netcdf atmos_month.198101-198112.aliq {
dimensions:
	time = UNLIMITED ; // (12 currently)
	pfull = 65 ;
	lat = 18 ;
	lon = 29 ;
	bnds = 2 ;
variables:
	float aliq(time, pfull, lat, lon) ;
		aliq:long_name = "Cloud fraction for large-scale liquid clouds" ;
		aliq:units = "dimensionless" ;
		aliq:_FillValue = -999.f ;
		aliq:missing_value = -999.f ;
		aliq:cell_methods = "time: mean" ;
		aliq:interp_method = "conserve_order2" ;
	double lat(lat) ;
		lat:standard_name = "latitude" ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_N" ;
		lat:axis = "Y" ;
		lat:bounds = "lat_bnds" ;
	double lat_bnds(lat, bnds) ;
	double lon(lon) ;
		lon:standard_name = "longitude" ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_E" ;
		lon:axis = "X" ;
		lon:bounds = "lon_bnds" ;
	double lon_bnds(lon, bnds) ;
	double pfull(pfull) ;
		pfull:standard_name = "air_pressure" ;
		pfull:long_name = "ref full pressure level" ;
		pfull:units = "mb" ;
		pfull:positive = "down" ;
		pfull:axis = "Z" ;
	double time(time) ;
		time:standard_name = "time" ;
		time:long_name = "time" ;
		time:bounds = "time_bnds" ;
		time:units = "days since 1979-01-01 00:00:00" ;
		time:calendar = "standard" ;
		time:axis = "T" ;
	double time_bnds(time, bnds) ;

// global attributes:
		:CDI = "Climate Data Interface version 2.4.4 (https://mpimet.mpg.de/cdi)" ;
		:Conventions = "CF-1.6" ;
		:title = "c96L65_am5f9d8r0_amip" ;
		:associated_files = "area: 19810101.grid_spec.nc" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
		:code_release_version = "2024.05" ;
		:git_hash = "5d306c05d9fe755cab04eedc8fd3de0d3c8355a0" ;
		:creationtime = "Mon Aug 11 19:59:00 2025" ;
		:hostname = "pp030" ;
		:history = "Mon Aug 11 16:17:05 2025: ncks -d lat,,,10 -d lon,,,10 atmos_month.198101-198112.aliq.nc reduced/atmos_month.198101-198112.aliq.nc\n",
			"Mon Aug 11 20:01:59 2025: cdo --history splitname 19810101.atmos_month.nc /home/Chris.Blanton/cylc-run/c96L65_am5f9d8r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run1/share/cycle/19810101T0000Z/split/regrid-xy/180_288.conserve_order2/19810101.atmos_month.\n",
			"fregrid --debug --standard_dimension --input_mosaic C96_mosaic.nc --input_dir /home/Chris.Blanton/cylc-run/c96L65_am5f9d8r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run1/share/cycle/19810101T0000Z/history/native --input_file 19810101.atmos_month --associated_file_dir /home/Chris.Blanton/cylc-run/c96L65_am5f9d8r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run1/share/cycle/19810101T0000Z/history/native --interp_method conserve_order2 --remap_file fregrid_remap_file_288_by_180.nc --nlon 288 --nlat 180 --scalar_field (**please see the field list in this file**) --output_file 19810101.atmos_month.nc" ;
		:CDO = "Climate Data Operators version 2.4.4 (https://mpimet.mpg.de/cdo)" ;
		:NCO = "netCDF Operators version 5.2.4 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco, Citation = 10.1016/j.envsoft.2008.03.004)" ;
data:

 aliq =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, -1.472766e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0.0006937876, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, -8.859464e-05, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0.007136224, 0.0001577576, 0, 0, 0, 0, 0, -1.934287e-05, 
    -9.565108e-07, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.872052e-05, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -4.39346e-05, -3.514404e-06, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -5.89307e-05, 0, 0, 3.978134e-06, 
    1.433759e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5.737614e-05, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, -1.724464e-07, 0.0120936, 0.0004463191, 0.000384264, 0, 0, 0, 0, 
    -8.537336e-06, 0.001258448, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -1.797572e-07, 0.001935643, 0.0003208703, 0, 0, 0,
  0, 0, -7.593926e-05, 0, 0.0001279515, 0, 0, 0, 0, 0, -5.277625e-05, 0, 0, 
    -6.375406e-05, -7.130552e-05, 0, 0, 0, 0, 0, 0, 0, 0, -4.231636e-07, 
    -3.574631e-10, -6.428992e-06, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0.0001190557, 0, 0, 0, 0.00031364, 0, -3.150605e-06, 
    1.414177e-05, 2.346066e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -7.097018e-06, 
    0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -5.039759e-05, 0.000228828, -3.142492e-06, 
    0, 0, 0.0002450024, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0.0004138202, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 9.926651e-05, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, -6.786352e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, -2.365432e-05, 0, -6.278254e-05, 0, 0,
  0, 0, -2.372363e-06, 0.02026818, 0.001227456, 0.001033425, -1.157516e-05, 
    0, 0, 0, -2.165174e-05, 0.003007225, -8.829799e-06, 0, 0, 0.0006000041, 
    -4.310576e-05, 6.075205e-06, 0, 0, 0, 0, 0, -5.392714e-07, 0.003088146, 
    0.0006935885, 0, 0, 0,
  0, 0, 3.441025e-06, 0, 0.0002308062, -3.376196e-05, 0, -0.000115214, 0, 0, 
    -9.187769e-05, 0, 0, -0.0001240168, -0.0001623784, 0.001692293, 0, 0, 0, 
    0, 0, 0, 0, -5.094277e-07, 0.0001457498, 0.0008252626, 0, 0, 0,
  0, 0, 0, 0, 0, -3.060938e-05, 0.0003255876, 0, 0, 1.243717e-05, 0.00166861, 
    0, 0.0006809267, 0.003407551, 0.002485566, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -4.001729e-06, -0.0001087688, 0, 0, 0,
  0, 0, 0, 0, 0, -2.305948e-05, 0, -6.103253e-06, 0, 0, -1.039713e-05, 
    0.0003604303, 0.0005862248, -1.226047e-05, 0, 0, 0.001640084, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0.003895391, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.001767339, 9.611149e-06, -1.21479e-05, 0, 0,
  0, 0, 0, 0, 0, 0, -9.331234e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0007865487, 
    0, -9.656748e-08, 0, 0, 0, 0, 0, 0.0001054962, -4.307667e-06, 
    0.0002252894, 0, 0,
  0, -3.13268e-05, -6.99511e-06, 0.0236889, 0.00157677, 0.004546942, 
    0.002003013, 0, 0, 0, -5.687013e-05, 0.00460363, -4.234822e-05, 
    0.0007572575, 0, 0.002668777, 0.0009593158, 0.0001680763, 0, 0, 0, 0, 0, 
    -5.972016e-06, 0.005633588, 0.002749736, 0, 0, 0,
  0, 0, 0.0005426285, -2.190082e-05, 0.0003485135, -7.051691e-05, 0, 
    -0.0002545489, 0, 0.0006650368, 0.0005717356, 0, -3.382835e-05, 
    -0.0002402301, 5.663486e-05, 0.002710611, -8.049917e-05, 0, 0, 0, 0, 0, 
    0, -1.328726e-05, 0.001382987, 0.00461814, 0, 0, 0,
  0, 0, 0, 0, 0, -9.29965e-05, 0.001354316, 0, -1.636023e-05, 0.0004603316, 
    0.003628717, 0, 0.005512783, 0.01574906, 0.01003844, -8.736784e-07, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.0001590806, -0.0002878008, 0, 0, 0,
  0, 0, 0, 0, 0, -8.11657e-05, 0, -4.174154e-05, 0, 0, -6.238277e-05, 
    0.001166105, 0.0008541506, -4.109742e-05, 0, -6.523454e-05, 0.002835321, 
    0, 0, 0, -1.421617e-05, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0.008343992, 0.0009114528, 0.001293845, 0, 0, 0, 0, 0, 0, 
    0.0001186547, 0, 0, 0, 0, 0, 0.0001673138, 0, 0, 0, 0, 0, 0.003162335, 
    0.001763347, 0.0002885991, 0, 0,
  0, 0, 0, 0, -7.451049e-05, -1.985206e-05, 0.005834769, 0, 0, 0, 0, 0, 
    0.000115252, 0, 0, -0.000195142, 0.004592948, -3.601257e-05, 
    -1.976732e-06, 0, 0, 0, 0, 0, 0.0002671952, -3.825757e-05, 0.00095856, 0, 0,
  0, 0.001403227, -8.484682e-06, 0.03453449, 0.004358964, 0.00992227, 
    0.00293378, 0, 0, 0, -0.0001001887, 0.01137423, 0.0002316539, 
    0.001314371, -2.042933e-05, 0.003830547, 0.001833382, 0.001799615, 
    0.001198491, 0, 0, 0, 0, -2.244666e-05, 0.01153202, 0.004415341, 
    -0.000113542, 0, 0,
  0, 0, 0.001012981, 4.447171e-05, 0.004288474, -4.104213e-06, 0.0003300337, 
    -0.0003901352, -1.499152e-05, 0.00300333, 0.001408786, 0, 8.265091e-06, 
    -0.0004672056, 0.002186738, 0.004287825, 0.0004291568, 0, 0, 0, 0, 0, 0, 
    -4.750135e-05, 0.003624529, 0.006640737, 0, 0, 0,
  0, 0, 0, 0, 0, 0.0004759502, 0.005797949, 6.639506e-06, 0.0004267685, 
    0.003989522, 0.01056721, 0.00042667, 0.008837565, 0.03232576, 0.01561988, 
    6.585116e-07, 0, 0, 0, 0, 0, 0, 0, 0, 0.0005661941, 0.001399894, 
    -1.689127e-05, 0, 0,
  0, 0, 0, 0, 0, -0.0002123437, 0, -0.0001803223, 0, 0, -0.0001724206, 
    0.002401567, 0.004640458, -5.344467e-05, -4.441674e-07, -0.0002618187, 
    0.006661501, -3.703219e-05, 0, -0.0001269492, 0.001463384, 0, 0, 0, 0, 0, 
    0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -9.211511e-06, -1.177576e-05, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, -3.316615e-05, 0, 0,
  0, 0, 0, 0.01310097, 0.0113409, 0.008312942, -3.819955e-05, 0.002299483, 0, 
    0.0001201431, 0, 0, 0.005629091, 0.000388413, 0, 0, 0, 0, 0.003485399, 0, 
    0, 0, 0, 0, 0.005253637, 0.004673911, 0.003746452, -7.115138e-06, 0,
  0, 0, -1.917401e-05, 0, 0.0004353519, -0.0006069292, 0.01200313, 0, 0, 0, 
    0, 0, 0.0004212857, 0, 0, 0.001695487, 0.006106403, -0.0001219719, 
    -2.134405e-05, 0, 0, 0, 0, 0, 0.001110418, 0.001039847, 0.00417747, 0, 0,
  0, 0.003336641, -8.73846e-05, 0.04866827, 0.01341496, 0.01768745, 
    0.009253288, 0, 0, 0, 0.0005603529, 0.02351537, 0.004446823, 0.001463429, 
    0.001500841, 0.0128781, 0.007622715, 0.006022552, 0.005467784, 0, 0, 0, 
    0, -3.825188e-05, 0.01888363, 0.005431178, 0.0002662464, 0, 0,
  0, 0.0004644131, 0.003997237, 0.00025983, 0.00791211, 0.0004561273, 
    0.001968146, -0.0003264459, -0.0001421912, 0.01134325, 0.003345656, 
    0.0007105229, 0.0004461732, 0.0007172734, 0.008137452, 0.004958616, 
    0.001935303, 0, 0, 0, 0, 0, 0, -8.124049e-05, 0.005854319, 0.0110364, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0.004009644, 0.01566105, 0.0004899393, 0.003861605, 
    0.01121365, 0.01817426, 0.001457157, 0.01399198, 0.05014511, 0.02152356, 
    1.913014e-08, 0, -4.807275e-05, 0, 0, -8.936544e-07, 0, 0, 0.0003648845, 
    0.0006408141, 0.007684371, 0.003400384, 0, 0,
  0, 0, 0, 0, -3.401454e-06, -0.000113326, 0, -0.0004218694, 0, 0, 
    0.0009016446, 0.005724819, 0.005649653, -0.0001322669, -3.154476e-05, 
    0.0004898475, 0.01676273, -0.0001559818, 0, -0.0002728934, 0.009169892, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    9.353714e-05, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -7.071937e-07, 0, 
    0.001158037, 0, -3.504581e-05, 0, 0, 0, 0, -4.404982e-06, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0.004774701, -1.19835e-05, 0.00380255, 0.00187045, 0, 0, 0, 
    0, 0.002683101, 0.002026333, 7.519333e-05, 0, 0, 0, 0.001508933, 0, 
    -1.266803e-06, 0, 0, 0, -3.671107e-05, 0.002388553, 0.0002982862, 0,
  0, 0, 0, 0.02100735, 0.01735664, 0.01312139, -0.0001526283, 0.004565664, 0, 
    0.003242472, 0, 0, 0.01192366, 0.003227046, 0, 2.374666e-06, 0.001054564, 
    -1.077092e-06, 0.02122932, -2.061595e-05, 0, -1.078302e-05, 0, 0, 
    0.0103673, 0.0146275, 0.01618539, -0.0001100378, 2.404269e-05,
  0, 0, 3.002381e-05, 0.001461118, 0.008869933, 0.007403553, 0.02098964, 0, 
    0, 1.301702e-08, 0, -8.715606e-07, 0.007065765, -3.282185e-05, 0, 
    0.009343321, 0.01208156, 0.0001330633, 0.001982456, 0, 0, 0, 0, 0, 
    0.01161033, 0.01175133, 0.01746604, 0, 0,
  0, 0.006143352, 0.0007313354, 0.05984046, 0.03555498, 0.02079896, 
    0.02284367, -7.635032e-06, 0, 0.0002540428, 0.003502957, 0.05029972, 
    0.01701766, 0.005044236, 0.005081624, 0.03010322, 0.02448489, 0.01708013, 
    0.009266905, 0, 0, 0, 0, -0.0001217416, 0.03976383, 0.00826327, 
    0.003242386, 0, 0,
  0, 0.001784364, 0.005794324, 0.003403245, 0.02349189, 0.0009982365, 
    0.002903386, 0.002972277, 0.00218567, 0.02231615, 0.007534591, 
    0.003360709, 0.00304671, 0.009635886, 0.02047818, 0.005892657, 
    0.01063241, 6.743719e-05, 0, 0, 0, 0, 0, 0.0003418043, 0.008788079, 
    0.02900005, 0, 0, 0,
  0, 0, 0, 0, 0, 0.01700131, 0.04441232, 0.003796361, 0.005545372, 
    0.02142588, 0.02897047, 0.003228472, 0.02145994, 0.08135524, 0.03402657, 
    6.169694e-06, 0, 0.0001234066, 0, 0, 0.0009081399, 0, -6.254966e-06, 
    0.001741957, 0.0004856199, 0.0199373, 0.009567134, 0, 0,
  0, 0, 0, 0, -0.00010417, 0.0006322098, 0, -2.473929e-05, 0, -8.667788e-06, 
    0.008576692, 0.01077471, 0.008941866, -0.0005190152, -0.0001739135, 
    0.00323487, 0.02698927, 0.004875037, 0, 0.001490941, 0.02245595, 0, 0, 0, 
    0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2.127526e-05, -3.142502e-05, 0, 0, 0, 
    -2.669262e-09, 0, 0, 0, 0, 0, 0, 0, 0.0008783058, -3.694812e-05, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.649374e-05, -2.430194e-06, 
    -4.385501e-09, 0, 0, 0.0008822044, 9.831617e-05, 0.005540906, 0, 
    0.00178945, 0, 0, 0, 0, -9.322792e-05, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001049165, 0.0005638892, 0, 
    -1.840591e-05, 0, 0, 0, 0.0006953641, -6.707195e-06, 0.001338171, 
    0.0002594438, -5.350614e-05, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -5.272202e-06, 0, 0, 0, 
    0, 0, 0, 0.0004015631, 0, -2.615859e-05, 0.0001054159, -1.208865e-05,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.040673e-09, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, -9.118078e-05, -2.862776e-05, 1.306333e-05, 0, 
    -7.512318e-10, 0, -3.250487e-05, 0, -8.689047e-05, 7.855488e-06, 0, 0, 0, 
    0, 0, 0, -2.173987e-05, 0, 0, 0, 0, 0, 0,
  0.003775821, 0, -2.239995e-06, 0, -4.741815e-06, 0.01232739, 2.637732e-05, 
    0.004316423, 0.004000438, -2.595611e-06, 0, 0, -1.825239e-05, 0.0186237, 
    0.003556376, 0.002584276, 0, 0, 0, 0.005272747, 0, 0.0004052112, 
    -7.469972e-05, 0, -3.478156e-08, 0.002142431, 0.005364846, 0.002797511, 
    0.002836286,
  -5.334283e-06, -1.826933e-05, 0, 0.02694618, 0.02094475, 0.01834189, 
    0.001727972, 0.005279781, -2.736284e-06, 0.005596489, -2.825068e-05, 
    0.0004777173, 0.0205015, 0.005086138, 0, 0.001584998, 0.008235758, 
    0.0002561485, 0.06829759, 0.0006783222, 0.0004776812, 0.0006316987, 0, 
    -1.312442e-05, 0.02246925, 0.03014934, 0.0353287, 0.0009351861, 
    0.000275635,
  0, -1.352292e-06, 0.001603873, 0.007447989, 0.02280378, 0.07205676, 
    0.02988904, 0.0001091174, -4.62637e-06, -7.178189e-07, 2.687274e-05, 
    -2.358455e-05, 0.01515508, -6.060786e-05, -1.313307e-08, 0.03102387, 
    0.01514308, 0.00530847, 0.02190731, -4.155102e-09, 0, 0, 0, 0, 
    0.02218226, 0.02987109, 0.0496699, -3.542416e-05, 0,
  0, 0.01121925, 0.006431811, 0.07661239, 0.0649745, 0.04699265, 0.05050655, 
    -0.0001294541, 0, 0.001744354, 0.01646071, 0.0954833, 0.04505311, 
    0.01290233, 0.01301502, 0.04069638, 0.04465448, 0.03302772, 0.01462508, 
    0, 0, -6.829149e-09, 0, 0.001181193, 0.09484513, 0.01063593, 0.005805835, 
    7.563836e-10, 0,
  0, 0.003969773, 0.01510022, 0.007269879, 0.0512012, 0.002195695, 0.0105931, 
    0.008038105, 0.004543005, 0.04208327, 0.01480628, 0.0151896, 0.01668875, 
    0.04126342, 0.05815561, 0.009954067, 0.02278836, 0.0001475489, 0, 0, 0, 
    0, 0, 0.0140139, 0.03353172, 0.05121136, -3.224164e-05, 0, 0,
  0, 0, -5.095349e-08, 2.592755e-06, -1.143332e-05, 0.04551544, 0.07753197, 
    0.005418638, 0.01613259, 0.03479406, 0.04395759, 0.01306514, 0.05413692, 
    0.1218652, 0.04281069, 0.0005317921, -3.610844e-08, 0.003343555, 0, 
    -7.224759e-08, 0.004774262, 0, 0.0008740409, 0.003295067, 0.001769906, 
    0.03619261, 0.01892219, 0, 0,
  -7.438752e-10, 0, 0, 0, 0.002047405, 0.006390009, -1.494058e-05, 
    0.003285361, -1.027751e-09, 3.151296e-05, 0.02385082, 0.04320751, 
    0.02195149, -0.0006354773, 0.000285962, 0.005662038, 0.04372184, 
    0.0148491, -1.353741e-06, 0.01031053, 0.04346411, 0, 0, -2.953643e-06, 0, 
    -2.564089e-08, -1.839989e-08, -3.865485e-07, -2.838055e-07,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.341348e-08, 0.001455614, 0.000851315, 0, 
    0, -1.080794e-10, 5.755079e-05, 0.002132244, 0.0004081314, -4.458086e-05, 
    0.002542594, 0, -0.000167908, 0, 0.005294443, 0.0001363259, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -9.036691e-05, -3.328565e-05, 
    -7.346646e-08, 1.197493e-07, 0.0005240929, 0.003682107, 0.01167168, 
    0.005919587, -1.748958e-06, 0.004428219, 0, 0, 0, 0, -0.0002594323, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -3.876234e-05, 0, 0.0006380586, 
    0.004068388, 0.002441155, 0.002266529, 0.001557072, 0, 0, -1.426018e-05, 
    0.00289713, 0.001061005, 0.005171843, 0.003322755, 0.001774215, 
    -1.745764e-05, 0,
  9.268554e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0009990215, 
    0.002678119, -2.575988e-05, 0, 0, 0, 0, -7.342242e-05, 0.002103144, 0, 
    0.0002865368, 0.002270219, 0.0007227496,
  0, -2.028044e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, -8.975259e-06, 0.002104853, 0.003172275, 0.003435694, 
    2.659268e-09, 5.122827e-05, 0, 0.001047963, -5.432886e-05, 0.0007983134, 
    0.0005218203, -0.000179285, 3.456122e-06, 0, 0, 0, 0, -6.00745e-05, 
    -5.712815e-05, 9.826575e-06, 0, 0, 0, 0,
  0.01203215, 0.000356448, -1.490361e-05, 0.0002766738, -0.0001308635, 
    0.03169787, 0.007034674, 0.006495763, 0.005613881, 0.004639222, 
    3.42595e-08, 0, 0.001159279, 0.04801995, 0.01020103, 0.006529465, 0, 
    -4.695986e-06, 0.002339396, 0.01804963, 0.009131851, 0.001015495, 
    0.00148378, 9.653436e-06, -4.743964e-06, 0.005902924, 0.009826377, 
    0.01431904, 0.018087,
  -8.331646e-05, 0.002215663, 7.709112e-06, 0.03446693, 0.03018813, 
    0.02567615, 0.01072633, 0.0071927, -0.0001791763, 0.007321812, 
    0.001395558, 0.003904324, 0.03796054, 0.01160851, 0.003465195, 
    0.006279265, 0.01488165, 0.006281551, 0.1125222, 0.01073406, 0.003152344, 
    0.001278707, 0.002227412, -3.601648e-05, 0.03464513, 0.05093595, 
    0.07314702, 0.01118767, 0.001656536,
  8.021953e-10, 5.515552e-05, 0.00773015, 0.02649207, 0.04847687, 0.1279398, 
    0.04291745, -8.277635e-05, 0.0006490864, 0.001627349, 0.001072384, 
    0.001208221, 0.02811266, 0.002607381, -6.915052e-05, 0.05470745, 
    0.0215055, 0.03141592, 0.07769007, 9.240015e-05, -6.978538e-05, 0, 0, 
    0.0001192944, 0.04283146, 0.05319962, 0.09754746, 0.0003053289, 
    -2.746952e-05,
  -7.7116e-07, 0.03146377, 0.03455766, 0.1544031, 0.1233964, 0.1575836, 
    0.106167, 0.005106352, -8.351501e-06, 0.008904575, 0.1267895, 0.1790003, 
    0.1619013, 0.0392766, 0.06831612, 0.1503412, 0.08413578, 0.05913828, 
    0.02074838, 0, -1.360808e-09, 0.0005420878, -7.794224e-09, 0.08319446, 
    0.2942149, 0.02112926, 0.008217817, -1.39316e-06, -1.669656e-08,
  3.108985e-07, 0.004647116, 0.02970248, 0.03458147, 0.1025682, 0.0368831, 
    0.04646416, 0.01619126, 0.01362201, 0.2177871, 0.08691826, 0.1430999, 
    0.1742764, 0.182881, 0.1853265, 0.06715754, 0.04165149, 0.0001535261, 
    0.0002740034, 7.592602e-05, 0, 0, 0.0002936813, 0.09904308, 0.1640193, 
    0.1055483, 0.002139203, -8.472322e-05, -1.993498e-08,
  -4.150072e-07, 7.201622e-07, 0.0001180591, -7.024221e-06, 1.120684e-05, 
    0.07106906, 0.1296269, 0.02811882, 0.05125472, 0.09627852, 0.1222451, 
    0.220801, 0.2057013, 0.2257328, 0.07554416, 0.004730452, 7.900484e-06, 
    0.01425083, 2.698982e-05, -1.805309e-06, 0.009530252, 4.190802e-08, 
    0.00829498, 0.01707816, 0.01335725, 0.06451581, 0.02761064, 0.0009765837, 
    3.679689e-07,
  -1.985681e-07, 0, 3.131167e-06, 0, 0.003781159, 0.01453479, 0.001177786, 
    0.01798749, -5.819021e-06, 0.005603249, 0.0759339, 0.1077302, 0.1009812, 
    0.02103982, 0.01314709, 0.007230566, 0.05550738, 0.02587015, 0.002457242, 
    0.02176694, 0.06045169, -2.277951e-07, -1.419884e-06, -2.230744e-05, 
    -4.096269e-06, 0.0009141212, 3.773435e-05, 0.0005696948, 0.0003007717,
  0, 0, 0, 2.866587e-08, 0, -2.904148e-08, -8.263175e-08, -3.621132e-08, 
    5.12783e-09, 2.566236e-07, 2.166035e-05, 0.02842462, 0.02638166, 
    1.155001e-05, 6.692876e-08, 9.485501e-07, 0.005562369, 0.01387784, 
    0.009669516, 0.00367193, 0.009627955, -4.769392e-06, 0.003124028, 0, 
    0.008080781, 0.004392048, 0, 9.655383e-05, -1.894124e-06,
  0, 0, 0, 0, 0, -4.571862e-11, 0, 0, 0, 8.890161e-09, 7.810972e-09, 
    -0.000125783, 0.0005833131, -1.405138e-05, 0.0001223563, 0.01456002, 
    0.009783264, 0.05007845, 0.01098977, -7.368993e-05, 0.009603413, 
    -0.0002157454, 0.001773418, -2.169592e-05, 0.000178539, 0.002824774, 
    4.155655e-06, 0, 0,
  4.641454e-06, 0, 0, 0.0001209519, 0, 0.0001787238, 0, 0, 0, 0, 0, 
    -8.56643e-06, 0.0001787818, 3.022761e-06, 0.004278152, 0.01154316, 
    0.007354361, 0.01752597, 0.003757715, 0.001002582, 0, 0.001224974, 
    0.009688654, 0.007463632, 0.007592422, 0.02096287, 0.01708155, 
    0.002217557, 0,
  5.802617e-05, 0.0004680644, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.004552902, 0.004125135, 0.0008484893, 0, 0, 0, 0, -4.260655e-05, 
    0.007463396, -6.264427e-05, 0.0003077422, 0.005571609, 0.00609199,
  0, 0.00268936, -4.224376e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.336789e-05,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.231614e-09, -3.926427e-11, 0, 0, 0, -0.0001310068, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0.006773925, 0.02454262, 0.02474549, 0.01574767, 
    0.0006204383, 0.001564584, 0, 0.003872872, 0.001059093, 0.01903298, 
    0.006157985, 0.001747728, 0.002719917, 0, 0, 0, 0, 0.003918799, 
    0.002132919, 0.004243432, 0.000688815, -5.068947e-05, 0.001751286, 
    0.0009734884,
  0.02254268, 0.002512562, 2.584921e-05, 0.001796013, 0.00685026, 0.06218086, 
    0.03809151, 0.04601912, 0.01728846, 0.02370491, 0.002097689, 
    5.374186e-06, 0.006668529, 0.09200621, 0.04171348, 0.02183605, 
    0.01722821, 0.01429236, 0.006543625, 0.02544905, 0.04640838, 0.009328437, 
    0.01656695, 0.003412892, 0.002624061, 0.01245155, 0.01318641, 0.02665683, 
    0.02475643,
  0.005604093, 0.01215185, 0.01150751, 0.04630484, 0.03876365, 0.06205237, 
    0.02831501, 0.02249293, 0.00335013, 0.02121203, 0.03091356, 0.01861826, 
    0.06477618, 0.05330922, 0.007639065, 0.01636259, 0.02318224, 0.01358438, 
    0.1835824, 0.06254981, 0.02876352, 0.00522513, 0.005568639, 
    -5.420125e-05, 0.04681161, 0.07642047, 0.1197054, 0.08468258, 0.02670659,
  0.003892707, 0.008996943, 0.05713688, 0.06100444, 0.07841541, 0.1905846, 
    0.1066078, 0.05093957, 0.03899869, 0.01086302, 0.009374445, 0.0303454, 
    0.06899671, 0.06104574, 0.0541306, 0.08958953, 0.1177155, 0.1823837, 
    0.2757882, 0.02377033, 0.0001422885, -1.198575e-06, 8.195287e-07, 
    0.009290141, 0.09612636, 0.1946311, 0.2336903, 0.02939088, 0.00185796,
  0.005244854, 0.157799, 0.1962769, 0.1608305, 0.1177836, 0.2347573, 
    0.1690866, 0.01811129, 7.298877e-07, 0.006007098, 0.1602535, 0.1934121, 
    0.163162, 0.1226345, 0.1276545, 0.1833818, 0.2057683, 0.1609031, 
    0.1316695, 2.194121e-05, 0.0002174145, 0.0004127744, 0.01763044, 
    0.1030342, 0.2899089, 0.1631083, 0.09690564, 0.0199775, 0.01257749,
  1.732021e-06, 0.0294521, 0.4153571, 0.1879035, 0.2654786, 0.1299326, 
    0.1292371, 0.03508735, 0.03253857, 0.241343, 0.09117135, 0.125832, 
    0.1377777, 0.1569574, 0.1716778, 0.07176399, 0.07606979, 0.009831319, 
    0.03362156, 0.004039351, -1.943716e-05, 2.236618e-05, 0.02601274, 
    0.432949, 0.3414966, 0.3074886, 0.1107134, 0.01527612, 0.02257853,
  3.993801e-05, 0.0005071213, 0.01022552, 0.03070433, 0.07563778, 0.2190185, 
    0.2386861, 0.1792135, 0.2008659, 0.3385437, 0.1920212, 0.2593484, 
    0.1841837, 0.1829828, 0.08361938, 0.008722214, 3.52209e-05, 0.0104471, 
    0.01116161, -3.127459e-06, 0.01196881, 3.251772e-05, 0.01662351, 
    0.2940246, 0.3031207, 0.3114732, 0.1200387, 0.02404417, 0.0300636,
  0.000129922, 4.457946e-07, 0.0001003385, -5.933606e-06, 0.006644789, 
    0.04661812, 0.008373838, 0.04889345, 0.002353814, 0.05471371, 0.09296131, 
    0.1038937, 0.08123355, 0.01340003, 0.003927086, 0.02368852, 0.09301914, 
    0.04387987, 0.0312519, 0.1282623, 0.1364271, 0.00945678, 0.0007176852, 
    0.002816236, 8.417852e-05, 0.001365092, 0.006111573, 0.03113176, 
    0.002196635,
  0.001333827, -3.228941e-07, -2.797852e-09, 2.443535e-06, 2.925046e-05, 
    5.723219e-05, -2.254877e-06, 2.418391e-06, 4.635017e-06, 1.068571e-05, 
    0.0004421529, 0.02510022, 0.027534, -5.337135e-06, 3.076015e-08, 
    0.0003139854, 0.02552854, 0.0739129, 0.02702237, 0.02876778, 0.1710181, 
    0.0004290416, 0.01725524, -2.959908e-08, 0.01526706, 0.01363989, 
    -0.0002720555, 0.004587225, 0.0002284737,
  0, 0, -2.623557e-08, 0.0001191761, -7.282798e-10, 1.94753e-08, 
    5.132816e-06, 0, 0, -7.502568e-07, -3.467864e-07, 0.0001982915, 
    0.004862449, -0.0002087023, 0.006929643, 0.02550044, 0.0196723, 
    0.09248762, 0.02064144, 0.002988294, 0.0198727, 0.01501345, 0.004087123, 
    0.0009846182, 0.0008984674, 0.01025091, 0.001036443, 0, 0.0003575785,
  0.00556625, 1.407152e-05, 1.905069e-07, 0.0008840006, -0.0002714233, 
    0.001420512, 0, 0, 0, 0, 0, 0.002816436, 0.002185069, 0.000507538, 
    0.009313163, 0.02219998, 0.04840734, 0.03671532, 0.009859761, 
    0.003340215, -1.604962e-05, 0.005522246, 0.01643788, 0.01940546, 
    0.01584872, 0.06067151, 0.04946744, 0.005147845, 0,
  0.004232762, 0.002517835, 0.0001874412, -8.842124e-06, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, -0.0001085819, 0.01212902, 0.008109676, 0.004188624, 
    0.001031322, 9.798616e-06, 0, 0, 0.00159343, 0.009409712, 0.001983877, 
    0.0006337698, 0.01395968, 0.01602577,
  0.00133043, 0.004802465, 2.395793e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, -1.079624e-05, 0, 0, 0, 0, 0, 0, 0, -6.747637e-05, 0, 
    -1.243259e-05, 0.0009709443,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4.685735e-06, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, -3.712872e-06, -0.0001236117, -1.517668e-05, 0, 0, 0, 
    0.0009781772, 0.0007444242, -5.68851e-06, -6.884235e-05, -6.606482e-09, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0.001381248, 0, 0, -1.76293e-06, -5.522649e-09, 0.01526785, 0.04046519, 
    0.03671639, 0.03522722, 0.0172668, 0.003389082, -1.716411e-06, 
    0.007210842, 0.00508914, 0.05864865, 0.06060015, 0.0441196, 0.01518574, 
    5.510731e-07, -2.333996e-05, 0, -1.658519e-05, 0.008843338, 0.01147432, 
    0.005753796, 0.002409897, 0.0009110237, 0.00320268, 0.002478006,
  0.05682894, 0.01038677, 0.01273028, 0.03727345, 0.07935446, 0.09614035, 
    0.07237422, 0.06077516, 0.05093296, 0.04517907, 0.009862567, 
    0.0008899994, 0.02388245, 0.1770928, 0.1195334, 0.08483155, 0.05703197, 
    0.04913766, 0.03640194, 0.0501197, 0.09714194, 0.06691672, 0.05036891, 
    0.01776046, 0.007336917, 0.02582597, 0.02878914, 0.06264652, 0.08298013,
  0.03870872, 0.03644352, 0.03789353, 0.07593803, 0.05897193, 0.06428856, 
    0.04390886, 0.05296196, 0.08360235, 0.05159455, 0.06235039, 0.07587483, 
    0.1348288, 0.09414775, 0.06795686, 0.03527344, 0.1036795, 0.02764825, 
    0.2051809, 0.1627643, 0.06200589, 0.0465758, 0.05545735, 0.002497717, 
    0.06970222, 0.1077221, 0.1713175, 0.1603874, 0.1080052,
  0.003035873, 0.00886144, 0.07230106, 0.05442462, 0.0908476, 0.2305381, 
    0.1406468, 0.05917778, 0.04042524, 0.01363621, 0.04148106, 0.05604595, 
    0.09716136, 0.09020898, 0.05514388, 0.1286359, 0.112733, 0.1888221, 
    0.3242805, 0.0553594, 0.08781893, 0.01270689, -2.567565e-06, 0.01161106, 
    0.09637916, 0.1930626, 0.2751842, 0.06988736, 0.02603749,
  0.001602846, 0.1202938, 0.1567702, 0.1385624, 0.1033709, 0.1916392, 
    0.1388915, 0.01406421, 3.326378e-05, 0.005435197, 0.1509505, 0.1726616, 
    0.1412539, 0.07840252, 0.1082394, 0.1576535, 0.1578987, 0.1518383, 
    0.09801902, 0.03300954, 0.004367235, 3.26806e-06, 0.002886835, 
    0.07482085, 0.2601114, 0.1320114, 0.06213473, 0.02395083, 0.04653858,
  1.894973e-07, 0.02285075, 0.353305, 0.1359638, 0.2389819, 0.08634994, 
    0.08801851, 0.02816044, 0.02382492, 0.2165867, 0.07064032, 0.09355163, 
    0.08961657, 0.1270129, 0.1517441, 0.05020826, 0.07314952, 0.001443896, 
    0.03189474, 0.01923367, -5.292174e-05, 5.607643e-06, 0.01039429, 
    0.3908093, 0.2832932, 0.2758065, 0.08675138, 0.01419431, 0.01942129,
  9.131953e-05, 5.564308e-05, 0.0006053066, 0.02475976, 0.04251753, 
    0.1512281, 0.2296216, 0.1470839, 0.1497067, 0.2816469, 0.1605553, 
    0.19729, 0.1504738, 0.1587718, 0.07359811, 0.006064822, 1.275454e-05, 
    0.002300295, 0.000520304, 4.133948e-05, 0.01194321, 0.0001600141, 
    0.01180269, 0.1688883, 0.2436138, 0.2696271, 0.08280738, 0.03963266, 
    0.0264168,
  0.01350747, 5.60606e-08, 1.55568e-05, 2.02413e-05, 0.001788685, 0.02603629, 
    0.007310153, 0.03887458, 0.001218633, 0.04009973, 0.07901103, 0.07765058, 
    0.05869503, 0.004328528, 0.0006292803, 0.01903849, 0.08586059, 
    0.03821492, 0.01721424, 0.08683626, 0.1054842, 0.003756811, 0.0005173651, 
    0.001507455, 0.0003327856, 0.0001497095, 0.01013199, 0.0870407, 0.131944,
  0.2713069, -0.0002243583, 1.280098e-06, 3.614755e-07, 3.370392e-06, 
    8.681436e-06, -8.689428e-07, 6.304266e-07, 1.86426e-06, 6.040432e-06, 
    4.154801e-05, 0.02005694, 0.02474599, 3.31491e-05, 1.637883e-07, 
    0.0001639732, 0.06658026, 0.1326862, 0.04535594, 0.1244272, 0.1740091, 
    -0.00031894, 0.01299589, -0.0001522736, 0.04882473, 0.02887307, 
    0.004299774, 0.04538925, 0.1513913,
  0.0001312322, 0.01250198, -1.252331e-06, 0.001834659, -1.252957e-07, 
    1.582094e-07, 7.188086e-06, 0, -1.819207e-11, 0.000134319, 0.0003284685, 
    0.001496926, 0.02667378, 0.001702915, 0.02641468, 0.04412932, 0.04012486, 
    0.1796153, 0.08495101, 0.02944921, 0.03800171, 0.08329735, 0.05283988, 
    0.06281251, 0.06777333, 0.05545194, 0.03410217, 0.0007438951, 0.002385894,
  0.01054885, 0.00143114, 0.0006953864, 0.003121686, 0.0003941773, 
    0.002272293, 0, 0, 0, 0, 0, 0.003888419, 0.01006362, 0.0067644, 
    0.0221287, 0.05594184, 0.1159491, 0.06468219, 0.04376764, 0.01038661, 
    -9.407415e-05, 0.01309516, 0.0446574, 0.0456784, 0.02980464, 0.08720861, 
    0.1106383, 0.03538521, 5.019725e-05,
  0.01802394, 0.00499346, 0.005552012, -1.955189e-05, -1.23467e-05, 0, 0, 0, 
    0, 0, 0, 0, 0, -9.839135e-06, -5.824923e-05, 0.001065996, 0.02340906, 
    0.01661674, 0.019673, 0.001616357, 0.0007233225, 0, 0, 0.003224134, 
    0.01391889, 0.005158602, 0.01180112, 0.04027255, 0.04188689,
  0.007831194, 0.006301747, 0.001224648, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -5.725734e-07, 2.133233e-06, -3.676295e-05, 5.285657e-05, 0.0001073314, 
    0, 0, 0, 0, 0, -1.3032e-05, 0.000334684, 0.0003530348, -0.0001637208, 
    0.005553123,
  0, -2.387045e-05, -9.292571e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -6.09016e-05, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001460483, -0.000204613, 
    -8.684158e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, -2.094802e-05, 0.001519886, -0.0001740563, -2.1403e-12, 
    0, -1.781093e-05, 0.005728921, 0.01569007, 0.0181354, 0.01178518, 
    0.009848853, 0.001863858, -2.117054e-06, 0, 0.009749125, 0, 0, 0, 0, 0, 
    0, 0, 0,
  0.01022074, 0.01269521, 0.005026861, -1.095647e-05, -3.072524e-07, 
    0.02331711, 0.05603605, 0.07069675, 0.08730489, 0.03998548, 0.009699055, 
    4.926926e-05, 0.01251665, 0.03465175, 0.09863457, 0.08310396, 0.09449287, 
    0.03847938, 0.02284629, 0.006715277, 0.02165268, 0.02125505, 0.02464789, 
    0.04275549, 0.0652453, 0.07321236, 0.03765222, 0.03016854, 0.02413306,
  0.1269676, 0.08031644, 0.073892, 0.0994412, 0.1502282, 0.1527813, 
    0.09952842, 0.08853927, 0.127405, 0.09793165, 0.04997296, 0.04886565, 
    0.09996824, 0.2422149, 0.1556107, 0.1445504, 0.09704566, 0.09310381, 
    0.09809729, 0.1120852, 0.1306096, 0.1384097, 0.211778, 0.07954045, 
    0.05191074, 0.08001195, 0.08197767, 0.08937176, 0.1347069,
  0.04189242, 0.033982, 0.04329761, 0.09446825, 0.06266331, 0.09292472, 
    0.06365192, 0.07452529, 0.08134088, 0.0605134, 0.08505106, 0.1117512, 
    0.1436067, 0.1174195, 0.09294804, 0.0431013, 0.1073072, 0.07026164, 
    0.2205248, 0.1728635, 0.05896817, 0.1217533, 0.07619336, 0.02749366, 
    0.09697272, 0.1352549, 0.1740222, 0.1502117, 0.09884398,
  0.009696648, 0.002812177, 0.05128835, 0.03464642, 0.08066268, 0.2220096, 
    0.1208763, 0.05378814, 0.02733734, 0.01702301, 0.03878348, 0.05879448, 
    0.1027803, 0.07649504, 0.04109647, 0.1001351, 0.08808511, 0.1631047, 
    0.3191808, 0.04152419, 0.06462161, 0.006586591, 2.999495e-07, 0.02995723, 
    0.09073683, 0.1725192, 0.2395412, 0.05554786, 0.01065589,
  0.005420617, 0.0880663, 0.136735, 0.1303135, 0.1089723, 0.1586128, 
    0.1260691, 0.009085932, 1.685743e-05, 0.005847581, 0.1570206, 0.1835489, 
    0.1351256, 0.05483442, 0.08166556, 0.1497566, 0.1459492, 0.1442186, 
    0.07672188, 0.0104646, 1.694625e-06, 0.000222966, 5.114722e-05, 
    0.05439366, 0.2322351, 0.1094015, 0.03403975, 0.02479054, 0.008197327,
  6.808895e-08, 0.02535148, 0.2646917, 0.1186356, 0.2080935, 0.06774958, 
    0.06832162, 0.02725734, 0.02105001, 0.1874036, 0.0636135, 0.07553228, 
    0.07025775, 0.1095785, 0.1513138, 0.04581213, 0.07369271, 0.001340589, 
    0.01209441, 0.008264643, -5.105408e-07, 1.937825e-06, 0.002827353, 
    0.3711676, 0.2520883, 0.2565442, 0.04615155, 0.01547611, 0.00335645,
  6.026412e-05, 1.963943e-05, 0.000399277, 0.005000314, 0.0118175, 0.1127477, 
    0.2194472, 0.122358, 0.1330753, 0.2650694, 0.1472185, 0.1590682, 
    0.1377315, 0.1470838, 0.07035638, 0.007708883, 1.530057e-05, 
    0.0003415324, 2.494443e-05, 6.744125e-05, 0.01735901, 2.560536e-05, 
    0.01305908, 0.1209204, 0.2056924, 0.2392277, 0.07114813, 0.04372857, 
    0.008855509,
  0.007856682, -1.603627e-09, 2.364574e-06, 0.0001055578, 0.001208425, 
    0.01557906, 0.002371991, 0.02814403, 0.002002514, 0.0324077, 0.07326768, 
    0.06894633, 0.0479339, 0.0003519482, 0.0004083498, 0.01336661, 
    0.06814043, 0.04419138, 0.02065844, 0.05623014, 0.095368, 0.003437769, 
    0.0003951395, 0.0009220954, 0.0004790583, 0.004091548, 0.020743, 
    0.1143657, 0.1050831,
  0.1487075, 7.452771e-05, 7.77734e-07, -3.085108e-08, 4.057503e-07, 
    1.764201e-06, 1.545318e-06, 5.688393e-07, 7.64127e-07, 4.636297e-06, 
    7.32375e-05, 0.01495505, 0.01433455, 3.112302e-06, 7.855795e-07, 
    0.001142776, 0.07951406, 0.1127469, 0.03876263, 0.1298463, 0.1048169, 
    -0.0002068371, 0.01095952, -6.09591e-06, 0.03329638, 0.04428667, 
    0.01714558, 0.05088494, 0.1956146,
  0.05579667, 0.03361699, -0.0001984141, 0.001193334, 3.44128e-05, 
    2.282449e-07, 0.0006406457, 0, -1.330619e-10, 0.004159353, 0.008033542, 
    0.01642848, 0.04457306, 0.02130838, 0.05409827, 0.06638233, 0.06017192, 
    0.2160651, 0.1023291, 0.07281277, 0.09501536, 0.1028052, 0.05428482, 
    0.04937416, 0.04284739, 0.09702241, 0.09782062, 0.03829809, 0.05806496,
  0.01902692, 0.007138094, 0.007428088, 0.01944833, 0.010147, 0.004071186, 
    -1.016489e-05, 0, 0, 0, -2.30073e-05, 0.00640501, 0.01287309, 0.02177551, 
    0.03922687, 0.09148255, 0.2119401, 0.1240914, 0.1041128, 0.04235707, 
    0.003852593, 0.04275132, 0.1185368, 0.1154409, 0.1010627, 0.1485993, 
    0.2099515, 0.178936, 0.02799852,
  0.07317155, 0.01184026, 0.0161658, 0.000725739, 0.00128419, 0, 0, 0, 0, 0, 
    0, 0, -3.295198e-05, 0.0001572819, 0.00915064, 0.00794714, 0.07325523, 
    0.08709042, 0.0398738, 0.003510793, 0.003421257, -6.318767e-06, 
    0.0005030842, 0.008165153, 0.02810503, 0.01539928, 0.04325801, 
    0.09602103, 0.1049397,
  0.0170477, 0.01124074, 0.003406085, 0.0001422856, 0.001755144, 
    -1.119886e-05, 0, 0, 0, 0, 0, 0, 0, 0, 2.80954e-05, 0.002876251, 
    0.007824379, 0.02112759, 0.001859933, 0.0001332076, 0, 0, 0, 0, 
    -0.0001484273, 0.001604565, 0.007525651, -0.0003218949, 0.01092147,
  0, 0.0003668278, 0.00185304, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.00031015, 
    -5.131786e-05, 0, 0.0007612183, -1.943678e-05, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0004146623, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -6.679932e-08, 0.01894299, 
    -5.10399e-05, -1.047863e-05, 2.892278e-06, 0, 0, 0, 0, 0, 0, 0, 
    -3.052446e-07, -3.440611e-08, 0, 0, 0,
  0, -1.208752e-06, 8.338256e-07, 0, 0, 0, -0.0001004592, 0.005327963, 
    0.001251801, -0.000357624, -3.168731e-12, -0.0003098361, 0.0139383, 
    0.08294717, 0.05800816, 0.02777438, 0.03395649, 0.01493519, 0.006051308, 
    9.211505e-05, 0.0193309, 0.01026131, 0.005212478, 0.02058313, 0.01540541, 
    -0.0001587255, -2.788224e-08, -2.182003e-05, 0,
  0.04768727, 0.03291542, 0.01467724, 0.003292762, 0.001837781, 0.04041864, 
    0.08514721, 0.1035699, 0.1311441, 0.07342725, 0.04259824, 0.008197422, 
    0.09776584, 0.1015732, 0.1030396, 0.1523055, 0.1236526, 0.09356006, 
    0.07154165, 0.0872073, 0.06809786, 0.06695744, 0.08288211, 0.1130808, 
    0.1282751, 0.1602906, 0.09888974, 0.09181093, 0.09433959,
  0.1571725, 0.1128467, 0.1332958, 0.156067, 0.1826607, 0.1741528, 0.1459415, 
    0.1469004, 0.1322204, 0.1588563, 0.127509, 0.1395591, 0.1412146, 
    0.2663444, 0.1507836, 0.1158562, 0.1083549, 0.130403, 0.1361548, 
    0.1312247, 0.1333608, 0.1733705, 0.2461849, 0.1388591, 0.09531962, 
    0.1072852, 0.08359398, 0.1099573, 0.1809457,
  0.03349487, 0.02700391, 0.03460466, 0.09305855, 0.04852497, 0.08528119, 
    0.05245565, 0.0599716, 0.07209174, 0.04957032, 0.08681362, 0.1147158, 
    0.1194662, 0.1025345, 0.09375943, 0.02387655, 0.09511453, 0.06637896, 
    0.2132069, 0.1862913, 0.06047965, 0.1023433, 0.07328766, 0.03358731, 
    0.1010411, 0.1208324, 0.1541184, 0.124444, 0.07973366,
  0.002538095, 0.001393598, 0.038309, 0.02627986, 0.06669085, 0.1810726, 
    0.1064908, 0.04974696, 0.01777259, 0.02711558, 0.03958572, 0.05740731, 
    0.09251616, 0.06117585, 0.02640168, 0.08702293, 0.09211794, 0.1274465, 
    0.3179278, 0.03639607, 0.04651258, 0.008469651, 7.630677e-08, 0.01555244, 
    0.08418294, 0.1506855, 0.2106118, 0.04557024, 0.0007562643,
  0.001827674, 0.06086854, 0.1050909, 0.1103855, 0.1012133, 0.1403111, 
    0.1216656, 0.006201338, 1.277335e-05, 0.005764608, 0.13923, 0.1752185, 
    0.135855, 0.05561027, 0.07512284, 0.1490535, 0.1313396, 0.1499135, 
    0.07343055, 0.008063006, -1.07591e-05, 1.348804e-05, -8.88628e-06, 
    0.04280441, 0.1945796, 0.1062956, 0.02631005, 0.008740344, 0.0001574133,
  7.193273e-07, 0.03084224, 0.184894, 0.09008903, 0.1519934, 0.05312254, 
    0.05231691, 0.03165369, 0.01912901, 0.1661181, 0.07438446, 0.06106569, 
    0.06012757, 0.08235543, 0.1528968, 0.02797025, 0.06283977, 0.003217683, 
    0.01034201, 0.004136559, 1.169024e-07, 8.357748e-07, 0.0005092583, 
    0.3098339, 0.2260507, 0.2238256, 0.0250928, 0.01310563, 5.024691e-05,
  -8.233917e-06, 6.46498e-06, 0.0002695355, 0.0009521538, 0.007843152, 
    0.09520546, 0.2240674, 0.08741703, 0.116244, 0.2382303, 0.1283574, 
    0.1292203, 0.1220159, 0.1503317, 0.06743645, 0.01039277, -2.997976e-05, 
    -0.0001598745, -2.983344e-05, -8.652201e-05, 0.0190291, 1.101584e-06, 
    0.01160785, 0.1073233, 0.1631282, 0.2601483, 0.06517702, 0.0301703, 
    0.001709284,
  0.0001421425, -5.365635e-11, 3.774828e-06, 4.383277e-05, 0.001495745, 
    0.009229846, 0.0005937148, 0.02480824, 0.00293273, 0.03031851, 
    0.06644114, 0.06320854, 0.04495573, 0.0009108894, 0.0004493483, 
    0.02611266, 0.05648172, 0.04243857, 0.03772491, 0.04946834, 0.08194681, 
    0.002673226, 0.0003955232, 0.0005726583, 0.001874278, 0.009615221, 
    0.02425627, 0.0958917, 0.09230081,
  0.04172825, -1.634304e-05, 1.592723e-07, -3.549932e-06, 4.305281e-07, 
    9.236032e-07, 5.299461e-06, 1.975318e-07, 5.089944e-07, -1.944102e-07, 
    7.191558e-05, 0.01257705, 0.02268366, -0.0001388665, 2.26602e-06, 
    0.006516857, 0.07091773, 0.07151096, 0.02739002, 0.107428, 0.05856609, 
    -3.799998e-05, 0.01083878, 1.856579e-05, 0.01514618, 0.04758601, 
    0.01600773, 0.09418299, 0.1822937,
  0.07196916, 0.0403709, 0.004316023, 0.003115881, 0.002264044, 1.623212e-05, 
    -0.0002483314, 0, 5.182291e-08, 0.01874592, 0.02321219, 0.06421766, 
    0.06238202, 0.07571969, 0.08737866, 0.0760185, 0.06080247, 0.2141499, 
    0.07696642, 0.0598792, 0.1243384, 0.0877817, 0.05698002, 0.02915496, 
    0.03695067, 0.06491794, 0.0708343, 0.03391542, 0.1145969,
  0.1023923, 0.04644817, 0.03886136, 0.04626894, 0.02825685, 0.01112107, 
    -0.0003871954, -1.820045e-06, 0, -3.47186e-07, 0.0003200784, 0.0171574, 
    0.02157896, 0.04773221, 0.07085085, 0.1359524, 0.2618804, 0.1888584, 
    0.1031393, 0.0836809, 0.01157211, 0.06623624, 0.1611669, 0.1775272, 
    0.1439601, 0.2237341, 0.2380294, 0.2331327, 0.124907,
  0.1546056, 0.05533228, 0.02886798, 0.008778653, 0.008749752, 0.006100637, 
    0, 0, 0, 0, 0, -1.082954e-05, 0.004278195, 0.001822112, 0.02019213, 
    0.07696846, 0.1974212, 0.1381295, 0.05332363, 0.02452218, 0.01153669, 
    0.02209058, 0.01618589, 0.03701784, 0.06578673, 0.06128384, 0.09176568, 
    0.1633484, 0.2366484,
  0.060693, 0.02244757, 0.01990044, 0.01216523, 0.01202122, -9.846173e-05, 
    0.0002045749, 0.003011281, 0, 0, 0, 0, 0, -0.0003387446, 0.01160298, 
    0.03131232, 0.07126741, 0.1180546, 0.01566948, 0.007900309, 0.007155339, 
    0.006736171, -1.240174e-06, 0, 0.002332962, 0.01150515, 0.03027446, 
    0.03481798, 0.04819056,
  1.118989e-05, 0.002281186, 0.008960692, 0.005979644, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 6.560043e-06, 0.01149653, -0.0002206859, 0.00250378, 0.0180024, 
    0.02609048, 0.002722215, 0, 0, 0, 0, -1.598415e-06, 0, 0, 0.0007986298, 
    9.79632e-05,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -8.47421e-06, 
    2.182474e-06, -1.051329e-05, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0002712897, 0.02856788, -0.00139728, 
    0.002239134, 0.009130533, 0.0002341481, 0.001445759, 0, 0, 0, 
    0.003304824, 0.03479387, 0.007211681, -0.0006098681, -4.476236e-05, 0, 0,
  0.008948452, -1.95731e-07, 0.01421306, 0.00252565, 0, 0, 0.00469787, 
    0.012324, 0.007559337, 0.001802493, 6.662113e-05, 0.006517565, 
    0.01468628, 0.1271848, 0.1039853, 0.06679514, 0.06870665, 0.07218429, 
    0.03005586, 0.0775413, 0.1299452, 0.08233406, 0.08893979, 0.04216377, 
    0.06901208, 0.07705209, 0.04578838, 0.02737562, 0.06253741,
  0.1174558, 0.08087785, 0.09236108, 0.1008474, 0.06715108, 0.1055362, 
    0.1380844, 0.1396873, 0.1807959, 0.1055774, 0.08476131, 0.086991, 
    0.1863905, 0.1911163, 0.1806869, 0.1797978, 0.1544196, 0.1176709, 
    0.1470138, 0.1433658, 0.110782, 0.09792089, 0.1344851, 0.2348438, 
    0.2362703, 0.2243691, 0.1745673, 0.1710481, 0.2095492,
  0.1875777, 0.1353581, 0.1506199, 0.1576552, 0.1990405, 0.1841405, 
    0.1428798, 0.1417309, 0.1328791, 0.1413115, 0.1267216, 0.1485842, 
    0.1230979, 0.2515277, 0.1489314, 0.1068696, 0.1013475, 0.1290146, 
    0.1257052, 0.1262319, 0.1366824, 0.1754884, 0.2306544, 0.1683617, 
    0.1085022, 0.1088688, 0.1128657, 0.09473003, 0.1972151,
  0.03060295, 0.02284357, 0.02722498, 0.09811207, 0.04395803, 0.07875302, 
    0.04356898, 0.05197647, 0.0502567, 0.03287702, 0.07701915, 0.08935894, 
    0.1050521, 0.08310612, 0.08315071, 0.01459724, 0.08849315, 0.06761593, 
    0.1935328, 0.1729522, 0.05286004, 0.08470494, 0.06904238, 0.03014928, 
    0.1000277, 0.09904088, 0.1512396, 0.1243143, 0.06632338,
  0.0006657527, 0.00134094, 0.03971684, 0.01680039, 0.05834969, 0.1352754, 
    0.08015272, 0.04667072, 0.008436249, 0.04684046, 0.02687163, 0.05890673, 
    0.07899159, 0.05280272, 0.01213306, 0.08355673, 0.0957247, 0.1056708, 
    0.3228114, 0.03240211, 0.03938675, 0.002934483, -1.706467e-07, 
    0.001563694, 0.06756268, 0.1282603, 0.1877867, 0.0329543, 3.645925e-05,
  0.0003336435, 0.04509489, 0.08076622, 0.1025918, 0.09785534, 0.1009861, 
    0.1060525, 0.007832205, 1.607912e-05, 0.004975153, 0.1218427, 0.1730061, 
    0.146235, 0.0525274, 0.06703336, 0.146275, 0.1317293, 0.1571932, 
    0.05975179, 0.0060547, 1.223385e-05, 1.693836e-06, -2.718511e-05, 
    0.03188634, 0.1607053, 0.1014542, 0.01274607, 2.410054e-05, 4.617554e-05,
  5.98392e-07, 0.02856663, 0.1127408, 0.07158168, 0.1018739, 0.03222083, 
    0.04154377, 0.03381774, 0.019793, 0.135768, 0.07013933, 0.04224327, 
    0.03930552, 0.06131275, 0.151918, 0.02526274, 0.0511056, 0.004188421, 
    0.009629672, 0.0001973502, 1.527197e-08, 5.675762e-07, 8.513006e-05, 
    0.2227071, 0.218494, 0.1919376, 0.01247654, 0.004383417, 4.586484e-06,
  -3.775859e-06, 1.977543e-06, 0.0002466077, 0.00051562, 0.004138271, 
    0.09421816, 0.1920551, 0.05252605, 0.09639662, 0.2176859, 0.1040417, 
    0.09445549, 0.1196872, 0.1499107, 0.06175427, 0.02715999, -0.0001611657, 
    0.0009180461, -0.0001544849, -7.66817e-05, 0.007205622, 7.672448e-08, 
    0.01270868, 0.1004598, 0.1047352, 0.2964052, 0.05501286, 0.01428652, 
    0.0006567467,
  1.809683e-05, 0, 7.73704e-06, 1.7297e-05, 0.002070686, 0.008582518, 
    0.001142858, 0.02365424, 0.002462099, 0.01303318, 0.05483389, 0.05646519, 
    0.05204536, 0.0006449683, 0.0005589204, 0.02925765, 0.06211329, 
    0.02819758, 0.04958313, 0.03555365, 0.06752237, 0.002354505, 
    0.0003999221, 0.0006340318, 0.002623149, 0.02627428, 0.03893929, 
    0.04365138, 0.07137553,
  0.009856525, -8.059467e-08, -3.91846e-10, -5.489707e-06, 1.594632e-07, 
    1.015544e-06, 2.490182e-05, 1.533516e-07, 3.831843e-06, 0.001247544, 
    0.0001675755, 0.01148627, 0.01776396, 3.490859e-06, 0.0003475132, 
    0.004780125, 0.06500071, 0.0305911, 0.0300682, 0.09654405, 0.03174379, 
    -3.825191e-06, 0.008719378, 1.997456e-05, 0.009253986, 0.05029973, 
    0.008354214, 0.08880276, 0.1329219,
  0.06933151, 0.02946466, 0.005977524, 0.01510991, 0.008161823, 4.3213e-05, 
    -0.0001668446, -5.375812e-07, 1.971172e-06, 0.07195333, 0.03885343, 
    0.08898628, 0.09873264, 0.100468, 0.06935201, 0.08903876, 0.05820107, 
    0.1994945, 0.05719977, 0.03514792, 0.1333401, 0.07807968, 0.04491226, 
    0.02937062, 0.0161315, 0.03804097, 0.03115086, 0.02507321, 0.1004468,
  0.1387353, 0.07043774, 0.0700729, 0.08329749, 0.05321188, 0.04994346, 
    0.001300407, 0.02223819, 2.681932e-05, 2.898362e-07, 0.01300655, 
    0.03176766, 0.03489893, 0.06335851, 0.1144594, 0.1460486, 0.2542813, 
    0.1924665, 0.1232445, 0.08953927, 0.03621264, 0.07238063, 0.1804021, 
    0.1735352, 0.1586214, 0.239519, 0.2356506, 0.2259072, 0.1347273,
  0.204898, 0.1372862, 0.06843045, 0.05653971, 0.06080473, 0.07382565, 
    0.02325076, 0, 0, -7.443777e-07, 0, 0.003218286, 0.02851502, 0.03726176, 
    0.08274105, 0.1392235, 0.2265546, 0.1320368, 0.05494736, 0.05027814, 
    0.02685402, 0.03619949, 0.02659487, 0.06891771, 0.07164999, 0.123192, 
    0.1161395, 0.2081768, 0.2984906,
  0.1266991, 0.06946625, 0.04143334, 0.03967643, 0.02684791, 0.01754535, 
    0.04746721, 0.04743768, 0.003876944, 9.211231e-05, 0, 0, -0.0008806228, 
    0.007561696, 0.05397872, 0.156202, 0.1955214, 0.2103717, 0.07007177, 
    0.03198112, 0.01987313, 0.01211436, 0.009228847, -1.287645e-05, 
    0.02343583, 0.05320389, 0.06873782, 0.1247189, 0.1305632,
  0.007404166, 0.01731408, 0.01694827, 0.01055442, 0.0004106294, 
    5.671614e-05, 0, 0, 0, 0, -5.474297e-09, 0, 0, 0.02308637, 0.02884199, 
    0.01864851, 0.08500641, 0.06226465, 0.07225677, 0.07296739, 0.00922839, 
    5.162027e-05, 0, 0, 0.0003772168, -6.383141e-06, 0, 0.001226496, 
    0.005193345,
  -1.988511e-07, 7.189078e-05, -1.905217e-08, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0001173974, 0.006865011, 0.00662177, 0.009211863, 0.01534035, 
    0.009315367, 2.970758e-05, -3.390612e-05, -3.362648e-06, 0, 0, 0, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0.0002184297, 0.005142181, 0.006470133, 
    0.02551256, 0.0198163, 0.09075433, 0.1321057, 0.06746123, 0.0434448, 
    0.01483453, -0.0005295214, -7.012729e-05, 0.02656828, 0.1185067, 
    0.05816685, -0.003449008, -0.0002198048, -6.491474e-05, 0,
  0.080253, 0.1128969, 0.07545514, 0.08155107, -0.0003483316, 0.0004003279, 
    0.08099213, 0.01948839, 0.008167316, 0.002705709, 0.01349988, 0.01978138, 
    0.07980127, 0.1714393, 0.1541914, 0.09552287, 0.1254947, 0.1200207, 
    0.1042998, 0.237173, 0.2393353, 0.160512, 0.2286139, 0.131272, 0.1842338, 
    0.1674587, 0.07106242, 0.07701563, 0.143446,
  0.1901245, 0.147134, 0.1846578, 0.185416, 0.1230706, 0.1396614, 0.1846599, 
    0.2083591, 0.2250209, 0.1552925, 0.1265779, 0.1347726, 0.2434042, 
    0.2164798, 0.1780186, 0.1691959, 0.1799211, 0.1080374, 0.1786088, 
    0.1714337, 0.1183242, 0.1704619, 0.1755581, 0.2403188, 0.2320331, 
    0.2214751, 0.1834201, 0.2360739, 0.2806433,
  0.1861578, 0.1594248, 0.153208, 0.1650479, 0.2132308, 0.2066906, 0.1385132, 
    0.1229224, 0.1164633, 0.1468448, 0.1251361, 0.1361587, 0.111016, 
    0.2306368, 0.1378617, 0.1063692, 0.0944737, 0.1198626, 0.1122659, 
    0.1260748, 0.1622564, 0.1646446, 0.221881, 0.1597599, 0.108094, 
    0.1000431, 0.1039837, 0.08610913, 0.2083054,
  0.04497431, 0.02255534, 0.03125124, 0.09636318, 0.03411239, 0.05883122, 
    0.03630774, 0.04414273, 0.03612502, 0.02120987, 0.07231946, 0.08033322, 
    0.09282171, 0.07497238, 0.0818548, 0.010464, 0.09487507, 0.07161321, 
    0.1717149, 0.1760045, 0.05301567, 0.07139247, 0.05212228, 0.03361698, 
    0.1020507, 0.08914629, 0.1362705, 0.1413033, 0.058608,
  0.000320261, 0.0002011234, 0.04374275, 0.01034939, 0.04875661, 0.1151286, 
    0.05347845, 0.04470561, 0.00682143, 0.04068518, 0.02202022, 0.05138215, 
    0.07245331, 0.03500276, 0.008140325, 0.08431824, 0.08826023, 0.07904779, 
    0.2717591, 0.01437734, 0.03717257, -3.842718e-05, -8.873079e-08, 
    0.0002409882, 0.05761098, 0.1165846, 0.1701065, 0.02181594, 6.607668e-05,
  0.002905587, 0.04068293, 0.05611377, 0.08206888, 0.09340061, 0.06475592, 
    0.0910501, 0.01038754, 2.35888e-05, 0.01120406, 0.0986903, 0.1728027, 
    0.1523029, 0.03721568, 0.04495986, 0.1491466, 0.1189796, 0.1635164, 
    0.04886403, 0.004236388, 7.119197e-06, 2.31153e-07, 9.58005e-06, 
    0.02112514, 0.1407381, 0.07379648, 0.004658367, 8.296992e-06, 7.163213e-07,
  9.326278e-07, 0.02667939, 0.08480005, 0.05766101, 0.08786748, 0.01955548, 
    0.03378323, 0.03070582, 0.02073727, 0.1240966, 0.06650522, 0.02995484, 
    0.03084528, 0.04870582, 0.1506909, 0.02323026, 0.03443851, 0.008007701, 
    0.01016696, 0.0001563842, -2.790461e-09, 7.546653e-07, 1.568759e-05, 
    0.1842074, 0.2019194, 0.1555724, 0.002698562, -0.0001055329, 1.328979e-06,
  -3.185445e-06, 5.404106e-07, 0.0001937165, 0.00035747, 0.003222791, 
    0.1005219, 0.1802963, 0.0323239, 0.07957868, 0.1884467, 0.09240997, 
    0.07870027, 0.1036212, 0.1475104, 0.06459355, 0.01942482, 0.0002531656, 
    0.009019909, -9.752491e-05, -2.902199e-05, 6.625619e-05, 8.157281e-08, 
    0.02984555, 0.09359927, 0.094257, 0.3198678, 0.04748216, 0.00363623, 
    0.0001244653,
  5.180762e-06, 0, 4.566747e-06, 5.344717e-06, 0.006702391, 0.01247369, 
    0.001826888, 0.04251461, 0.00167459, 0.005628082, 0.04406136, 0.05749241, 
    0.05642305, 0.001530976, 0.0004583307, 0.02062835, 0.06069023, 
    0.03217672, 0.05852102, 0.02547265, 0.06718627, 0.002198858, 
    0.0008827235, 0.0004495702, 0.01699564, 0.04575293, 0.01028315, 
    0.006461705, 0.08104965,
  0.001226488, 5.479976e-08, 4.041218e-09, -2.926866e-06, 3.320482e-07, 
    3.041955e-07, -0.0001852608, 1.238527e-07, 5.606831e-05, 0.01557408, 
    0.002322946, 0.01197017, 0.01674137, 4.215914e-05, 0.01163528, 
    0.0007894131, 0.06397083, 0.01725159, 0.01083596, 0.1306807, 0.01927869, 
    5.271384e-06, 0.004052117, 2.051273e-05, 0.0101167, 0.04309712, 
    0.0004698836, 0.05835095, 0.09422402,
  0.03141557, 0.01458382, 0.01188257, 0.01714601, 0.005611674, 2.010423e-05, 
    -8.933738e-05, 2.724407e-06, 2.897026e-06, 0.1246189, 0.05644168, 
    0.09324771, 0.1243323, 0.1352196, 0.08673582, 0.1022393, 0.05578292, 
    0.1911066, 0.05382732, 0.02074496, 0.1184572, 0.06828207, 0.05269016, 
    0.03475795, 0.01543365, 0.03163616, 0.02195719, 0.011725, 0.0711532,
  0.1244224, 0.05616147, 0.07236107, 0.1407321, 0.1136994, 0.0763322, 
    0.01477755, 0.05889842, 0.01046141, -0.0002074239, 0.05726684, 
    0.07545766, 0.08448731, 0.1059411, 0.152034, 0.1548391, 0.2476646, 
    0.2070769, 0.1132479, 0.1061, 0.05097887, 0.08796413, 0.1801995, 
    0.1660535, 0.1676973, 0.2389156, 0.2381195, 0.1962123, 0.125089,
  0.2307091, 0.1774088, 0.1343204, 0.131289, 0.1980808, 0.2148012, 0.0655402, 
    -6.096192e-05, 6.693145e-05, 0.0004609837, -2.789435e-07, 0.01153479, 
    0.04640349, 0.08456387, 0.1715053, 0.1784859, 0.2259272, 0.1359751, 
    0.08124492, 0.06891193, 0.03265052, 0.08066881, 0.07233271, 0.07958591, 
    0.1108395, 0.1395202, 0.1224366, 0.2130679, 0.3019433,
  0.1814139, 0.1343259, 0.09315227, 0.09970444, 0.1147359, 0.1262642, 
    0.2048206, 0.123764, 0.0708212, 0.02514772, 1.52316e-07, -6.707918e-05, 
    0.01222455, 0.04030292, 0.137501, 0.2454586, 0.2535696, 0.2571983, 
    0.1565655, 0.06086805, 0.05050991, 0.05949065, 0.04833655, 0.01115112, 
    0.06491765, 0.1098897, 0.1377862, 0.1796189, 0.1685933,
  0.05037462, 0.0787728, 0.05760653, 0.06213605, 0.02210415, 0.01147803, 
    0.009131555, 0.01838506, 0.009937459, 0.006465934, 6.539698e-05, 
    -2.688243e-05, 0.02138407, 0.03632726, 0.04516046, 0.06731702, 0.1308467, 
    0.09853123, 0.09735611, 0.1235405, 0.07431669, 0.004144541, 0, 
    -4.71866e-05, 0.005316881, 1.325786e-05, -4.333002e-07, 0.008286336, 
    0.03190907,
  0.0002306163, 0.005471081, 1.199799e-06, -0.0001412099, 0, 0, 0, 0, 0, 0, 
    0, 0, -0.0001145903, 0.01291522, 0.02559573, 0.02875206, 0.0340785, 
    0.03077631, 0.02449643, 0.009651441, 0.0003626339, -1.335783e-05, 0, 0, 
    0, 0, 0, 0, -6.556245e-05,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.008833406, 0.010794, 0.01415368, 
    0.04715635, 0.02415616, 0.09773054, 0.1553831, 0.192149, 0.1268664, 
    0.03707774, 0.05217016, 0.01579833, 0.1212069, 0.1512659, 0.09014225, 
    0.01101924, 0.0149466, 0.003499964, 0,
  0.1330335, 0.2276006, 0.222768, 0.1681449, -0.00279696, -0.003357538, 
    0.1746503, 0.03035748, 0.009639248, 0.02030393, 0.02771709, 0.01682729, 
    0.1391535, 0.182974, 0.1729876, 0.1124013, 0.1542729, 0.1281555, 
    0.1254859, 0.3069713, 0.3315439, 0.25195, 0.3058115, 0.2386662, 
    0.2823145, 0.2314879, 0.1180156, 0.09889606, 0.2811433,
  0.2163139, 0.2054773, 0.2631762, 0.2441564, 0.1908574, 0.1781282, 
    0.2010652, 0.2090953, 0.2704383, 0.1813764, 0.1681506, 0.1687139, 
    0.2392926, 0.238904, 0.1713063, 0.1581525, 0.187423, 0.1076674, 
    0.1776723, 0.1853645, 0.1530797, 0.2166938, 0.2265262, 0.2359004, 
    0.2378639, 0.2243431, 0.190717, 0.2546127, 0.3087812,
  0.1820008, 0.1708661, 0.1448418, 0.1609676, 0.2041135, 0.2165361, 
    0.1396687, 0.1110541, 0.1154551, 0.134268, 0.1383148, 0.1260111, 
    0.127449, 0.2168498, 0.145229, 0.1023134, 0.09822536, 0.1008306, 
    0.09857883, 0.1192999, 0.1536895, 0.1622755, 0.2112425, 0.1692404, 
    0.1050917, 0.100308, 0.1099371, 0.08489253, 0.1988062,
  0.04667055, 0.01613284, 0.02213426, 0.09327117, 0.03138801, 0.04441627, 
    0.03373656, 0.04419231, 0.04030256, 0.01502097, 0.08188727, 0.07819179, 
    0.08495462, 0.06011476, 0.07474693, 0.01071881, 0.1015842, 0.07436715, 
    0.1623186, 0.1552528, 0.04062956, 0.06021557, 0.05647452, 0.03257349, 
    0.1080042, 0.08118923, 0.1189305, 0.1297113, 0.07506286,
  0.0002465664, -1.814566e-05, 0.05480651, 0.01691058, 0.03473878, 0.12416, 
    0.03915223, 0.03859287, 0.004414236, 0.03369321, 0.02641366, 0.04684752, 
    0.06710925, 0.02523274, 0.01140012, 0.06427919, 0.07511821, 0.07001941, 
    0.2556091, 0.00582417, 0.03349444, -0.0001928586, -5.288014e-07, 
    0.0002283961, 0.04767513, 0.1011097, 0.1469883, 0.01382186, 5.199979e-05,
  0.0005863875, 0.03250863, 0.04768951, 0.08065712, 0.09197903, 0.04244584, 
    0.079276, 0.00537783, 1.076866e-05, 0.032801, 0.08092201, 0.1679368, 
    0.1656714, 0.04057319, 0.0331011, 0.1436867, 0.1248216, 0.154322, 
    0.04697124, 0.00355462, 1.222746e-05, 8.134548e-08, 8.228335e-06, 
    0.017648, 0.1281565, 0.06073204, 0.001954895, 2.433335e-06, 3.936331e-07,
  1.433475e-06, 0.02922702, 0.09260257, 0.05096681, 0.07611638, 0.01490692, 
    0.02848773, 0.02797115, 0.02035879, 0.1179293, 0.06330408, 0.02820502, 
    0.02563407, 0.04346525, 0.1469477, 0.02764944, 0.02518238, 0.01231492, 
    0.01322324, 9.121685e-05, 2.113583e-08, 2.463658e-06, 1.271069e-05, 
    0.1352623, 0.2081493, 0.1261328, 0.001595963, -1.175303e-05, 1.103339e-07,
  3.211844e-05, 4.484005e-07, 0.0001420174, 0.0003083677, 0.003185635, 
    0.1057694, 0.1475859, 0.01845951, 0.0736729, 0.1849383, 0.08932178, 
    0.06863124, 0.0910008, 0.1400111, 0.06367141, 0.003960155, 0.004237215, 
    -0.00023935, -1.137294e-05, -2.88733e-05, -2.39758e-06, 1.684424e-07, 
    0.05486024, 0.07981444, 0.1102891, 0.2970451, 0.0407512, 0.002282239, 
    0.000822442,
  6.907839e-07, 0, 1.805338e-06, 2.765431e-06, 0.0153579, 0.02154687, 
    0.001512253, 0.06385274, 0.001033528, 0.01083992, 0.04008691, 0.06573299, 
    0.06039826, 0.005583642, 0.003105096, 0.0206888, 0.06326861, 0.01997288, 
    0.07618062, 0.02271336, 0.06721734, 0.002095079, 0.0008425035, 
    0.0003049008, 0.003928398, 0.02670025, 0.008766513, 0.006194737, 
    0.07861434,
  -6.792972e-05, 2.77668e-09, -2.944591e-11, -2.616102e-06, 5.382885e-07, 
    1.008698e-05, -1.53423e-05, 2.062287e-05, 2.937529e-05, 0.01758794, 
    0.004712136, 0.01875847, 0.01586859, 1.801902e-05, 0.002742061, 
    0.004673965, 0.07471427, 0.01718917, 0.003337645, 0.1159538, 0.01201396, 
    2.041126e-05, 0.002288762, 1.926236e-05, 0.008966641, 0.04764632, 
    2.914688e-06, 0.05459129, 0.07527576,
  0.006223164, 0.001822419, 0.01284786, 0.02120616, 0.007759923, 
    0.0003862199, -4.618259e-05, 1.176098e-06, 0.001535996, 0.1615226, 
    0.08112403, 0.1204032, 0.1112564, 0.1193545, 0.1143436, 0.1021543, 
    0.05878432, 0.173148, 0.04167427, 0.0135941, 0.1124754, 0.05677161, 
    0.04471508, 0.05065152, 0.01550279, 0.03279524, 0.01965355, 0.01998185, 
    0.05518726,
  0.09341865, 0.03546939, 0.06672415, 0.2100132, 0.144351, 0.09090945, 
    0.04333058, 0.1110312, 0.06889295, 0.02933931, 0.07439648, 0.07470234, 
    0.1061365, 0.1214158, 0.147164, 0.1802199, 0.2543462, 0.2139399, 
    0.115774, 0.1225752, 0.06349328, 0.1251344, 0.1809354, 0.1766888, 
    0.1844571, 0.2490725, 0.2219498, 0.1678865, 0.1033,
  0.2475666, 0.185893, 0.1650716, 0.1600562, 0.2147976, 0.2358993, 0.1453504, 
    -0.001092833, 0.0007868984, 0.007907785, 0.02154904, 0.06162916, 
    0.1133254, 0.1334212, 0.2416462, 0.2645984, 0.221766, 0.1611042, 
    0.1271854, 0.08076621, 0.04861959, 0.1434304, 0.1839114, 0.1517363, 
    0.1585847, 0.1487655, 0.1534667, 0.2075119, 0.2817401,
  0.2365475, 0.14838, 0.1655979, 0.1874719, 0.1626432, 0.1907048, 0.2909647, 
    0.2232141, 0.1587039, 0.1132872, 0.004965775, 0.008842945, 0.02340901, 
    0.1133614, 0.1892768, 0.2802075, 0.2917428, 0.3002928, 0.1688541, 
    0.09041351, 0.1109421, 0.1233273, 0.07198242, 0.04508498, 0.1605244, 
    0.1765583, 0.1761771, 0.2038025, 0.1787587,
  0.1218274, 0.1600803, 0.1043652, 0.1186334, 0.134623, 0.1028075, 
    0.09211352, 0.06992839, 0.03442088, 0.03055098, 0.004542231, 0.001794913, 
    0.04312173, 0.06358334, 0.09324218, 0.09378013, 0.1667627, 0.1887096, 
    0.211074, 0.178139, 0.09055731, 0.04369767, 0.00317509, -0.001518846, 
    0.02926907, 3.321049e-06, -0.0001038256, 0.02762208, 0.07754157,
  0.04512226, 0.05296092, 0.04727905, 0.05586072, 0.0308379, 0.006555973, 
    0.004760303, 0.007094484, 0.0005250319, 1.1837e-05, 0, -0.0001584126, 
    0.008814365, 0.02302264, 0.03472364, 0.03718466, 0.03898189, 0.03789801, 
    0.03699452, 0.01811258, 0.01043932, 1.756505e-05, -2.403833e-10, 0, 0, 0, 
    -8.781481e-06, -0.001734326, 0.02316126,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -0.0003252596, -0.0003252596, -0.0003252596, -0.0003252596, 
    -0.0003252596, -0.0003252596, -0.0003252596, 0,
  -4.491342e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0.006690585, 0.01316396, 0.01714539, 
    0.009417224, 0.06760813, 0.03143923, 0.09590505, 0.1498353, 0.210777, 
    0.1945749, 0.1095003, 0.1159764, 0.1045811, 0.1309356, 0.1150232, 
    0.06152285, 0.0006305941, 0.04104248, 0.06843889, 0.000836756,
  0.126917, 0.2359067, 0.187609, 0.1546195, -0.0009673594, 0.008917241, 
    0.2110392, 0.06539234, 0.02814951, 0.09271673, 0.08052239, 0.1097952, 
    0.1628917, 0.1612277, 0.1591447, 0.1241513, 0.2039279, 0.1682277, 
    0.1426141, 0.3017446, 0.3604554, 0.2664358, 0.327222, 0.264436, 
    0.2894198, 0.2298008, 0.1455347, 0.1232229, 0.2737918,
  0.2410995, 0.2022423, 0.259777, 0.2480405, 0.2019003, 0.2103326, 0.2116807, 
    0.2137995, 0.2430234, 0.1969844, 0.2011141, 0.1740638, 0.2314934, 
    0.260455, 0.1703628, 0.1844062, 0.1899849, 0.1169533, 0.1932684, 
    0.2040409, 0.1838392, 0.2654507, 0.2492028, 0.2257775, 0.236599, 
    0.2299535, 0.2229394, 0.2672477, 0.3019446,
  0.177455, 0.1682421, 0.1369393, 0.1522594, 0.2151131, 0.2099914, 0.1317797, 
    0.1016355, 0.09974582, 0.1094885, 0.1256465, 0.1383341, 0.12088, 
    0.2103035, 0.141768, 0.08539449, 0.08366026, 0.0855217, 0.101751, 
    0.1253713, 0.1488211, 0.1714562, 0.2059202, 0.1637418, 0.09664965, 
    0.08919665, 0.09749153, 0.07038393, 0.1813135,
  0.05074384, 0.01290179, 0.01307527, 0.09029699, 0.0247807, 0.03536151, 
    0.03600957, 0.04582474, 0.03012648, 0.008758071, 0.07599609, 0.07536082, 
    0.07483309, 0.05759985, 0.06069512, 0.008133982, 0.06662113, 0.06445876, 
    0.1736273, 0.1510992, 0.03767795, 0.06228885, 0.04722461, 0.0251281, 
    0.1048186, 0.0801703, 0.09928502, 0.1069091, 0.06634081,
  0.0002239293, 9.592959e-05, 0.07727938, 0.01278242, 0.02397122, 0.1218233, 
    0.03448349, 0.0369329, 0.002424332, 0.03329801, 0.0266966, 0.03331854, 
    0.06078405, 0.01459227, 0.01460398, 0.06688534, 0.04813778, 0.06488635, 
    0.2323206, 0.004492214, 0.02951591, -0.0002215534, -1.519403e-06, 
    6.475712e-05, 0.04006291, 0.07432707, 0.1383885, 0.006846305, 0.0002895068,
  4.873324e-06, 0.02366174, 0.04612464, 0.08877917, 0.0930155, 0.03439375, 
    0.0796687, 0.003957338, 5.470294e-07, 0.03532331, 0.05450535, 0.153417, 
    0.1650471, 0.02798946, 0.02822388, 0.1258095, 0.1324943, 0.1466434, 
    0.04672029, 0.003046836, 6.425412e-07, -1.560263e-08, 5.897034e-06, 
    0.01513079, 0.1302152, 0.05589116, 0.001429377, 7.206864e-07, 3.502191e-08,
  1.583743e-05, 0.04188247, 0.1158843, 0.05618775, 0.0629244, 0.01366558, 
    0.02597165, 0.02246399, 0.01453516, 0.1139111, 0.06982949, 0.03289984, 
    0.03026356, 0.04303388, 0.144249, 0.03848604, 0.02575117, 0.01610398, 
    0.004172175, 0.0002148861, 8.119168e-08, 3.069651e-06, 8.567001e-05, 
    0.1091193, 0.2251637, 0.1194642, 0.001406805, 0.0001808156, 3.96414e-08,
  0.001755526, 9.743048e-06, 0.003518339, 0.0008481337, 0.003285421, 
    0.1125828, 0.1367421, 0.01085764, 0.07752983, 0.1740493, 0.08268198, 
    0.06671266, 0.08710214, 0.1361826, 0.06171715, 0.001674245, 0.009972041, 
    0.0003727115, -5.909116e-06, -1.574788e-05, 1.024323e-09, -8.190796e-08, 
    0.08325458, 0.07009739, 0.09831415, 0.2615705, 0.03735512, 0.003244852, 
    0.00676385,
  1.212371e-08, -3.438229e-11, 1.414113e-06, 2.225372e-06, 0.02134643, 
    0.03765145, 0.006707634, 0.0671098, 0.00133871, 0.01836652, 0.0345363, 
    0.06390991, 0.07067671, 0.009715367, 0.004535399, 0.01626673, 0.06608216, 
    0.0104427, 0.06730033, 0.02577055, 0.06052542, 0.002837421, 0.001897539, 
    0.001089674, 0.005748575, 0.00933629, 0.0004789219, 0.002147959, 
    0.06664917,
  3.640747e-06, -8.602333e-10, 0, -1.658856e-06, 2.210257e-06, 0.0004533943, 
    0.006677674, 0.006961318, -3.158122e-05, 0.01963462, 0.01104982, 
    0.02634631, 0.01541189, 7.188214e-06, 0.0001260081, 0.000763542, 
    0.07244349, 0.01039492, 0.002310442, 0.113047, 0.007768149, 3.201434e-05, 
    0.006926946, 4.761232e-05, 0.009544309, 0.05030935, 2.134002e-06, 
    0.03684437, 0.02802448,
  -8.423194e-05, 0.0002221792, 0.01567629, 0.01433976, 0.01528222, 
    0.0001542552, -4.110194e-05, 5.319035e-07, 0.006530334, 0.1690456, 
    0.08994681, 0.1184669, 0.07683095, 0.08698829, 0.1379838, 0.09645559, 
    0.06694888, 0.1734264, 0.03861113, 0.01340155, 0.1091921, 0.05681729, 
    0.05818019, 0.05441253, 0.02058607, 0.03188815, 0.01702538, 0.01810878, 
    0.04018071,
  0.07349216, 0.02058551, 0.07735463, 0.2738421, 0.1295911, 0.1062216, 
    0.08109844, 0.1277987, 0.08031515, 0.06987753, 0.06664881, 0.1046338, 
    0.1203249, 0.1317564, 0.1580214, 0.1991978, 0.2414511, 0.2089692, 
    0.0905502, 0.1629791, 0.1074857, 0.1245368, 0.1873683, 0.1818112, 
    0.1740424, 0.2405228, 0.2023054, 0.1426083, 0.088181,
  0.2504942, 0.2140189, 0.163649, 0.1807369, 0.1919139, 0.2505841, 0.1596168, 
    0.009248109, 0.02799198, 0.01954834, 0.04619742, 0.1266502, 0.1886168, 
    0.1424969, 0.2815585, 0.2805096, 0.2343705, 0.1726405, 0.1342434, 
    0.104061, 0.08322504, 0.1583408, 0.224535, 0.1904275, 0.1918458, 
    0.1898964, 0.177684, 0.2105712, 0.2637876,
  0.250834, 0.1430317, 0.1996533, 0.2424213, 0.2026545, 0.1999907, 0.3236437, 
    0.2961156, 0.2170912, 0.1738293, 0.03855283, 0.03476032, 0.04160442, 
    0.1740971, 0.2544195, 0.2919441, 0.3004209, 0.3362272, 0.1681091, 
    0.1246463, 0.1872739, 0.1662297, 0.1136385, 0.2170281, 0.2049722, 
    0.2245951, 0.1986799, 0.2088457, 0.2153884,
  0.2184, 0.1867362, 0.13374, 0.1658692, 0.1721367, 0.1731357, 0.2105965, 
    0.1796939, 0.1158184, 0.07376242, 0.04088377, 0.05107839, 0.06951115, 
    0.0983488, 0.1068619, 0.1198596, 0.2151966, 0.2229015, 0.2592924, 
    0.2128925, 0.09800895, 0.06443159, 0.02114438, -0.007995868, 0.07599087, 
    0.001571618, 4.698954e-05, 0.07532481, 0.123362,
  0.1431598, 0.1470371, 0.1001946, 0.1246108, 0.04087848, 0.009005902, 
    0.0125996, 0.01580887, 0.03084298, 0.02391816, 0.001427231, 0.00385366, 
    0.03919973, 0.06396806, 0.06894058, 0.05756338, 0.06026801, 0.06291304, 
    0.06419186, 0.02572918, 0.02017826, 0.02438577, -0.0001621823, 
    -6.119063e-05, -0.0008517188, -3.057616e-05, -0.001914287, 0.006983805, 
    0.1306621,
  0.02296697, 0.02169413, 0.0204213, 0.01914847, 0.01787563, 0.0166028, 
    0.01532997, 0.01983974, 0.02017077, 0.0205018, 0.02083283, 0.02116385, 
    0.02149488, 0.02182591, 0.02204191, 0.02394352, 0.02584513, 0.02774675, 
    0.02964836, 0.03154998, 0.03345159, 0.02894863, 0.02798882, 0.02702901, 
    0.0260692, 0.0251094, 0.02414959, 0.02318978, 0.02398524,
  0.0009700851, -9.700741e-06, 0, 0, 0, 0, 0, 0, 0.000325851, 0.01469388, 
    0.01609581, 0.01530689, 0.01145026, 0.05876083, 0.04140523, 0.08550776, 
    0.1513492, 0.2288949, 0.216778, 0.1529602, 0.1490283, 0.1367859, 
    0.142322, 0.08260369, 0.02567876, -0.004816513, 0.03210609, 0.1417359, 
    0.04270904,
  0.1470665, 0.2336357, 0.1761532, 0.1466709, 0.05096289, 0.06720813, 
    0.2181682, 0.1629097, 0.131548, 0.1741046, 0.1157834, 0.1752711, 
    0.1565509, 0.154528, 0.1465048, 0.1505371, 0.2256893, 0.2561896, 
    0.1582054, 0.3086103, 0.3963121, 0.3374277, 0.327448, 0.2843391, 
    0.2978097, 0.2331191, 0.1229859, 0.1152772, 0.2593803,
  0.2451607, 0.1924436, 0.2434172, 0.2468799, 0.2285621, 0.2083581, 
    0.2290478, 0.238404, 0.2674409, 0.2357504, 0.2221371, 0.1999094, 
    0.2275805, 0.2469577, 0.1996275, 0.1695253, 0.1671844, 0.1145151, 
    0.1865961, 0.2232447, 0.193412, 0.270171, 0.2443101, 0.2367586, 
    0.2442758, 0.2232358, 0.2296244, 0.2625294, 0.2955818,
  0.1804047, 0.1707986, 0.1434935, 0.1579218, 0.2105832, 0.2263543, 0.144844, 
    0.09155868, 0.1002273, 0.1278944, 0.1418239, 0.1542395, 0.1338013, 
    0.2151333, 0.1453166, 0.07571535, 0.08046787, 0.09209502, 0.07843459, 
    0.1291226, 0.1475439, 0.1762141, 0.1824197, 0.157938, 0.09862509, 
    0.08701777, 0.1016108, 0.07504977, 0.1686816,
  0.04615583, 0.01386822, 0.007909376, 0.08605126, 0.02118213, 0.02677357, 
    0.03062589, 0.04437212, 0.03576237, 0.009286615, 0.05640493, 0.06768717, 
    0.07052955, 0.06340691, 0.05219838, 0.007517256, 0.05856711, 0.08265281, 
    0.1855144, 0.1363408, 0.03355128, 0.05752557, 0.03789789, 0.0212043, 
    0.09511767, 0.0821059, 0.08807197, 0.08999994, 0.05953212,
  0.001270082, 0.002275199, 0.1106876, 0.008006195, 0.02204, 0.1224046, 
    0.03313932, 0.03688578, 0.0003173522, 0.03336561, 0.01463647, 0.01827125, 
    0.06367903, 0.005957636, 0.01873685, 0.07173647, 0.0616864, 0.06374568, 
    0.1920289, 0.00510511, 0.02247057, -0.0002254802, -4.423924e-07, 
    -9.296503e-06, 0.03220065, 0.0659207, 0.1425689, 0.003872673, 0.0004297463,
  2.808072e-06, 0.02625304, 0.06014733, 0.09582491, 0.1096247, 0.04156987, 
    0.07397567, 0.0004746862, 2.281481e-06, 0.05097235, 0.05125298, 
    0.1449289, 0.1720407, 0.04331194, 0.03344727, 0.1525103, 0.1596539, 
    0.1517062, 0.04044816, 0.002563181, -3.581992e-06, 9.289655e-09, 
    1.160447e-05, 0.01178921, 0.1481605, 0.04516026, 0.00171669, 
    1.860419e-06, 3.687952e-08,
  0.008153216, 0.07901878, 0.1396994, 0.08902854, 0.06801074, 0.01420509, 
    0.0275769, 0.02508119, 0.01352153, 0.1172784, 0.08253504, 0.04406851, 
    0.05026228, 0.04516486, 0.1361358, 0.04426598, 0.03557584, 0.01782589, 
    0.00207798, 0.0007428648, 3.18979e-08, 3.064863e-06, 0.0004465605, 
    0.1011812, 0.249071, 0.1376225, 0.003713737, 2.492801e-05, 5.148221e-06,
  0.07842527, 0.00176186, 0.04063419, 0.003898271, 0.003774588, 0.1079755, 
    0.1351283, 0.007227638, 0.05700586, 0.17191, 0.09667412, 0.07664061, 
    0.08626942, 0.13019, 0.06334369, 0.00244596, 0.003339942, -7.489946e-05, 
    0.001545362, -8.219162e-06, 4.982321e-05, -3.711598e-07, 0.08497915, 
    0.07308844, 0.1083488, 0.2151705, 0.03722394, 0.005932624, 0.02187113,
  -3.78966e-06, 9.754132e-10, 1.100775e-06, 1.971635e-05, 0.03171183, 
    0.03657148, 0.01290745, 0.06485271, 0.001469353, 0.02662087, 0.03384032, 
    0.06144319, 0.08256436, 0.01133498, 0.004825624, 0.01998427, 0.06068068, 
    0.008176161, 0.05515104, 0.03220883, 0.0606471, 0.005279381, 0.005665178, 
    0.003728849, 0.005642406, 0.001479863, 0.001264138, 0.0001518029, 
    0.0440152,
  2.887013e-06, -4.93566e-09, 0, 8.4736e-06, 2.286357e-06, 0.00122825, 
    0.01199932, 0.001599292, -1.733107e-05, 0.03887017, 0.01895985, 
    0.03478717, 0.01557463, -3.694348e-06, 6.536137e-06, 0.0009303333, 
    0.05917145, 0.004380157, 0.006072089, 0.08809378, 0.006764506, 
    0.0008735463, 0.007634802, 0.000109265, 0.01645036, 0.05566968, 
    8.676252e-07, 0.01354515, 0.01346787,
  0.0009781154, 8.345916e-05, 0.01698424, 0.01746897, 0.02443589, 
    8.994031e-05, 0.000195489, -2.413031e-06, 0.02654909, 0.1736665, 
    0.08649825, 0.08749655, 0.06369726, 0.08206221, 0.140548, 0.08329611, 
    0.06390947, 0.1629598, 0.02567917, 0.006154258, 0.1100769, 0.05793128, 
    0.06867883, 0.05120201, 0.02027657, 0.03381464, 0.01593837, 0.008709989, 
    0.02991857,
  0.06588754, 0.01468405, 0.1034856, 0.322736, 0.1076923, 0.1001404, 
    0.1509735, 0.1134969, 0.07377183, 0.07296313, 0.06023807, 0.1227577, 
    0.1301547, 0.133091, 0.1640451, 0.1819441, 0.2241215, 0.2199285, 
    0.0888657, 0.1953998, 0.1426524, 0.1164305, 0.179852, 0.18397, 0.1681609, 
    0.2247667, 0.1765454, 0.1232569, 0.0675616,
  0.194048, 0.2035401, 0.1666495, 0.1686576, 0.1704085, 0.2447835, 0.1946443, 
    0.08764961, 0.0923097, 0.05000776, 0.06628408, 0.1589702, 0.2284224, 
    0.163322, 0.301223, 0.2816572, 0.2209142, 0.1705164, 0.1052936, 
    0.1413655, 0.1259298, 0.1577909, 0.2579626, 0.2498089, 0.2066408, 
    0.2168815, 0.189479, 0.2029844, 0.2616958,
  0.2361608, 0.1403136, 0.195749, 0.2510622, 0.2323045, 0.2796362, 0.3246506, 
    0.3336025, 0.2492217, 0.2184599, 0.109502, 0.05729191, 0.07413885, 
    0.2045893, 0.3052821, 0.3316523, 0.3277961, 0.3601055, 0.2162955, 
    0.1494544, 0.1898246, 0.2120791, 0.1737806, 0.2687394, 0.2095672, 
    0.3045791, 0.2511663, 0.2336199, 0.2240358,
  0.2591861, 0.2663525, 0.1465486, 0.1981331, 0.1629078, 0.2101743, 
    0.2510613, 0.2496662, 0.1764245, 0.1007081, 0.03830114, 0.09536308, 
    0.1262469, 0.1452557, 0.1179992, 0.1529564, 0.2594762, 0.2743073, 
    0.2901722, 0.2294871, 0.09596581, 0.06958158, 0.05609242, 0.0364947, 
    0.1008413, 0.01809723, -0.001078844, 0.1494975, 0.1649975,
  0.226321, 0.2154141, 0.1467234, 0.1640055, 0.09652393, 0.04527127, 
    0.06296804, 0.06560215, 0.06206479, 0.05819248, 0.0374199, 0.02119086, 
    0.05565365, 0.1143212, 0.1613071, 0.1816848, 0.1543707, 0.1143091, 
    0.1168976, 0.08990213, 0.04953251, 0.04054143, 0.008428883, -0.003082468, 
    0.0008985535, -0.0003167414, -0.01042328, 0.1159317, 0.2384861,
  0.03809136, 0.03797016, 0.03784896, 0.03772775, 0.03760655, 0.03748535, 
    0.03736415, 0.04379889, 0.04448894, 0.04517899, 0.04586904, 0.04655909, 
    0.04724914, 0.04793919, 0.04843481, 0.04833822, 0.04824163, 0.04814504, 
    0.04804845, 0.04795187, 0.04785528, 0.04310247, 0.0426302, 0.04215794, 
    0.04168568, 0.04121342, 0.04074116, 0.0402689, 0.03818832,
  0.06700874, -0.002116767, -2.805523e-05, -1.523818e-08, 0.0001742398, 
    -0.0004867392, 0, -7.599677e-07, 0.009229839, 0.01934232, 0.01425858, 
    0.0343443, 0.02757425, 0.05811846, 0.07737096, 0.09059855, 0.1551468, 
    0.2694305, 0.2550188, 0.1871418, 0.1715637, 0.1880421, 0.2075698, 
    0.05325089, 0.01117674, -0.004566818, 0.04182236, 0.1790955, 0.1056587,
  0.1615234, 0.2159404, 0.1959132, 0.136779, 0.08214076, 0.1178836, 
    0.2326718, 0.2596834, 0.2427866, 0.1844078, 0.2436968, 0.2217512, 
    0.1685929, 0.1561061, 0.1432548, 0.2124133, 0.2560101, 0.2750143, 
    0.209709, 0.2995285, 0.4182869, 0.3497798, 0.3539845, 0.3290251, 
    0.3241038, 0.2659577, 0.1055999, 0.1452404, 0.2845886,
  0.2676133, 0.2347362, 0.2626843, 0.2877809, 0.2558682, 0.2199151, 
    0.2199776, 0.2537692, 0.2790006, 0.2638428, 0.2326867, 0.2281148, 
    0.236687, 0.2434357, 0.1861935, 0.1651143, 0.176618, 0.1612509, 
    0.2068086, 0.2317175, 0.2795376, 0.285847, 0.2373552, 0.2473787, 
    0.2321294, 0.2147013, 0.2390287, 0.2978165, 0.3018087,
  0.1817732, 0.1598419, 0.1856885, 0.1996152, 0.2243535, 0.2211762, 
    0.1380763, 0.08185484, 0.08708166, 0.1319026, 0.1562397, 0.1666101, 
    0.1211628, 0.1954114, 0.1467546, 0.07276665, 0.07426535, 0.09134466, 
    0.09329902, 0.1289747, 0.1570437, 0.1838118, 0.1814984, 0.152257, 
    0.1028446, 0.08265225, 0.09930308, 0.09463301, 0.1873877,
  0.04787433, 0.01304103, 0.008225916, 0.08095711, 0.01251253, 0.02649118, 
    0.03346149, 0.04052131, 0.03525326, 0.008672126, 0.04105095, 0.06097278, 
    0.07249244, 0.07001782, 0.04008832, 0.00782068, 0.06192713, 0.07693023, 
    0.1974085, 0.1492887, 0.02954496, 0.05682343, 0.0343884, 0.01733945, 
    0.0851064, 0.08672097, 0.08336248, 0.0797655, 0.05596794,
  0.002712063, 0.0002073452, 0.1370639, 0.005318033, 0.02241919, 0.1161622, 
    0.03143598, 0.04247596, 3.521209e-06, 0.02926034, 0.03263129, 0.01910261, 
    0.06087669, 0.006480112, 0.02368202, 0.06954525, 0.05517176, 0.06500391, 
    0.1620477, 0.007873432, 0.0232728, -0.0001564221, -3.065285e-08, 
    -7.929372e-06, 0.0297566, 0.06828339, 0.1545519, 0.0059791, 0.0001135367,
  7.117134e-06, 0.03805278, 0.07843509, 0.1070058, 0.1288115, 0.05497532, 
    0.0903905, 0.0003265293, 2.406041e-06, 0.0693532, 0.05944805, 0.1464864, 
    0.1861278, 0.04510152, 0.04120228, 0.2042467, 0.1775301, 0.1622076, 
    0.03413296, 0.002533877, 1.300006e-05, 8.467085e-08, 2.00924e-05, 
    0.009571313, 0.1754729, 0.04828841, 0.003089054, 2.183756e-06, 
    3.612107e-07,
  0.03172995, 0.1364212, 0.1949784, 0.1259468, 0.08535923, 0.0180206, 
    0.031772, 0.02250244, 0.02290055, 0.1434506, 0.09072586, 0.06694407, 
    0.07671727, 0.06405017, 0.152515, 0.0524152, 0.05019544, 0.01609496, 
    0.002480198, 0.001142839, 6.912869e-07, 9.789691e-06, 7.617777e-05, 
    0.1159318, 0.297949, 0.1596724, 0.007982007, 3.932333e-05, 0.0001160811,
  0.1415934, 0.03702936, 0.06894857, 0.005897279, 0.008198106, 0.1049198, 
    0.1379691, 0.008718109, 0.04975433, 0.1956775, 0.1095985, 0.08866749, 
    0.101709, 0.135608, 0.06152738, 0.002248991, 0.00228214, -0.0007156255, 
    0.0001341047, -4.861849e-06, 0.01360699, 0.001370076, 0.07510597, 
    0.06335308, 0.1048975, 0.1950243, 0.04390806, 0.004002516, 0.02224722,
  -0.0001218546, 2.86389e-07, 0.0001102344, 0.000101017, 0.04088053, 
    0.03828107, 0.02235444, 0.06918795, 0.002896619, 0.043614, 0.04431294, 
    0.07554451, 0.09140267, 0.01570678, 0.009594603, 0.02333238, 0.0617416, 
    0.001584581, 0.05099998, 0.03919993, 0.06107837, 0.004041051, 
    0.007526946, 0.003318181, 0.004231764, 0.0006060963, 0.0007169094, 
    -5.577347e-05, 0.02602912,
  1.31912e-06, -4.519618e-10, 0, 0.0001351679, 1.7302e-06, 0.0008424222, 
    0.01554083, 0.001268256, 8.487699e-06, 0.02854662, 0.02356891, 
    0.03865166, 0.02617176, 8.154882e-05, -1.722038e-05, 0.00116683, 
    0.05376637, 0.003378043, 0.001122958, 0.07932647, 0.0221737, 0.008914982, 
    0.01017167, 0.0005004551, 0.01860829, 0.05679394, 3.276066e-06, 
    0.001638362, 0.02477657,
  9.069997e-05, -1.934546e-05, 0.02180249, 0.01462758, 0.0325436, 
    0.000127185, 0.00160782, -4.775494e-05, 0.07055377, 0.1686515, 
    0.07362198, 0.06969832, 0.06851615, 0.08845302, 0.1465607, 0.09207741, 
    0.06878756, 0.1450909, 0.01674508, 0.00629525, 0.107922, 0.07503283, 
    0.07457465, 0.05520288, 0.02271676, 0.03877749, 0.02073873, 0.009631124, 
    0.02201713,
  0.05125468, 0.01185401, 0.1235155, 0.3208141, 0.09969783, 0.09496054, 
    0.1805325, 0.1004073, 0.06159605, 0.06416278, 0.05662416, 0.1233681, 
    0.1286364, 0.1345137, 0.1836831, 0.1987713, 0.2255116, 0.2357297, 
    0.1003057, 0.2015143, 0.1722649, 0.1089701, 0.1900747, 0.1824688, 
    0.1790217, 0.2170826, 0.1756627, 0.1180636, 0.07417194,
  0.1798071, 0.1962074, 0.1683301, 0.169656, 0.1539438, 0.2396073, 0.201598, 
    0.1442057, 0.152444, 0.06032437, 0.0721641, 0.1954553, 0.2397081, 
    0.156416, 0.2995067, 0.2632582, 0.1980338, 0.1487036, 0.09251229, 
    0.1445405, 0.1346131, 0.1495909, 0.3012407, 0.2743412, 0.1999809, 
    0.2259866, 0.1934681, 0.196216, 0.2593142,
  0.2266356, 0.1444092, 0.1977233, 0.2982885, 0.217093, 0.2597426, 0.327607, 
    0.3600301, 0.2957483, 0.2998997, 0.1572353, 0.1135341, 0.1405642, 
    0.2214686, 0.3462806, 0.3329431, 0.3264431, 0.3557533, 0.2208965, 
    0.2105888, 0.2071986, 0.2295194, 0.2208335, 0.3079181, 0.2414392, 
    0.3405182, 0.2391163, 0.2153279, 0.2279623,
  0.2741548, 0.2619944, 0.2049821, 0.2304066, 0.1687199, 0.2437316, 
    0.2779389, 0.2994347, 0.2709199, 0.2350376, 0.07836158, 0.1747293, 
    0.205847, 0.1910608, 0.146344, 0.1744117, 0.2772515, 0.2897549, 
    0.2819147, 0.2247164, 0.1190201, 0.08407696, 0.06492411, 0.04714456, 
    0.1593472, 0.04647313, -0.001393051, 0.1706184, 0.1732981,
  0.225715, 0.2480897, 0.1717364, 0.1968724, 0.1360952, 0.09019466, 
    0.1167036, 0.1382114, 0.09218463, 0.0757094, 0.04855043, 0.06553848, 
    0.1066162, 0.1415966, 0.2308079, 0.238127, 0.1859211, 0.1137799, 
    0.1220489, 0.1112804, 0.09382381, 0.06858084, 0.062367, -0.0008637134, 
    0.02703919, 0.005761165, -0.004868314, 0.2348048, 0.2406419,
  0.07488589, 0.07580532, 0.07672475, 0.07764418, 0.0785636, 0.07948303, 
    0.08040246, 0.08182472, 0.08026912, 0.07871352, 0.07715791, 0.07560232, 
    0.07404672, 0.07249112, 0.04868697, 0.04946999, 0.050253, 0.05103602, 
    0.05181903, 0.05260205, 0.05338506, 0.08801804, 0.08787121, 0.08772437, 
    0.08757752, 0.08743069, 0.08728384, 0.087137, 0.07415035,
  0.1655094, 0.03911929, -0.002195228, -6.044349e-06, 0.0009469087, 
    0.001018556, -0.000782294, -0.0003900543, 0.01362049, 0.02225146, 
    0.04130077, 0.04294284, 0.06084031, 0.08144593, 0.1126199, 0.1890032, 
    0.1671163, 0.2875903, 0.2752092, 0.2114429, 0.1752005, 0.2051217, 
    0.2011482, 0.02291062, 0.004946683, -0.004983597, 0.05760048, 0.2308547, 
    0.1136641,
  0.1455798, 0.1946623, 0.2257879, 0.1462861, 0.08124382, 0.1392823, 
    0.2513666, 0.3235807, 0.2549191, 0.1872218, 0.2504503, 0.2321713, 
    0.1486085, 0.1754004, 0.1632836, 0.217322, 0.2755971, 0.3048345, 
    0.1825207, 0.3556991, 0.423368, 0.364043, 0.3322841, 0.3464463, 
    0.3153774, 0.2611887, 0.1214221, 0.2283991, 0.2934546,
  0.2994342, 0.3077338, 0.2582619, 0.3262627, 0.3117699, 0.2545491, 
    0.2500393, 0.3114457, 0.2740583, 0.2908344, 0.2529199, 0.2526167, 
    0.2543809, 0.252573, 0.1771382, 0.1482271, 0.1868315, 0.1568952, 
    0.2207242, 0.2687415, 0.2716452, 0.2868434, 0.2667924, 0.2375839, 
    0.2482585, 0.2657254, 0.237571, 0.2844616, 0.3006271,
  0.1642869, 0.1704608, 0.2099286, 0.2079288, 0.2230507, 0.2214549, 
    0.1490648, 0.09068334, 0.07601511, 0.1273577, 0.1325314, 0.1873848, 
    0.1209277, 0.1909206, 0.1451234, 0.08953045, 0.06772566, 0.09502451, 
    0.1062288, 0.1355956, 0.1610438, 0.1955174, 0.1554544, 0.1417185, 
    0.1049301, 0.09746751, 0.0963474, 0.1081337, 0.151029,
  0.05099023, 0.009170922, 0.01437122, 0.08755667, 0.01347949, 0.03868686, 
    0.03344865, 0.04071367, 0.04704555, 0.006067082, 0.0316393, 0.06322515, 
    0.08325439, 0.08529178, 0.0512111, 0.006420743, 0.05141571, 0.0722549, 
    0.2144366, 0.1612272, 0.03169401, 0.06032791, 0.0168181, 0.02912812, 
    0.07185588, 0.1111251, 0.09319598, 0.07976034, 0.0638747,
  0.005134639, 0.0005108197, 0.1366112, 0.00539582, 0.0252783, 0.09967799, 
    0.02962489, 0.04230307, -6.433285e-05, 0.01900851, 0.02384944, 
    0.02375682, 0.06345171, 0.004887918, 0.02358049, 0.07713358, 0.05182806, 
    0.08686297, 0.1497951, 0.00785411, 0.02790178, 0.0002411045, 
    6.678491e-08, 0.0001276725, 0.04666176, 0.08058239, 0.1834291, 
    0.01772753, 0.0002076822,
  -1.431556e-05, 0.05762372, 0.09741092, 0.1179228, 0.1452398, 0.06992593, 
    0.1102358, 0.0007945456, 1.590089e-06, 0.07024787, 0.0721015, 0.1606029, 
    0.1818657, 0.04575231, 0.0410303, 0.2485968, 0.2033281, 0.1829261, 
    0.0307574, 0.00364572, 7.804819e-05, 1.120248e-07, 1.179497e-05, 
    0.007001376, 0.2062648, 0.05989208, 0.005955546, 2.92368e-08, 4.269107e-07,
  0.02549121, 0.1286867, 0.2679767, 0.1671157, 0.09790049, 0.02784187, 
    0.0373124, 0.02282917, 0.02332173, 0.1813079, 0.1031782, 0.07649089, 
    0.09541527, 0.07565545, 0.1484339, 0.05319589, 0.05651207, 0.01926075, 
    0.003582946, 0.0007759667, 3.8669e-07, 5.577313e-05, 0.0001805792, 
    0.1467065, 0.3482571, 0.1932586, 0.01024546, 5.70607e-05, 9.78396e-05,
  0.1601563, 0.0557454, 0.08893199, 0.01352076, 0.009933317, 0.09912633, 
    0.1346691, 0.0174849, 0.06964666, 0.2190479, 0.1302657, 0.1085647, 
    0.1059986, 0.1412001, 0.07348399, 0.002101385, 0.007709443, 
    -0.0005013265, -4.194945e-05, -3.752803e-05, 0.001487214, 0.01610448, 
    0.0943606, 0.07613939, 0.149191, 0.2007258, 0.05099407, 0.003137814, 
    0.04377972,
  -1.065432e-05, 2.775686e-06, 0.0009349539, 0.002016881, 0.04646853, 
    0.03935714, 0.02609254, 0.07821337, 0.005794421, 0.05147925, 0.04631463, 
    0.08507121, 0.08918453, 0.01771688, 0.02182694, 0.03451518, 0.06701738, 
    0.002229155, 0.04573862, 0.04362765, 0.06753313, 0.007671795, 0.01133726, 
    0.004440323, 0.004530916, 0.003283921, -1.188829e-06, 1.226839e-05, 
    0.02106167,
  2.001836e-06, 4.962977e-07, -4.82641e-11, 0.001896553, 4.176015e-07, 
    2.789623e-06, 0.01713791, 0.01624775, 0.0001157087, 0.03081987, 
    0.02728796, 0.05989252, 0.03852491, -2.410659e-06, 0.0005439214, 
    0.001519733, 0.05681393, 0.00394867, 0.001531406, 0.08334335, 0.04910281, 
    0.02642104, 0.02560163, 0.001909631, 0.02264052, 0.0701001, 4.741238e-06, 
    0.003532808, 0.0488543,
  3.612368e-06, -3.666079e-06, 0.02440899, 0.01586293, 0.03777093, 
    0.00255175, 0.001812091, 6.078454e-05, 0.1198134, 0.159349, 0.07258788, 
    0.0655179, 0.06503775, 0.0969854, 0.1436142, 0.1037985, 0.07094332, 
    0.1306109, 0.01641843, 0.01460889, 0.1050893, 0.08864414, 0.07454295, 
    0.05838621, 0.031875, 0.05100689, 0.02802959, 0.004138308, 0.04329229,
  0.0291031, 0.00828233, 0.1394226, 0.3254248, 0.09402428, 0.08455294, 
    0.1881402, 0.08363265, 0.05002069, 0.04885221, 0.04980761, 0.1135975, 
    0.1197795, 0.1416164, 0.2177488, 0.2055253, 0.2212862, 0.2215263, 
    0.09668653, 0.1914753, 0.1846972, 0.1088677, 0.1824398, 0.1618148, 
    0.1720371, 0.2119698, 0.1767529, 0.1102334, 0.07015505,
  0.1866259, 0.2041492, 0.1603788, 0.1535422, 0.1344571, 0.2224305, 
    0.1887192, 0.178343, 0.160705, 0.05806622, 0.07738329, 0.2072062, 
    0.2349951, 0.1582645, 0.3002598, 0.2595164, 0.1780834, 0.1496201, 
    0.08667537, 0.1273429, 0.1527594, 0.1337315, 0.3286845, 0.3286214, 
    0.2308098, 0.221815, 0.1906226, 0.1907747, 0.235687,
  0.2240812, 0.1467783, 0.2086359, 0.3220859, 0.2237998, 0.2684638, 
    0.3291491, 0.3555366, 0.3092624, 0.3569933, 0.1815385, 0.1149544, 
    0.1441748, 0.2417017, 0.3825119, 0.3452537, 0.3218261, 0.3594121, 
    0.2309686, 0.2220787, 0.2118017, 0.2287657, 0.2035618, 0.3491522, 
    0.2663588, 0.3823791, 0.2601198, 0.2144413, 0.2492591,
  0.2542658, 0.2184418, 0.1883169, 0.210998, 0.1946429, 0.2740409, 0.2773771, 
    0.3419269, 0.30922, 0.2842765, 0.1066059, 0.1932359, 0.2032051, 0.213332, 
    0.1360466, 0.1529445, 0.3060839, 0.2929683, 0.2573502, 0.203694, 
    0.1307551, 0.1094475, 0.07534919, 0.07386328, 0.1697217, 0.08030545, 
    0.01710501, 0.1990215, 0.1677332,
  0.2126245, 0.2388243, 0.2260815, 0.232146, 0.2026079, 0.1615855, 0.167774, 
    0.1821997, 0.1348453, 0.1231497, 0.1625991, 0.1458308, 0.1294505, 
    0.2002507, 0.2784401, 0.2545168, 0.2518737, 0.1572326, 0.1341778, 
    0.1109068, 0.09704809, 0.1607668, 0.1456892, 0.04181151, 0.06934274, 
    0.01546086, 0.08978442, 0.2883634, 0.2257819,
  0.06676793, 0.06918348, 0.07159902, 0.07401457, 0.07643011, 0.07884566, 
    0.0812612, 0.08234894, 0.08538918, 0.08842944, 0.09146969, 0.09450994, 
    0.09755019, 0.1005904, 0.106934, 0.1069954, 0.1070569, 0.1071183, 
    0.1071797, 0.1072411, 0.1073025, 0.1020845, 0.09656728, 0.09105007, 
    0.08553284, 0.08001563, 0.07449841, 0.06898119, 0.06483549,
  0.1666038, 0.09632391, 0.02008725, 0.0002769304, 0.004431889, 0.002232981, 
    -0.0005397892, 0.01043795, 0.02486699, 0.1096328, 0.06439686, 0.05701457, 
    0.06428157, 0.1218027, 0.1554894, 0.1635819, 0.1882309, 0.3225642, 
    0.3200866, 0.2503216, 0.1874873, 0.2190688, 0.2042419, 0.005906682, 
    0.004970141, -0.001547754, 0.08328877, 0.2692035, 0.1184008,
  0.1722044, 0.1831038, 0.2429018, 0.166071, 0.09113974, 0.1600168, 
    0.2592411, 0.3405371, 0.303099, 0.2167312, 0.2594096, 0.2382415, 
    0.1632498, 0.1804416, 0.2245801, 0.2450228, 0.3223482, 0.3618801, 
    0.2012757, 0.3461074, 0.421149, 0.4381615, 0.3578915, 0.347929, 
    0.2872396, 0.2002481, 0.1035908, 0.2176128, 0.2577813,
  0.3050974, 0.3515529, 0.273958, 0.414219, 0.3419111, 0.248099, 0.2602169, 
    0.2952822, 0.2690804, 0.2713926, 0.2203773, 0.246436, 0.2463488, 
    0.2602892, 0.1689903, 0.1779581, 0.1993373, 0.2127888, 0.2598681, 
    0.2788137, 0.2522727, 0.2507814, 0.2103946, 0.2245389, 0.2208398, 
    0.24406, 0.2297618, 0.252884, 0.2872166,
  0.224015, 0.1932806, 0.2480963, 0.2272701, 0.2403374, 0.232598, 0.1284632, 
    0.09538449, 0.08167763, 0.123823, 0.1552436, 0.1723704, 0.1276152, 
    0.1896131, 0.1384406, 0.09722453, 0.07475821, 0.09828956, 0.1065261, 
    0.1377902, 0.1693909, 0.2084923, 0.1453849, 0.1495505, 0.1128009, 
    0.0916787, 0.09924959, 0.1182148, 0.1777969,
  0.0590514, 0.007634294, 0.02008161, 0.0890739, 0.02088811, 0.04435395, 
    0.04098965, 0.04507167, 0.05553244, 0.002913671, 0.02610103, 0.0684013, 
    0.09260022, 0.08530378, 0.05426139, 0.008051851, 0.05113149, 0.08811899, 
    0.2195314, 0.1664866, 0.03641648, 0.05812661, 0.0123509, 0.02184326, 
    0.06789922, 0.1292997, 0.1033056, 0.08806325, 0.07586994,
  0.006813414, 0.004805761, 0.1384957, 0.02274327, 0.02559296, 0.0881062, 
    0.03659473, 0.05316469, 8.650573e-06, 0.005074202, 0.007738451, 
    0.03383667, 0.07410157, 0.004518854, 0.03037124, 0.1058298, 0.05389721, 
    0.1050086, 0.1449753, 0.008820035, 0.03124945, 0.0005054965, 
    5.792413e-07, 0.000675682, 0.07152397, 0.09312888, 0.1842609, 0.02095333, 
    0.001235074,
  0.001916265, 0.07331746, 0.1409594, 0.09704486, 0.1270538, 0.05382936, 
    0.09969218, 0.003704059, 6.146884e-07, 0.04694447, 0.07368708, 0.1684232, 
    0.1593412, 0.03550485, 0.04536294, 0.2467533, 0.2193141, 0.1803214, 
    0.02865344, 0.006321633, 0.0001357204, 1.809235e-07, 5.807859e-06, 
    0.0006822113, 0.1912085, 0.08662624, 0.01024957, -5.904191e-06, 
    2.401297e-07,
  0.002092152, 0.04789196, 0.3407015, 0.178087, 0.08111935, 0.03578197, 
    0.03633499, 0.03342351, 0.01627628, 0.1457827, 0.09743449, 0.04500821, 
    0.07263371, 0.06111022, 0.1122946, 0.05309707, 0.05301547, 0.01702979, 
    0.003068962, 0.0007866661, 5.604467e-08, 8.516496e-06, 9.370301e-05, 
    0.1605975, 0.3490432, 0.222514, 0.008460688, 0.0001614302, 0.006490735,
  0.1166, 0.1046378, 0.06041952, 0.02142248, 0.01224161, 0.09491877, 
    0.1361185, 0.01995468, 0.08127686, 0.2581648, 0.1223253, 0.088213, 
    0.08158936, 0.1295018, 0.0762701, 0.002755521, 0.0110137, -0.0004010891, 
    -1.822192e-05, 5.802278e-05, 0.0007092311, 0.06651459, 0.1270839, 
    0.09486702, 0.149115, 0.1827255, 0.05098118, 0.003260744, 0.05381751,
  2.92141e-07, 7.418731e-05, 0.0006521019, 0.03424929, 0.04430746, 
    0.02460953, 0.0327054, 0.06705, 0.01139203, 0.04919651, 0.05718983, 
    0.07710302, 0.07733995, 0.02099039, 0.03992634, 0.02566882, 0.06750469, 
    0.007410541, 0.04496171, 0.044564, 0.07195379, 0.009059415, 0.02025687, 
    0.008579046, 0.005925893, 0.002345054, 0.0001483515, -8.399607e-05, 
    0.02535833,
  3.867787e-06, 1.085862e-06, 3.167215e-10, 0.002875712, 9.466992e-07, 
    2.355632e-07, 0.02765338, 0.02253434, 0.000231072, 0.04766236, 
    0.02581276, 0.07463957, 0.0299725, 1.353331e-05, 0.001342624, 
    0.002481018, 0.06210269, 0.006890415, 0.0001323701, 0.1209179, 
    0.05908505, 0.04200923, 0.02439906, 0.004683778, 0.03135899, 0.08086934, 
    7.260762e-06, 0.002446759, 0.05107804,
  -1.929057e-05, 1.189968e-06, 0.01770964, 0.01380931, 0.05098195, 
    0.003739693, 0.002207872, 0.0003711558, 0.1434329, 0.1478024, 0.07828269, 
    0.06990758, 0.06235902, 0.1284403, 0.1350719, 0.09710626, 0.06809777, 
    0.1201573, 0.01834407, 0.0200939, 0.09452194, 0.09120688, 0.08032245, 
    0.04474055, 0.03598941, 0.07113089, 0.03207671, 0.007578512, 0.04487718,
  0.0265921, 0.006441454, 0.1491826, 0.3355065, 0.109996, 0.07844316, 
    0.2002652, 0.06597862, 0.03957572, 0.04904275, 0.04739637, 0.10374, 
    0.1211354, 0.1500618, 0.2187232, 0.2055568, 0.2094454, 0.2135765, 
    0.08493436, 0.194615, 0.1938349, 0.09990392, 0.2153577, 0.1612826, 
    0.1646341, 0.2062556, 0.1876866, 0.1018176, 0.05671624,
  0.1724554, 0.1889832, 0.165475, 0.1488736, 0.1325432, 0.2267556, 0.1828104, 
    0.1826193, 0.1797606, 0.04812019, 0.07421716, 0.1901144, 0.2302964, 
    0.1554849, 0.3041489, 0.2489728, 0.1656705, 0.1448485, 0.08867806, 
    0.121366, 0.1755642, 0.1757075, 0.3248204, 0.3229237, 0.2552686, 
    0.2129212, 0.1786297, 0.1839895, 0.2267243,
  0.2223528, 0.159659, 0.2460206, 0.3443816, 0.2131509, 0.2736176, 0.3092788, 
    0.3357698, 0.3023224, 0.38487, 0.1769219, 0.1260384, 0.1439644, 
    0.2625588, 0.3762615, 0.3232638, 0.294906, 0.3516252, 0.2306623, 
    0.2114253, 0.2249781, 0.2358243, 0.2661448, 0.3876658, 0.2570555, 
    0.3658559, 0.2940918, 0.2367063, 0.2504884,
  0.2694739, 0.2176912, 0.1967342, 0.2383914, 0.2187493, 0.2910482, 
    0.2921088, 0.3564642, 0.3272808, 0.2952143, 0.1464674, 0.1893712, 
    0.2041527, 0.2073267, 0.1267711, 0.1507154, 0.2978199, 0.2910305, 
    0.2039383, 0.1967695, 0.1174413, 0.1312545, 0.08205742, 0.1199125, 
    0.1630699, 0.142667, 0.03043935, 0.2193841, 0.1632476,
  0.1869224, 0.2319211, 0.2185379, 0.2403851, 0.2096718, 0.1594562, 
    0.1628232, 0.1918942, 0.1519784, 0.1384136, 0.1888514, 0.1832285, 
    0.1450381, 0.2133953, 0.2872928, 0.2964521, 0.2599886, 0.1528143, 
    0.1272704, 0.1015557, 0.1022572, 0.1977243, 0.2002384, 0.04199034, 
    0.07479598, 0.06425337, 0.1762602, 0.2836207, 0.2213718,
  0.04636255, 0.05091704, 0.05547153, 0.06002602, 0.06458051, 0.069135, 
    0.07368949, 0.08832121, 0.0957183, 0.1031154, 0.1105125, 0.1179096, 
    0.1253067, 0.1327038, 0.1522309, 0.1485088, 0.1447868, 0.1410647, 
    0.1373427, 0.1336207, 0.1298987, 0.09334355, 0.08511399, 0.07688444, 
    0.06865489, 0.06042534, 0.05219579, 0.04396624, 0.04271896,
  0.1564192, 0.1190029, 0.04933016, 0.02114604, 0.0119794, 0.0384131, 
    0.06573766, 0.08669979, 0.1880226, 0.2085327, 0.119125, 0.04618651, 
    0.06296001, 0.1541163, 0.2122802, 0.283447, 0.166394, 0.3586856, 
    0.2742024, 0.2794311, 0.2197946, 0.2617297, 0.1928905, 0.006133667, 
    0.01157107, 0.04046717, 0.07918394, 0.2318075, 0.1183413,
  0.1680184, 0.1865493, 0.2596527, 0.1986227, 0.109736, 0.1790098, 0.2960904, 
    0.337687, 0.2997101, 0.2602492, 0.254746, 0.2304787, 0.1823407, 
    0.1571058, 0.2362681, 0.2393972, 0.2926064, 0.3537682, 0.2366032, 
    0.4557706, 0.4507198, 0.4329666, 0.3078437, 0.3468957, 0.2516387, 
    0.1949964, 0.1303472, 0.2861436, 0.3257783,
  0.3236667, 0.340821, 0.2886424, 0.4078039, 0.3726152, 0.2845697, 0.2589881, 
    0.3434716, 0.2507022, 0.3520158, 0.3104037, 0.2944422, 0.2741885, 
    0.2807105, 0.2144984, 0.1707137, 0.1815764, 0.166266, 0.2613782, 
    0.2610728, 0.2476617, 0.2755476, 0.225596, 0.2393552, 0.2609703, 
    0.230023, 0.2471845, 0.3128465, 0.3258871,
  0.2018831, 0.2065071, 0.2214849, 0.2335714, 0.2255507, 0.2289385, 
    0.1373356, 0.09118553, 0.1033786, 0.1272798, 0.1585927, 0.1603895, 
    0.1319201, 0.1968899, 0.1519823, 0.1042638, 0.07106154, 0.1130133, 
    0.1090783, 0.1372831, 0.2037048, 0.2205468, 0.1647991, 0.1551186, 
    0.1033088, 0.1229614, 0.1181475, 0.1245503, 0.1761283,
  0.05873837, 0.008186776, 0.01932593, 0.09177685, 0.02389111, 0.04296333, 
    0.05200246, 0.06017088, 0.02190248, 0.001981432, 0.0227928, 0.06850969, 
    0.1025427, 0.1012042, 0.06908366, 0.02062911, 0.05706968, 0.06655648, 
    0.2092559, 0.1714475, 0.04981731, 0.06110613, 0.01062813, 0.01611761, 
    0.0666025, 0.1399009, 0.1105099, 0.1012462, 0.08841947,
  0.01160098, 0.006068198, 0.141949, 0.03057665, 0.02215813, 0.07790339, 
    0.04154161, 0.02534018, 1.466599e-05, 0.001247982, 0.0004876083, 
    0.02285096, 0.08564074, 0.01741771, 0.03536794, 0.1006967, 0.0544941, 
    0.111309, 0.1301109, 0.01469049, 0.03338342, 0.001323359, 1.077047e-06, 
    0.003851952, 0.0652619, 0.07569721, 0.1747225, 0.02978351, 0.004082859,
  0.0007834738, 0.06438642, 0.1600779, 0.08472367, 0.1048337, 0.04835239, 
    0.07739464, 0.001171576, 4.528951e-07, 0.03492301, 0.0564738, 0.1377762, 
    0.1572825, 0.03313165, 0.04512671, 0.2344391, 0.1919165, 0.1665924, 
    0.02605611, 0.009516073, 0.0001673496, -1.741731e-08, 2.944487e-06, 
    0.0003453274, 0.1448825, 0.104046, 0.02446227, 8.441633e-05, 1.241533e-07,
  2.519382e-06, 0.01471908, 0.3818663, 0.1281018, 0.07638645, 0.0347465, 
    0.03438554, 0.04132566, 0.009107078, 0.1218597, 0.08591132, 0.03569456, 
    0.06106333, 0.05817046, 0.1105137, 0.05973463, 0.0529009, 0.01950855, 
    0.004002003, 0.001308253, 5.173271e-08, 1.87712e-06, 2.88373e-05, 
    0.1077057, 0.2468247, 0.1737566, 0.01557786, 0.0002475725, 0.0002768705,
  0.04491765, 0.03855392, 0.04820703, 0.02608003, 0.01262757, 0.09536052, 
    0.1341759, 0.022654, 0.06744125, 0.2456751, 0.1182779, 0.06721065, 
    0.06342693, 0.1044409, 0.06995829, 0.003623851, 0.01824316, 
    -0.0003789036, -3.861256e-06, 0.00174772, 9.190003e-05, 0.04917572, 
    0.1515596, 0.06481598, 0.1122504, 0.1495619, 0.05363351, 0.006578053, 
    0.02809341,
  2.587333e-07, 2.60608e-06, 2.406038e-05, 0.1507722, 0.0396424, 0.02316713, 
    0.03280723, 0.05614952, 0.01776446, 0.0522586, 0.07593454, 0.07316907, 
    0.07174355, 0.03031164, 0.04799515, 0.0217782, 0.05517562, 0.01140987, 
    0.04962935, 0.04585785, 0.06636262, 0.02208526, 0.03521104, 0.01395115, 
    0.01021127, 0.001124513, 1.808395e-05, -0.0001521058, 0.03613413,
  1.994681e-06, 1.074455e-06, 1.756571e-09, 0.00440163, 0.003017694, 
    2.152955e-07, 0.04113914, 0.03409744, 0.0004902122, 0.04169328, 
    0.02551703, 0.06867627, 0.02328662, 0.0001670076, 0.003482168, 
    0.00427006, 0.05179088, 0.006587454, 0.001118275, 0.1067771, 0.03926329, 
    0.05205704, 0.01076424, 0.01231762, 0.03906227, 0.08106395, 5.798645e-05, 
    0.004229348, 0.04159173,
  -2.077273e-06, 2.187885e-06, 0.01939269, 0.01344038, 0.06862134, 
    0.004282289, 0.005047261, 0.004344792, 0.1626565, 0.1430974, 0.06375514, 
    0.0730556, 0.07855944, 0.1496076, 0.1326161, 0.09722864, 0.06746483, 
    0.1071956, 0.02253299, 0.02595093, 0.0817057, 0.07386597, 0.0930176, 
    0.05038212, 0.05935255, 0.07700263, 0.0336211, 0.01386446, 0.05215322,
  0.02604751, 0.00747336, 0.1580215, 0.3490702, 0.1201145, 0.06768377, 
    0.206538, 0.05867624, 0.0243423, 0.05555346, 0.04643831, 0.1053666, 
    0.1247443, 0.1604845, 0.2102461, 0.2061365, 0.2027305, 0.2142476, 
    0.1070299, 0.1883163, 0.2037854, 0.1119206, 0.2090706, 0.1663684, 
    0.1681841, 0.2179168, 0.2119917, 0.1008147, 0.04700178,
  0.185456, 0.210713, 0.1500216, 0.2275672, 0.1291815, 0.2203968, 0.1922092, 
    0.1795021, 0.1884681, 0.03643108, 0.05833866, 0.1744476, 0.2319937, 
    0.1826819, 0.3492546, 0.2700447, 0.1615281, 0.1465388, 0.08491018, 
    0.1339075, 0.2096411, 0.2006172, 0.3224108, 0.3112218, 0.2689256, 
    0.195603, 0.1782943, 0.1833038, 0.2243176,
  0.2489472, 0.1788881, 0.2388507, 0.305797, 0.2311941, 0.2770316, 0.2966268, 
    0.3394856, 0.2939425, 0.3676158, 0.1663686, 0.1175378, 0.1515211, 
    0.3156846, 0.4431048, 0.3180477, 0.2982619, 0.348226, 0.2186715, 
    0.2124961, 0.2151111, 0.2344019, 0.2862025, 0.3938736, 0.2765308, 
    0.3288276, 0.30615, 0.255647, 0.2358114,
  0.2786484, 0.2118153, 0.2000444, 0.2240128, 0.2110745, 0.2886723, 
    0.2868362, 0.3781513, 0.3343984, 0.2903768, 0.1788047, 0.1820847, 
    0.221005, 0.2013052, 0.1271855, 0.1583174, 0.3005137, 0.2844445, 
    0.1841035, 0.2163768, 0.111632, 0.1385312, 0.1010752, 0.1170491, 
    0.1597862, 0.238578, 0.05402385, 0.2421891, 0.1631598,
  0.1892894, 0.2304564, 0.1939931, 0.2129874, 0.1957117, 0.1663373, 
    0.1726752, 0.2351825, 0.2040866, 0.1799559, 0.2193677, 0.1830731, 
    0.1778259, 0.2112024, 0.2663243, 0.2684098, 0.2165227, 0.1426072, 
    0.1026271, 0.1123, 0.1201398, 0.2044238, 0.2013344, 0.04190604, 
    0.06672636, 0.06556269, 0.2325995, 0.277292, 0.2151298,
  0.03815215, 0.04370495, 0.04925775, 0.05481055, 0.06036334, 0.06591614, 
    0.07146894, 0.1006148, 0.1084965, 0.1163782, 0.1242599, 0.1321416, 
    0.1400232, 0.1479049, 0.1436778, 0.1393464, 0.1350149, 0.1306835, 
    0.1263521, 0.1220206, 0.1176892, 0.09102042, 0.08191738, 0.07281432, 
    0.06371128, 0.05460823, 0.04550518, 0.03640213, 0.03370991,
  0.1479255, 0.1209658, 0.1003359, 0.06759905, 0.06146624, 0.1089905, 
    0.1374907, 0.1857693, 0.1917482, 0.1895148, 0.08569284, 0.05616511, 
    0.09537951, 0.1182891, 0.1199385, 0.1653954, 0.2076752, 0.3255993, 
    0.29218, 0.2131736, 0.2155842, 0.2487866, 0.1855994, 0.0105156, 
    0.01472101, 0.05966963, 0.08263852, 0.1571436, 0.130851,
  0.2784761, 0.2992199, 0.1642722, 0.1811413, 0.1381662, 0.2355754, 
    0.2917787, 0.3507098, 0.2993472, 0.2851381, 0.2562228, 0.213828, 
    0.2240829, 0.1816635, 0.2173919, 0.3080906, 0.3053904, 0.3527225, 
    0.261592, 0.4839778, 0.5024377, 0.4337628, 0.3341796, 0.4314943, 
    0.3015004, 0.2172754, 0.1537719, 0.2260952, 0.2579228,
  0.3313066, 0.3507972, 0.4456265, 0.492603, 0.4182687, 0.3031326, 0.2761486, 
    0.3375911, 0.2738776, 0.4496047, 0.3665369, 0.3469701, 0.2836956, 
    0.3032588, 0.23839, 0.2033141, 0.2616165, 0.2262795, 0.2885267, 
    0.2975486, 0.2765286, 0.2588258, 0.239839, 0.2392491, 0.2353931, 
    0.1785454, 0.2337651, 0.2730613, 0.2815441,
  0.2081047, 0.2128004, 0.2854175, 0.2841569, 0.2423656, 0.2371362, 
    0.1454774, 0.1019675, 0.1135591, 0.1466094, 0.1959867, 0.1650662, 
    0.1672458, 0.1906462, 0.1747232, 0.1354224, 0.08989581, 0.1188934, 
    0.1257303, 0.1394055, 0.2304021, 0.2085405, 0.1752477, 0.1686538, 
    0.09687321, 0.1202212, 0.1263755, 0.1500509, 0.1755318,
  0.06677199, 0.01735813, 0.02849536, 0.1101923, 0.03240474, 0.04259422, 
    0.08092433, 0.1197238, 0.01394761, 0.002401486, 0.02865168, 0.06670272, 
    0.1059505, 0.108136, 0.08934217, 0.03936777, 0.0660441, 0.07679864, 
    0.1930464, 0.1504667, 0.05774401, 0.07046688, 0.02190593, 0.01988724, 
    0.06469113, 0.1447432, 0.1109803, 0.1001759, 0.09625331,
  0.01231977, 0.009547364, 0.1325593, 0.02708842, 0.02033454, 0.06532659, 
    0.04834294, 0.04668976, 1.341908e-05, 0.0001350183, -1.365721e-06, 
    0.009258963, 0.08609135, 0.02340811, 0.03431247, 0.08082492, 0.06972282, 
    0.1194962, 0.0871155, 0.01737143, 0.02257767, 0.005954892, 4.239236e-06, 
    0.003170648, 0.05682005, 0.06464158, 0.1748165, 0.03325313, 0.00746713,
  0.0005000128, 0.04364632, 0.1486558, 0.07707323, 0.1028108, 0.0490111, 
    0.0611956, 0.001673374, 1.244852e-06, 0.02546616, 0.04787065, 0.1352083, 
    0.1584312, 0.03426262, 0.04285651, 0.21491, 0.1717223, 0.1526369, 
    0.02701461, 0.02203269, 0.001335501, 0.0001789603, 1.167184e-06, 
    9.489764e-05, 0.1345723, 0.09199452, 0.04340059, 0.004420025, 3.394561e-06,
  -1.326843e-06, 0.01653186, 0.3432137, 0.08874987, 0.07001077, 0.03051494, 
    0.03387217, 0.041748, 0.01138531, 0.1041999, 0.07228903, 0.0283892, 
    0.05661145, 0.0513573, 0.1091897, 0.07374705, 0.05576274, 0.01746243, 
    0.008589709, 0.001833754, 5.214354e-08, 1.907419e-07, 6.323972e-06, 
    0.1028133, 0.2050994, 0.1279459, 0.02944342, 0.0002807842, 3.790437e-06,
  0.01931017, 0.01117296, 0.03851847, 0.05659272, 0.0153634, 0.1084507, 
    0.1358797, 0.02792387, 0.07639036, 0.2296546, 0.1110025, 0.05686563, 
    0.05860466, 0.09631453, 0.06556118, 0.003777954, 0.0177104, 
    -0.0004314342, 7.048564e-06, 0.0004579613, 0.00103288, 0.04342347, 
    0.1447377, 0.06113504, 0.1089906, 0.1317407, 0.05451712, 0.01621516, 
    0.02344335,
  1.33136e-07, 4.172374e-07, 1.968012e-05, 0.1963886, 0.04298356, 0.03555231, 
    0.03710767, 0.05529261, 0.03284758, 0.06355209, 0.08629835, 0.07958246, 
    0.06538622, 0.03792008, 0.05232859, 0.0277022, 0.04240936, 0.01089831, 
    0.03794638, 0.04711855, 0.06148065, 0.02739785, 0.05481831, 0.02337595, 
    0.03494633, 0.001370417, 9.178041e-06, 3.408298e-05, 0.03775334,
  1.408316e-06, 4.686893e-07, 6.567531e-10, 0.0110415, 0.03243378, 
    3.471126e-08, 0.04934887, 0.04713237, 0.004788955, 0.03356921, 
    0.03674185, 0.08557986, 0.0216392, 0.002029943, 0.0104347, 0.007597727, 
    0.04460616, 0.003891184, 0.002628405, 0.09502132, 0.01907927, 0.0623895, 
    0.006794206, 0.04283649, 0.04677582, 0.07892902, 0.0005248755, 
    0.002633143, 0.03460165,
  4.086269e-06, 1.371509e-06, 0.03439281, 0.02364553, 0.08573807, 
    0.007641859, 0.008456751, 0.0093623, 0.1817971, 0.1449655, 0.05657828, 
    0.1037499, 0.08303365, 0.1426565, 0.1220262, 0.1281133, 0.06950335, 
    0.1162589, 0.03243591, 0.03541972, 0.07361589, 0.06269513, 0.1038416, 
    0.05367811, 0.08730456, 0.08387333, 0.03973348, 0.01791819, 0.05333636,
  0.03677914, 0.01277454, 0.1620015, 0.3719418, 0.130441, 0.06533578, 
    0.2068284, 0.05199313, 0.0157251, 0.04774228, 0.03756498, 0.1031151, 
    0.1361749, 0.1927174, 0.2079062, 0.1990621, 0.2008684, 0.2058198, 
    0.1241699, 0.1892932, 0.2119169, 0.09826328, 0.1669438, 0.1539637, 
    0.1794188, 0.216534, 0.2196376, 0.1185095, 0.04058933,
  0.2128194, 0.2540875, 0.1793835, 0.2643247, 0.1205915, 0.2244957, 
    0.1765947, 0.1753261, 0.1691741, 0.03285972, 0.03391313, 0.1825096, 
    0.2250905, 0.1889718, 0.3331816, 0.2604981, 0.171637, 0.1548482, 
    0.09319877, 0.1504969, 0.1877163, 0.2024235, 0.3372377, 0.3388465, 
    0.2621948, 0.1849859, 0.1943818, 0.1828617, 0.2250934,
  0.2478331, 0.1773901, 0.3026501, 0.3130207, 0.269298, 0.2983055, 0.3062835, 
    0.3228319, 0.3034139, 0.4111356, 0.1768624, 0.1064108, 0.1728714, 
    0.2865482, 0.4581052, 0.3084273, 0.3203119, 0.3681409, 0.2253579, 
    0.2364782, 0.213148, 0.2118187, 0.263858, 0.3923551, 0.289553, 0.3312066, 
    0.3261544, 0.2616341, 0.2424355,
  0.2831326, 0.2435409, 0.2007233, 0.228125, 0.2146584, 0.3034233, 0.2776417, 
    0.399005, 0.346516, 0.2834793, 0.1828548, 0.1621549, 0.2133987, 
    0.1811404, 0.118714, 0.1186639, 0.3046023, 0.3026297, 0.1864562, 
    0.2422833, 0.129435, 0.1610567, 0.1184542, 0.1081079, 0.161502, 
    0.3074465, 0.1021804, 0.2651824, 0.1689463,
  0.1784895, 0.2517179, 0.2101902, 0.2659054, 0.2035916, 0.1575346, 
    0.2016582, 0.2490204, 0.1943142, 0.1676269, 0.217696, 0.1673883, 
    0.1752423, 0.2132749, 0.2570902, 0.2474536, 0.1911659, 0.128363, 
    0.08879177, 0.1201119, 0.1277124, 0.2035487, 0.1863903, 0.04461996, 
    0.05173483, 0.1162122, 0.2420011, 0.2659828, 0.2063806,
  0.04313901, 0.04795041, 0.05276182, 0.05757323, 0.06238464, 0.06719604, 
    0.07200745, 0.1002263, 0.1078436, 0.115461, 0.1230784, 0.1306957, 
    0.1383131, 0.1459305, 0.1600332, 0.1585507, 0.1570682, 0.1555857, 
    0.1541032, 0.1526207, 0.1511381, 0.108793, 0.09784669, 0.08690042, 
    0.07595415, 0.06500789, 0.05406162, 0.04311535, 0.03928988,
  0.1471429, 0.1154234, 0.08325859, 0.08779299, 0.128087, 0.2370825, 
    0.249563, 0.221829, 0.2146639, 0.2061987, 0.09048703, 0.09193125, 
    0.09545822, 0.08752573, 0.05333912, 0.1903336, 0.2144108, 0.2725341, 
    0.2376108, 0.1986455, 0.2086312, 0.2537494, 0.1619296, 0.06780565, 
    0.1009955, 0.149742, 0.04501764, 0.1106927, 0.1367955,
  0.2134129, 0.3048175, 0.1967411, 0.1642482, 0.1603865, 0.3088025, 
    0.2640958, 0.3658695, 0.2945846, 0.32419, 0.271563, 0.2064218, 0.1737764, 
    0.1708866, 0.2173809, 0.3639733, 0.2396402, 0.3613837, 0.2349646, 
    0.3937709, 0.4613776, 0.4579975, 0.3506403, 0.4758401, 0.2151723, 
    0.2226027, 0.1636565, 0.1942425, 0.2648542,
  0.3355843, 0.4136544, 0.3822647, 0.435703, 0.4517723, 0.382621, 0.3197154, 
    0.3324298, 0.2801973, 0.3244831, 0.387143, 0.3524439, 0.34231, 0.3073271, 
    0.249524, 0.2004543, 0.2688293, 0.2469153, 0.3119977, 0.3466507, 
    0.2889554, 0.2391783, 0.2269052, 0.2752781, 0.2926982, 0.1951221, 
    0.2732603, 0.3130358, 0.2895144,
  0.2341931, 0.2554357, 0.2977963, 0.2702729, 0.2402797, 0.2329479, 
    0.1504108, 0.1193364, 0.1426861, 0.1348054, 0.2094069, 0.1819481, 
    0.1854295, 0.1877362, 0.162126, 0.1196241, 0.1075234, 0.1264616, 
    0.1419728, 0.1743059, 0.2020478, 0.2294439, 0.1895409, 0.1853623, 
    0.07138443, 0.1061846, 0.1495147, 0.1344292, 0.1983069,
  0.06802858, 0.03364183, 0.03281781, 0.132896, 0.05567037, 0.03963193, 
    0.1078132, 0.1366046, 0.02667404, 0.002410934, 0.03396484, 0.06849363, 
    0.1071484, 0.1174817, 0.1073193, 0.04805699, 0.07513991, 0.1054436, 
    0.1840658, 0.1442323, 0.06656534, 0.06943376, 0.03107519, 0.02852213, 
    0.06066553, 0.1389066, 0.09964365, 0.1045708, 0.08899922,
  0.01193882, 0.009427506, 0.135465, 0.01931158, 0.02355761, 0.06655388, 
    0.0574991, 0.04996518, 4.62775e-05, -1.207333e-05, -3.831954e-05, 
    0.003571898, 0.0864455, 0.02798584, 0.03875633, 0.0651514, 0.06658101, 
    0.1221332, 0.07480556, 0.02642019, 0.01957018, 0.01877536, -4.315368e-06, 
    0.0002419282, 0.0485103, 0.06718241, 0.1542911, 0.04015952, 0.01589195,
  0.003900865, 0.0311873, 0.159297, 0.07932921, 0.1033562, 0.05454284, 
    0.06115615, 0.005518233, 0.0001416698, 0.02128497, 0.03589302, 0.127313, 
    0.1542175, 0.03313249, 0.04119154, 0.1806445, 0.1512272, 0.1436148, 
    0.02896265, 0.04378147, 0.01994149, 0.01058116, 3.33428e-07, 
    1.006183e-05, 0.1263609, 0.09057575, 0.05765409, 0.03892175, 0.002366767,
  4.052711e-06, 0.01788426, 0.344963, 0.06124798, 0.05641131, 0.02893524, 
    0.03596244, 0.03993241, 0.01468689, 0.09568095, 0.06485409, 0.02396915, 
    0.06367362, 0.04351008, 0.09446266, 0.06828019, 0.04841801, 0.02465351, 
    0.01797713, 0.007328177, -5.869516e-06, 8.768116e-07, -2.699443e-07, 
    0.1018981, 0.1799799, 0.1033036, 0.02858276, 0.000851839, 9.5562e-06,
  0.009691188, 0.007427421, 0.01664775, 0.07642769, 0.02118576, 0.1205367, 
    0.1477955, 0.02948067, 0.1051368, 0.2186201, 0.09789427, 0.05072483, 
    0.05399926, 0.09918601, 0.0625599, 0.00608996, 0.01850719, -0.0003978935, 
    0.0004745599, 0.0019361, 0.002159058, 0.04509307, 0.1230436, 0.06502192, 
    0.1122057, 0.1196268, 0.04894855, 0.0208124, 0.02293538,
  4.812372e-08, 1.243552e-07, -4.941318e-06, 0.1211477, 0.05803182, 
    0.04142212, 0.04685382, 0.04271204, 0.04472923, 0.0729, 0.09279997, 
    0.08406466, 0.06468023, 0.04752839, 0.05094773, 0.03396408, 0.03992774, 
    0.01514111, 0.0407222, 0.04712622, 0.05918382, 0.03038907, 0.07630023, 
    0.0315629, 0.04209807, 0.003841665, 2.668363e-05, -1.101133e-05, 
    0.03123312,
  1.639189e-06, 8.980626e-08, -8.272828e-07, 0.02631133, 0.001048635, 
    6.146513e-06, 0.04396813, 0.0562984, 0.02081659, 0.05014805, 0.09305936, 
    0.08520287, 0.0373553, 0.00743893, 0.02444822, 0.01337308, 0.04879335, 
    0.009790263, 0.006564801, 0.08889443, 0.004543141, 0.09792326, 
    0.01080165, 0.05953602, 0.06283468, 0.07252564, 0.002256842, 0.002955257, 
    0.02482976,
  4.858206e-06, -7.318097e-05, 0.03724163, 0.03090523, 0.08907459, 
    0.01120063, 0.002034255, 0.01130184, 0.1846007, 0.1345835, 0.05320163, 
    0.1391351, 0.09497033, 0.1388079, 0.1190544, 0.1422483, 0.09010311, 
    0.1190065, 0.054325, 0.03931333, 0.06636477, 0.05900685, 0.1145079, 
    0.06448188, 0.08794685, 0.07948729, 0.0402427, 0.02739754, 0.03652965,
  0.03302725, 0.02456896, 0.1515038, 0.3958747, 0.1440818, 0.08152931, 
    0.2054885, 0.0406462, 0.01025678, 0.0346665, 0.03389569, 0.111553, 
    0.1513897, 0.2046259, 0.2191647, 0.1973602, 0.2038665, 0.193646, 
    0.1373443, 0.1899314, 0.2067878, 0.0912863, 0.1491521, 0.1557775, 
    0.2098679, 0.2143274, 0.2314356, 0.1517906, 0.05953078,
  0.2367983, 0.2788066, 0.1951797, 0.2873721, 0.1285804, 0.2012302, 
    0.1603753, 0.1791348, 0.1452667, 0.02707786, 0.01836258, 0.2003506, 
    0.278853, 0.2562682, 0.3508328, 0.2942377, 0.16231, 0.1750826, 
    0.09621009, 0.1781723, 0.1806535, 0.180466, 0.2883376, 0.3422821, 
    0.256202, 0.2307947, 0.2164048, 0.1835772, 0.2358188,
  0.2414021, 0.1710763, 0.2738682, 0.2882674, 0.2574304, 0.3025423, 
    0.3211245, 0.3154222, 0.2922001, 0.4152224, 0.2173871, 0.08851418, 
    0.207408, 0.2688412, 0.4391693, 0.2908333, 0.3185681, 0.3689824, 
    0.2270745, 0.2082159, 0.178301, 0.2254797, 0.2543099, 0.3577679, 
    0.2874682, 0.3486065, 0.3314869, 0.2647345, 0.2553129,
  0.2823807, 0.2869658, 0.179779, 0.3166776, 0.3036698, 0.2829834, 0.2590097, 
    0.4031059, 0.3505748, 0.2827092, 0.1845493, 0.1634611, 0.2066078, 
    0.1941621, 0.09540451, 0.1145424, 0.2946725, 0.2985267, 0.2301981, 
    0.1997875, 0.1932562, 0.1472854, 0.1231683, 0.1060792, 0.1785173, 
    0.3895253, 0.1382521, 0.2910056, 0.2004076,
  0.1596985, 0.2128875, 0.1975848, 0.2613043, 0.1718934, 0.1558774, 
    0.2021611, 0.2835094, 0.1943239, 0.1647647, 0.1992918, 0.1610836, 
    0.1769592, 0.2164117, 0.2446064, 0.2292696, 0.179779, 0.1124436, 
    0.07841717, 0.1554316, 0.1445892, 0.1901709, 0.1909173, 0.05048364, 
    0.04432348, 0.121594, 0.245144, 0.2456072, 0.1831709,
  0.02838382, 0.03280894, 0.03723406, 0.04165919, 0.04608431, 0.05050944, 
    0.05493456, 0.08603474, 0.09322954, 0.1004243, 0.1076191, 0.1148139, 
    0.1220087, 0.1292035, 0.1399237, 0.1380192, 0.1361148, 0.1342104, 
    0.1323059, 0.1304015, 0.1284971, 0.07980661, 0.07009112, 0.06037563, 
    0.05066015, 0.04094466, 0.03122917, 0.02151368, 0.02484372,
  0.156526, 0.1384603, 0.08720683, 0.08259605, 0.1438297, 0.2694138, 
    0.292828, 0.2327532, 0.2187762, 0.247786, 0.109183, 0.08661935, 
    0.09440725, 0.02135051, 0.02382163, 0.07774719, 0.1043385, 0.1932136, 
    0.1692968, 0.1837655, 0.2304762, 0.2189973, 0.1528479, 0.02666691, 
    0.2028385, 0.2654713, 0.1381306, 0.1206043, 0.1581055,
  0.1304656, 0.1582567, 0.1493654, 0.1794456, 0.1408045, 0.3561797, 
    0.2530911, 0.3784778, 0.3081481, 0.3245194, 0.2761832, 0.1805744, 
    0.2047363, 0.1444166, 0.2176814, 0.3078249, 0.2999102, 0.33813, 
    0.2225838, 0.3271168, 0.3459898, 0.3825317, 0.4083745, 0.4793751, 
    0.1688136, 0.1622336, 0.2011077, 0.2127777, 0.3031,
  0.3376417, 0.4058074, 0.3117507, 0.3696671, 0.3420419, 0.2848943, 
    0.3169922, 0.3343218, 0.2617244, 0.3186511, 0.3170518, 0.337068, 
    0.3234273, 0.299753, 0.2359829, 0.1920472, 0.2422545, 0.2220839, 
    0.3001357, 0.3377009, 0.2670387, 0.2278622, 0.2428131, 0.2712646, 
    0.2739963, 0.1948607, 0.2779715, 0.2934377, 0.2972218,
  0.2217022, 0.2656694, 0.2768276, 0.2495218, 0.2579494, 0.2506015, 
    0.1716653, 0.125506, 0.1526427, 0.1630472, 0.2458457, 0.2129495, 
    0.2022686, 0.1860527, 0.1472994, 0.1244823, 0.09730717, 0.1465614, 
    0.1309244, 0.2052334, 0.2070821, 0.2039199, 0.2217819, 0.1765409, 
    0.07939473, 0.1063017, 0.1232834, 0.1285386, 0.2037005,
  0.08874545, 0.06840724, 0.04681251, 0.1464273, 0.0803552, 0.05194298, 
    0.1054728, 0.1032746, 0.02237015, 0.000782975, 0.03572125, 0.08075496, 
    0.108035, 0.1344722, 0.1362827, 0.07026257, 0.09190524, 0.1267967, 
    0.1745851, 0.1613624, 0.08116839, 0.0724223, 0.05905892, 0.03465282, 
    0.05172741, 0.1339931, 0.1073188, 0.1005063, 0.10227,
  0.01034501, 0.001026537, 0.1224121, 0.01521446, 0.03061986, 0.06573088, 
    0.06991663, 0.07132046, 0.000122832, 3.679227e-07, -0.0002378726, 
    0.0007116707, 0.07045529, 0.0304816, 0.05020013, 0.07409575, 0.07087067, 
    0.1314278, 0.07361796, 0.03706649, 0.03797222, 0.04332943, 0.002507879, 
    1.168159e-05, 0.04133033, 0.06355488, 0.1468974, 0.05738308, 0.0276424,
  0.003584852, 0.01879257, 0.1867259, 0.08135588, 0.09667419, 0.06082043, 
    0.07467224, 0.00697116, 0.004001345, 0.0273564, 0.03242166, 0.09882466, 
    0.1478855, 0.03840961, 0.04050069, 0.1393922, 0.1328333, 0.124289, 
    0.02637625, 0.04659385, 0.06926162, 0.03611684, -1.251558e-05, 
    5.920092e-05, 0.1185303, 0.08575106, 0.0334502, 0.07043555, 0.0239877,
  0.0008965685, 0.02077418, 0.3349177, 0.05183986, 0.04357874, 0.02375364, 
    0.03782149, 0.03828588, 0.01639865, 0.08479724, 0.06152181, 0.01930263, 
    0.05685597, 0.03496476, 0.07217639, 0.05705304, 0.03879419, 0.02056366, 
    0.02130084, 0.0177793, -0.0001512233, 0.0001219761, 1.796858e-06, 
    0.08847807, 0.1500438, 0.08632017, 0.02682324, 0.002706615, 0.000737351,
  0.004283424, 0.01061667, 0.00427008, 0.05458628, 0.02879265, 0.1202991, 
    0.1464875, 0.02847138, 0.1209866, 0.2233122, 0.09191611, 0.04210158, 
    0.04184672, 0.08595654, 0.0600018, 0.01041204, 0.02207139, 0.01240868, 
    0.001856587, 0.001797439, 0.01120062, 0.03171391, 0.09085, 0.07041413, 
    0.1120728, 0.1048991, 0.04182762, 0.02569588, 0.02379333,
  1.306017e-08, 2.885438e-08, -1.38953e-07, 0.06245732, 0.0633862, 
    0.05914776, 0.06449872, 0.03852313, 0.04130668, 0.07988768, 0.0988607, 
    0.07875038, 0.06131287, 0.05320064, 0.05141659, 0.03716808, 0.04090893, 
    0.02068966, 0.04723438, 0.04458472, 0.05460146, 0.03422111, 0.1143367, 
    0.03195746, 0.03338195, 0.01080729, 0.0003405146, 0.0001473421, 0.02543047,
  1.902425e-06, 2.400945e-08, -9.178122e-05, 0.05445088, -1.116267e-05, 
    0.001371572, 0.05137252, 0.05645778, 0.04545947, 0.1368779, 0.1117527, 
    0.09244288, 0.04710775, 0.02121067, 0.04792622, 0.01777366, 0.04988033, 
    0.01806283, 0.01141742, 0.08466343, 0.0009629357, 0.1455539, 0.01831985, 
    0.06966009, 0.06270697, 0.07485876, 0.01288305, 0.007715529, 0.01212734,
  6.639771e-06, 0.0007405287, 0.05789826, 0.03316603, 0.08113809, 0.0120874, 
    -0.0006051441, 0.01121156, 0.1677899, 0.1139806, 0.0815751, 0.1742471, 
    0.1217282, 0.1423545, 0.124533, 0.158792, 0.1099753, 0.106387, 
    0.08129416, 0.03493593, 0.08392751, 0.04427698, 0.1309783, 0.1020942, 
    0.09211725, 0.09019212, 0.05148383, 0.02908212, 0.0291835,
  0.04315514, 0.06108448, 0.1370117, 0.4360479, 0.1671324, 0.08469803, 
    0.1950919, 0.03380526, 0.005969508, 0.03119913, 0.03098398, 0.1565422, 
    0.1881744, 0.2142857, 0.2386514, 0.2108212, 0.2037721, 0.1786103, 
    0.1566742, 0.2051537, 0.1996247, 0.1120284, 0.1591699, 0.1744819, 
    0.2746286, 0.2264527, 0.2376052, 0.158129, 0.06002674,
  0.2075908, 0.288205, 0.2208142, 0.2197265, 0.1560662, 0.177788, 0.14891, 
    0.1807491, 0.1232129, 0.02252592, 0.0146009, 0.2104608, 0.3558055, 
    0.3508894, 0.3710145, 0.3225752, 0.1741148, 0.1964174, 0.1029829, 
    0.2115432, 0.2203051, 0.191084, 0.2635005, 0.3389256, 0.2542086, 
    0.2814201, 0.2177938, 0.2093348, 0.2512378,
  0.2360805, 0.1964085, 0.2384967, 0.2695375, 0.2582162, 0.2779691, 
    0.3065086, 0.3286389, 0.2916711, 0.3877427, 0.2306838, 0.07607361, 
    0.2124862, 0.2634557, 0.4483389, 0.252088, 0.3052597, 0.3744823, 
    0.2414619, 0.171772, 0.1801163, 0.2406134, 0.3066483, 0.3261448, 
    0.2818308, 0.3332114, 0.3528053, 0.2748003, 0.2428513,
  0.298331, 0.3232296, 0.1906135, 0.3410341, 0.2637371, 0.2833107, 0.2909034, 
    0.435169, 0.3516114, 0.2777691, 0.1862335, 0.1671828, 0.2080306, 
    0.214024, 0.1049737, 0.1047696, 0.3066977, 0.3074249, 0.2665567, 
    0.1861363, 0.2074524, 0.168048, 0.1310305, 0.1031649, 0.203855, 
    0.4267418, 0.152584, 0.2679381, 0.239501,
  0.1855396, 0.1974288, 0.2293974, 0.2881769, 0.2219016, 0.2102471, 
    0.2144484, 0.260499, 0.173224, 0.1955101, 0.1838987, 0.1822139, 
    0.2090356, 0.2504446, 0.235164, 0.2198181, 0.1825321, 0.111797, 
    0.09981754, 0.1680836, 0.1761621, 0.2151163, 0.1936962, 0.04339243, 
    0.05278134, 0.1036198, 0.2679854, 0.2747115, 0.2236067,
  0.01250187, 0.01664344, 0.02078501, 0.02492658, 0.02906815, 0.03320972, 
    0.03735129, 0.07491489, 0.08108246, 0.08725002, 0.09341758, 0.09958514, 
    0.1057527, 0.1119203, 0.1252989, 0.1232799, 0.1212609, 0.1192419, 
    0.1172229, 0.1152038, 0.1131848, 0.06858487, 0.06029474, 0.05200461, 
    0.04371448, 0.03542435, 0.02713422, 0.01884409, 0.009188617,
  0.1523077, 0.1374102, 0.09571946, 0.07108313, 0.1674342, 0.2826901, 
    0.3005965, 0.2445621, 0.2216648, 0.2407615, 0.1532508, 0.09494039, 
    0.1197843, 0.001916072, 0.1262103, 0.06404095, 0.1547353, 0.1659153, 
    0.1608444, 0.1640504, 0.2405418, 0.2245385, 0.1522655, 0.0767808, 
    0.2760775, 0.2290696, 0.05293286, 0.1016031, 0.2002714,
  0.1836055, 0.1796128, 0.1690653, 0.1014117, 0.1624694, 0.3541366, 
    0.2023522, 0.384359, 0.3208659, 0.2937927, 0.3014053, 0.1940877, 
    0.2044688, 0.1534699, 0.2563842, 0.3671042, 0.3144801, 0.3281015, 
    0.2056552, 0.3549773, 0.3849514, 0.3649594, 0.2803618, 0.4800907, 
    0.1503523, 0.1560918, 0.2003749, 0.3697711, 0.3450359,
  0.3579414, 0.4267775, 0.3442522, 0.3596736, 0.3198142, 0.2947102, 
    0.3583679, 0.343588, 0.3238208, 0.3572682, 0.3347389, 0.3090007, 
    0.2901076, 0.3261411, 0.2611983, 0.2021606, 0.2527299, 0.2355858, 
    0.3176822, 0.3753366, 0.2843635, 0.2354675, 0.279506, 0.2964348, 
    0.2929884, 0.1980164, 0.2818896, 0.3394901, 0.34216,
  0.2678378, 0.2985987, 0.271189, 0.2778758, 0.2742055, 0.2649385, 0.190183, 
    0.1607586, 0.1593813, 0.1823829, 0.2846797, 0.2314384, 0.2326768, 
    0.2032088, 0.1404375, 0.13331, 0.1204392, 0.206994, 0.1609645, 0.2660222, 
    0.226582, 0.2336647, 0.2452061, 0.165198, 0.06651511, 0.1154407, 
    0.1202381, 0.1444807, 0.238067,
  0.1386184, 0.1060135, 0.092791, 0.2020922, 0.1269403, 0.1009388, 0.12817, 
    0.129306, 0.04626457, 0.003549196, 0.05265213, 0.1238965, 0.1076821, 
    0.1329239, 0.1533816, 0.08748158, 0.1150284, 0.1535166, 0.1903743, 
    0.1837885, 0.1105983, 0.09692461, 0.1396624, 0.03981093, 0.04691776, 
    0.1372419, 0.1156149, 0.1005837, 0.1199532,
  0.03219904, 0.00380839, 0.1297243, 0.03039216, 0.03985194, 0.07062241, 
    0.08255842, 0.07997843, 0.0102955, 3.272327e-07, -0.0001468889, 
    -6.107332e-06, 0.07393109, 0.08553118, 0.06324678, 0.07837441, 
    0.07605642, 0.1621298, 0.0670242, 0.04561966, 0.07086254, 0.05948518, 
    0.026562, -2.828297e-05, 0.04139759, 0.05689277, 0.1402946, 0.06319503, 
    0.0508393,
  0.01748804, 0.02527803, 0.1877194, 0.08387319, 0.08913612, 0.05934633, 
    0.06790005, 0.01497681, 0.01368091, 0.04839328, 0.02877609, 0.07868554, 
    0.1258713, 0.03438907, 0.03879279, 0.1128569, 0.1208295, 0.1070435, 
    0.02538612, 0.03100868, 0.07547205, 0.07189203, 0.001317187, 
    0.0002350267, 0.1236474, 0.09810222, 0.02630864, 0.05006883, 0.06355812,
  0.01057766, 0.01649489, 0.3047338, 0.05076953, 0.03489883, 0.02179204, 
    0.03541126, 0.04328826, 0.01937339, 0.07234304, 0.06497788, 0.01601477, 
    0.05458625, 0.02852643, 0.05276607, 0.03884815, 0.03342277, 0.01962896, 
    0.02016989, 0.0362269, 0.009884449, 0.004718903, 0.0001677465, 
    0.07926258, 0.1174338, 0.07119285, 0.03117649, 0.004842915, 0.006045558,
  0.005533406, 0.01260303, 0.002156494, 0.03883374, 0.02605428, 0.09993733, 
    0.134216, 0.02510215, 0.1106089, 0.2337932, 0.0865438, 0.03199543, 
    0.03367704, 0.07279532, 0.05890618, 0.01442299, 0.02447712, 0.01887087, 
    0.005479794, 0.002739379, 0.01477362, 0.02945662, 0.05602524, 0.07369272, 
    0.09578012, 0.09045532, 0.03813222, 0.02436426, 0.02002836,
  3.679181e-09, 8.285866e-09, 1.563038e-08, 0.02639502, 0.09573945, 
    0.08831863, 0.06690106, 0.04332374, 0.06199627, 0.07088742, 0.1040154, 
    0.07393926, 0.05334246, 0.05659771, 0.05096157, 0.03921131, 0.03895959, 
    0.02465387, 0.0528104, 0.03989252, 0.04270139, 0.02383944, 0.1406168, 
    0.03470861, 0.03087694, 0.02090416, 0.007031674, 9.974078e-05, 0.02005734,
  6.506774e-07, 8.333149e-09, 0.0009257719, 0.06256389, -2.003137e-05, 
    0.04686096, 0.0539808, 0.06341256, 0.06718194, 0.2189305, 0.1122847, 
    0.1259914, 0.06231421, 0.04072481, 0.08575591, 0.0429617, 0.04513332, 
    0.03503432, 0.03364132, 0.0771499, 0.0006315839, 0.1801622, 0.02103279, 
    0.05970716, 0.06115568, 0.07372079, 0.05369153, 0.01968948, 0.001654423,
  4.299367e-06, 0.004091553, 0.08628905, 0.04620408, 0.0793177, 0.005974504, 
    -0.0006383361, 0.01160057, 0.1546221, 0.1005486, 0.1553912, 0.2251362, 
    0.1383988, 0.1536623, 0.1516134, 0.1827987, 0.1184551, 0.09492587, 
    0.128368, 0.04907117, 0.1089211, 0.0567971, 0.1188829, 0.1488235, 
    0.1096249, 0.1070522, 0.06519512, 0.03747987, 0.0218247,
  0.04293137, 0.05883026, 0.1265424, 0.444956, 0.1530191, 0.09166306, 
    0.1721908, 0.02195019, 0.008573901, 0.03233677, 0.03111907, 0.2639959, 
    0.2784631, 0.1957208, 0.2314641, 0.2435732, 0.2315427, 0.180265, 
    0.213162, 0.2289837, 0.2311133, 0.1328299, 0.190075, 0.2440992, 
    0.3498008, 0.2321902, 0.2815446, 0.1860582, 0.06939648,
  0.2140564, 0.265346, 0.274835, 0.2117474, 0.1460136, 0.1970774, 0.1580616, 
    0.177164, 0.1140838, 0.01990243, 0.02139596, 0.2009272, 0.44713, 
    0.4199205, 0.393039, 0.3425777, 0.2115237, 0.2322186, 0.1288546, 
    0.2096188, 0.228369, 0.2169938, 0.2921579, 0.3208185, 0.30399, 0.3412917, 
    0.2298881, 0.21831, 0.2561604,
  0.2416181, 0.1790064, 0.2597195, 0.2878399, 0.2756378, 0.2507275, 0.351608, 
    0.3384143, 0.2975365, 0.4093087, 0.2549196, 0.06357256, 0.204819, 
    0.2955868, 0.462106, 0.2528944, 0.3288588, 0.3941112, 0.2694201, 
    0.1554243, 0.1973043, 0.2681874, 0.2830149, 0.3406669, 0.3133213, 
    0.3079183, 0.3538356, 0.299897, 0.241284,
  0.3514604, 0.3436061, 0.2654279, 0.2938073, 0.273313, 0.3315898, 0.3230041, 
    0.4541564, 0.3652199, 0.3300999, 0.1886037, 0.1673775, 0.2095442, 
    0.2557842, 0.1094, 0.1007001, 0.3226927, 0.3316779, 0.2633435, 0.1916551, 
    0.2266726, 0.18217, 0.1440554, 0.0886335, 0.1829574, 0.4389194, 
    0.1679611, 0.2563126, 0.2982826,
  0.223918, 0.1975764, 0.2360576, 0.2987718, 0.2352368, 0.2309062, 0.2060738, 
    0.2407793, 0.1661807, 0.2100078, 0.191183, 0.1858982, 0.2148532, 
    0.2663358, 0.2274458, 0.2286697, 0.2103569, 0.1372481, 0.1500652, 
    0.1862546, 0.1869482, 0.2366342, 0.1702662, 0.03732179, 0.0614826, 
    0.0869068, 0.2902814, 0.3104995, 0.3278887,
  0.001425399, 0.005074626, 0.008723853, 0.01237308, 0.01602231, 0.01967154, 
    0.02332076, 0.05926349, 0.06529163, 0.07131977, 0.07734791, 0.08337605, 
    0.08940419, 0.09543233, 0.107362, 0.1045275, 0.1016931, 0.0988586, 
    0.09602413, 0.09318966, 0.0903552, 0.05041086, 0.04356796, 0.03672506, 
    0.02988216, 0.02303926, 0.01619636, 0.009353467, -0.001493983,
  0.1776326, 0.1497964, 0.1499573, 0.07000459, 0.2175092, 0.2981783, 
    0.3250598, 0.2842628, 0.2471856, 0.2747665, 0.1340571, 0.1048109, 
    0.1311947, 0.005279536, 0.1071331, 0.1410291, 0.1361133, 0.1730611, 
    0.205823, 0.1432931, 0.2529723, 0.2324782, 0.2097425, 0.1037677, 
    0.1739237, 0.1503834, 0.09989546, 0.1305787, 0.2178718,
  0.2753192, 0.1972383, 0.169045, 0.1125855, 0.1660011, 0.3539755, 0.1804133, 
    0.3544737, 0.337125, 0.2729782, 0.3058067, 0.1919261, 0.2470873, 
    0.1766789, 0.3332073, 0.4362299, 0.3156651, 0.414358, 0.3076608, 
    0.3944651, 0.4627787, 0.4955675, 0.2910834, 0.4736483, 0.133596, 
    0.161078, 0.2959864, 0.3735709, 0.3896347,
  0.433752, 0.4262303, 0.3570924, 0.4493787, 0.3794606, 0.3629104, 0.3457685, 
    0.4198439, 0.3645076, 0.4220856, 0.3643534, 0.404391, 0.3293742, 
    0.3507358, 0.3408485, 0.2820114, 0.2996669, 0.287103, 0.3747194, 
    0.4033403, 0.3256003, 0.2883944, 0.3266295, 0.3641829, 0.4278666, 
    0.3262988, 0.3151196, 0.3272074, 0.3902837,
  0.345973, 0.3307698, 0.3651109, 0.3390653, 0.3018567, 0.3147859, 0.2240035, 
    0.2352527, 0.1790795, 0.2092753, 0.3264215, 0.2730361, 0.2773383, 
    0.2123889, 0.1352653, 0.2147555, 0.1380741, 0.2528106, 0.2049353, 
    0.3023319, 0.2946377, 0.2819045, 0.2856135, 0.1449409, 0.05917437, 
    0.1247404, 0.1559529, 0.1866234, 0.2848725,
  0.195218, 0.1504789, 0.1945396, 0.2569321, 0.2042793, 0.2019933, 0.1903659, 
    0.20197, 0.05878041, 0.05653476, 0.09023492, 0.1515487, 0.09952103, 
    0.1553935, 0.1878289, 0.1296085, 0.1787378, 0.173502, 0.2159523, 
    0.2359453, 0.1384916, 0.1525308, 0.1881856, 0.04107305, 0.05588773, 
    0.151978, 0.136043, 0.1237839, 0.1604841,
  0.09392664, 0.02468424, 0.1249757, 0.05678598, 0.05335151, 0.09596179, 
    0.09295961, 0.1045114, 0.02725391, 4.449671e-06, -0.0001357251, 
    3.451157e-05, 0.05931618, 0.09414794, 0.07616306, 0.09881, 0.08127371, 
    0.161515, 0.07153133, 0.04920071, 0.07274972, 0.06408771, 0.1055747, 
    -3.304529e-05, 0.04641311, 0.0641955, 0.1391961, 0.06796013, 0.0736969,
  0.06030316, 0.01993083, 0.1585869, 0.0748735, 0.07418475, 0.0555534, 
    0.05402697, 0.04799976, 0.0292945, 0.05328904, 0.02623636, 0.06294507, 
    0.112429, 0.03519747, 0.04211466, 0.1007177, 0.1155123, 0.09439903, 
    0.0294147, 0.03076668, 0.05525645, 0.1917079, 0.02506675, 0.0002896886, 
    0.1158057, 0.1174489, 0.03140453, 0.04897063, 0.08794333,
  0.01847326, 0.01340252, 0.2623849, 0.05394097, 0.0324992, 0.02363219, 
    0.03290547, 0.05391585, 0.03153332, 0.06010322, 0.07128967, 0.01572236, 
    0.05401538, 0.02670819, 0.04125196, 0.03145796, 0.0337579, 0.02675405, 
    0.02584962, 0.03050872, 0.05202017, 0.04390389, 0.006558903, 0.07170682, 
    0.09325157, 0.05877138, 0.04537306, 0.02544133, 0.02751759,
  0.03344292, 0.02643687, 0.001732014, 0.02517439, 0.02484789, 0.08031817, 
    0.1153781, 0.02641571, 0.1249578, 0.2257596, 0.07504372, 0.02718874, 
    0.03011654, 0.0652604, 0.05321768, 0.01614425, 0.02796716, 0.00871906, 
    0.008705839, 0.01174115, 0.04901693, 0.02648852, 0.03465215, 0.06740966, 
    0.07974618, 0.07721019, 0.03816318, 0.02607874, 0.02704006,
  8.312026e-10, 1.929766e-09, 3.697661e-09, 0.01168024, 0.156636, 0.1337027, 
    0.04468401, 0.1019108, 0.06999076, 0.08228333, 0.1076725, 0.06815569, 
    0.0478728, 0.06235782, 0.06724279, 0.03778159, 0.03901425, 0.03246982, 
    0.05621928, 0.03718751, 0.03628009, 0.02232068, 0.1452323, 0.04431462, 
    0.03436647, 0.03440172, 0.01434127, -7.273973e-05, 0.01533281,
  1.11913e-07, 2.871196e-09, 0.001067421, 0.0610975, 1.328174e-06, 
    0.08763276, 0.04408043, 0.07602677, 0.05217149, 0.2672367, 0.1563149, 
    0.1837047, 0.1397513, 0.08353138, 0.1626589, 0.07870142, 0.05670731, 
    0.05371037, 0.0618336, 0.1225903, 0.000661269, 0.2395633, 0.06577861, 
    0.07470022, 0.06490336, 0.06985689, 0.1186382, 0.02641471, -4.954671e-05,
  2.007744e-06, 0.03088723, 0.1488609, 0.06750309, 0.08250726, 0.001934549, 
    -0.0006521951, 0.009365547, 0.1294626, 0.09481368, 0.2157395, 0.2262453, 
    0.1356475, 0.1482173, 0.1463355, 0.1834372, 0.1317251, 0.1829391, 
    0.1129258, 0.1237868, 0.1144024, 0.09769451, 0.09403612, 0.250925, 
    0.1104547, 0.1280192, 0.09808496, 0.04295504, 0.02043575,
  0.038615, 0.05132223, 0.1366635, 0.4444714, 0.155017, 0.0960772, 0.1473341, 
    0.009567199, 0.003144711, 0.03382054, 0.04784517, 0.3219213, 0.2903352, 
    0.1672775, 0.1891424, 0.2474854, 0.240785, 0.1963224, 0.2337509, 
    0.231254, 0.2632157, 0.1180408, 0.2214485, 0.25021, 0.3710442, 0.2878518, 
    0.262028, 0.1969565, 0.09282997,
  0.2409965, 0.3137372, 0.2974009, 0.2850561, 0.1984396, 0.2323446, 
    0.1852083, 0.1894225, 0.1038905, 0.02377001, 0.04104636, 0.2256941, 
    0.4228458, 0.2875811, 0.3699581, 0.3938012, 0.2280569, 0.2616824, 
    0.1244932, 0.2191128, 0.2279044, 0.2370439, 0.3208934, 0.3185216, 
    0.3675939, 0.3556158, 0.2168778, 0.2212194, 0.2773838,
  0.3240536, 0.1633791, 0.2786929, 0.2991106, 0.3004948, 0.2943679, 
    0.4073265, 0.3602564, 0.3275054, 0.4238708, 0.2637194, 0.0662085, 
    0.1972194, 0.3907227, 0.4950124, 0.2640882, 0.381085, 0.4090923, 
    0.2606263, 0.1633397, 0.2156943, 0.2756967, 0.2725848, 0.3701779, 
    0.4257346, 0.2847274, 0.3400445, 0.2748922, 0.2525145,
  0.3577509, 0.3495133, 0.2729388, 0.2900012, 0.296934, 0.3676478, 0.3337572, 
    0.478341, 0.3951858, 0.368911, 0.2071385, 0.1717982, 0.2443039, 
    0.2709997, 0.1355778, 0.1485704, 0.3717747, 0.3261057, 0.2587982, 
    0.2122959, 0.2297894, 0.1976854, 0.1610093, 0.0823108, 0.1617043, 
    0.4485592, 0.172979, 0.2475739, 0.3600287,
  0.222105, 0.2319533, 0.2538243, 0.3007513, 0.2089821, 0.2306509, 0.2340615, 
    0.2367157, 0.1827223, 0.2328285, 0.231773, 0.1789615, 0.2087745, 
    0.2502181, 0.2128415, 0.2481877, 0.2178137, 0.1201382, 0.1230636, 
    0.1807287, 0.1823931, 0.2261446, 0.1791677, 0.03082622, 0.05687734, 
    0.04984339, 0.3180917, 0.3498394, 0.3175268,
  0.05075943, 0.05286239, 0.05496535, 0.05706832, 0.05917128, 0.06127425, 
    0.06337721, 0.08919532, 0.09398523, 0.09877514, 0.1035651, 0.108355, 
    0.1131449, 0.1179348, 0.1056252, 0.1016167, 0.09760825, 0.09359977, 
    0.0895913, 0.08558282, 0.08157435, 0.04392844, 0.04104404, 0.03815963, 
    0.03527524, 0.03239083, 0.02950643, 0.02662203, 0.04907705,
  0.2353781, 0.1482287, 0.1834535, 0.08912367, 0.2939041, 0.3327465, 
    0.3643856, 0.2985277, 0.2091427, 0.2772418, 0.1883624, 0.1618715, 
    0.1696052, 0.006310094, 0.1033097, 0.06972757, 0.1461746, 0.1935607, 
    0.1899861, 0.2105579, 0.3430134, 0.2476472, 0.2582476, 0.1788797, 
    0.1074284, 0.1466773, 0.07379979, 0.1725612, 0.230857,
  0.2770969, 0.1754026, 0.1859083, 0.126776, 0.2071001, 0.394569, 0.1610665, 
    0.32832, 0.3581696, 0.3287185, 0.3062105, 0.28416, 0.2816854, 0.2277894, 
    0.3480713, 0.4969979, 0.4622438, 0.5377866, 0.3718194, 0.4563427, 
    0.4867023, 0.4879284, 0.3287733, 0.4763011, 0.1445566, 0.3269796, 
    0.4743708, 0.3512797, 0.4482411,
  0.4708691, 0.4689113, 0.3648576, 0.4964382, 0.4292649, 0.4283349, 
    0.3935279, 0.4905508, 0.4666118, 0.4704117, 0.4575117, 0.4323708, 
    0.4390967, 0.433441, 0.3824615, 0.3821077, 0.3871253, 0.3662599, 
    0.4841495, 0.4070559, 0.364264, 0.3387284, 0.3311343, 0.3905855, 
    0.4462638, 0.3776088, 0.4275101, 0.456179, 0.456401,
  0.3874041, 0.4148745, 0.4782853, 0.3805958, 0.3500086, 0.3381198, 
    0.2591082, 0.2983697, 0.2411203, 0.2542999, 0.3401723, 0.3925336, 
    0.2616455, 0.213923, 0.1541302, 0.2755078, 0.1414344, 0.2393076, 
    0.2673984, 0.2604891, 0.2609712, 0.2953629, 0.3374221, 0.1387512, 
    0.06281335, 0.1687324, 0.2349166, 0.2758344, 0.3238686,
  0.2285688, 0.2090121, 0.1849535, 0.2170071, 0.2382071, 0.2411924, 
    0.2562404, 0.2828816, 0.1131856, 0.1406693, 0.2014903, 0.1494172, 
    0.07941955, 0.2057529, 0.2278899, 0.2276749, 0.3082123, 0.2327142, 
    0.2800578, 0.2636028, 0.148833, 0.2358948, 0.2437516, 0.04416025, 
    0.07587602, 0.1771803, 0.2018258, 0.2118275, 0.2370948,
  0.1132982, 0.04361816, 0.09716252, 0.139827, 0.07903302, 0.09110309, 
    0.1493964, 0.1624346, 0.1497405, 0.0001642739, 0.001014664, 1.80763e-05, 
    0.04424281, 0.09280542, 0.08881388, 0.1257614, 0.1626382, 0.1575933, 
    0.09982558, 0.09021696, 0.07451619, 0.1110839, 0.2367587, -6.574931e-05, 
    0.04462912, 0.0684552, 0.144256, 0.06620767, 0.1039743,
  0.1771055, 0.02296265, 0.1344694, 0.08036976, 0.07530002, 0.05992319, 
    0.06259585, 0.1183612, 0.05906755, 0.06534383, 0.02284221, 0.04956895, 
    0.08732288, 0.03709726, 0.07031281, 0.09533831, 0.1368518, 0.09519294, 
    0.0409525, 0.04128973, 0.05296594, 0.2426151, 0.1882688, 0.0003770092, 
    0.07207845, 0.1055326, 0.04420691, 0.05035727, 0.1135388,
  0.06860995, 0.01746175, 0.2204355, 0.04685776, 0.03423028, 0.0295366, 
    0.03779751, 0.05980028, 0.04147778, 0.05518482, 0.06807043, 0.0193438, 
    0.04941446, 0.03809232, 0.05965132, 0.03578358, 0.04648983, 0.0643023, 
    0.07206435, 0.05671436, 0.07098975, 0.09408896, 0.04799283, 0.05712545, 
    0.08315211, 0.04130731, 0.07471718, 0.05613229, 0.08953178,
  0.01725357, 0.02811725, 0.001155235, 0.01471536, 0.03721964, 0.09408294, 
    0.1224961, 0.03852451, 0.128805, 0.2192796, 0.06994841, 0.03044408, 
    0.03143331, 0.06551582, 0.06654844, 0.04693392, 0.02929244, 0.005348834, 
    0.01799234, 0.01967033, 0.04937321, 0.0610173, 0.03268724, 0.0500222, 
    0.06748823, 0.06242454, 0.0422551, 0.03344577, 0.0150444,
  1.594358e-10, 6.173511e-10, 8.943751e-10, 0.001159335, 0.1764658, 
    0.1182385, 0.01902899, 0.1366939, 0.08393215, 0.06044216, 0.1171195, 
    0.07343632, 0.04861977, 0.04913426, 0.06226778, 0.06579226, 0.05141962, 
    0.04189918, 0.05857775, 0.0370609, 0.04521749, 0.02730769, 0.177844, 
    0.05076664, 0.04993861, 0.09299207, 0.2403818, 0.01889838, 0.01606865,
  2.635949e-08, -9.539816e-08, 0.0002921258, 0.01772932, -1.607772e-07, 
    0.02887199, 0.03642787, 0.06026021, 0.02597317, 0.3866374, 0.1861881, 
    0.2725025, 0.1572709, 0.1191401, 0.145021, 0.1378357, 0.06664735, 
    0.0556214, 0.141016, 0.2351228, 0.003667557, 0.2858233, 0.08641668, 
    0.07012779, 0.08723734, 0.09241475, 0.2120592, 0.01807347, -1.35784e-05,
  1.305838e-06, 0.08532279, 0.2117147, 0.09605375, 0.08502977, -0.000202108, 
    -0.0005238657, 0.005299374, 0.101694, 0.07733832, 0.2922529, 0.1442274, 
    0.108479, 0.1034018, 0.1054534, 0.1719696, 0.1598194, 0.1777249, 
    0.07040797, 0.09604038, 0.1297828, 0.1807749, 0.1512537, 0.2461138, 
    0.1153193, 0.1361966, 0.1538008, 0.07441476, 0.01758521,
  0.04380242, 0.09469544, 0.1446958, 0.4433329, 0.1395106, 0.08089694, 
    0.1291772, 0.003937118, 0.0007118253, 0.03000075, 0.05872501, 0.2337742, 
    0.1794053, 0.1160601, 0.1714533, 0.2419807, 0.2802141, 0.2431454, 
    0.2073264, 0.2311713, 0.2792082, 0.1187616, 0.2522699, 0.214896, 
    0.3202077, 0.2281555, 0.2480061, 0.2065352, 0.1218895,
  0.2870193, 0.3680744, 0.3145362, 0.3042659, 0.2896672, 0.2518316, 0.218177, 
    0.2116059, 0.1036467, 0.03388271, 0.05121377, 0.2512743, 0.2840119, 
    0.1517351, 0.3143125, 0.409303, 0.2974402, 0.2840495, 0.1509008, 
    0.2358875, 0.2766872, 0.272773, 0.3737246, 0.3494571, 0.4059577, 
    0.2977695, 0.1612351, 0.1773217, 0.2918089,
  0.2961352, 0.1643259, 0.3216152, 0.3364694, 0.3378192, 0.3329446, 
    0.4391394, 0.3935798, 0.3327225, 0.4615084, 0.3318501, 0.08608902, 
    0.1861431, 0.3867175, 0.5883346, 0.3029633, 0.4407327, 0.4374412, 
    0.2671578, 0.1594208, 0.2435118, 0.2819276, 0.246246, 0.3775703, 
    0.5734996, 0.2152301, 0.2406069, 0.2183879, 0.2238886,
  0.2940034, 0.2425672, 0.2534173, 0.2702847, 0.3522979, 0.3662694, 0.354958, 
    0.547716, 0.4129714, 0.4019565, 0.2355496, 0.1532832, 0.2826798, 
    0.3242334, 0.2143153, 0.1692155, 0.3787479, 0.3567485, 0.3004318, 
    0.2586473, 0.220069, 0.2121009, 0.1626894, 0.07486851, 0.129639, 
    0.4486934, 0.1749431, 0.2079499, 0.4291826,
  0.202638, 0.2083941, 0.2280776, 0.289629, 0.2202629, 0.2694342, 0.3337056, 
    0.3095962, 0.2520759, 0.2829036, 0.2434596, 0.1842626, 0.222716, 
    0.2646092, 0.190466, 0.2615138, 0.1851371, 0.1052394, 0.1403787, 
    0.1868015, 0.1848938, 0.212734, 0.1659273, 0.03001578, 0.05504981, 
    0.04018784, 0.3457501, 0.3707489, 0.3650993,
  0.1081508, 0.108836, 0.1095212, 0.1102065, 0.1108917, 0.1115769, 0.1122622, 
    0.1296141, 0.132938, 0.1362618, 0.1395857, 0.1429096, 0.1462334, 
    0.1495573, 0.1418996, 0.1400679, 0.1382363, 0.1364047, 0.1345731, 
    0.1327414, 0.1309098, 0.1169836, 0.1148061, 0.1126286, 0.1104512, 
    0.1082737, 0.1060963, 0.1039188, 0.1076026,
  0.3321565, 0.2291835, 0.2357639, 0.145242, 0.3704091, 0.3767069, 0.4125096, 
    0.3388168, 0.2525619, 0.3202173, 0.2795219, 0.2599894, 0.195424, 
    0.01066566, 0.1297324, 0.06700802, 0.1441536, 0.2100655, 0.1757122, 
    0.1940458, 0.3785779, 0.3425128, 0.312758, 0.2529452, 0.1152508, 
    0.2375655, 0.02947634, 0.1349279, 0.2473344,
  0.2645388, 0.1698841, 0.2094889, 0.1385417, 0.2116173, 0.4399353, 
    0.1583628, 0.3292156, 0.3860775, 0.3735027, 0.2863823, 0.4263869, 
    0.2615968, 0.2747844, 0.4329282, 0.5793296, 0.5257403, 0.6304175, 
    0.4122012, 0.4398986, 0.4982527, 0.5172911, 0.4219907, 0.5167941, 
    0.138563, 0.4355132, 0.465959, 0.3752044, 0.3795577,
  0.5765298, 0.513265, 0.419876, 0.4887469, 0.4756352, 0.4275429, 0.446961, 
    0.5015794, 0.4725097, 0.5086724, 0.4920582, 0.4157156, 0.4913008, 
    0.4932779, 0.3747631, 0.3859439, 0.4614866, 0.4938286, 0.5010027, 
    0.3794964, 0.3513962, 0.3437906, 0.3940723, 0.4470358, 0.3882002, 
    0.4231548, 0.5264162, 0.5527555, 0.5210297,
  0.4039776, 0.4772771, 0.4809364, 0.3399437, 0.3755823, 0.4020346, 
    0.3173873, 0.36198, 0.3213581, 0.3132927, 0.3402063, 0.3402815, 0.306361, 
    0.2708828, 0.1780468, 0.3486694, 0.2461423, 0.2808444, 0.3678114, 
    0.3345298, 0.2338145, 0.342131, 0.3573273, 0.1389563, 0.1228311, 
    0.1922263, 0.3502655, 0.3736154, 0.3487783,
  0.2768908, 0.2762353, 0.1346309, 0.1986593, 0.1524299, 0.2232392, 
    0.2687052, 0.4165708, 0.3348776, 0.2605353, 0.3322124, 0.103009, 
    0.05391398, 0.1829108, 0.2232185, 0.2726555, 0.2930855, 0.2705117, 
    0.3313923, 0.2722891, 0.2461293, 0.3094015, 0.2444726, 0.05813703, 
    0.08992752, 0.1790339, 0.2228736, 0.2804244, 0.2618953,
  0.1460531, 0.1117362, 0.07630174, 0.1233439, 0.0747312, 0.1165928, 
    0.1072336, 0.2190667, 0.1891306, 0.004773745, 0.0003697313, 5.205699e-06, 
    0.02477813, 0.09047123, 0.09349022, 0.1258894, 0.1616877, 0.153422, 
    0.09830751, 0.1190816, 0.09321255, 0.1281588, 0.3149402, 0.008046932, 
    0.04460836, 0.06791682, 0.163556, 0.09146081, 0.1535829,
  0.3146642, 0.04075781, 0.1125174, 0.07936686, 0.05005342, 0.08375514, 
    0.08715024, 0.1543662, 0.3152551, 0.07143644, 0.02297194, 0.03812432, 
    0.09222969, 0.05200593, 0.07211986, 0.08098333, 0.1135172, 0.08842839, 
    0.05854508, 0.05101664, 0.04787058, 0.1510123, 0.6564403, 0.005273261, 
    0.05304327, 0.0827304, 0.07266644, 0.03597775, 0.09055481,
  0.1886684, 0.04390883, 0.1759179, 0.04590237, 0.03982947, 0.0545557, 
    0.07474902, 0.09702586, 0.1004151, 0.0802291, 0.05050675, 0.1061995, 
    0.04417282, 0.0903669, 0.04822495, 0.04001627, 0.06560527, 0.1069276, 
    0.03829598, 0.08910783, 0.1604407, 0.2213512, 0.1930401, 0.03976491, 
    0.06283265, 0.02998509, 0.07013004, 0.1571276, 0.1678264,
  0.03014329, 0.01889887, 0.0004215432, 0.009574563, 0.06150838, 0.1498774, 
    0.09698371, 0.04864517, 0.1185683, 0.2125515, 0.06733789, 0.03796529, 
    0.04881324, 0.07907635, 0.08028463, 0.05788763, 0.04363243, 0.008730039, 
    0.01865087, 0.03889037, 0.05679836, 0.07569991, 0.05541519, 0.02975831, 
    0.03878987, 0.06060733, 0.04799176, 0.04281278, 0.023082,
  4.192775e-11, 2.734621e-10, -9.423367e-12, -0.005226656, 0.2036336, 
    0.09912299, 0.004720317, 0.1454832, 0.09342024, 0.06769338, 0.1003545, 
    0.075518, 0.03797764, 0.03729673, 0.04588426, 0.07119748, 0.05504786, 
    0.06706619, 0.06616869, 0.04541245, 0.04827207, 0.04419667, 0.2834337, 
    0.06330948, 0.03925437, 0.03260557, 0.06133644, 0.04282993, 0.01494282,
  9.469931e-09, -9.848189e-06, 0.0003240925, 0.00529334, -3.02319e-08, 
    0.007522086, 0.0281235, 0.04061333, 0.01896887, 0.3732227, 0.1114341, 
    0.1805761, 0.1060356, 0.07855707, 0.06026552, 0.084438, 0.1908827, 
    0.04952473, 0.1410485, 0.2718613, 0.003699267, 0.3124454, 0.1395586, 
    0.03804874, 0.04508405, 0.05492944, 0.09246186, 0.01841906, -6.726669e-07,
  0.0001149718, 0.0769074, 0.1381545, 0.05107513, 0.08760152, -0.0005196102, 
    -0.0003282699, 0.001915529, 0.0730514, 0.0719779, 0.2334768, 0.09308667, 
    0.06645369, 0.07452751, 0.07677786, 0.1838356, 0.1940564, 0.1263393, 
    0.1357504, 0.05773063, 0.1585264, 0.1949729, 0.1561054, 0.1926449, 
    0.1125838, 0.09971917, 0.15749, 0.1168684, 0.01581143,
  0.05650184, 0.08704171, 0.088971, 0.4548653, 0.1097779, 0.1301266, 
    0.1190479, 0.002678027, -0.0001274299, 0.01753254, 0.06859894, 
    0.09708545, 0.1031025, 0.09464249, 0.1327894, 0.1882987, 0.2663241, 
    0.2569301, 0.198945, 0.2587948, 0.2746561, 0.1170081, 0.2615247, 
    0.1797937, 0.2129497, 0.1859471, 0.2255954, 0.1831736, 0.1654357,
  0.3427733, 0.3918454, 0.2934498, 0.3130061, 0.3113849, 0.243681, 0.2309665, 
    0.2356809, 0.1054185, 0.05007358, 0.06574667, 0.2616505, 0.1328789, 
    0.05388259, 0.250537, 0.3994816, 0.3236499, 0.3138746, 0.2138813, 
    0.2722505, 0.2823861, 0.2722909, 0.4085537, 0.4464665, 0.4798709, 
    0.2399411, 0.1432904, 0.1941183, 0.3026128,
  0.2313623, 0.1591429, 0.3902082, 0.4024817, 0.3334147, 0.37587, 0.5485941, 
    0.4893282, 0.4168922, 0.4866807, 0.420993, 0.1145008, 0.1901264, 
    0.2903228, 0.6271048, 0.327989, 0.4792341, 0.4769081, 0.2794471, 
    0.1792722, 0.292441, 0.3114877, 0.2655615, 0.3640002, 0.6421503, 
    0.1617231, 0.1820814, 0.1660559, 0.2056081,
  0.1876972, 0.1680134, 0.2095667, 0.2477182, 0.40756, 0.3181582, 0.3860811, 
    0.6267157, 0.3959241, 0.4379235, 0.2764725, 0.1822791, 0.3175853, 
    0.3266342, 0.2950446, 0.198703, 0.3901213, 0.3790967, 0.3358256, 
    0.3308239, 0.2081782, 0.2457831, 0.1774051, 0.07612323, 0.1056634, 
    0.429359, 0.1712417, 0.1650229, 0.3113239,
  0.1906898, 0.2140182, 0.2848981, 0.3177617, 0.2790696, 0.327697, 0.4048784, 
    0.3945211, 0.3197018, 0.3011336, 0.2683143, 0.2172966, 0.2327606, 
    0.3048387, 0.2202132, 0.263595, 0.1771091, 0.1325618, 0.1992524, 
    0.2564108, 0.185082, 0.2209319, 0.1714599, 0.04071628, 0.05662148, 
    0.04179319, 0.3462565, 0.3891636, 0.4794558,
  0.1397576, 0.1457741, 0.1517905, 0.1578069, 0.1638233, 0.1698398, 
    0.1758562, 0.168293, 0.1683028, 0.1683127, 0.1683225, 0.1683323, 
    0.1683421, 0.1683519, 0.1827906, 0.1809546, 0.1791187, 0.1772828, 
    0.1754468, 0.1736109, 0.171775, 0.128392, 0.1242017, 0.1200114, 0.115821, 
    0.1116307, 0.1074404, 0.1032501, 0.1349445,
  0.3102934, 0.2428513, 0.2437631, 0.2025868, 0.4525647, 0.353281, 0.369888, 
    0.3197167, 0.3030646, 0.3724521, 0.249491, 0.236425, 0.1985892, 
    0.01461169, 0.112912, 0.1206764, 0.1377616, 0.3008106, 0.1977225, 
    0.1146414, 0.31629, 0.3153097, 0.272831, 0.199617, 0.09764093, 0.2075886, 
    0.1285257, 0.1232438, 0.2134563,
  0.2076293, 0.1307598, 0.2085423, 0.1110211, 0.1274355, 0.3854536, 
    0.1489735, 0.2803098, 0.3220419, 0.275611, 0.2370619, 0.3413931, 
    0.2034854, 0.3340116, 0.5522504, 0.5824564, 0.5077302, 0.5916082, 
    0.4321422, 0.5022013, 0.556532, 0.5275006, 0.5028599, 0.554599, 
    0.1839933, 0.4741388, 0.3136361, 0.3002791, 0.3044003,
  0.5538445, 0.4891154, 0.3835477, 0.4815866, 0.5265614, 0.4529497, 0.54426, 
    0.5030594, 0.4808243, 0.5258806, 0.4722239, 0.437338, 0.4633819, 
    0.4617676, 0.350916, 0.3896847, 0.4931409, 0.554144, 0.4764771, 
    0.3397773, 0.3347692, 0.3106887, 0.3848129, 0.4152212, 0.3923248, 
    0.3736056, 0.5220037, 0.5766249, 0.4725035,
  0.4154803, 0.4709761, 0.4260608, 0.3266343, 0.3703834, 0.4112506, 
    0.3365844, 0.4561443, 0.4505966, 0.3664891, 0.2929989, 0.2182847, 
    0.2515874, 0.2334581, 0.1982456, 0.3454324, 0.3323179, 0.388033, 
    0.372325, 0.3414103, 0.2395552, 0.3206443, 0.3272386, 0.1262046, 
    0.07998662, 0.2151803, 0.398035, 0.4295473, 0.3742504,
  0.303422, 0.2604578, 0.09229585, 0.1734312, 0.1061182, 0.2075558, 
    0.2364766, 0.4221897, 0.4102374, 0.3697976, 0.1993667, 0.07247643, 
    0.05873353, 0.1387609, 0.2256217, 0.210231, 0.1537095, 0.1968933, 
    0.3255246, 0.3573258, 0.2960998, 0.2786296, 0.2289285, 0.07213905, 
    0.07169459, 0.1949665, 0.2174437, 0.3183464, 0.2396818,
  0.1615678, 0.2288809, 0.06773629, 0.05911447, 0.05462082, 0.04646805, 
    0.06802151, 0.1102819, 0.2535179, 0.003182461, 0.0001818312, 
    5.524489e-07, 0.02004654, 0.03641371, 0.0964854, 0.07158916, 0.1181865, 
    0.1503486, 0.1223026, 0.0510058, 0.0726343, 0.08912013, 0.1683636, 
    0.02322071, 0.03514122, 0.07692482, 0.1439058, 0.02942878, 0.0660559,
  0.1630533, 0.07199777, 0.08423321, 0.09488663, 0.02408909, 0.05597212, 
    0.06074952, 0.06952151, 0.3062912, 0.145257, 0.01986192, 0.02737566, 
    0.06615555, 0.03935502, 0.0607407, 0.05910172, 0.08144771, 0.06411247, 
    0.01662168, 0.01146982, 0.02446597, 0.0419981, 0.3822699, 0.2009027, 
    0.04192733, 0.06968595, 0.01749566, 0.006620708, 0.03816885,
  0.2199879, 0.1285325, 0.1420964, 0.05098519, 0.03604059, 0.1037216, 
    0.05094579, 0.04975929, 0.05818517, 0.04604654, 0.03588818, 0.03397736, 
    0.04087433, 0.02419611, 0.01972231, 0.01819481, 0.02709917, 0.02220159, 
    0.005590671, 0.02362606, 0.05586415, 0.183269, 0.4224688, 0.02553074, 
    0.04839585, 0.01820389, 0.01132957, 0.06178605, 0.1793421,
  0.009371196, 0.01258476, 0.0001048373, 0.004341567, 0.03923498, 0.07809256, 
    0.08327622, 0.02438757, 0.06593727, 0.1571569, 0.04110371, 0.03836203, 
    0.05527038, 0.05246178, 0.04490704, 0.038528, 0.04312948, 0.01459844, 
    0.01123116, 0.0399894, 0.1219754, 0.1264304, 0.1307594, 0.01729356, 
    0.01837534, 0.05779641, 0.02235153, 0.01030198, 0.08176943,
  2.837052e-11, 1.743695e-10, -1.58441e-10, -0.006638091, 0.1674593, 
    0.04105854, -0.003912979, 0.0465824, 0.01821465, 0.04069439, 0.0824182, 
    0.04025179, 0.02322982, 0.01950001, 0.01506886, 0.0302578, 0.0296181, 
    0.03441771, 0.06571423, 0.07183979, 0.02787512, 0.03397952, 0.3956802, 
    0.1173634, 0.006367474, 0.005721065, 0.01889584, 0.009978526, 0.01336462,
  6.843734e-09, -2.657761e-05, 0.005426623, 0.001318559, -2.124869e-08, 
    0.002396452, 0.02592776, 0.01962137, 0.01477346, 0.3265952, 0.07367696, 
    0.09574331, 0.05359968, 0.02945899, 0.03455543, 0.02702872, 0.06515664, 
    0.03212697, 0.06974428, 0.1826779, 0.01387113, 0.3053971, 0.03869881, 
    0.012567, 0.01941067, 0.02539708, 0.02627121, 0.004059664, 8.486725e-08,
  0.001503522, 0.06061138, 0.05604748, 0.02721726, 0.08664569, -3.094238e-05, 
    -0.0002960188, 0.001161549, 0.04753374, 0.130148, 0.1650149, 0.06883767, 
    0.04301775, 0.064698, 0.07565712, 0.166355, 0.1971686, 0.0786475, 
    0.1237539, 0.05628059, 0.1669046, 0.2329016, 0.1207616, 0.1842104, 
    0.09176251, 0.09621004, 0.1129777, 0.05462996, 0.01584846,
  0.0624652, 0.05335226, 0.05569495, 0.4531938, 0.07304437, 0.1151052, 
    0.103659, 0.002660508, -0.0002266463, 0.01319186, 0.08690174, 0.04352263, 
    0.0706473, 0.07510883, 0.09966358, 0.1693912, 0.2451439, 0.2240759, 
    0.1474193, 0.2787005, 0.246085, 0.1046321, 0.2595763, 0.1453799, 
    0.1457928, 0.1447362, 0.1998461, 0.2759859, 0.2150919,
  0.3321376, 0.344169, 0.2726243, 0.4000334, 0.3272303, 0.2812088, 0.2299645, 
    0.2505296, 0.1014548, 0.0516842, 0.0529734, 0.2586884, 0.05646074, 
    0.02200811, 0.2175184, 0.4063798, 0.3950628, 0.3924381, 0.2290776, 
    0.2960165, 0.3111911, 0.249807, 0.4008881, 0.5077251, 0.4542622, 
    0.1847247, 0.1406531, 0.1893188, 0.2927708,
  0.2006331, 0.1631729, 0.4694067, 0.4553096, 0.3754463, 0.3826075, 
    0.6543645, 0.5309609, 0.4198326, 0.533787, 0.478191, 0.1594504, 
    0.1985772, 0.2315785, 0.5610921, 0.3006641, 0.4951245, 0.4638358, 
    0.2798373, 0.1949171, 0.3493467, 0.3205637, 0.2865202, 0.3744815, 
    0.5570045, 0.1117463, 0.1482192, 0.130998, 0.1734383,
  0.130355, 0.1147203, 0.2032271, 0.2234956, 0.4659409, 0.3694827, 0.4382447, 
    0.6934637, 0.3765735, 0.4529083, 0.3337067, 0.2365618, 0.4025473, 
    0.3545235, 0.3176721, 0.2498783, 0.4112876, 0.3750393, 0.3692632, 
    0.383916, 0.2238587, 0.2808739, 0.2419444, 0.09118661, 0.08999836, 
    0.4269198, 0.179429, 0.1212795, 0.2100816,
  0.2345076, 0.252353, 0.354419, 0.3437511, 0.2791408, 0.3534441, 0.4518006, 
    0.4455548, 0.3466216, 0.3595953, 0.336224, 0.2847851, 0.2637118, 
    0.3471868, 0.2853398, 0.3112567, 0.2093711, 0.1907173, 0.2362726, 
    0.319618, 0.2365129, 0.2348187, 0.1751646, 0.06592643, 0.06598522, 
    0.04680116, 0.319144, 0.409345, 0.6019003,
  0.2326029, 0.2407883, 0.2489737, 0.2571591, 0.2653445, 0.2735299, 
    0.2817152, 0.2294762, 0.2287535, 0.2280308, 0.2273082, 0.2265855, 
    0.2258628, 0.2251401, 0.2953192, 0.2937223, 0.2921254, 0.2905285, 
    0.2889317, 0.2873348, 0.2857379, 0.2062374, 0.2003716, 0.1945057, 
    0.1886399, 0.182774, 0.1769082, 0.1710424, 0.2260546,
  0.2703567, 0.2392209, 0.1917105, 0.1559191, 0.3452987, 0.2563963, 0.322483, 
    0.3000764, 0.2759842, 0.3528494, 0.2126867, 0.1362577, 0.1610178, 
    0.01204871, 0.1026892, 0.2452114, 0.1732977, 0.3418076, 0.1754573, 
    0.06320761, 0.2177505, 0.2235972, 0.2433917, 0.1153857, 0.1862981, 
    0.1524104, 0.180368, 0.05525115, 0.1835922,
  0.1643085, 0.08946786, 0.1305468, 0.09935269, 0.07454412, 0.2956772, 
    0.1474904, 0.2178633, 0.2314079, 0.2163898, 0.1632797, 0.2321369, 
    0.1341031, 0.2852134, 0.534756, 0.5439631, 0.4826754, 0.5165966, 
    0.3952764, 0.5180239, 0.6038564, 0.5423111, 0.5608445, 0.5995002, 
    0.2387265, 0.4342526, 0.2551895, 0.239142, 0.2754145,
  0.4297345, 0.4343569, 0.3519854, 0.4448309, 0.5522934, 0.4726856, 
    0.5322217, 0.4957118, 0.4602244, 0.4572126, 0.3964157, 0.4423824, 
    0.4878082, 0.4486174, 0.4148056, 0.4275129, 0.50555, 0.5257145, 
    0.4378722, 0.3149674, 0.2816286, 0.2727685, 0.3579307, 0.3636909, 
    0.3814385, 0.3849274, 0.5482954, 0.5637606, 0.4085208,
  0.4175981, 0.4146928, 0.3900528, 0.3371123, 0.3736838, 0.393025, 0.3469167, 
    0.4111433, 0.4378505, 0.3602393, 0.232931, 0.1481957, 0.2201274, 
    0.2393662, 0.2199796, 0.3639769, 0.3805, 0.4034055, 0.2992122, 0.2952939, 
    0.2396137, 0.3115053, 0.2981513, 0.1078956, 0.08252517, 0.2824848, 
    0.4403414, 0.4246118, 0.3693848,
  0.2867761, 0.2002561, 0.05088958, 0.1519054, 0.0845901, 0.1536261, 
    0.2242385, 0.3417294, 0.2732514, 0.2135759, 0.07303648, 0.03993464, 
    0.05418774, 0.1822264, 0.223256, 0.1166321, 0.08533491, 0.1510126, 
    0.3404302, 0.407561, 0.3025198, 0.2285614, 0.1662512, 0.0846543, 
    0.05599929, 0.1923315, 0.2687935, 0.3119836, 0.2578354,
  0.05608821, 0.1190332, 0.05327721, 0.01847248, 0.01570845, 0.01893747, 
    0.04257793, 0.06531657, 0.135556, 0.007832022, -5.780725e-05, 
    -5.569768e-07, 0.01687556, 0.01329655, 0.05706426, 0.04142629, 
    0.09984291, 0.1185796, 0.09048609, 0.009338059, 0.02976016, 0.02590489, 
    0.064542, 0.04241987, 0.02658743, 0.03653419, 0.08415941, 0.007146407, 
    0.01503114,
  0.04655554, 0.1019054, 0.06741504, 0.02417231, 0.006722455, 0.03547602, 
    0.05513794, 0.01206831, 0.1234728, 0.1542043, 0.01585494, 0.02244441, 
    0.0328609, 0.008414362, 0.01191248, 0.0462501, 0.05088594, 0.03582234, 
    0.001253556, 0.0007773564, 0.002323042, 0.009201718, 0.1323204, 
    0.1314467, 0.03412825, 0.05902273, 0.003199406, 0.0002878328, 0.006392129,
  0.09128591, 0.04625848, 0.1164313, 0.04927246, 0.01059977, 0.01276298, 
    0.01120402, 0.01113529, 0.01023348, 0.01532086, 0.02034426, 0.005946368, 
    0.01032377, 0.005004616, 0.008770283, 0.002577826, 0.002804532, 
    0.00528064, 0.0004338768, 0.004571219, 0.01412875, 0.04281569, 0.1108355, 
    0.02339441, 0.04267861, 0.01599549, -0.0005242905, 0.01421111, 0.04873219,
  0.001611007, 0.01060632, 4.560054e-05, 0.00260996, 0.01009327, 0.03593107, 
    0.06541785, 0.003122719, 0.04390394, 0.09779444, 0.0217509, 0.0131232, 
    0.01865324, 0.03729178, 0.0215999, 0.005140074, 0.0232524, 0.009170556, 
    0.004093145, 0.01773796, 0.07969045, 0.2312827, 0.358055, 0.01343585, 
    0.01040951, 0.04699568, 0.006800184, 0.0003086162, 0.01899877,
  2.439697e-11, 1.442777e-10, -1.675012e-10, -0.001348706, 0.08242447, 
    0.01050187, -0.007030174, 0.009221556, 0.004215439, 0.02142784, 
    0.05779057, 0.01629101, 0.01477439, 0.009299473, 0.003303655, 0.01033306, 
    0.01377658, 0.009066463, 0.02895164, 0.03374886, 0.00679643, 0.008395236, 
    0.4258231, 0.1236336, -0.0001031969, 0.001630573, 0.006365533, 
    0.00396047, 0.01513095,
  6.399459e-09, -9.448462e-06, 0.003717198, 0.0007424523, -4.098173e-08, 
    0.001114093, 0.02218171, 0.01085807, 0.01343462, 0.2423585, 0.04249002, 
    0.05242377, 0.01503013, 0.007763021, 0.005684251, 0.01042562, 0.02257499, 
    0.02069302, 0.03840126, 0.125922, 0.02557215, 0.2408075, 0.009559801, 
    -2.066016e-05, 0.008486997, 0.008149221, 0.01044516, 0.001118269, 
    -1.88541e-07,
  0.004424268, 0.04089702, 0.03386045, 0.02005167, 0.08155292, 0.0005349752, 
    -0.0002724281, 0.0005309758, 0.03248531, 0.09621286, 0.1231351, 
    0.04995797, 0.03410149, 0.0576985, 0.065339, 0.1554988, 0.2000833, 
    0.06105644, 0.09926338, 0.04479535, 0.1513947, 0.2538906, 0.09344987, 
    0.1246326, 0.07091615, 0.05739975, 0.03768661, 0.01779943, 0.01477805,
  0.05748168, 0.04493124, 0.03269804, 0.4200364, 0.04349389, 0.1031825, 
    0.09140213, 0.002298617, -0.0001834925, 0.01170609, 0.1016579, 
    0.02427618, 0.05260281, 0.05713926, 0.07826598, 0.1563398, 0.2503259, 
    0.1818046, 0.108424, 0.2823396, 0.231097, 0.09767218, 0.2414045, 
    0.1355778, 0.1004556, 0.1067842, 0.148641, 0.2723032, 0.2336446,
  0.3338998, 0.3191086, 0.2621473, 0.4495803, 0.2847647, 0.3031451, 
    0.2121835, 0.2508117, 0.107443, 0.05309336, 0.05147686, 0.291079, 
    0.02885672, 0.006562176, 0.1848704, 0.3919528, 0.4201312, 0.3337147, 
    0.2421285, 0.3351651, 0.2936567, 0.2823476, 0.3966773, 0.5183191, 
    0.3717132, 0.1596448, 0.1187657, 0.1483101, 0.2990001,
  0.1724201, 0.1964343, 0.4940015, 0.4932784, 0.4441996, 0.4034238, 
    0.6837319, 0.5792004, 0.4597562, 0.5724487, 0.513372, 0.2112487, 
    0.2293535, 0.2106536, 0.4861736, 0.3051111, 0.5420467, 0.4435522, 
    0.2785095, 0.2060605, 0.4728458, 0.3344646, 0.3281552, 0.3050648, 
    0.500816, 0.08130285, 0.120027, 0.1003301, 0.1317683,
  0.09982904, 0.08378454, 0.1925919, 0.1796774, 0.4387791, 0.4526857, 
    0.525215, 0.6647149, 0.338883, 0.4759196, 0.4353266, 0.3125379, 
    0.4445593, 0.3957458, 0.3190063, 0.2880512, 0.455658, 0.3554924, 
    0.3676543, 0.4327989, 0.2351078, 0.3399622, 0.3120672, 0.1156074, 
    0.0888102, 0.4162871, 0.1956342, 0.08394498, 0.1517951,
  0.3001789, 0.2767681, 0.4419152, 0.3917933, 0.3413406, 0.4432125, 
    0.5253904, 0.4770038, 0.3862617, 0.4456927, 0.3847726, 0.3389803, 
    0.3232651, 0.4024963, 0.338886, 0.3611099, 0.2652068, 0.2439592, 
    0.2888348, 0.3438228, 0.2887171, 0.2459735, 0.1728017, 0.1028129, 
    0.08113808, 0.05750811, 0.2920796, 0.3930982, 0.7047072,
  0.2384491, 0.2508228, 0.2631966, 0.2755704, 0.2879442, 0.300318, 0.3126918, 
    0.3296503, 0.3285989, 0.3275474, 0.326496, 0.3254446, 0.3243932, 
    0.3233418, 0.3635581, 0.3591779, 0.3547977, 0.3504174, 0.3460372, 
    0.341657, 0.3372768, 0.2843947, 0.2774525, 0.2705103, 0.2635681, 
    0.256626, 0.2496838, 0.2427416, 0.22855,
  0.2067465, 0.1889161, 0.1276865, 0.09239559, 0.219465, 0.1838335, 
    0.2622164, 0.30461, 0.2619474, 0.280666, 0.1244263, 0.06330593, 
    0.1099066, 0.01012248, 0.06500705, 0.2083375, 0.1756943, 0.3144599, 
    0.1208157, 0.03084257, 0.1431904, 0.151385, 0.210642, 0.0516462, 
    0.1391602, 0.1026352, 0.1665034, 0.05216754, 0.1229044,
  0.1473176, 0.07781967, 0.08141544, 0.06273817, 0.04759566, 0.2227701, 
    0.1346206, 0.1591167, 0.1646958, 0.1566676, 0.09904096, 0.1745314, 
    0.0892808, 0.2675606, 0.4712633, 0.5039573, 0.449892, 0.4531814, 
    0.3214028, 0.5326753, 0.5895545, 0.5188149, 0.5463876, 0.6525884, 
    0.2733219, 0.3611495, 0.2504848, 0.1863012, 0.2143008,
  0.3499593, 0.376878, 0.2875976, 0.4097559, 0.4902994, 0.4295956, 0.4597642, 
    0.4243765, 0.3960081, 0.3813722, 0.3335886, 0.3882176, 0.5163196, 
    0.4309255, 0.4012673, 0.4249818, 0.4759091, 0.5080279, 0.4308401, 
    0.2608864, 0.248618, 0.2277093, 0.2794004, 0.2980869, 0.3550422, 
    0.3952218, 0.5602787, 0.5235324, 0.3734587,
  0.3516697, 0.3646425, 0.3560099, 0.3158953, 0.3818898, 0.3851242, 
    0.3356903, 0.3585849, 0.3563353, 0.3091335, 0.1669938, 0.1054715, 
    0.1869672, 0.2469596, 0.3060484, 0.400054, 0.3463848, 0.3389801, 
    0.222346, 0.2442948, 0.2090155, 0.2756726, 0.2701171, 0.0803901, 
    0.1064751, 0.3479576, 0.4069508, 0.3707254, 0.3425638,
  0.213598, 0.1280275, 0.02408275, 0.1452185, 0.06392851, 0.09771301, 
    0.1892177, 0.3023283, 0.2287365, 0.1025309, 0.031531, 0.0245467, 
    0.049308, 0.1680512, 0.2369165, 0.07124049, 0.05611761, 0.1200951, 
    0.2975681, 0.3362072, 0.2394179, 0.1726084, 0.1005518, 0.09501031, 
    0.05095645, 0.1481507, 0.2900292, 0.2779295, 0.196988,
  0.02206396, 0.05438351, 0.04450269, 0.006520645, 0.00576854, 0.007440238, 
    0.02589634, 0.04027953, 0.06692714, 0.01139689, -2.876603e-05, 
    -2.161225e-07, 0.01430375, 0.004982127, 0.04648007, 0.01943053, 
    0.07249062, 0.09192057, 0.05050586, 0.002159859, 0.01043544, 0.005393001, 
    0.02068291, 0.03769237, 0.01835084, 0.01786102, 0.04676269, 0.001738186, 
    0.004051213,
  0.01380393, 0.112173, 0.05068376, 0.005647237, -0.001338792, 0.01110693, 
    0.01310992, 0.00470657, 0.05241764, 0.06509164, 0.01328148, 0.02553077, 
    0.01187434, 0.003052728, 0.002397008, 0.02955605, 0.01898251, 0.0236593, 
    0.0002207106, 0.0001512513, 0.0008204434, 0.002923556, 0.04168963, 
    0.04435226, 0.02641185, 0.05412471, 0.001120186, 2.96223e-05, 0.001234695,
  0.03343289, 0.01038991, 0.1063411, 0.03704529, 0.005661305, 0.002719347, 
    0.001239729, 0.003016212, 0.00204971, 0.002724323, 0.01207265, 
    0.001181103, 0.002096627, 0.0007009272, 0.003477459, 0.0002781673, 
    0.0005648449, 0.002275191, 0.0001776901, 0.00183293, 0.004785698, 
    0.01544301, 0.04301495, 0.0197511, 0.03331975, 0.01289485, -0.0006935851, 
    0.005263616, 0.0173547,
  0.0002618092, 0.01127154, 5.595651e-05, 0.002801446, 0.001200454, 
    0.0236436, 0.04546672, 0.0002394439, 0.03154675, 0.08707883, 0.01028415, 
    0.00429224, 0.005846494, 0.02367672, 0.01478187, 0.0009318964, 
    0.009282122, 0.001847515, 9.28215e-05, 0.002101904, 0.0218439, 0.0896248, 
    0.1284823, 0.0117156, 0.005554446, 0.02862471, 0.002123068, 4.881366e-05, 
    0.008467252,
  2.370196e-11, 1.371054e-10, -1.602421e-10, 0.002693182, 0.04381752, 
    0.002677567, -0.006347644, 0.002890098, 0.001226911, 0.006376897, 
    0.02544013, 0.005195545, 0.004683945, 0.006202711, 0.0009559571, 
    0.001883379, 0.006562174, 0.0006463235, 0.005903981, 0.006524095, 
    0.001341503, 0.0008252913, 0.3724348, 0.09825961, -1.886599e-05, 
    0.0007243862, 0.002980409, 0.002075001, 0.0157154,
  6.173748e-09, -3.844972e-06, 0.0009462585, 0.0005316113, 2.485082e-09, 
    0.0006879995, 0.02047355, 0.005597307, 0.0157852, 0.1679102, 0.01983986, 
    0.02548181, 0.002945316, 0.002387387, 0.001483571, 0.004572794, 
    0.008594586, 0.01524905, 0.03677306, 0.0612073, 0.005632824, 0.1833235, 
    0.003999772, -0.002110512, 0.002633946, 0.002759141, 0.005445265, 
    0.0003051214, -3.369558e-05,
  0.002150204, 0.02525845, 0.02634367, 0.01655706, 0.07671613, 0.0004076563, 
    -0.000288383, 0.0002688723, 0.02065052, 0.0747845, 0.09536184, 
    0.03161044, 0.03094397, 0.04168272, 0.04717963, 0.1449007, 0.1635162, 
    0.03433082, 0.07387377, 0.02534105, 0.1234717, 0.2131431, 0.08958466, 
    0.06056765, 0.05090405, 0.03405809, 0.01417823, 0.00748953, 0.01176952,
  0.04447735, 0.08138754, 0.02048196, 0.3731199, 0.02474284, 0.1042981, 
    0.08492348, 0.001298351, -0.0001427938, 0.01074602, 0.115057, 0.01648654, 
    0.0393103, 0.04401996, 0.05822324, 0.1410129, 0.2478288, 0.1515571, 
    0.07281001, 0.2586627, 0.2196549, 0.09380419, 0.2133267, 0.1193599, 
    0.06792036, 0.07438997, 0.09994569, 0.1901802, 0.1891091,
  0.2979604, 0.2799172, 0.2161449, 0.4038148, 0.2739104, 0.3124463, 
    0.1861356, 0.2274834, 0.1025718, 0.05895578, 0.05246279, 0.3414564, 
    0.01720602, 0.002465225, 0.155549, 0.3390972, 0.3747815, 0.2726079, 
    0.1595266, 0.3452681, 0.2392137, 0.270941, 0.3494823, 0.5687039, 
    0.2953991, 0.1420121, 0.08663829, 0.09461305, 0.2556539,
  0.1203288, 0.2267557, 0.5128424, 0.4934072, 0.4823152, 0.3970289, 
    0.6817477, 0.6093453, 0.5048524, 0.5753536, 0.5764052, 0.2945561, 
    0.263828, 0.1908998, 0.4331284, 0.3418206, 0.5843964, 0.4118641, 
    0.2764115, 0.2203185, 0.5823197, 0.3282033, 0.3395261, 0.2762476, 
    0.4576408, 0.05971602, 0.1008591, 0.06740218, 0.09893711,
  0.07441172, 0.06743009, 0.1940628, 0.1323982, 0.3996371, 0.4862352, 
    0.6210789, 0.633838, 0.2650275, 0.5633671, 0.5036303, 0.376789, 0.51998, 
    0.4626299, 0.3718371, 0.3061502, 0.4373415, 0.3041383, 0.3396634, 
    0.4130993, 0.2388729, 0.4425506, 0.3405911, 0.1690982, 0.08747917, 
    0.366778, 0.2080901, 0.05538331, 0.1252775,
  0.4030785, 0.2939436, 0.4762437, 0.4163496, 0.3771003, 0.4756544, 
    0.5733254, 0.5231866, 0.5090712, 0.5645455, 0.4670294, 0.4194714, 
    0.4063439, 0.4715135, 0.4099214, 0.4323594, 0.368149, 0.3311188, 
    0.3545678, 0.4306714, 0.3821888, 0.2528482, 0.1854926, 0.1858479, 
    0.1012337, 0.05996971, 0.230274, 0.3547798, 0.6646941,
  0.2435669, 0.2561018, 0.2686368, 0.2811718, 0.2937067, 0.3062417, 
    0.3187767, 0.3036354, 0.3030933, 0.3025512, 0.302009, 0.3014669, 
    0.3009247, 0.3003826, 0.3485139, 0.3418142, 0.3351147, 0.3284151, 
    0.3217155, 0.3150159, 0.3083163, 0.2837895, 0.2784962, 0.273203, 
    0.2679098, 0.2626165, 0.2573233, 0.25203, 0.2335389,
  0.1352055, 0.1311978, 0.08436626, 0.08074537, 0.1395578, 0.1311299, 
    0.2006218, 0.2475188, 0.2150795, 0.2146808, 0.0723101, 0.04019647, 
    0.07769109, 0.01082886, 0.04524548, 0.1409674, 0.1545153, 0.2730308, 
    0.0757755, 0.01186492, 0.09778354, 0.133179, 0.1666401, 0.04324534, 
    0.1168924, 0.07853876, 0.1177836, 0.03952203, 0.09369016,
  0.1129565, 0.07035527, 0.05214044, 0.03858766, 0.03226892, 0.1589366, 
    0.1148635, 0.1116087, 0.1231355, 0.1180981, 0.06732113, 0.1373181, 
    0.06713724, 0.220093, 0.39943, 0.4454089, 0.3353637, 0.4003106, 0.260872, 
    0.4883225, 0.4970595, 0.4675523, 0.473115, 0.6422781, 0.263295, 
    0.3033272, 0.206034, 0.1451162, 0.1836877,
  0.2946045, 0.3205494, 0.2525842, 0.3549241, 0.3896573, 0.3398576, 
    0.3819884, 0.338308, 0.3315548, 0.3160207, 0.2578644, 0.3243175, 
    0.4815783, 0.3765181, 0.3371574, 0.3738799, 0.4308315, 0.4475585, 
    0.3732275, 0.214562, 0.2038097, 0.167916, 0.1941822, 0.2098632, 0.303644, 
    0.3800908, 0.5446199, 0.4628893, 0.3089022,
  0.2847624, 0.2881568, 0.3000273, 0.2570032, 0.3393641, 0.326741, 0.2869199, 
    0.2984994, 0.2772887, 0.2324877, 0.1146467, 0.06250849, 0.1527703, 
    0.2183191, 0.310274, 0.3883164, 0.2752358, 0.2659893, 0.1559881, 
    0.1900106, 0.1611151, 0.2253103, 0.2281551, 0.05913256, 0.1022665, 
    0.3275498, 0.3460462, 0.2970374, 0.2842653,
  0.1502679, 0.07397353, 0.012385, 0.1263539, 0.05150959, 0.06330029, 
    0.1546105, 0.267099, 0.1867909, 0.05615739, 0.01697811, 0.01667718, 
    0.04587777, 0.1166623, 0.2141871, 0.03183345, 0.03340453, 0.0960501, 
    0.2675264, 0.267065, 0.1478082, 0.1090825, 0.05178254, 0.09553425, 
    0.05686186, 0.1093172, 0.2299724, 0.2156205, 0.1268233,
  0.01011193, 0.02528839, 0.03066964, 0.003464049, 0.002040696, 0.002419475, 
    0.009699835, 0.02611881, 0.02698311, 0.01000469, -1.164823e-05, 
    -5.670341e-08, 0.009445534, 0.001753705, 0.01766634, 0.008235374, 
    0.05124459, 0.06338461, 0.03049801, 0.001122877, 0.002715535, 
    0.002473357, 0.01088256, 0.01924999, 0.01194693, 0.007295088, 0.02854027, 
    0.001022441, 0.002216259,
  0.006083902, 0.09048975, 0.03387632, 0.001822722, -0.001979997, 
    0.003320187, 0.005590104, 0.002654027, 0.02711774, 0.02848862, 
    0.007828712, 0.01693197, 0.002809333, 0.0008862827, 0.001069873, 
    0.01507149, 0.00616904, 0.01394982, 0.0001026977, 7.738172e-05, 
    0.0004700436, 0.001401385, 0.0170502, 0.02485693, 0.02337709, 0.04220995, 
    0.000560421, 1.10935e-05, 0.000609312,
  0.01623791, 0.003670483, 0.09504499, 0.02738966, 0.00377204, 0.00114859, 
    0.0002761196, 0.001153519, 0.000913811, 0.0002453018, 0.005590984, 
    0.0005575673, 0.00043966, 0.0002160604, 0.001758308, 6.148264e-05, 
    0.0003107224, 0.001370242, 9.891285e-05, 0.001060632, 0.002625463, 
    0.008298766, 0.02301028, 0.01601653, 0.02709978, 0.01297552, 
    -0.0001260411, 0.002806033, 0.00876665,
  0.0001306039, 0.007337795, 2.966281e-05, 0.001685692, 0.0003784137, 
    0.01370342, 0.02030509, 8.840856e-05, 0.03859744, 0.0849264, 0.004544502, 
    0.001483185, 0.004030963, 0.01417308, 0.01175813, 0.0004371147, 
    0.004881629, 0.000125074, 2.682291e-05, 0.0005722504, 0.004384866, 
    0.02801171, 0.05579435, 0.0116972, 0.002409476, 0.01373533, 0.0007467894, 
    1.991585e-05, 0.004504553,
  2.345832e-11, 1.3469e-10, -1.534504e-10, 0.003156848, 0.02508149, 
    0.0008179647, -0.005285476, 0.001566152, 0.0006733173, 0.0008646712, 
    0.01143939, 0.001225082, 0.002041136, 0.003160753, 0.0003613743, 
    0.0004875814, 0.002423581, 0.0002051584, 0.001577399, 0.001920999, 
    0.000434393, 0.0001766709, 0.2827191, 0.07335889, -2.968253e-06, 
    0.0004069931, 0.001738174, 0.00132608, 0.01603176,
  6.102977e-09, -2.000251e-06, 0.0003349576, 0.0003390517, 1.869964e-08, 
    0.0004881948, 0.02034861, 0.002523005, 0.01696447, 0.1006171, 0.00835121, 
    0.01269377, 0.001117009, 0.00100278, 0.0008133174, 0.002005627, 
    0.003563439, 0.006923519, 0.0293054, 0.0237614, 0.002326131, 0.1352941, 
    0.002352082, -0.001814865, 0.0009523312, 0.001006272, 0.003449315, 
    0.0001621055, -2.336769e-05,
  0.0008542086, 0.01972338, 0.01805784, 0.01260589, 0.06862663, 0.0002777592, 
    -0.0002807126, 0.0001501826, 0.01336582, 0.06164746, 0.0769943, 
    0.01781751, 0.01825905, 0.02519875, 0.02942622, 0.112741, 0.1195417, 
    0.01791297, 0.03865177, 0.01527542, 0.1048096, 0.1770966, 0.08151923, 
    0.02660949, 0.0319343, 0.02029327, 0.007344343, 0.004360763, 0.008310923,
  0.02896762, 0.06712648, 0.01405043, 0.3285584, 0.01574298, 0.08928754, 
    0.08237857, 0.0004207904, -0.0001164732, 0.01112994, 0.1139593, 
    0.01263422, 0.02873333, 0.03216911, 0.038124, 0.1160831, 0.2118832, 
    0.1285755, 0.05038291, 0.2381536, 0.2049527, 0.08824761, 0.1877602, 
    0.1017436, 0.0466861, 0.04755645, 0.05934775, 0.1060476, 0.128714,
  0.22663, 0.2563533, 0.1637381, 0.3204497, 0.2423932, 0.2762111, 0.1580819, 
    0.2007681, 0.08970334, 0.07303872, 0.04550306, 0.3902262, 0.009268295, 
    0.001445141, 0.1245247, 0.288443, 0.3228178, 0.2068223, 0.09934151, 
    0.338354, 0.1799589, 0.1926597, 0.2897691, 0.6092577, 0.2438431, 
    0.1245454, 0.06492034, 0.06434553, 0.1959249,
  0.07072251, 0.2300042, 0.4978323, 0.4625086, 0.4649551, 0.3292024, 
    0.6150083, 0.5640911, 0.4886541, 0.5445836, 0.6357296, 0.3729562, 
    0.2965125, 0.193159, 0.3787875, 0.3368356, 0.6097283, 0.3708863, 
    0.2636001, 0.2342262, 0.6795564, 0.3264147, 0.3178381, 0.2720399, 
    0.42659, 0.04486819, 0.08169391, 0.04337858, 0.07399724,
  0.05715376, 0.05385556, 0.2011272, 0.09749385, 0.3563551, 0.4757568, 
    0.6168917, 0.5875009, 0.2443181, 0.6046849, 0.6260018, 0.4078904, 
    0.6572987, 0.5047293, 0.3853652, 0.2674925, 0.4113525, 0.2535643, 
    0.3220228, 0.3830296, 0.2918628, 0.5546584, 0.4587953, 0.2492339, 
    0.1063753, 0.3042271, 0.2265937, 0.0406442, 0.09623962,
  0.4006471, 0.2715266, 0.4792227, 0.4221292, 0.4855745, 0.5680909, 0.632723, 
    0.6126333, 0.6753454, 0.6515203, 0.6049443, 0.6110742, 0.5581488, 
    0.5531567, 0.4926128, 0.4581293, 0.4454349, 0.4421098, 0.4396425, 
    0.5108321, 0.4448987, 0.2743344, 0.1904665, 0.280258, 0.08823483, 
    0.06058107, 0.1799093, 0.2875812, 0.6047097,
  0.1939361, 0.2054376, 0.2169391, 0.2284407, 0.2399422, 0.2514437, 
    0.2629452, 0.2229484, 0.2250546, 0.2271608, 0.229267, 0.2313732, 
    0.2334794, 0.2355856, 0.2907313, 0.2808788, 0.2710263, 0.2611739, 
    0.2513214, 0.241469, 0.2316165, 0.2070268, 0.2032716, 0.1995163, 
    0.195761, 0.1920058, 0.1882505, 0.1844952, 0.1847349,
  0.09318246, 0.08330628, 0.05786098, 0.05914129, 0.1131926, 0.088846, 
    0.1543332, 0.1979289, 0.1820699, 0.1678172, 0.04949972, 0.0237444, 
    0.04320429, 0.005028029, 0.02943651, 0.07911559, 0.1186048, 0.2268115, 
    0.05665376, 0.005523042, 0.06581439, 0.09900672, 0.1257753, 0.03823926, 
    0.1172633, 0.06430503, 0.07505065, 0.03044618, 0.06881544,
  0.07341527, 0.05272507, 0.03064364, 0.02427879, 0.02344304, 0.120589, 
    0.09629665, 0.07904025, 0.09567774, 0.1023466, 0.04930749, 0.1096973, 
    0.05204032, 0.1716079, 0.3269227, 0.3569558, 0.2647596, 0.3185746, 
    0.1897141, 0.3577362, 0.3630691, 0.3919779, 0.4178877, 0.5685008, 
    0.2247641, 0.2433696, 0.1558542, 0.1080151, 0.1480162,
  0.2238262, 0.2422427, 0.1947821, 0.2769584, 0.3033714, 0.2529353, 0.28596, 
    0.2632568, 0.2633751, 0.2507108, 0.1933348, 0.247272, 0.384019, 
    0.2891399, 0.2555582, 0.2938105, 0.3638978, 0.3695171, 0.3042571, 
    0.1591993, 0.1410386, 0.1124627, 0.1233982, 0.1245762, 0.2333384, 
    0.3191192, 0.4528299, 0.3664898, 0.2310177,
  0.2262817, 0.2146429, 0.2187614, 0.1916823, 0.2743865, 0.2646146, 
    0.2182851, 0.2223383, 0.2165211, 0.157414, 0.06905822, 0.03229456, 
    0.1144929, 0.1662676, 0.263141, 0.2881934, 0.1965136, 0.1778452, 
    0.09660509, 0.1426573, 0.1115132, 0.1600148, 0.1782999, 0.04361562, 
    0.07793579, 0.3052332, 0.2876548, 0.2334935, 0.2220803,
  0.09727342, 0.03982665, 0.007027458, 0.09194702, 0.03714159, 0.03646592, 
    0.1086209, 0.2187263, 0.1437964, 0.03559886, 0.01085483, 0.01016719, 
    0.03897914, 0.07855133, 0.1870007, 0.01391308, 0.0166864, 0.07581097, 
    0.2364766, 0.2001286, 0.08381362, 0.05522015, 0.02452701, 0.09011167, 
    0.05485506, 0.07782498, 0.1448064, 0.1267882, 0.07246935,
  0.006243449, 0.0121078, 0.01505757, 0.002017248, 0.001090113, 0.00110314, 
    0.003082217, 0.01596177, 0.01453824, 0.006422805, -6.932511e-06, 
    -1.134508e-08, 0.005104386, 0.0007840516, 0.004200388, 0.003535151, 
    0.02746204, 0.04088429, 0.01652149, 0.0007152572, 0.001415286, 
    0.001636921, 0.00731696, 0.01312282, 0.007805148, 0.003261378, 
    0.01448768, 0.0006572413, 0.001509867,
  0.003765013, 0.059152, 0.02011524, 0.0010141, -0.001578505, 0.001271506, 
    0.002045627, 0.001770407, 0.01695008, 0.01507218, 0.003514678, 
    0.009111314, 0.0008617736, 0.000447139, 0.0006374434, 0.00519002, 
    0.001765848, 0.005727247, 6.621497e-05, 5.181165e-05, 0.0003213824, 
    0.000846205, 0.009187474, 0.01678054, 0.0161316, 0.03088038, 
    0.0003492991, 6.087512e-06, 0.0003862055,
  0.01012919, 0.001839609, 0.08704486, 0.02514558, 0.002268091, 0.0006450976, 
    0.0001853573, 0.0004048585, 0.0006004397, 2.918931e-05, 0.002556083, 
    0.0003601148, 0.0002158792, 0.0001523391, 0.0008157221, 4.145193e-05, 
    0.0002142376, 0.0009477047, 6.585752e-05, 0.0007194597, 0.00171603, 
    0.005468198, 0.01510812, 0.01345052, 0.02256303, 0.009802991, 
    -1.665455e-05, 0.001802168, 0.005516019,
  8.449828e-05, 0.005607462, 1.364863e-05, 0.0007234684, 0.0002001836, 
    0.006844402, 0.008646803, 5.18731e-05, 0.04008381, 0.07737208, 
    0.001885067, 0.0006210056, 0.001911039, 0.006195008, 0.006902496, 
    0.0002662258, 0.001711257, 6.924149e-05, 1.364839e-05, 0.0003139853, 
    0.001868865, 0.01450682, 0.03109929, 0.01114552, 0.001568333, 
    0.006164897, 0.0002360593, 1.203324e-05, 0.002714308,
  2.376115e-11, 1.329689e-10, -1.487927e-10, 0.002707758, 0.01386302, 
    0.0004670978, -0.003565137, 0.001103922, 0.0003325892, 0.0001718328, 
    0.00537165, 0.0004152717, 0.0008899747, 0.001585583, 0.0002175017, 
    0.0002018813, 0.0006490039, 0.0001198098, 0.0006268431, 0.001011139, 
    0.0001502693, 0.0001008301, 0.2231296, 0.05384166, -1.279091e-06, 
    0.0002683538, 0.001182895, 0.0009515259, 0.01455051,
  6.105228e-09, -1.211899e-06, 0.0001978611, 0.0002443218, -6.786487e-08, 
    0.0003783728, 0.01803136, 0.001226458, 0.01543695, 0.0621983, 
    0.003631497, 0.007899399, 0.0007174914, 0.0006545191, 0.0005513891, 
    0.00129179, 0.002109981, 0.001562646, 0.02171332, 0.0114339, 0.001241361, 
    0.09877703, 0.001607087, -0.001573493, 0.0005686948, 0.0005157262, 
    0.002468772, 0.0001046597, -1.581368e-05,
  0.0005204588, 0.01589302, 0.01104867, 0.008086486, 0.06178443, 
    0.0002578591, -0.0002290372, 0.0003487153, 0.01195744, 0.04490714, 
    0.05779626, 0.00963967, 0.009760236, 0.01316338, 0.01625863, 0.07560797, 
    0.07218525, 0.008507127, 0.0204304, 0.009127872, 0.08260816, 0.1405344, 
    0.07235045, 0.01498285, 0.01770405, 0.01006827, 0.004533904, 0.003029906, 
    0.005816382,
  0.02028977, 0.05959593, 0.009869994, 0.2893803, 0.01086634, 0.07000658, 
    0.07625637, 0.0007611934, -9.45889e-05, 0.01576524, 0.09967488, 
    0.00936054, 0.02018168, 0.0219891, 0.02391613, 0.08670994, 0.1537045, 
    0.09691803, 0.02980375, 0.2137607, 0.1786329, 0.07674775, 0.165173, 
    0.08410326, 0.03121553, 0.03012298, 0.03268875, 0.05182913, 0.08044104,
  0.1738917, 0.2218356, 0.1403461, 0.25434, 0.2009025, 0.225987, 0.1334734, 
    0.1808941, 0.08784971, 0.08922666, 0.03418665, 0.3946354, 0.006166744, 
    0.0009915789, 0.0961491, 0.2268731, 0.2578854, 0.1457649, 0.06703622, 
    0.329901, 0.1300295, 0.131763, 0.2490449, 0.6123612, 0.2022254, 0.107894, 
    0.04670028, 0.0420297, 0.1382145,
  0.04348379, 0.2560402, 0.4633368, 0.3862279, 0.479212, 0.2652831, 
    0.5161396, 0.4394627, 0.4573348, 0.4381097, 0.5878317, 0.4381615, 
    0.3331023, 0.1859209, 0.3288962, 0.2982854, 0.6129325, 0.33374, 
    0.2559597, 0.236572, 0.6760221, 0.3789459, 0.247108, 0.2791311, 
    0.4047671, 0.03423723, 0.0605753, 0.03066384, 0.05346438,
  0.04346424, 0.04141099, 0.2416904, 0.07691456, 0.3038315, 0.4301206, 
    0.5942079, 0.4946169, 0.3243334, 0.7118826, 0.6958402, 0.3649912, 
    0.754539, 0.4683577, 0.3600662, 0.2280008, 0.3484769, 0.2192302, 
    0.3086995, 0.370268, 0.3004926, 0.5967808, 0.5990182, 0.3868369, 
    0.1358359, 0.2485946, 0.2606911, 0.02518052, 0.07483906,
  0.4036355, 0.246892, 0.4180525, 0.3887611, 0.5325235, 0.5780653, 0.5785046, 
    0.5475838, 0.6140092, 0.6290413, 0.5424159, 0.6500645, 0.6369518, 
    0.5500247, 0.4502012, 0.3854533, 0.3875321, 0.4481282, 0.4348089, 
    0.4549421, 0.4831296, 0.258214, 0.1942086, 0.3584469, 0.04741001, 
    0.06453745, 0.1630043, 0.2587419, 0.5273525,
  0.1153693, 0.1234577, 0.1315461, 0.1396345, 0.1477229, 0.1558113, 
    0.1638997, 0.143607, 0.1463773, 0.1491476, 0.1519179, 0.1546882, 
    0.1574585, 0.1602288, 0.2031896, 0.1955205, 0.1878514, 0.1801824, 
    0.1725133, 0.1648442, 0.1571752, 0.1206204, 0.1174307, 0.1142411, 
    0.1110514, 0.1078618, 0.1046721, 0.1014825, 0.1088986,
  0.07297079, 0.06063513, 0.04276587, 0.06499421, 0.09134517, 0.06706244, 
    0.1065464, 0.1690217, 0.1487356, 0.1415384, 0.04349769, 0.01727917, 
    0.02761297, 0.00361315, 0.02073997, 0.05716909, 0.08625933, 0.1951279, 
    0.04818879, 0.003797988, 0.04842959, 0.08027848, 0.09457503, 0.03480605, 
    0.1106893, 0.0551505, 0.05661726, 0.02765578, 0.06347953,
  0.04762994, 0.03848719, 0.02336758, 0.01790771, 0.01930314, 0.09760476, 
    0.08346388, 0.06373075, 0.07895727, 0.09350018, 0.03930907, 0.09124281, 
    0.0452148, 0.1441806, 0.2521363, 0.2778205, 0.2126956, 0.2490097, 
    0.1492966, 0.2661847, 0.2770944, 0.3076435, 0.3440531, 0.4842285, 
    0.1986422, 0.1969029, 0.1190389, 0.08216731, 0.1088418,
  0.1726931, 0.181423, 0.1490087, 0.2173577, 0.2417195, 0.1980923, 0.2278731, 
    0.2073303, 0.2117888, 0.2077502, 0.1635062, 0.192617, 0.3053108, 
    0.2226114, 0.190344, 0.2294578, 0.2952655, 0.298798, 0.2482145, 
    0.1169522, 0.1035739, 0.07739003, 0.08470687, 0.08024389, 0.1751143, 
    0.2515928, 0.3598219, 0.2877111, 0.176918,
  0.1757717, 0.1636127, 0.1590592, 0.1479868, 0.2293415, 0.2348286, 
    0.1761521, 0.1754777, 0.1742211, 0.1156251, 0.04193829, 0.02007476, 
    0.07992811, 0.1187414, 0.2148102, 0.20909, 0.1359986, 0.1162618, 
    0.06473757, 0.1125885, 0.07993861, 0.1167827, 0.140172, 0.03505418, 
    0.05861695, 0.2556697, 0.234833, 0.1866972, 0.1842587,
  0.06559845, 0.02359238, 0.005181186, 0.05935885, 0.02434389, 0.02162999, 
    0.07057671, 0.1683822, 0.09677184, 0.02614696, 0.008059318, 0.004685419, 
    0.03006416, 0.04955728, 0.1631851, 0.008221094, 0.009022492, 0.05457557, 
    0.1745205, 0.1470925, 0.04905437, 0.0288, 0.01408273, 0.08931885, 
    0.04198491, 0.05666758, 0.09249929, 0.08233008, 0.04472832,
  0.004538088, 0.007339655, 0.009968591, 0.001360125, 0.0007570775, 
    0.0007508591, 0.001579331, 0.009282348, 0.01036756, 0.004770534, 
    -4.971839e-06, -1.45714e-09, 0.004713827, 0.0004841439, 0.001898051, 
    0.001940406, 0.01609092, 0.0224837, 0.009763899, 0.0005499737, 
    0.0009579547, 0.001246584, 0.005593679, 0.009412325, 0.006069887, 
    0.001679922, 0.007579976, 0.0004695703, 0.00115716,
  0.00271781, 0.04298159, 0.01089476, 0.0007429261, -0.001213527, 
    0.0006758782, 0.00100805, 0.001314805, 0.01220269, 0.01029291, 
    0.001597059, 0.004534213, 0.0004903363, 0.0003262683, 0.0004498543, 
    0.002170062, 0.0006365556, 0.002391334, 4.855657e-05, 3.901609e-05, 
    0.0002468286, 0.0005952406, 0.006035704, 0.0127826, 0.01061838, 
    0.02280718, 0.0002557566, 2.900649e-06, 0.0002804986,
  0.007334639, 0.001195985, 0.07398115, 0.03026127, 0.001321068, 
    0.0004447917, 0.0001219504, 0.0001763981, 0.000445919, 0.0001097289, 
    0.001631863, 0.0002639869, 0.0001656461, 0.0001287024, 0.0004360033, 
    3.43424e-05, 0.0001629083, 0.0007266619, 4.931045e-05, 0.0005476, 
    0.00127632, 0.004085098, 0.01127802, 0.01654977, 0.0176815, 0.008009577, 
    -6.542669e-05, 0.001321844, 0.003984917,
  6.389843e-05, 0.005687174, -3.183111e-05, 0.0004719755, 0.0001329262, 
    0.003568509, 0.004019212, 3.792866e-05, 0.04398786, 0.07668175, 
    0.0008918997, 0.0003423215, 0.0009817124, 0.002912238, 0.003283326, 
    0.0001851347, 0.0007435363, 4.393133e-05, 8.928042e-06, 0.0002098997, 
    0.001143562, 0.009563102, 0.02032913, 0.01185664, 0.002335423, 
    0.002874044, 0.0001333431, 8.393262e-06, 0.001930193,
  2.487473e-11, 1.331355e-10, -1.451869e-10, 0.0051201, 0.008823706, 
    0.0003296211, -0.002346733, 0.0008684886, 1.656969e-05, 0.0001016094, 
    0.002982205, 0.0002035979, 0.0003746975, 0.0006892406, 0.0001560418, 
    0.0001596896, 0.0001856382, 8.499243e-05, 0.0003960845, 0.0006554121, 
    8.117451e-05, 7.049302e-05, 0.1702529, 0.03559374, -9.002905e-07, 
    0.0002014401, 0.0008937217, 0.0007506495, 0.01050091,
  6.180161e-09, -8.469219e-07, 0.0001447566, 0.0001997094, -2.008414e-06, 
    0.0003143082, 0.01547946, 0.0008924787, 0.013349, 0.04355002, 
    0.002212308, 0.004903132, 0.0005456505, 0.0005121467, 0.0004218966, 
    0.0009952413, 0.00153393, 0.0008746196, 0.01293684, 0.007242827, 
    0.000895453, 0.07899579, 0.001231109, -0.001217038, 0.0002985692, 
    0.0003611807, 0.001943607, 7.726259e-05, -2.405877e-05,
  0.0003751268, 0.01374072, 0.007516098, 0.00528895, 0.05834991, 
    0.0002937968, -0.0002499985, 0.001194727, 0.01365951, 0.03154804, 
    0.04462206, 0.005475304, 0.005078264, 0.006601118, 0.009639882, 
    0.04801909, 0.04797403, 0.00488922, 0.01331524, 0.006535455, 0.07554589, 
    0.1135347, 0.05926785, 0.01003839, 0.009824688, 0.005455076, 0.003307331, 
    0.002352589, 0.005540021,
  0.01506503, 0.05490785, 0.007502506, 0.2636001, 0.008729818, 0.05902772, 
    0.06807697, 0.004788124, -7.384707e-05, 0.02845838, 0.09701405, 
    0.007212781, 0.01576937, 0.01596394, 0.01654787, 0.0626266, 0.1048351, 
    0.06939861, 0.0175386, 0.1922055, 0.1638596, 0.06920798, 0.155901, 
    0.07794162, 0.02252606, 0.02016757, 0.02054207, 0.02874915, 0.05541036,
  0.1329692, 0.1981643, 0.1365946, 0.2187161, 0.1777995, 0.1910656, 
    0.1163361, 0.194574, 0.1308661, 0.08711258, 0.02875896, 0.3852546, 
    0.004657034, 0.0007651211, 0.07633228, 0.1762809, 0.2043588, 0.1138129, 
    0.05129834, 0.3178014, 0.1054128, 0.1003287, 0.2215801, 0.5876383, 
    0.1803762, 0.09350871, 0.03488667, 0.03004839, 0.0984914,
  0.03089939, 0.3059183, 0.4295053, 0.3412724, 0.4752034, 0.2405419, 
    0.4283874, 0.3560008, 0.3749983, 0.3615608, 0.5178275, 0.5435721, 
    0.3956611, 0.2081967, 0.2923568, 0.2669199, 0.6013112, 0.3031884, 
    0.2965145, 0.2581641, 0.6178692, 0.433318, 0.1705762, 0.2400109, 
    0.3910023, 0.02917564, 0.0466943, 0.02434418, 0.03885964,
  0.03542721, 0.0329208, 0.3177902, 0.06522933, 0.2628425, 0.3545643, 
    0.566937, 0.4452648, 0.4229727, 0.7536872, 0.7532952, 0.3663914, 
    0.6745138, 0.3324836, 0.3143999, 0.2155863, 0.2940865, 0.1929929, 
    0.2722721, 0.2616306, 0.2901556, 0.5418071, 0.5098698, 0.4312653, 
    0.1459078, 0.1907726, 0.3023854, 0.02625921, 0.06203751,
  0.3400968, 0.237281, 0.354729, 0.3029151, 0.4137706, 0.4758334, 0.4165767, 
    0.3191842, 0.4521648, 0.4238626, 0.3339257, 0.4108237, 0.4184541, 
    0.3539873, 0.2945841, 0.2422164, 0.2649513, 0.3378752, 0.2679171, 
    0.2859998, 0.3379076, 0.2220759, 0.2475915, 0.3883034, 0.05976139, 
    0.04753751, 0.1553637, 0.2238358, 0.3990099,
  0.07150491, 0.07684118, 0.08217745, 0.08751372, 0.09285, 0.09818628, 
    0.1035225, 0.09442618, 0.09744594, 0.1004657, 0.1034855, 0.1065052, 
    0.109525, 0.1125447, 0.1475483, 0.1418978, 0.1362472, 0.1305966, 
    0.1249461, 0.1192955, 0.1136449, 0.0837395, 0.08103403, 0.07832856, 
    0.0756231, 0.07291763, 0.07021217, 0.0675067, 0.06723588,
  0.07309344, 0.05491544, 0.05156107, 0.1023467, 0.1097082, 0.05460025, 
    0.08810288, 0.155142, 0.1590969, 0.1338156, 0.04318388, 0.01340918, 
    0.02006847, 0.003001909, 0.01917542, 0.05371434, 0.0713019, 0.1798886, 
    0.04422211, 0.006239702, 0.04123161, 0.07035262, 0.07670388, 0.03250555, 
    0.1089655, 0.04979134, 0.05126306, 0.02549431, 0.06948458,
  0.03766056, 0.03311595, 0.02122986, 0.016897, 0.01690236, 0.08927576, 
    0.07799713, 0.06220961, 0.07987246, 0.08650562, 0.03461768, 0.09418587, 
    0.04431367, 0.1354341, 0.2083847, 0.2308013, 0.1740399, 0.2122963, 
    0.1276767, 0.2257636, 0.2346663, 0.2583616, 0.3019754, 0.4256939, 
    0.1843578, 0.1678512, 0.09783858, 0.0698472, 0.08502784,
  0.144897, 0.1509651, 0.1167411, 0.1810895, 0.2057299, 0.1649753, 0.196531, 
    0.1757641, 0.183196, 0.1776841, 0.1420667, 0.156644, 0.2540388, 
    0.1768219, 0.1466456, 0.1880412, 0.2450793, 0.2576752, 0.2120834, 
    0.09394005, 0.08748455, 0.05960479, 0.06488878, 0.06215246, 0.1364044, 
    0.2029821, 0.3001576, 0.2385328, 0.1490115,
  0.146904, 0.1375151, 0.1277194, 0.1205205, 0.1934453, 0.1910785, 0.1488239, 
    0.1448823, 0.1483991, 0.09563632, 0.03052008, 0.0151154, 0.06082197, 
    0.08341859, 0.1685373, 0.167436, 0.09412386, 0.08287246, 0.04951447, 
    0.08746783, 0.06138553, 0.08473426, 0.1098123, 0.03611395, 0.04755383, 
    0.2090865, 0.19098, 0.1571123, 0.1560512,
  0.04935063, 0.01697258, 0.003515996, 0.03728418, 0.01622162, 0.01523597, 
    0.04652094, 0.1262633, 0.06756192, 0.02188745, 0.006668814, 0.003308501, 
    0.02268623, 0.0323694, 0.1599056, 0.006016159, 0.006593172, 0.04090628, 
    0.1220872, 0.09887224, 0.03360002, 0.01723805, 0.00931086, 0.09213042, 
    0.03258096, 0.04107222, 0.06889605, 0.06191033, 0.03171071,
  0.003723332, 0.005387414, 0.01163789, 0.001153395, 0.0006309514, 
    0.0006128044, 0.001138077, 0.005352319, 0.008483408, 0.00390806, 
    -3.96238e-06, 3.363122e-09, 0.007949654, 0.0003741242, 0.001352388, 
    0.001396006, 0.01137582, 0.01211716, 0.005256006, 0.0004536018, 
    0.0007629926, 0.00104099, 0.004613419, 0.007668879, 0.0162326, 
    0.001187366, 0.004770741, 0.0003855023, 0.0009750421,
  0.002227657, 0.03398215, 0.007324877, 0.0006033372, -0.00113644, 
    0.0004691435, 0.0006660681, 0.001101708, 0.009954152, 0.008170331, 
    0.0008621717, 0.003078249, 0.0003715579, 0.0002678007, 0.0003659263, 
    0.001255776, 0.0003938783, 0.001322914, 3.974127e-05, 3.248774e-05, 
    0.0002078509, 0.0004768389, 0.004708142, 0.01008151, 0.02917205, 
    0.06341805, 0.0002105905, 2.25514e-06, 0.0002285785,
  0.00596242, 0.000813131, 0.1029882, 0.1000621, 0.0008720883, 0.0003463792, 
    9.536924e-05, 0.0001294618, 0.0003691137, 9.209873e-05, 0.001291522, 
    0.0002147895, 0.0001470276, 0.0001102019, 0.0003161818, 2.920777e-05, 
    0.0001363677, 0.0006060147, 4.058825e-05, 0.0004634578, 0.001064128, 
    0.003395363, 0.009323569, 0.1312222, 0.05665366, 0.04840311, 
    -2.179092e-05, 0.001094953, 0.003244342,
  4.324339e-05, 0.0303524, 0.0003987002, 0.001211003, 0.0001049497, 
    0.002451174, 0.002696406, 3.172516e-05, 0.08319874, 0.1096744, 
    0.0006088094, 0.0002463633, 0.0007179244, 0.001764126, 0.002112234, 
    0.000151671, 0.00045381, 3.551585e-05, 7.340808e-06, 0.00016715, 
    0.0008413383, 0.007275453, 0.01565911, 0.06504031, 0.02878517, 
    0.001804391, 0.0001032962, 6.924911e-06, 0.001568285,
  2.519292e-11, 1.332698e-10, -1.423364e-10, 0.007447142, 0.006615931, 
    0.0002705811, -0.001525533, 0.0007451908, -0.000255989, 7.774537e-05, 
    0.001849561, 0.0001408091, 0.0002432792, 0.0003952651, 0.0001285175, 
    0.0001377366, 0.0001088024, 7.084961e-05, 0.0003084603, 0.0005063663, 
    6.190487e-05, 6.158793e-05, 0.178442, 0.02911383, -7.033553e-07, 
    0.0001821246, 0.0007683189, 0.0006495543, 0.007559663,
  6.234825e-09, -6.93369e-07, 0.0001127331, 0.0001794525, -2.713229e-07, 
    0.0002796821, 0.01296353, 0.0007209735, 0.01424557, 0.03172095, 
    0.001605857, 0.003357874, 0.0004615724, 0.0004418796, 0.000359274, 
    0.0008502725, 0.00125909, 0.0006279206, 0.008172469, 0.005586036, 
    0.0007286429, 0.06963179, 0.001052939, -0.001195231, 0.0002283995, 
    0.0002926892, 0.001679366, 6.449522e-05, -1.61879e-05,
  0.00030103, 0.01199558, 0.005755065, 0.005399416, 0.0568726, 0.000217798, 
    -0.0003039745, 0.01639981, 0.02668128, 0.02709293, 0.03587633, 
    0.004054532, 0.003270523, 0.004151965, 0.006631164, 0.03341126, 
    0.03355177, 0.003314461, 0.009897043, 0.005065285, 0.06840123, 0.1026656, 
    0.06308807, 0.007599085, 0.006409192, 0.003606592, 0.002756497, 
    0.002004958, 0.005491617,
  0.01332428, 0.05136697, 0.006137342, 0.2619282, 0.007918259, 0.05296953, 
    0.06450523, 0.01121099, -6.362188e-05, 0.04097392, 0.1110807, 
    0.006266539, 0.01379943, 0.01235033, 0.01342491, 0.04820286, 0.0804977, 
    0.05073863, 0.01272818, 0.1910579, 0.1745468, 0.06514709, 0.1546744, 
    0.07312559, 0.01890938, 0.01625811, 0.01486187, 0.01880636, 0.04592867,
  0.1164654, 0.2041964, 0.1670765, 0.208846, 0.1621392, 0.1773849, 0.1083, 
    0.2907343, 0.235439, 0.1019277, 0.03681328, 0.4280832, 0.003994955, 
    0.0006761463, 0.06495535, 0.1448453, 0.1671618, 0.09677552, 0.04332203, 
    0.3397819, 0.1018067, 0.1105389, 0.233268, 0.5835962, 0.1791893, 
    0.08419238, 0.02921597, 0.02403733, 0.07816183,
  0.02536537, 0.43221, 0.4244689, 0.3391972, 0.5400905, 0.2803599, 0.4142415, 
    0.3517584, 0.4519415, 0.4127656, 0.5031287, 0.6251554, 0.4944218, 
    0.2596453, 0.277893, 0.2538287, 0.6167944, 0.3103979, 0.3888462, 
    0.3370017, 0.5828839, 0.5054484, 0.139432, 0.2535251, 0.3858695, 
    0.03096939, 0.03978384, 0.0215184, 0.03207372,
  0.03100325, 0.02808558, 0.4015341, 0.0569714, 0.2474532, 0.3263193, 
    0.4985603, 0.4405281, 0.54878, 0.6810784, 0.7727576, 0.5138268, 
    0.4748471, 0.2717897, 0.2619521, 0.1964921, 0.2728159, 0.2239839, 
    0.2417414, 0.2062122, 0.2511518, 0.4492812, 0.3825325, 0.4510917, 
    0.1099739, 0.1470963, 0.3479586, 0.02804905, 0.05600245,
  0.2989557, 0.2199288, 0.3371213, 0.2621923, 0.3201458, 0.4018629, 
    0.3354977, 0.2568425, 0.3478339, 0.3258116, 0.225693, 0.2633515, 
    0.2808408, 0.2681332, 0.225125, 0.1944945, 0.214542, 0.2502576, 
    0.1553519, 0.1847539, 0.2484573, 0.2012062, 0.2807632, 0.4521835, 
    0.08337008, 0.06902114, 0.1333292, 0.2247162, 0.3305343,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -5.411817e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2.164727e-05, 0, 0.0002055592, 0, 
    0.0001886555, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.305299e-06, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, -3.355794e-06, 0, 0, 0, 0, 0, 0, 0, -3.788272e-05, 0, 0.0003083388, 
    0, 0.003046372, 0, 0, 0, 0, 0, 0, 0, 0, -6.883334e-06, -2.098926e-05, 
    -3.034003e-05, 0, 0, 0,
  0, 0, 0, 0, 2.619012e-05, 0, 0, 0, 0, 0, 0, 0, -3.761071e-06, 0, 
    0.001257751, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -2.587943e-06, 0, 0, 0,
  0, -2.204198e-05, 7.845841e-06, 0, -4.410226e-05, 0, 0, 0, 0, 0, 0, 
    -3.74637e-06, 0, 0, -1.887482e-05, -1.567366e-05, 0, 0, 0, 0, 0, 0, 0, 0, 
    -8.605624e-05, 0, 0, 0, 0,
  0, 0, -1.829965e-05, -5.380213e-07, -7.121686e-05, 0, 0, 0, 0, 0, 
    -0.0001177985, -9.494125e-06, 0.0003823341, 0, 0.005744819, 0.0005043011, 
    -5.206281e-06, 0, 0, 0, 0, 0, 0, 0.0002274138, 0.000573748, -5.80938e-05, 
    0, 0, 0,
  0, 0, 0, 0, 8.913322e-05, -3.037261e-08, 0, 0, 0, 0, 0, 0, -1.382865e-05, 
    0, 0.001234856, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2.321504e-05, 0, 0, 0, 0, 0, 0, 0, 
    0.0002067014, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, -9.846931e-06, 0, 0, 0, 0, 0, 0, -3.264982e-08, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, -7.704073e-05, 0, 0, 0,
  0, -3.708341e-05, 1.257235e-05, 0, 0.0008627046, 0, 0, 0, 0, -7.637327e-05, 
    0.0009609844, -4.749408e-05, 0, 1.446114e-05, -6.034203e-05, 
    -0.0001905254, -0.0001286665, 0, 0, 0, 0, 0, 0, 0, 0.000957779, 0, 0, 0, 0,
  0, -1.730894e-05, 4.034965e-05, -1.076043e-06, -0.000206784, 0, 0, 0, 0, 0, 
    -0.0003256857, -2.373531e-05, 0.001285338, 0, 0.009510338, 0.005873011, 
    -7.753933e-05, 0, 0, 0, 0, 0, 0, 0.0002402589, 0.002055614, 
    -0.0001021359, 0, 0, 0,
  0, 0, 0, 0, -9.546314e-05, -3.922419e-05, 0, 0.001939925, 0.0001822327, 0, 
    0, 0, -3.660685e-05, 3.302647e-05, 0.00302186, 7.750856e-05, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.0003210028, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0008179464, -2.126973e-05, -5.971547e-06, 
    0, 0, 0, 0, 0, 0.0005625795, -6.601838e-05, -3.391533e-05, 0, 0, 0, 0, 0, 
    0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, -8.772076e-06, 0, 0.0001818331, 0, 0, 0, 0, 0, 0, 0, 0, 
    -7.457583e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -3.008e-07, 0, 0, 0,
  0, 0, 0, 0, 0.0001744413, 0, 0, 0, 0, 0, 0, -6.529964e-08, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, -0.0001051216, -3.501155e-06, 0, 0,
  0, -8.518782e-05, 0.0005686621, 0, 0.002149958, 0, 0, 0, 0, 0.0006684253, 
    0.002198623, -0.0001616019, 0, 0.002932171, -0.0003104772, -0.0002700041, 
    0.001263337, 0, 0, 0, 0, 0, 0, 0, 0.003843983, -4.988793e-05, 0, 0, 0,
  0, -4.327235e-05, 0.002678841, -2.211369e-06, -4.720793e-05, 8.998202e-06, 
    0, 0, 0, 0, -0.0005098439, -3.586598e-05, 0.002431631, -0.000231297, 
    0.0201702, 0.00769698, -8.04275e-05, 0, 0, 0, 0, 0, 0, 0.005057122, 
    0.003035691, -0.0001516381, 0, 0, 0,
  0, 0, 0, 0, 0.004836143, -0.0001117378, -7.7178e-05, 0.003483181, 
    0.0003686855, 0, 0, 0, -0.0001458485, 0.0006570484, 0.004998479, 
    9.698674e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.00242975, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.003507685, -9.627608e-05, 0.002349882, 0, 
    0, 0, -3.662099e-05, 0, 0.001353344, 0.0009397238, 0.000250668, 0, 0, 0, 
    0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.613279e-10, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, -2.89054e-05, 0, 0.002022218, 0, 0, 0, 0, 0, 0, 0.0003833752, 0, 
    0.0009604525, -9.79977e-07, 0, 0, 0, 0, 0, 0, 0, 0, 0, -3.560461e-05, 0, 
    0, 0,
  0, 0, 0.0001313514, 0, 0.001062501, 0, 0, 0, 0, 0, 0, -8.191415e-06, 0, 0, 
    0.002920393, 0, -0.0001348043, -1.411167e-05, 0, 0, 0, 0, 0, 0, 0, 
    -0.0002092977, -3.30609e-05, 0, 0,
  0, -0.0001636711, 0.001748721, 0, 0.007112237, 0, 0, 0, 0, 0.002087721, 
    0.009561258, 0.0007410301, 0, 0.009415463, -0.0009209231, 0.001013529, 
    0.01336929, 0, 0, 0, 0, 0, 0, 0, 0.005451963, -0.0002140499, 0, 0, 0,
  0, -0.0001038536, 0.009504644, -6.432496e-06, 0.001228527, 1.677747e-05, 0, 
    0, 0, 0, -0.0003767808, 0.0002219216, 0.004363848, 0.0001572723, 
    0.04123167, 0.02108771, 0.000798827, 0, 0, 0, 0, 0, 0, 0.005896872, 
    0.007598687, 0.0007556813, 0, 0, 0,
  0, 0, 0, 0, 0.01809419, 0.002207413, 0.0001038868, 0.007735374, 
    0.002143939, -8.921206e-06, 0, -5.201483e-05, -0.0001920927, 0.001878354, 
    0.005610707, 4.999844e-05, 0, 0, -1.662938e-05, -9.51632e-08, 0, 0, 0, 0, 
    -2.979329e-10, 0.006716309, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, -9.494938e-05, 0.006880656, -2.106987e-05, 
    0.006310261, 0, -5.958201e-06, 0, -0.0001087368, 0, 0.004594787, 
    0.002815763, 0.002690571, -3.49759e-05, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0.0001524975, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, -3.733483e-05, -0.000123488, 0, 0, 0, 0, 0.0001916344, 0, 
    0, -1.582747e-07, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, -8.199934e-05, 0, 0.004334837, 0.000622252, 0.0008433596, 0, 0, 0, 
    -9.113525e-06, 0.002534018, 0, 0.003492155, 0.0009109825, 0, 0, 
    0.0001146481, -2.283354e-05, 0, 0, 0, 0, 0.001203725, 0.003692332, 0, 0, 0,
  0, 0, 0.0005232688, 0, 0.004233647, -1.091244e-05, 0, 0, 0, 0, 0, 
    -0.0001072365, 0, 0, 0.006494161, 0, 7.790307e-05, -3.312892e-05, 
    -1.757072e-06, 0.0003457669, 0, 0, 0, 0, 6.509421e-05, 0.004340635, 
    0.002272922, 0, 0,
  0, 0.0002212933, 0.003479674, -1.021829e-05, 0.01973913, 0, 0, 0, 0, 
    0.007722528, 0.02591678, 0.003186967, 0, 0.01504243, 0.004605784, 
    0.005486692, 0.02407812, -1.246363e-06, 0, 0, 0, 0, 0, 0, 0.009311444, 
    0.0007238901, -1.635368e-05, 0, 0,
  0, -0.0002378636, 0.02144559, -3.454688e-06, 0.00528594, 3.161917e-05, 0, 
    0, 0, 0.0001222261, 0.002087893, 0.00156732, 0.004872798, 0.002239809, 
    0.07635342, 0.04449753, 0.001015226, 0, 0, 0, 0, 0, 0, 0.009966062, 
    0.01559706, 0.002045607, 0, 0, 0,
  0, 0, 0, 0, 0.02876141, 0.009442593, 4.673827e-05, 0.01036226, 0.007361908, 
    0.0002193589, -5.322453e-06, 2.456397e-05, 0.0006015901, 0.005235968, 
    0.009140308, 0.003785818, 0, 0, -9.372171e-05, -1.022424e-06, 0, 0, 0, 0, 
    0.0002716395, 0.01583454, 0, 0, 0,
  0, 0, 0, 0, 0, -6.004461e-06, 0, 0, 0, -0.0001660465, 0.01256623, 
    0.001972324, 0.01146572, -1.085057e-05, -2.166481e-05, 0, 2.600949e-05, 
    0.0001458515, 0.01380934, 0.004045996, 0.004124697, -0.0001365346, 0, 0, 
    0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.934141e-05, 0, 0, 0, 0, 0, 
    -0.0003024316, 0, -4.79251e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, -6.339394e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -1.493165e-05, 0, -1.974749e-05, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 5.912656e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.0004690716,
  0, 0, 0, -1.367418e-05, 0.0001131214, 0, 0.002888317, 0.004277149, 
    -2.251256e-05, 0, 0, -5.778927e-06, 0.00946449, -1.007419e-06, 0, 
    0.001166816, 0, 0, 0, 0, 0.0005620924, -1.194809e-05, 0, 4.37516e-06, 0, 
    0.0006894576, 0.001140498, 0, 0,
  0, 0, 0, -0.0002023822, -0.0001742535, 0.0167493, 0.00470407, 0.001547253, 
    0, 0, -1.474446e-06, 0.003667439, 0.00881574, 0.0002007215, 0.01761441, 
    0.009835673, 0.0005177873, -8.994566e-06, 0.007854253, 0.001564228, 
    -4.797883e-05, 0, 0, 0, 0.003042853, 0.01898532, -4.774523e-05, 
    0.0002062982, 0.0002026607,
  0, 0, 0.001825667, -3.03979e-05, 0.009718906, 0.003173212, 0.006073666, 0, 
    0, 0, -3.093643e-05, 0.0008707286, 0, 0, 0.01565668, 2.940392e-06, 
    0.001158487, 0.004778305, 6.524626e-05, 0.0004235032, 0, 0, 0, 0, 
    0.0005774384, 0.01475851, 0.006041005, 0.001114965, 0,
  0, 0.000304795, 0.007954234, -2.982141e-05, 0.0628543, 0, 0, 0, 0, 
    0.01379201, 0.03681504, 0.009047956, 0.0001313323, 0.0206563, 0.01738952, 
    0.01153957, 0.04410361, 0.0001420093, -1.894541e-05, 0, 0, 0, 0, 
    -2.349529e-07, 0.01602075, 0.002659546, -0.0002244154, 0, 0,
  0, -0.0005354402, 0.04083, 0.0002921523, 0.01405207, 0.0002428889, 0, 
    -4.311789e-09, 0, 8.463093e-05, 0.004475083, 0.006461367, 0.01425874, 
    0.01711176, 0.1208765, 0.06621881, 0.002736933, 0, 1.322215e-08, 
    1.815113e-05, 0, 0, 0, 0.01809363, 0.03941113, 0.003392377, 
    -2.140535e-05, 0, 0,
  0, 0, -3.44033e-06, 0, 0.0488857, 0.01894327, 0.003022105, 0.01481655, 
    0.01672203, 0.005823737, -1.596736e-05, 0.001395385, 0.01313026, 
    0.01681657, 0.02308582, 0.005432924, -5.619211e-06, 0, -0.0001016396, 
    -1.675642e-06, 3.289904e-05, 0, -2.431804e-11, 0, 0.002246579, 
    0.03048799, 0, 0, 0,
  0, 0, 0, 0, -1.605816e-05, -3.183215e-05, -1.873466e-05, 0, 0, 
    -0.0003035782, 0.03882091, 0.005846588, 0.02142661, -5.533993e-05, 
    -4.323841e-05, 0, 0.001442336, 0.01096376, 0.03157244, 0.008585386, 
    0.007237005, 0.000299134, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0004271441, 0.0001421168, -9.0417e-08, 0, 
    0, 0, -1.514636e-06, 0.004345967, 0, -0.0001406288, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, -0.0001402356, 4.051666e-07, 0, 0, 0, 
    -1.588982e-08, 0, 0, 0, -4.460104e-07, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -3.102881e-06, 0, 0, 0, -5.736999e-06, 0, 
    0, 0, 0, 0, 0, -2.569346e-05, 1.963125e-06, 0.0005531273, 0, 0.001398927, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8.581055e-05, 0, 0, 0, 
    0, 0, 0, 0, 0, -1.022649e-06, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, -2.983965e-07, 0, 0, 0, 0.0004398928, 0, 7.709936e-05, 0, 0, 0, 0, 
    0, 0, 9.698882e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001259913,
  0.0006791758, 0.0004848015, -9.010217e-06, 0.001022816, 0.002066508, 
    0.003334102, 0.01271961, 0.0126281, 0.002441818, 0, 0, -0.0001335913, 
    0.01972413, 0.003636717, -4.343123e-05, 0.02117185, 0.001239826, 
    -6.248232e-06, 0, -5.983756e-08, 0.003063046, -0.0001117415, 0.001474302, 
    0.001102474, 0, 0.01455349, 0.004093632, 0.006124422, 0.002499427,
  0.0004341056, -1.477604e-08, 0.001421848, 0.0009904578, 0.002803102, 
    0.02946606, 0.01298876, 0.006377836, 0, 0, 0.00140978, 0.03267098, 
    0.01404136, 0.005203616, 0.02579325, 0.03513251, 0.003824327, 
    0.0009813826, 0.0197228, 0.009178149, -0.0002583792, 0, 0, 0, 
    0.006730125, 0.04281167, 0.00567891, 0.00411927, 0.004430027,
  0, 0, 0.003956989, -9.604978e-05, 0.01226328, 0.008593735, 0.01650999, 
    -3.221673e-07, 0, 0, 0.001166245, 0.003806479, -1.50341e-11, 
    -2.615089e-06, 0.05362194, 0.002055658, 0.005437112, 0.02697904, 
    0.002053184, 0.0004354845, 0, 0, 0, 0, 0.001600357, 0.01973057, 
    0.01441913, 0.01035842, 0,
  0, 0.007375711, 0.01865592, 9.43769e-05, 0.126311, 0, 0, -5.974359e-11, 0, 
    0.02357842, 0.05131254, 0.0316243, 0.0005881288, 0.05090746, 0.06812733, 
    0.02715004, 0.06431433, 0.001386528, 0.0008322662, 0, 0, -1.923023e-09, 
    0, -9.860679e-06, 0.04757254, 0.0133185, 0.0004350391, 0, 0,
  0, 8.525419e-05, 0.0773503, 0.002190161, 0.025558, 0.000305338, 
    -7.733657e-06, -9.888948e-06, -9.47586e-06, 0.001676356, 0.00796672, 
    0.02212799, 0.03177129, 0.1116473, 0.2006532, 0.08099023, 0.006698556, 
    -3.933087e-06, 3.665068e-07, 8.373832e-05, 0, 0, 3.129363e-09, 
    0.04041985, 0.1043211, 0.01805886, 0.0001330054, 0, 0,
  0, 0, -2.069667e-05, 0.00035544, 0.07911566, 0.03796713, 0.005766421, 
    0.02506853, 0.04892775, 0.008732835, 8.067803e-05, 0.003678867, 
    0.02616047, 0.06081526, 0.03522874, 0.00967632, -0.0001186007, 
    4.087287e-07, 0.0007094232, -1.590486e-05, 0.004261067, 0, 6.686582e-10, 
    2.094273e-05, 0.005947823, 0.0521461, 0.0007335815, 0, 0,
  0, 0, 0, -1.326699e-06, 0.0005521991, -9.383606e-05, -0.0001202708, 
    -4.163472e-06, 2.850877e-06, 7.41792e-05, 0.08137145, 0.0215707, 
    0.03466106, 0.003760609, -9.210064e-05, 0, 0.003030494, 0.03484144, 
    0.05050503, 0.02555477, 0.01744978, 0.008184843, 0, 0, 0, -1.2738e-07, 
    -4.91628e-22, -1.212931e-08, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0.000320491, 0.006339565, 0.002138555, 
    0.000269691, -8.162412e-06, 1.054545e-07, -1.675503e-07, 0.009223685, 
    0.01826597, -0.0002331416, 0.002990636, 1.256642e-05, 0.0006932949, 0, 0, 
    0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, -0.0003352475, 4.422517e-05, -4.099304e-08, 0, 
    0, 0.0004258379, -1.540956e-05, -5.393908e-05, -1.879939e-05, 
    0.0001851952, -3.951803e-08, 0, 0, -4.248953e-05, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.005042839, -1.070153e-06, 0, 0, 0, 
    -6.926712e-05, 0, -8.526948e-06, 0, 0, 0, 0, 0.003557879, 0.004966138, 
    0.006803643, 0, 0.006927068, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5.895911e-05, 0, 0, 0, 
    0, 0, 0, -3.895425e-05, 0, 0.0003063882, -6.371976e-06, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  -2.888441e-05, 0, 0, -2.217327e-05, 0.0006193545, 0, 0, 0.001841748, 
    0.001914409, 0.001422811, 0, 0, 0, 0, 8.029348e-05, -1.122122e-05, 
    0.0002353499, 0.0007518224, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.002831605,
  0.004900619, 0.003889616, 0.0007222082, 0.004971705, 0.01298604, 
    0.01700126, 0.02691013, 0.03119455, 0.00769662, 0.0004267017, 0, 
    0.00108825, 0.02621461, 0.0101679, 0.0002606212, 0.03508247, 0.003639604, 
    0.001276822, -2.924868e-07, 0.0006180527, 0.01191483, 0.01476941, 
    0.006880469, 0.002453078, -2.815916e-07, 0.03056456, 0.008159772, 
    0.01932796, 0.01336127,
  0.003699846, -4.324634e-05, 0.003998808, 0.007578952, 0.01093776, 
    0.04347589, 0.01541115, 0.01203761, 1.178028e-07, -3.173579e-10, 
    0.007627747, 0.0576126, 0.02067137, 0.008833398, 0.0565801, 0.1039933, 
    0.01109081, 0.01695427, 0.04643936, 0.02871964, 8.091995e-05, 
    -3.760363e-06, 0.001001351, 0, 0.008529303, 0.06015984, 0.02052509, 
    0.009713956, 0.006999327,
  0, -4.419994e-07, 0.008483251, 0.007596141, 0.01752124, 0.02258971, 
    0.02303525, 0.0003230185, 0, -2.265077e-09, 0.02307926, 0.01437456, 
    0.001290363, 0.001145513, 0.1449073, 0.02071023, 0.0168133, 0.0641297, 
    0.009469093, 0.001666877, -8.870006e-05, -1.859043e-06, 0, 0, 0.0146787, 
    0.06557847, 0.02255021, 0.01531976, -5.104947e-07,
  7.604638e-07, 0.04120941, 0.06305702, 0.002044597, 0.2280278, 
    -4.253391e-06, -8.674409e-06, 0.0008619371, 4.261974e-06, 0.06802974, 
    0.1473403, 0.1867903, 0.01245188, 0.123649, 0.2518582, 0.1011743, 
    0.09309044, 0.01096297, 0.001987257, 0, 1.270615e-05, -8.171525e-05, 0, 
    0.0009720082, 0.2262402, 0.05048063, 0.00923691, 0, -4.268207e-08,
  2.366685e-07, -0.0004465393, 0.1531813, 0.01317301, 0.04428056, 
    0.001482981, 0.0003836028, -2.869274e-05, -2.848486e-05, 0.01977962, 
    0.03515016, 0.2063413, 0.192521, 0.3622388, 0.5170559, 0.1429812, 
    0.02702928, 0.004141601, 3.584547e-05, 0.005032141, 0.001155584, 0, 
    0.003098253, 0.160957, 0.3356265, 0.07604975, 3.583489e-05, 3.011743e-05, 0,
  -1.900338e-09, 0.0007061443, -7.368631e-05, 0.00174102, 0.1192872, 
    0.07541607, 0.01763067, 0.03763256, 0.116815, 0.05607331, 0.02224665, 
    0.06438944, 0.1222479, 0.3016421, 0.1195659, 0.03490274, 0.01143228, 
    0.0001528945, 0.006084788, -3.400235e-05, 0.008516719, 0, 1.751078e-06, 
    0.000822692, 0.0196884, 0.1138932, 0.0009842924, 0.001294008, 0,
  4.922578e-05, 0, 4.210171e-09, -1.647635e-05, 0.003749297, 0.0001214492, 
    -0.0001321845, -3.993464e-05, 7.576167e-06, 0.001828017, 0.1389005, 
    0.08424848, 0.05284208, 0.03690052, 0.0003377388, 0.0001854852, 
    0.00585204, 0.05028008, 0.06824112, 0.04247743, 0.02471165, 0.01916045, 
    -8.43443e-09, 1.069197e-06, 9.065793e-06, 0.0006052437, 0.0005690894, 
    2.668467e-06, 1.194279e-07,
  1.33437e-07, 0, 0, 0, -3.311015e-08, 4.192423e-08, -8.996619e-06, 0, 0, 
    0.0006418108, 0.01380742, 0.004039845, 0.002624214, -2.963976e-05, 
    0.000385129, -8.823432e-06, 0.02921009, 0.03951525, 0.01976335, 
    0.01148713, 0.001548205, 0.002821053, -6.602606e-06, -1.393604e-10, 
    -3.535983e-10, 0, 0, 0, 9.997381e-10,
  0, 0, 0, 0, -4.687213e-07, 1.400029e-06, -2.073041e-09, 0, 0, 0.003638391, 
    0.007018988, 0.0001495246, 0.004467545, 2.690365e-05, 0.01286008, 
    0.008685919, 0.008336734, 0.01722179, 0.004231209, -5.038129e-05, 
    -4.72745e-05, -1.97201e-06, -0.0001325785, 0.0009761456, 7.494345e-05, 
    5.105577e-06, 0.0005310205, 0.00263093, 0,
  0.0001006991, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01226187, 2.132087e-05, 
    2.783348e-06, 0.001898657, 7.517463e-06, 0.01478477, -9.930837e-05, 
    0.008416323, -6.435976e-06, 0, 0, 0, 0.009766797, 0.01901954, 0.01517856, 
    0.002633793, 0.01570447, 0.004136106, 1.533683e-05,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0006674352, 0.003445049, 
    0, 0, 0, 0, 0, 0, 0.0006303963, -3.936642e-05, 0.005403225, 0.00030827, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.001297346, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0.001098575, -2.724547e-08, 0, -2.603125e-05, 0.002470239, 0.003760824, 
    0.0004873776, 0.006788106, 0.004353661, 0.002867071, -1.621699e-05, 
    0.002798231, -1.239107e-05, -4.728504e-05, 0.00525, 6.320034e-05, 
    0.007890087, 0.004934, -0.0001447803, 0, 0, 0, 0.001207756, 
    -1.494226e-06, -1.735839e-05, -0.0001888003, -0.0001438787, 0.001272921, 
    0.00424495,
  0.01199305, 0.01326651, 0.004976539, 0.0148866, 0.02153966, 0.03372924, 
    0.03680836, 0.04314072, 0.02641841, 0.003960464, -7.542477e-05, 
    0.005826196, 0.03230171, 0.0259081, 0.007780053, 0.04976007, 0.01200518, 
    0.01209495, 8.50118e-05, 0.005812222, 0.02267191, 0.03692789, 0.01542496, 
    0.005125936, -6.33478e-05, 0.04430323, 0.03145695, 0.04310786, 0.03595288,
  0.01964346, 0.002998437, 0.006379841, 0.02320336, 0.02181162, 0.1377992, 
    0.06164619, 0.02975917, 0.004964491, 0.0027269, 0.01574946, 0.07804634, 
    0.05112247, 0.0223294, 0.1001586, 0.1977101, 0.0765844, 0.07771589, 
    0.07579617, 0.06700998, 0.01557577, 0.001048409, 0.003471339, 
    0.0003864197, 0.02033043, 0.1033816, 0.1048452, 0.06270313, 0.01350536,
  1.797171e-07, 7.087993e-06, 0.04936657, 0.05081982, 0.1091357, 0.1910045, 
    0.1182829, 0.04037271, 0.002327082, -5.128182e-05, 0.04245333, 
    0.03018238, 0.002071628, 0.009935747, 0.231985, 0.09543817, 0.1133583, 
    0.1748345, 0.1260465, 0.006693775, -0.0001750416, 0.04280309, 
    -8.096823e-06, -5.334294e-05, 0.05598814, 0.1798278, 0.1202667, 
    0.07256082, -0.0001030069,
  -1.506964e-06, 0.1502125, 0.2416747, 0.01546609, 0.2500316, 0.03758202, 
    0.005313839, 0.02416809, 3.111099e-06, 0.05419405, 0.1400899, 0.181324, 
    0.01960467, 0.1180485, 0.2120841, 0.1639504, 0.2024663, 0.1552648, 
    0.07161902, 1.293531e-06, 0.002185954, 0.02173482, 9.463181e-06, 
    0.003176797, 0.2374624, 0.2167869, 0.167786, 0.01941161, -2.157099e-06,
  0.004554207, 0.08063073, 0.547279, 0.133389, 0.09908686, 0.02288711, 
    0.05214839, 0.0006049352, 0.02135222, 0.0653101, 0.03688906, 0.2022766, 
    0.1439762, 0.3016632, 0.4624272, 0.1611137, 0.05699782, 0.04838118, 
    0.02638107, 0.01433843, 0.03211064, 4.955364e-07, 0.0440504, 0.4088044, 
    0.4499157, 0.3025897, 0.1821212, 0.07753924, 3.377612e-09,
  1.393611e-05, 0.03693893, 0.1209612, 0.07279558, 0.2168993, 0.3171855, 
    0.09373235, 0.1325538, 0.3303906, 0.2572908, 0.07610178, 0.1121249, 
    0.122885, 0.2663364, 0.08778492, 0.01942401, 0.00828691, 0.007034523, 
    0.0126673, 0.008335127, 0.01386007, 2.760787e-06, 3.705371e-06, 
    0.1558198, 0.1852766, 0.2385941, 0.1604761, 0.03064413, -4.741646e-06,
  0.0002190313, 4.254267e-06, 0.0001903057, -1.478893e-05, 0.02673538, 
    0.01009888, 0.005504407, 0.0001365966, 0.005167732, 0.06344812, 
    0.1779229, 0.07571298, 0.048829, 0.02513265, 5.144504e-05, 0.0001208692, 
    0.02668103, 0.1202106, 0.1963027, 0.1380832, 0.1261386, 0.03939017, 
    0.0001592764, 3.338696e-06, 6.541795e-06, 0.003700294, 0.002212298, 
    0.07825641, 0.000451015,
  3.26802e-05, 6.389278e-05, 3.614507e-10, 4.102625e-08, 7.375892e-06, 
    0.000132613, 0.0001877665, 0, 0, 0.0001075959, 0.03281474, 0.005757385, 
    0.01374387, 0.002513112, 0.009578724, -3.120253e-05, 0.04419163, 
    0.07111388, 0.1033452, 0.09036093, 0.1210033, 0.02889165, 0.004034833, 
    1.434907e-06, -6.320651e-07, 1.903093e-06, 1.11062e-06, -5.434062e-05, 
    3.881249e-05,
  0, -6.739661e-06, 0, 0, 0.0003071664, 0.001590365, -2.028742e-05, 0, 0, 
    0.01197505, 0.02206219, 0.02335635, 0.01290741, 0.01146228, 0.03357902, 
    0.02903728, 0.07145914, 0.04900904, 0.009600668, 0.006944931, 
    -0.0002005077, 0.02414108, 0.0196345, 0.01638376, 0.005849571, 
    0.00180668, 0.006644174, 0.00650145, -1.023609e-06,
  0.0180292, -9.185785e-10, 0, 0, 0, 0, 0, 0, 0, -2.486041e-06, 0.01732391, 
    0.006862944, 0.0009021315, 0.006644265, 0.0008457179, 0.04427641, 
    0.008513942, 0.02479338, 0.006531467, 0, 0, 0.0002519259, 0.01795719, 
    0.06496896, 0.04207335, 0.01826463, 0.02540589, 0.01356591, 0.01029121,
  -5.329653e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.009601e-05, 
    -4.476407e-05, 0, 0, 0.003497161, 0.009378632, 0.002384975, 0, 0, 0, 0, 
    -1.056942e-05, 0.001621789, 0.000374183, 0.01960672, 0.006162709, 
    -8.902974e-05,
  0, -2.64659e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, -1.365993e-05, 0.003161544, -1.622401e-05, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -6.108413e-05, -4.992158e-05, 
    0.001437047, -7.894189e-06, 0, 0, 0, 0, 0, -1.499046e-05, 0, 0, 0, 0, 0,
  0.00253432, 0.0002421149, 4.344661e-06, 4.505027e-05, 0.005985839, 
    0.008846561, 0.0004740669, 0.008849179, 0.006828503, 0.003497281, 
    -7.351697e-05, 0.004661578, -0.0001041583, 0.009053182, 0.01935771, 
    0.02513658, 0.03913943, 0.02255973, 0.007734384, -6.990698e-06, 
    -2.019868e-08, 0, 0.004684168, -8.356632e-05, 0.005094693, 0.004828003, 
    0.006749574, 0.006701171, 0.006339101,
  0.0434913, 0.03935817, 0.0465652, 0.05512681, 0.06044402, 0.1051675, 
    0.1346736, 0.07915524, 0.05341062, 0.03400053, 0.04044548, 0.04378543, 
    0.09601144, 0.06401011, 0.05503746, 0.1079523, 0.0824294, 0.04743214, 
    0.02192465, 0.0276592, 0.056832, 0.1060329, 0.06478079, 0.02108598, 
    0.01073413, 0.07116105, 0.05669356, 0.08774839, 0.091479,
  0.07134534, 0.03016225, 0.02736204, 0.06013344, 0.0600079, 0.1679326, 
    0.1035212, 0.1120262, 0.01897444, 0.02061371, 0.0377572, 0.112835, 
    0.09100204, 0.03975576, 0.1404227, 0.2483219, 0.09946969, 0.1599888, 
    0.1643969, 0.2056434, 0.1036375, 0.04592209, 0.03368589, 0.008120751, 
    0.0935532, 0.168663, 0.1644527, 0.1662142, 0.08584785,
  2.616819e-06, 1.431762e-05, 0.107485, 0.05408167, 0.09369113, 0.190993, 
    0.1192465, 0.05672863, 0.004454252, -0.000135879, 0.07111055, 0.04168819, 
    0.01792308, 0.01062189, 0.2419811, 0.1082238, 0.1666693, 0.2323442, 
    0.1709515, 0.1120286, 0.04823182, 0.006041581, 8.342806e-07, 
    0.0001802543, 0.07699787, 0.17242, 0.1379771, 0.1099145, 0.0009352767,
  6.753327e-06, 0.118471, 0.2032633, 0.01441253, 0.2160598, 0.01889998, 
    0.004652374, 0.02018137, 3.745635e-06, 0.03965195, 0.1462806, 0.1312166, 
    0.0106293, 0.1054636, 0.1861781, 0.1389649, 0.196251, 0.1020572, 
    0.08746952, 0.04507861, 0.02747907, 0.01204128, 6.722874e-06, 
    -1.00419e-06, 0.1869674, 0.2022809, 0.1787822, 0.005453383, 1.639339e-06,
  0.00253944, 0.04429205, 0.5126739, 0.1073608, 0.08441837, 0.009805275, 
    0.03130347, 0.0006925734, 0.009316475, 0.03851675, 0.0280384, 0.1675249, 
    0.111855, 0.2464746, 0.3946953, 0.1290619, 0.03425049, 0.04307147, 
    0.01861532, 0.01508033, 0.03628626, 8.672463e-08, 0.02560717, 0.3481098, 
    0.3822902, 0.2789527, 0.1480386, 0.02569285, 9.235533e-09,
  4.545124e-06, 0.01958719, 0.0556033, 0.0587641, 0.1824538, 0.2329928, 
    0.06394226, 0.09191661, 0.2723204, 0.2009026, 0.04582507, 0.07787045, 
    0.08120101, 0.2121233, 0.09423323, 0.0130217, 0.009363208, 0.005181363, 
    0.006445492, 0.003336451, 0.01616547, 1.638095e-06, 8.502921e-05, 
    0.06640791, 0.1386768, 0.2150756, 0.1142443, 0.01802942, 9.132374e-07,
  3.376161e-05, 4.041872e-06, 1.248706e-05, 0.0002386456, 0.02147632, 
    0.006012949, 0.000154207, 0.0002850109, 0.002403747, 0.03897543, 
    0.1625542, 0.05661758, 0.04298726, 0.01924166, -0.000116045, 
    3.521985e-05, 0.02857105, 0.124753, 0.1640638, 0.09475532, 0.08745287, 
    0.02789937, 6.879774e-05, -1.115668e-06, -2.597253e-05, 0.0003566771, 
    9.231658e-05, 0.08245328, 0.04288063,
  0.1154633, 0.003940414, -1.132698e-07, 6.445101e-07, 3.112909e-06, 
    4.397471e-05, 1.346612e-05, 0, 0, 0.0001190191, 0.03131723, 0.01473562, 
    0.02251377, 0.001020064, 0.01354731, 0.0002913106, 0.04100832, 0.1008078, 
    0.1441769, 0.09966088, 0.1211517, 0.03191114, 0.002966504, 0.0001138993, 
    -1.994645e-06, 2.898773e-07, 0.0001517283, 0.006215121, 0.06318755,
  -1.217875e-07, 0.001805252, -4.783177e-09, 0, 0.003500067, 0.005871588, 
    0.007520122, 0, 0, 0.03772298, 0.02286575, 0.03511195, 0.01476711, 
    0.02399118, 0.06247751, 0.09126998, 0.101802, 0.134737, 0.1015048, 
    0.04628988, 0.004875571, 0.1048828, 0.1574932, 0.1097925, 0.09490421, 
    0.06842887, 0.03124328, 0.01987786, -0.000280735,
  0.05720239, -5.768248e-05, 0, 0, -3.790512e-06, 0, -1.018853e-05, 0, 0, 
    -2.081152e-05, 0.02574265, 0.03107895, 0.01613719, 0.02384018, 
    0.00961335, 0.06673124, 0.02980949, 0.05360132, 0.02601204, -3.67764e-05, 
    -3.565684e-09, 0.01688184, 0.05368273, 0.1747123, 0.1552347, 0.1070949, 
    0.06698652, 0.03815929, 0.04977054,
  0.001323394, -1.719081e-05, -2.227888e-06, 0, 0, 0, 0, 0, 0, 0, 0, 
    -4.983593e-05, 0.004302337, 0.001244384, 0, 0.004106684, 0.01132216, 
    0.01810369, 0.0139764, -3.607842e-05, 0, 0, 0, -2.284858e-05, 
    0.004543275, 0.002806315, 0.04388615, 0.01289462, 0.002040659,
  -0.0001120217, 0.0005114767, -1.813522e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, -8.040287e-05, 0, 0, 0, 0, 0, 0, 0, 0.001564305, 0.007729678, 
    0.0006769554, 0.001156082,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.000160573, 6.249784e-06,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  -6.066007e-05, 0, 0, 0, -1.210607e-05, 0, 9.116585e-06, 0, 0, 0, 0, 0, 0, 
    0, 0.0009478896, 0.002056111, 0.004822288, 0.004438527, 0.0001118259, 0, 
    0, 0, 1.518125e-06, 0.001406771, 0, 0, 0, 0, -4.17549e-05,
  0.01680666, 0.03445403, 0.03790352, 0.0101993, 0.05462768, 0.06169257, 
    0.07177228, 0.03294463, 0.01181517, 0.005113327, 0.004779501, 
    0.007231446, -0.0004962074, 0.0564349, 0.08507208, 0.1327171, 0.1087297, 
    0.08986861, 0.0565464, 0.01079136, -2.380585e-06, -1.706349e-06, 
    0.004911171, 0.002292603, 0.03267447, 0.02029887, 0.02060586, 0.02838646, 
    0.01247955,
  0.1066999, 0.08115725, 0.09401473, 0.1515864, 0.2043405, 0.1918518, 
    0.1670371, 0.1586132, 0.1118973, 0.08337618, 0.07473359, 0.146044, 
    0.2086217, 0.1173581, 0.09095546, 0.1152073, 0.1157502, 0.08033755, 
    0.06906111, 0.07760869, 0.1240091, 0.2180419, 0.1863351, 0.06243093, 
    0.08373415, 0.1625561, 0.1128383, 0.1802007, 0.1767452,
  0.07635348, 0.03261979, 0.02457419, 0.06111467, 0.06155438, 0.1685036, 
    0.0852666, 0.135362, 0.01436353, 0.0199806, 0.03224147, 0.1042158, 
    0.08042991, 0.03540914, 0.1626654, 0.2795061, 0.08544241, 0.1519914, 
    0.1665563, 0.2038407, 0.1068482, 0.04364685, 0.01065664, 0.02579272, 
    0.09371883, 0.1705453, 0.1420158, 0.1815487, 0.09838901,
  4.01628e-05, 2.07516e-05, 0.1283423, 0.03976878, 0.06698482, 0.2259222, 
    0.1155269, 0.0421316, 0.001783492, 2.449783e-05, 0.0708396, 0.04479132, 
    0.01042031, 0.0131236, 0.2199667, 0.08279412, 0.1560122, 0.2206097, 
    0.1610655, 0.06262285, 0.0456115, 0.001391388, 4.94598e-07, 0.0009169796, 
    0.06937587, 0.1469259, 0.1213758, 0.0985148, 0.0004479175,
  1.05981e-05, 0.09518629, 0.1658558, 0.01325681, 0.1954532, 0.01528398, 
    0.00327671, 0.002225328, 4.335332e-06, 0.03540318, 0.163171, 0.09430461, 
    0.004771193, 0.1126167, 0.1830843, 0.1257268, 0.2049196, 0.07423872, 
    0.05036972, 0.02004352, 0.0131968, 0.001228898, 5.592743e-07, 
    -0.0003865111, 0.1542339, 0.1938383, 0.169019, 0.004046691, 2.074721e-05,
  0.0008537948, 0.02853084, 0.4515173, 0.1107797, 0.07670132, 0.01101869, 
    0.02489263, 0.002076236, 0.005305012, 0.03564834, 0.02836872, 0.1557847, 
    0.09583665, 0.2083512, 0.3462925, 0.1312876, 0.03111365, 0.009846192, 
    0.01149611, 0.01216809, 0.02096425, 1.063565e-07, 0.006241973, 0.3055434, 
    0.3544346, 0.2571977, 0.0920933, 0.005309338, 6.347816e-09,
  1.034765e-05, 0.01266243, 0.01757671, 0.03548796, 0.1548868, 0.1881122, 
    0.07701931, 0.07694755, 0.2376631, 0.1719919, 0.03560235, 0.05210271, 
    0.04903447, 0.1907344, 0.09754297, 0.009396399, 0.01685241, 0.02503382, 
    0.005490249, 0.004806027, 0.02013077, -5.163096e-08, -5.26235e-06, 
    0.02380656, 0.09728595, 0.2231222, 0.09260286, 0.0103739, 2.871573e-07,
  2.138473e-06, 1.04299e-06, 7.014191e-06, 7.766701e-05, 0.02195939, 
    0.004916307, -9.201899e-05, -4.180312e-05, 0.002504596, 0.02492133, 
    0.1550581, 0.04960554, 0.04565882, 0.01740421, -0.0002513368, 
    0.0001142794, 0.03537127, 0.121473, 0.1496346, 0.0883994, 0.07836399, 
    0.01280398, 0.004182823, 0.00039714, 3.752933e-05, 6.095652e-05, 
    1.173498e-05, 0.04120727, 0.03983464,
  0.09213194, 0.00598942, -6.461264e-06, -4.962775e-08, 1.67687e-06, 
    1.450698e-05, 4.82545e-06, -1.970482e-08, 0, 0.0004619118, 0.02619259, 
    0.02852438, 0.02195946, 0.00444682, 0.0234196, 0.001274426, 0.03262525, 
    0.09814414, 0.1435241, 0.06729908, 0.09336005, 0.01264498, 0.002033933, 
    0.000464007, 1.766771e-07, -1.58102e-05, 7.108646e-05, 0.02137101, 
    0.1805522,
  0.06067418, 0.02931917, 0.005579399, 2.472945e-08, 0.001347746, 0.02062527, 
    0.02045108, 0, 6.33292e-11, 0.08745504, 0.02703683, 0.04945077, 
    0.03960659, 0.06956736, 0.1231276, 0.167254, 0.1572155, 0.1821744, 
    0.1683057, 0.0402303, 0.01030543, 0.09873591, 0.1848206, 0.1079742, 
    0.09215861, 0.07225905, 0.1142818, 0.1132078, 0.02161572,
  0.1247002, 0.04019128, 0.0001276426, -9.044555e-08, -5.692055e-06, 
    -8.050765e-06, 3.802478e-05, 0, 0, -5.593851e-05, 0.04641066, 0.03875364, 
    0.03319914, 0.03592613, 0.03521062, 0.1427472, 0.1239227, 0.2854185, 
    0.1365103, 0.02844188, 0.0010958, 0.02259894, 0.1300496, 0.2335357, 
    0.235731, 0.2013026, 0.1256643, 0.06123124, 0.09412551,
  0.01471883, 0.001896786, 7.756909e-05, -3.590835e-05, 0, 0, 0, 0, 0, 0, 0, 
    -0.000121957, 0.008816889, 0.007999831, -1.207463e-05, 0.01167476, 
    0.02259414, 0.06908377, 0.08606727, 0.01080533, -2.643624e-05, 0, 
    -3.579837e-05, -0.0001870282, 0.01057035, 0.0140662, 0.07478786, 
    0.02158742, 0.02209738,
  0.001897691, 0.00418438, -3.023988e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, -1.731798e-05, 0.006362507, 0.0005695362, -3.142139e-05, 0, 0, 0, 0, 
    0, 0.005336212, 0.03056801, 0.01459135, 0.008279053,
  -5.616624e-05, 3.899467e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, -5.624735e-06, 0.001188783, 0.002753901,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0.01555033, 0.02404838, 0.02965324, 0.004099261, -4.412046e-05, 
    -0.0002899425, 0.003246516, -4.068814e-12, 0, 0, 0, 0, -8.776748e-06, 
    -1.477644e-05, 0.02239008, 0.05299681, 0.06547394, 0.03034887, 
    0.01546975, 0.007989069, -0.000411365, 0.006680305, 0.01531428, 
    0.01363022, 0.01774513, 0.01870269, 0.01171248, 0.005562576, 0.01774726,
  0.04600802, 0.08219954, 0.05545896, 0.07752567, 0.09482422, 0.09290355, 
    0.1475245, 0.1165565, 0.07114347, 0.04528359, 0.03926484, 0.03319157, 
    0.04672141, 0.1791539, 0.1518335, 0.1709465, 0.1543812, 0.1324272, 
    0.09392995, 0.0529171, 0.02446775, 0.009204728, 0.02353765, 0.0341243, 
    0.09742646, 0.08749076, 0.1003333, 0.06835444, 0.02598243,
  0.1486861, 0.1597006, 0.1499114, 0.1985497, 0.2079303, 0.1679458, 
    0.1532858, 0.1598918, 0.1791894, 0.14958, 0.1214748, 0.2181926, 
    0.1960379, 0.1178222, 0.08537458, 0.1188347, 0.113316, 0.1056974, 
    0.09586543, 0.1262621, 0.1476049, 0.2425208, 0.2034069, 0.1018795, 
    0.1158815, 0.1872849, 0.1431382, 0.1897069, 0.1848106,
  0.06523326, 0.029499, 0.02726303, 0.05902106, 0.06031405, 0.1538314, 
    0.09172776, 0.1370409, 0.01374, 0.02851216, 0.03218842, 0.09787297, 
    0.07958575, 0.02655502, 0.1494067, 0.233526, 0.08295996, 0.1345931, 
    0.1536512, 0.1939455, 0.09968874, 0.04006177, 0.004867172, 0.02728039, 
    0.09874687, 0.1458678, 0.1173693, 0.1634356, 0.08798472,
  4.255067e-07, 0.0001538389, 0.1232997, 0.04093439, 0.05301159, 0.2443116, 
    0.1149533, 0.0217536, 0.0002559886, -2.879867e-05, 0.06260308, 
    0.04117689, 0.01220227, 0.01798372, 0.1859888, 0.06244907, 0.143317, 
    0.2353126, 0.1640306, 0.05029624, 0.03853849, 0.0005588168, 6.430431e-07, 
    0.0008082928, 0.04587263, 0.1350909, 0.1182581, 0.1024333, 6.933921e-05,
  0.0002957623, 0.08388956, 0.1267775, 0.01061409, 0.1956417, 0.01241574, 
    0.002033674, 0.0003683573, 3.33959e-06, 0.02925352, 0.1748933, 
    0.06877875, 0.00428762, 0.1188204, 0.2017898, 0.1291154, 0.2215088, 
    0.05732141, 0.02698877, 0.01667933, 0.005342765, 0.01292401, 
    -3.588215e-08, -0.00021523, 0.1170619, 0.2132078, 0.163781, 0.0202764, 
    0.001748006,
  -9.131622e-06, 0.02007688, 0.4011906, 0.09897378, 0.06275578, 0.009538211, 
    0.0175262, 0.001521969, 0.003958859, 0.03335599, 0.02199562, 0.1427881, 
    0.08186336, 0.1665914, 0.3184074, 0.1329531, 0.03210821, 0.005357017, 
    0.01079389, 0.01177076, 0.0003299173, 7.258834e-08, 0.004812771, 
    0.2256369, 0.3144317, 0.2405261, 0.05950385, 0.0002550604, 2.695408e-09,
  2.171552e-06, 0.004699802, 0.005011504, 0.02413881, 0.1305831, 0.160332, 
    0.07285772, 0.06962144, 0.1999163, 0.1271023, 0.02865838, 0.04585877, 
    0.04300323, 0.1627402, 0.10542, 0.0118044, 0.02160703, 0.01425469, 
    0.006157451, 0.01148248, 0.02596088, 8.286226e-08, 6.00558e-06, 
    0.01312137, 0.08549444, 0.2328676, 0.08031195, 0.007499818, 1.134209e-07,
  5.870236e-07, 3.547e-09, 1.119598e-05, 0.0001789605, 0.02108822, 
    0.003345253, -1.282332e-05, 8.790957e-05, 0.001913635, 0.02524491, 
    0.1595457, 0.04523633, 0.04975853, 0.0161996, 0.0001284515, 8.086929e-05, 
    0.04553862, 0.1224619, 0.1275, 0.0891583, 0.07152745, 0.001346111, 
    0.003150229, 0.002899754, 0.000587462, -2.886274e-05, 1.508902e-05, 
    0.07226094, 0.01320572,
  0.1061496, 0.003476158, -2.328376e-06, -2.90008e-08, 1.920538e-06, 
    3.143752e-05, -9.542346e-06, -7.870873e-09, 0, 0.0002923773, 0.03143759, 
    0.02168578, 0.01134566, 0.0106848, 0.03531083, 0.00119257, 0.02680214, 
    0.1040369, 0.1429018, 0.06942695, 0.07842403, 0.01087415, 0.001871805, 
    0.0006819198, 6.411689e-06, 1.355322e-05, 0.0007807264, 0.02312487, 
    0.160174,
  0.06601619, 0.0296435, 0.003633546, 0.001831243, 0.0005529858, 0.03728916, 
    0.01537928, 0, -1.464852e-05, 0.1182631, 0.04090553, 0.05175488, 
    0.06728511, 0.08974252, 0.17192, 0.1767414, 0.1278215, 0.1901285, 
    0.109667, 0.02365066, 0.02165631, 0.08562405, 0.174963, 0.07300939, 
    0.05020631, 0.05311444, 0.1036767, 0.1409098, 0.07820846,
  0.1996221, 0.05827354, 0.03414123, 0.001888991, -7.098206e-05, 0.001642965, 
    0.0005283896, -3.162386e-05, 0.004364016, -2.105582e-05, 0.05913711, 
    0.05432453, 0.06358834, 0.05145734, 0.0662527, 0.2110183, 0.213003, 
    0.3040609, 0.1441434, 0.05287756, 0.00343192, 0.02954847, 0.1538836, 
    0.219643, 0.2176728, 0.2283849, 0.2380589, 0.1741103, 0.2274168,
  0.04724611, 0.02878089, 0.04349723, 0.007747357, 0, 0, 0, 0, 0, 0, 0, 
    0.0004156181, 0.01505981, 0.01066579, 0.00276651, 0.02068746, 0.06483501, 
    0.1984195, 0.2752199, 0.03269872, 0.005428181, 0, -0.0001031056, 
    0.005206978, 0.02980234, 0.03319975, 0.1509399, 0.09336243, 0.04155681,
  0.03639415, 0.02042107, 0.008819076, -5.254616e-05, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, -0.0002730699, 0.03670469, 0.007372799, 0.004528957, 
    -0.0001951414, 0, 0, 0, -2.358305e-06, 0.01066346, 0.07432985, 0.0568378, 
    0.03855593,
  0.01033318, 0.00779293, 0.001462772, -1.821531e-05, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, -1.523921e-05, 0.004879064, 0, 0, 0, 0, 0, 0, 0, 
    3.280762e-05, 0.006422426, 0.01039845,
  -4.292203e-07, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, -3.656517e-07,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0.0007709427, -0.000404293, 
    0.004011254, -9.638876e-06, 0, 0, 0, 0, 0.0002679545, -2.343636e-05, 0, 
    0, 0, 0,
  0.04345381, 0.06162491, 0.07234029, 0.04557911, 0.001738665, 0.003861066, 
    0.02347965, -4.621953e-06, 0, 0, 0, 0, -4.399728e-05, 0.05528932, 
    0.1067671, 0.126842, 0.1145516, 0.07007743, 0.02961183, 0.04607888, 
    0.07252816, 0.04257468, 0.03162295, 0.02196078, 0.01833544, 0.0273409, 
    0.0386391, 0.08869427, 0.02708006,
  0.08961838, 0.100546, 0.07088996, 0.1532024, 0.1548837, 0.1345136, 
    0.2029137, 0.1620913, 0.118133, 0.08665629, 0.1097511, 0.1119624, 
    0.1793942, 0.2645797, 0.1725459, 0.1741869, 0.1712596, 0.1629472, 
    0.1144061, 0.082994, 0.07765112, 0.06567533, 0.1208891, 0.1164625, 
    0.2143861, 0.1786916, 0.2151668, 0.1388064, 0.09173927,
  0.1478946, 0.1903127, 0.1606809, 0.1832199, 0.1996576, 0.154906, 0.1354761, 
    0.1456115, 0.1997949, 0.1998589, 0.157666, 0.2077453, 0.182889, 
    0.1212618, 0.08317351, 0.1332174, 0.1087544, 0.1164289, 0.1165555, 
    0.1364974, 0.1543635, 0.2365519, 0.2043362, 0.09909193, 0.1222165, 
    0.1836129, 0.1487159, 0.1713561, 0.1688329,
  0.0560069, 0.03154828, 0.03122145, 0.06248756, 0.052758, 0.1473393, 
    0.09445556, 0.1143665, 0.01921817, 0.01766434, 0.03870953, 0.1055037, 
    0.07336579, 0.02233598, 0.1478391, 0.2155387, 0.06911335, 0.1199703, 
    0.1364547, 0.1957458, 0.09841897, 0.04618183, 0.004005723, 0.01701382, 
    0.08329127, 0.1266459, 0.1018525, 0.137633, 0.07593728,
  1.205066e-06, 1.176173e-06, 0.131981, 0.02971901, 0.03144473, 0.2558453, 
    0.1048332, 0.007709116, 1.19566e-05, -9.807522e-06, 0.05997176, 
    0.02530173, 0.009051558, 0.02196132, 0.1863487, 0.02842388, 0.1426806, 
    0.2210848, 0.1506518, 0.04214432, 0.03181447, 0.0008925023, 7.257697e-08, 
    0.0001261295, 0.02704491, 0.1016194, 0.08427242, 0.1007492, 0.000165257,
  0.0004524596, 0.07508831, 0.09104077, 0.0089108, 0.1889154, 0.009348617, 
    0.001520481, 0.0001256437, 1.501605e-06, 0.02354969, 0.1576514, 
    0.04900719, 0.00212662, 0.1145843, 0.1918243, 0.1255372, 0.2128098, 
    0.03905614, 0.01442571, 0.01046275, 0.002767136, 0.005822148, 
    -4.455257e-08, 0.0006857964, 0.08292323, 0.2177918, 0.1490912, 
    0.02795821, 0.0008134953,
  1.775309e-06, 0.01526202, 0.3574424, 0.08658349, 0.04564152, 0.008479129, 
    0.0135164, 0.001471992, 0.003028359, 0.0234024, 0.01633018, 0.1123998, 
    0.06929256, 0.1237962, 0.2963163, 0.1311665, 0.03113968, 0.004749744, 
    0.006905198, 0.0121332, 7.227803e-06, 6.732775e-09, 0.005526646, 
    0.1567927, 0.2893984, 0.2226238, 0.03865134, 8.813858e-05, -7.161349e-09,
  1.258932e-06, 0.00309004, 0.004030975, 0.017924, 0.1503536, 0.1222505, 
    0.06373766, 0.06091382, 0.1578867, 0.0881082, 0.02300816, 0.02502279, 
    0.02911301, 0.1180765, 0.110747, 0.01021819, 0.01407921, 0.002569449, 
    0.005162263, 0.02109312, 0.02644219, -2.97257e-07, -4.131629e-06, 
    0.01105428, 0.0707649, 0.2582468, 0.05011058, 0.006406656, 1.340327e-08,
  1.55236e-07, -7.871323e-09, 8.869541e-06, 0.0005258448, 0.02760125, 
    0.004959425, 2.642468e-07, 5.295521e-05, 0.001896416, 0.02648947, 
    0.1676282, 0.04015353, 0.06259201, 0.01378258, 0.00073507, 0.0001038992, 
    0.06624557, 0.1076069, 0.12828, 0.1034794, 0.0707057, 0.002358607, 
    0.002025354, 0.001311203, 0.00225789, -2.556523e-06, 0.003002902, 
    0.1517233, 0.003211066,
  0.06452819, -1.676238e-05, -9.033341e-10, -7.946635e-09, 3.116172e-06, 
    0.002461898, -0.0001376651, -4.086038e-09, 0, 0.000174053, 0.04364478, 
    0.05176155, 0.01572176, 0.03528977, 0.02750075, 0.001240095, 0.02377201, 
    0.1145975, 0.1062781, 0.05891109, 0.07099994, 0.009710435, 0.001288607, 
    0.001113003, -2.988121e-06, -8.039369e-06, 9.649486e-05, 0.03121711, 
    0.1104045,
  0.06426088, 0.01858867, 0.0008501649, 0.00256486, 0.003667203, 0.03818959, 
    0.006637567, -1.206103e-09, 0.0008039675, 0.1384694, 0.04808335, 
    0.08528808, 0.07654508, 0.1013416, 0.182505, 0.1828995, 0.1233674, 
    0.1272249, 0.06424086, 0.006730254, 0.02040064, 0.07737403, 0.1365904, 
    0.05819497, 0.03819337, 0.04094982, 0.1003376, 0.0943253, 0.07690565,
  0.2382689, 0.07934432, 0.06136173, 0.01770016, 0.04638842, 0.03983207, 
    0.004525472, 0.04868015, 0.01201655, 0.01509813, 0.09306242, 0.1049146, 
    0.07847041, 0.09580136, 0.1124077, 0.2305152, 0.2290676, 0.271174, 
    0.09550924, 0.05196607, 0.007132059, 0.08097788, 0.1849358, 0.2158828, 
    0.236599, 0.2285773, 0.2310756, 0.1718737, 0.2180974,
  0.1657069, 0.09077744, 0.06822588, 0.04086389, 0.04884909, 0.00626165, 
    0.0001551991, 0, 0, 0, 0.009476209, 0.005950686, 0.02125193, 0.01220826, 
    0.01494378, 0.07668377, 0.1672356, 0.2460856, 0.3058828, 0.1459802, 
    0.04697851, 0.0005119853, -0.0004295562, 0.01580117, 0.03823441, 
    0.07910507, 0.1963312, 0.1205141, 0.08524975,
  0.1081074, 0.07378703, 0.04306041, 0.05026858, 0.007405974, 0.00539198, 
    -0.0001795104, 0, 0, 0, 0, 0, 0, 0, 0, 0.01286152, 0.03770316, 
    0.08603432, 0.03206836, 0.02654929, 0.01701104, -7.059468e-05, 0, 0, 
    4.952549e-05, 0.03940202, 0.1372058, 0.1976188, 0.114308,
  0.04639738, 0.04932653, 0.01177218, 0.009612613, -1.619323e-05, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.004064683, 0.01972334, 0.02572945, 0.02461868, 
    0.008283628, -7.443695e-08, 0, 0, 0, 1.490941e-05, -7.336414e-06, 
    0.03880762, 0.04806827,
  -0.0002164402, 0.0003332661, -2.759265e-07, -1.119046e-05, -4.56315e-06, 0, 
    0, 0, 0, 0, 0, 0, 2.278913e-06, 3.790778e-06, 1.189873e-08, 3.550772e-07, 
    -1.09704e-07, 9.761089e-07, 1.539481e-05, -8.204464e-09, 0, 0, 0, 0, 0, 
    0, 0, -7.316887e-05, -0.0002175627,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8.71173e-06, -0.0001683973, 
    0.01847435, 0.02515663, 0.01334775, 0.0008309372, -2.848234e-05, 0, 0, 
    0.00326515, 0.01130536, 0.01827985, 0.04197068, 0.02546823, 
    -0.0003522852, 0,
  0.1115076, 0.1588459, 0.2085181, 0.1178116, 0.002814982, 0.01543981, 
    0.03904865, -0.0004372266, -3.103436e-09, 0, -9.853776e-06, 0, 
    -0.004996756, 0.1795561, 0.1881783, 0.1797806, 0.179923, 0.1170079, 
    0.1371786, 0.1908164, 0.09087815, 0.05857716, 0.1684039, 0.1282731, 
    0.06598745, 0.04365486, 0.05466474, 0.2057892, 0.1134304,
  0.1758899, 0.1955946, 0.1573535, 0.2045205, 0.1923635, 0.1658807, 
    0.2165544, 0.2144333, 0.1588533, 0.1611147, 0.1875286, 0.2218411, 
    0.2296699, 0.2698574, 0.163365, 0.1619613, 0.1874563, 0.2143709, 
    0.1569607, 0.1655975, 0.1548988, 0.1612625, 0.1994645, 0.2076959, 
    0.2724633, 0.21975, 0.272804, 0.1754872, 0.1535726,
  0.1600048, 0.1769035, 0.1613336, 0.1835586, 0.1869073, 0.1429245, 
    0.1145681, 0.136488, 0.1859692, 0.2007647, 0.1884448, 0.1949519, 
    0.1617877, 0.124396, 0.07716238, 0.1319204, 0.09925539, 0.1209189, 
    0.1105911, 0.117075, 0.1564513, 0.223795, 0.2076833, 0.1029015, 
    0.09249634, 0.1813465, 0.132595, 0.1621855, 0.1578896,
  0.05253305, 0.02178534, 0.03702202, 0.06951141, 0.04190619, 0.1407257, 
    0.09401293, 0.108999, 0.01061629, 0.01015992, 0.03149386, 0.07948443, 
    0.07082133, 0.01551419, 0.1449192, 0.1838154, 0.04779239, 0.09876287, 
    0.1494559, 0.1946143, 0.1010708, 0.04148841, 0.005018292, 0.01165226, 
    0.06293438, 0.1130529, 0.1022727, 0.1272896, 0.07716887,
  6.692161e-07, 1.94733e-06, 0.1265371, 0.02864153, 0.02095174, 0.2401073, 
    0.0891756, 0.01026935, 4.60795e-06, -9.871989e-06, 0.0584062, 0.02007029, 
    0.005463346, 0.02308674, 0.2122831, 0.01653556, 0.1384427, 0.2063632, 
    0.1239539, 0.04438593, 0.009598438, 0.0005101761, 4.14931e-08, 
    -6.7521e-05, 0.01479484, 0.0811403, 0.06102777, 0.1052625, 0.0003272081,
  -1.327715e-05, 0.06588051, 0.06513292, 0.004400061, 0.2035852, 0.008887449, 
    0.0009940044, 3.330597e-05, 1.015127e-06, 0.01391854, 0.1457979, 
    0.03522761, 0.001677201, 0.09727885, 0.1787455, 0.1199585, 0.1855631, 
    0.03015373, 0.00851125, 0.007833818, 0.0006876678, 0.0001923492, 
    -1.542057e-08, 0.003077792, 0.06243958, 0.2405775, 0.09441447, 
    0.004402513, -1.621395e-05,
  2.221256e-05, 0.01909101, 0.2973716, 0.08064941, 0.03156951, 0.006380503, 
    0.01034934, 0.001682674, 0.002349373, 0.01291098, 0.01255285, 0.08476729, 
    0.06724686, 0.1136097, 0.2856417, 0.1152655, 0.02241088, 0.00414025, 
    0.004619803, 0.006456513, 1.871249e-06, 5.323795e-08, 0.005256872, 
    0.1151245, 0.2878351, 0.1952548, 0.01647712, 8.304819e-05, -3.558256e-07,
  1.296333e-05, 0.005631626, 0.004260588, 0.01337485, 0.1531236, 0.1101936, 
    0.0763756, 0.04848976, 0.1400561, 0.05458445, 0.01870095, 0.01393296, 
    0.0215186, 0.08627214, 0.1160304, 0.009944188, 0.02114794, 0.0005893871, 
    0.007075409, 0.03747238, 0.02214196, -1.280492e-06, 2.32318e-05, 
    0.01145364, 0.05565205, 0.2960492, 0.02228959, 0.004144148, 1.22321e-07,
  1.066078e-08, 2.419104e-08, 1.963876e-06, 0.0001992295, 0.01963032, 
    0.01360699, 1.890478e-05, -8.880575e-05, 0.001399341, 0.03138313, 
    0.1787189, 0.03573282, 0.06408138, 0.01265917, 0.01190394, 0.0004370684, 
    0.08988936, 0.09437707, 0.1281072, 0.1082722, 0.07547587, -0.0001918382, 
    0.001252845, 0.0008495812, 0.0110041, 3.110263e-08, -0.0002171797, 
    0.04214685, 0.0003552111,
  0.01710324, -9.191973e-05, 1.86319e-08, -2.71052e-09, 3.667596e-06, 
    0.00739552, -0.0001028835, -1.022849e-10, 0, 0.0002122991, 0.07227223, 
    0.07073523, 0.009316598, 0.04975472, 0.02993661, 0.000504642, 0.01506191, 
    0.1117549, 0.07816128, 0.04865075, 0.04658803, 0.005907248, 0.001229989, 
    0.0005995983, 2.59901e-06, -3.882269e-07, 0.0001586525, 0.03313967, 
    0.06343939,
  0.04632913, 0.008754423, -0.0001564074, 0.0012242, 0.008209772, 0.03658019, 
    0.006662307, -3.422126e-08, 0.004873668, 0.1637598, 0.06300512, 
    0.09919099, 0.07903568, 0.0952119, 0.1771443, 0.1793529, 0.09641597, 
    0.08404911, 0.03517338, 0.004895091, 0.01535509, 0.07318146, 0.118186, 
    0.04737746, 0.04273476, 0.03282602, 0.08579636, 0.07854344, 0.06932772,
  0.2353417, 0.08594539, 0.08354563, 0.04334568, 0.1226183, 0.119579, 
    0.01262328, 0.1124873, 0.09151961, 0.06603207, 0.1325286, 0.1246019, 
    0.09046327, 0.1450576, 0.1264931, 0.2359584, 0.2333828, 0.26177, 
    0.08278926, 0.04674425, 0.03866541, 0.1147249, 0.1764486, 0.2223559, 
    0.2531583, 0.2324845, 0.2207956, 0.1738452, 0.2170777,
  0.1511583, 0.1489515, 0.1090533, 0.08222365, 0.1692405, 0.1028513, 
    0.06749516, -2.41276e-05, -7.250142e-11, -0.0005539446, 0.02293044, 
    0.005581695, 0.02168254, 0.03240821, 0.09523757, 0.09453824, 0.2050072, 
    0.28399, 0.2922769, 0.2515882, 0.1066434, 0.05776533, 0.04308266, 
    0.02388653, 0.09637094, 0.1239486, 0.2101039, 0.1383147, 0.1040786,
  0.1838541, 0.1702045, 0.09619406, 0.08070479, 0.02975606, 0.004353271, 
    0.01212974, 0.0005776263, -1.651976e-05, 0, 0, 0, 0, 0, 0.001692521, 
    0.1338249, 0.09434242, 0.1319524, 0.07889625, 0.06057582, 0.02678593, 
    0.03003541, 0.02171368, 0, 0.003282302, 0.08051439, 0.2208003, 0.2255095, 
    0.1164124,
  0.1258257, 0.1435837, 0.05202019, 0.03393305, 0.01765537, 0.004734358, 
    -3.601797e-05, 0, 0, 0, 0, 0, -8.410969e-05, 6.175697e-05, 0.01200598, 
    0.002470271, 0.1048117, 0.08977558, 0.05573725, 0.05840494, 0.02864663, 
    -0.0002336831, -1.111019e-07, -2.686837e-07, 0.0009413795, 0.003153743, 
    -0.0003741011, 0.1033732, 0.1095078,
  0.01157044, 0.00236642, 0.0006182958, 0.001117046, 0.00166038, 
    -9.117562e-07, 0, 0, 0, 0, 0, -4.60277e-05, 0.002212325, -0.0001366838, 
    2.622603e-05, 0.00030927, 0.0007911464, 0.002893004, 0.0001231111, 
    -2.488236e-05, 9.069204e-07, -1.401834e-05, -2.321139e-05, -9.018049e-06, 
    -9.854689e-05, -2.348499e-06, -9.154344e-05, -0.002219931, 0.01889367,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.002146319, 0.06176692, 0.1476729, 
    0.2255351, 0.1692706, 0.02321781, 0.0004624558, -0.001302429, 
    -0.0006034104, 0.008364693, 0.04365582, 0.05681068, 0.1211849, 0.2142134, 
    -0.002334907, 0,
  0.1927157, 0.2518876, 0.3352248, 0.244837, 0.01693424, 0.02396732, 
    0.03714415, -0.001000021, -4.505634e-05, -0.0001486972, -9.078671e-05, 
    -0.0002612627, 0.07714675, 0.3683392, 0.2395102, 0.2231497, 0.2201371, 
    0.1782902, 0.183182, 0.183808, 0.09824079, 0.1503831, 0.3379265, 
    0.2312692, 0.2017314, 0.1084748, 0.08825025, 0.220155, 0.1205326,
  0.1927207, 0.2229331, 0.2001193, 0.2212997, 0.2214083, 0.1915226, 
    0.2295707, 0.2292526, 0.2160346, 0.2261291, 0.2303904, 0.2970316, 
    0.2755485, 0.2679825, 0.1654737, 0.1652631, 0.1901936, 0.2576364, 
    0.1770981, 0.2386758, 0.2464026, 0.2383158, 0.2457027, 0.2359024, 
    0.2815493, 0.2488146, 0.3187047, 0.191026, 0.1829863,
  0.161762, 0.1602659, 0.162011, 0.180302, 0.1644071, 0.1428584, 0.1084502, 
    0.1227722, 0.179873, 0.2077341, 0.191954, 0.2044131, 0.1294134, 
    0.1174264, 0.08180884, 0.1203992, 0.09964017, 0.1092519, 0.1053238, 
    0.114889, 0.1652805, 0.1954734, 0.218962, 0.1058741, 0.08936004, 
    0.1817577, 0.1332283, 0.1605224, 0.1686337,
  0.04304599, 0.01817378, 0.03452143, 0.08652234, 0.03106797, 0.1134066, 
    0.08764452, 0.09475245, 0.008724424, 0.006373994, 0.03583613, 0.07052103, 
    0.06157352, 0.00879131, 0.1470267, 0.1632618, 0.05232219, 0.08349956, 
    0.1247198, 0.1405941, 0.09667172, 0.04137763, 0.003289038, 0.01129887, 
    0.05572066, 0.1062511, 0.1019581, 0.118149, 0.05804716,
  5.867881e-07, 3.608131e-06, 0.1206426, 0.01939483, 0.01487321, 0.2153239, 
    0.08312106, 0.003578538, -4.112003e-07, 9.127047e-06, 0.06449441, 
    0.02234432, 0.009314636, 0.02374643, 0.2448951, 0.007951807, 0.1084089, 
    0.2056935, 0.1286362, 0.04034425, 0.007542246, 0.0002806451, 
    5.439346e-08, -0.000141687, 0.01107776, 0.09174466, 0.04877916, 
    0.06795939, 0.0002528328,
  0.0002926805, 0.0552869, 0.0456501, 0.003934176, 0.2173599, 0.007397375, 
    0.0009358443, 3.872001e-07, 3.384772e-06, 0.006638336, 0.1371725, 
    0.02742636, 0.001666174, 0.08547837, 0.1840763, 0.1113034, 0.1543445, 
    0.03069161, 0.006529888, 0.006131752, 0.000304746, 1.784464e-05, 
    -1.683307e-09, 0.004575226, 0.05632641, 0.2617256, 0.04974268, 
    0.005050303, -0.0001806495,
  1.050258e-05, 0.0342998, 0.2508439, 0.07974077, 0.02346701, 0.005722738, 
    0.009553482, 0.001655126, 0.00138966, 0.009710538, 0.009356812, 
    0.07233411, 0.07758544, 0.1209665, 0.2730787, 0.09736553, 0.01760928, 
    0.006627143, 0.003886743, 0.001208132, 1.19309e-07, 5.92573e-08, 
    0.005054665, 0.09308476, 0.3039793, 0.1978485, 0.01689168, 7.326463e-05, 
    -7.147909e-07,
  0.0001021721, 0.003751474, 0.005958163, 0.009532145, 0.1481057, 0.1043647, 
    0.1041611, 0.06110222, 0.119061, 0.03335423, 0.02709691, 0.01217934, 
    0.01394562, 0.06054469, 0.1112272, 0.01002755, 0.006502162, 0.0001337559, 
    0.01578218, 0.03704184, 0.01645059, 9.628895e-05, 0.001211131, 
    0.01013307, 0.06046567, 0.325371, 0.01405854, 0.003468982, 1.823275e-06,
  6.204109e-10, 5.929339e-08, 1.505823e-06, 0.0008372575, 0.02456167, 
    0.005673986, 5.368749e-05, -0.0001930211, 0.0008321677, 0.03204664, 
    0.1865743, 0.0418171, 0.07761564, 0.01676219, 0.01681511, 0.0005219614, 
    0.09970339, 0.08107913, 0.1309439, 0.1006958, 0.07855552, 3.223546e-05, 
    0.0007197857, 0.0009916257, 0.02782022, 2.675098e-06, -5.768135e-05, 
    0.01169127, 0.004008957,
  0.001304986, -7.645728e-05, 2.291514e-07, -4.458821e-09, 2.740619e-06, 
    0.002229987, 0.0002145764, -5.588431e-10, 1.071389e-10, 0.0008042088, 
    0.09258559, 0.09848654, 0.0002899667, 0.04477062, 0.02339672, 
    0.0003276479, 0.01707873, 0.09078581, 0.04041161, 0.03783737, 0.03421248, 
    0.005630842, 0.001676973, 0.0005607887, 1.512282e-06, 5.015882e-08, 
    0.0005434153, 0.02809173, 0.03418764,
  0.03979073, 0.002962428, -5.746727e-05, 0.005463439, 0.01069993, 
    0.03784704, 0.005696916, -2.210387e-05, 0.02151687, 0.2013492, 
    0.09264528, 0.1013745, 0.07777695, 0.09950982, 0.1362577, 0.1412391, 
    0.05990481, 0.07972096, 0.03157217, 0.001773341, 0.01124687, 0.06611077, 
    0.1262538, 0.05422382, 0.048032, 0.03312805, 0.07164805, 0.08733279, 
    0.0680054,
  0.2125691, 0.08422383, 0.07276948, 0.08996145, 0.130782, 0.158575, 
    0.03880907, 0.1679015, 0.1007419, 0.09971675, 0.1599832, 0.1257051, 
    0.1192254, 0.1433376, 0.1367226, 0.2426892, 0.2356979, 0.2650375, 
    0.09869896, 0.04935005, 0.06056646, 0.138785, 0.1594944, 0.2494507, 
    0.2347024, 0.2377962, 0.2002132, 0.1410924, 0.189895,
  0.1474796, 0.151976, 0.1028993, 0.09557641, 0.1950368, 0.143384, 0.1514778, 
    -0.0003440939, -7.514458e-05, 0.03627335, 0.04857863, 0.01430888, 
    0.05475651, 0.09258943, 0.1506699, 0.1204538, 0.2499723, 0.3241282, 
    0.2825823, 0.2752666, 0.1159009, 0.09115234, 0.1162141, 0.06037499, 
    0.1786461, 0.1739697, 0.2444032, 0.1663739, 0.1315069,
  0.2057357, 0.2193197, 0.1374777, 0.1338438, 0.09073485, 0.09366482, 
    0.1047544, 0.189964, 0.07555076, 0.01496008, 0.00248736, -1.993382e-05, 
    -1.454002e-05, -2.080684e-07, 0.04604405, 0.184273, 0.1302565, 0.212066, 
    0.1020693, 0.1090106, 0.04187388, 0.05224978, 0.03605193, 0.0001238503, 
    0.02022404, 0.1782778, 0.2747814, 0.2476619, 0.2004123,
  0.2239978, 0.1688028, 0.07828286, 0.06013944, 0.04225918, 0.04368911, 
    0.02969258, 0.03692275, 0.004557458, -1.449394e-06, 0, 0.001102181, 
    5.403285e-05, 0.004192195, 0.03814205, 0.06223897, 0.127835, 0.1029792, 
    0.06757307, 0.09915193, 0.0368574, 0.006541211, 3.635757e-05, 
    -0.0001456663, 0.03745926, 0.01662902, 0.01104532, 0.1736635, 0.1767191,
  0.07868433, 0.07828769, 0.06723275, 0.04269003, 0.03059296, 0.002760263, 
    0.00448035, 0.005393189, 0.001041376, 0.0001853726, -8.178193e-07, 
    -9.696427e-05, 0.005957793, -0.0006404522, 0.002669709, 0.01439458, 
    0.008903475, 0.04074172, 0.05273212, 0.03084435, 0.0197079, 0.01439339, 
    9.576733e-05, -0.0007858012, 0.001948949, -4.947616e-05, -0.003246387, 
    0.03481651, 0.07884162,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5.914359e-05, 0.06266651, 0.1323264, 
    0.2086042, 0.2355026, 0.2173484, 0.08631561, 0.02849887, 0.02162538, 
    0.009923371, 0.08528029, 0.05388136, 0.1057089, 0.1491368, 0.2544907, 
    0.2169343, 0.001599893,
  0.2310548, 0.3187627, 0.3725114, 0.2822961, 0.07524318, 0.07735145, 
    0.03131942, -0.002178882, -6.826951e-05, -0.0005773856, -0.0001722954, 
    -0.003036397, 0.2355133, 0.3655285, 0.2579941, 0.2272474, 0.2264978, 
    0.2011872, 0.2516777, 0.1722454, 0.09101167, 0.1587378, 0.3122152, 
    0.2542189, 0.2332537, 0.1319757, 0.1032406, 0.2219705, 0.1781671,
  0.2089287, 0.238849, 0.1977519, 0.2336925, 0.260676, 0.212925, 0.2258928, 
    0.2360681, 0.2320113, 0.254038, 0.2485628, 0.319391, 0.295441, 0.2715492, 
    0.167572, 0.1556842, 0.1887771, 0.2521574, 0.1926068, 0.257214, 0.259279, 
    0.2428542, 0.2378775, 0.2267042, 0.2652779, 0.2380597, 0.308053, 
    0.2003294, 0.2228415,
  0.1650968, 0.1514284, 0.1316895, 0.1845218, 0.1523583, 0.1270886, 
    0.07930908, 0.1144012, 0.1812879, 0.2247243, 0.1843087, 0.2127877, 
    0.1274295, 0.1156295, 0.09616277, 0.1141205, 0.09743822, 0.1138184, 
    0.1041221, 0.1130738, 0.1538487, 0.1977502, 0.1940846, 0.08786222, 
    0.09073278, 0.1775021, 0.1310909, 0.1609753, 0.1761123,
  0.04101915, 0.01388416, 0.02819969, 0.09602547, 0.02525163, 0.1032516, 
    0.0864851, 0.07746759, 0.0245982, 0.005625384, 0.04681804, 0.08009378, 
    0.05657949, 0.006259861, 0.145689, 0.1485928, 0.05019005, 0.07415529, 
    0.1187938, 0.1302651, 0.1007437, 0.05359313, 0.00208292, 0.01002949, 
    0.04449826, 0.1095634, 0.08081648, 0.1171726, 0.04914704,
  3.627849e-07, 6.24267e-06, 0.1228007, 0.01558951, 0.01503862, 0.1871004, 
    0.07031099, 0.004617148, 3.381408e-08, 2.285002e-05, 0.09728406, 
    0.02118754, 0.01028542, 0.03398255, 0.2328917, 0.005088445, 0.09772616, 
    0.1791871, 0.1039078, 0.03927405, 0.005604402, 0.0002810635, 
    -3.614804e-09, -6.218738e-05, 0.01186009, 0.08232431, 0.03693533, 
    0.04514058, -4.208225e-05,
  0.000147593, 0.05284451, 0.03660718, 0.004639216, 0.2107295, 0.007388729, 
    0.001163805, 7.364209e-07, 1.443407e-05, 0.007033479, 0.1378751, 
    0.02705212, 0.001898333, 0.0859113, 0.1840064, 0.103576, 0.1337895, 
    0.03743771, 0.005581131, 0.005381744, 5.934477e-07, 5.02368e-06, 
    2.289486e-09, 0.002941869, 0.06043156, 0.2916342, 0.01825556, 
    0.001052897, -7.550842e-05,
  0.001537904, 0.04010386, 0.2246977, 0.07581749, 0.02024442, 0.004598813, 
    0.009480591, 0.00142317, 0.001118226, 0.00864305, 0.01337586, 0.06515882, 
    0.1008073, 0.1156228, 0.2655844, 0.08263569, 0.0196876, 0.01103423, 
    0.003344867, 1.646874e-05, 7.60357e-09, 1.749908e-07, 0.004456066, 
    0.1100727, 0.3209656, 0.2061152, 0.01498903, 0.0001871696, 4.519729e-05,
  0.03623582, 0.005844483, 0.003953133, 0.00920083, 0.1365043, 0.08803514, 
    0.1130252, 0.09320375, 0.09268676, 0.02775834, 0.03902185, 0.01170203, 
    0.01055245, 0.04781219, 0.09458145, 0.00522722, 0.0008725971, 
    5.308562e-07, 0.03516365, 0.0343279, 0.01477623, 0.01485816, 0.02872494, 
    0.007963321, 0.04261173, 0.3345284, 0.01076894, 0.003948001, 0.00051655,
  2.112951e-08, 6.426819e-07, 1.595367e-06, 0.0005564994, 0.02777666, 
    0.001901813, 6.162214e-05, -0.0002626259, 0.0008375917, 0.03637366, 
    0.1983187, 0.05751568, 0.0748909, 0.02575251, 0.01524949, 0.008094823, 
    0.1061306, 0.08127016, 0.114408, 0.1125579, 0.07946527, 0.001089166, 
    0.0008170492, 0.001181829, 0.02362043, 0.0001783606, -0.0001569674, 
    0.008584859, 0.001794543,
  2.873598e-05, 5.595e-08, 2.151007e-07, -1.148782e-08, 1.683872e-06, 
    0.0003232248, 0.00132495, -1.067154e-08, 2.573013e-09, 0.006200377, 
    0.1167945, 0.09135562, 0.0004455947, 0.04048477, 0.01763877, 5.26599e-05, 
    0.02072213, 0.07609125, 0.04161566, 0.03022921, 0.02246479, 0.006517884, 
    0.002779227, 0.0003234555, -7.002251e-07, 2.374447e-08, 0.0005094177, 
    0.03459793, 0.00598719,
  0.02335103, 0.0005516573, -0.0003897473, 0.0101238, 0.01443424, 0.04070373, 
    0.003941095, -0.0002087338, 0.05102782, 0.2487511, 0.1205037, 0.070028, 
    0.06333192, 0.08215971, 0.1299324, 0.1108242, 0.04099144, 0.07237479, 
    0.04397083, 0.0002531419, 0.01165346, 0.0687733, 0.1228535, 0.04483401, 
    0.04671422, 0.0304872, 0.06046566, 0.09394772, 0.06013002,
  0.1880285, 0.07834245, 0.0648823, 0.1257519, 0.1275633, 0.1411261, 
    0.09308598, 0.1538678, 0.1109993, 0.09887557, 0.1579598, 0.1052755, 
    0.1152953, 0.1528517, 0.1581499, 0.2616898, 0.2199127, 0.2766912, 
    0.09515153, 0.04292107, 0.06464729, 0.1363145, 0.1680378, 0.251571, 
    0.2289056, 0.2331537, 0.1751324, 0.1302067, 0.1683377,
  0.1297007, 0.1496299, 0.1031998, 0.1045729, 0.2200999, 0.1616181, 
    0.1967975, 0.004760687, 0.0345648, 0.04232094, 0.07127629, 0.02473296, 
    0.07975346, 0.1386759, 0.2007407, 0.1693063, 0.2608937, 0.3294431, 
    0.2706833, 0.2808957, 0.1462298, 0.1384173, 0.1593393, 0.1414004, 
    0.2335667, 0.2129699, 0.2635649, 0.1945898, 0.1451624,
  0.190719, 0.2153825, 0.1508735, 0.2138306, 0.2022111, 0.126444, 0.1821817, 
    0.2486293, 0.2119423, 0.153825, 0.1498043, 0.001462632, -0.00153022, 
    0.02298034, 0.1826149, 0.2975934, 0.2191806, 0.320589, 0.1953204, 
    0.1627076, 0.08243363, 0.08264273, 0.09057996, 0.01875914, 0.1305157, 
    0.2731917, 0.3048313, 0.2788632, 0.2022721,
  0.2226462, 0.1916903, 0.09930138, 0.09489246, 0.06813325, 0.07144314, 
    0.04335628, 0.04505892, 0.02661978, 0.02411463, 0.005952199, 0.008926992, 
    0.0006415771, 0.01049059, 0.1161281, 0.1199505, 0.1840894, 0.1729496, 
    0.1178565, 0.1275318, 0.06506697, 0.009022661, 0.01042652, -0.001676382, 
    0.09377199, 0.05224832, 0.02315622, 0.2504612, 0.217118,
  0.1069303, 0.1300132, 0.1313448, 0.1057594, 0.08836047, 0.04944779, 
    0.04564784, 0.049635, 0.05052257, 0.01737889, 0.001157121, 0.006841244, 
    0.01656408, 0.0165884, 0.01450595, 0.04611859, 0.05935336, 0.06365821, 
    0.07712709, 0.09180863, 0.07273211, 0.03807135, 0.01401429, 
    -0.0004397092, 0.009202091, 0.002855461, 0.005106713, 0.06632781, 
    0.1617042,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -0.0001264613, -0.0001264613, -0.0001264613, -0.0001264613, 
    -0.0001264613, -0.0001264613, -0.0001264613, 0,
  0.004711038, -0.0001543938, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.000829988, 
    0.164201, 0.1799083, 0.2449349, 0.2011732, 0.1880823, 0.08031161, 
    0.0854435, 0.05133956, 0.05394008, 0.1439866, 0.07947135, 0.1238249, 
    0.1643423, 0.292046, 0.2577158, 0.08688121,
  0.2804509, 0.3638048, 0.3363892, 0.2689809, 0.1585415, 0.1275494, 
    0.02227163, -0.0006346811, -0.002289173, 0.03524105, 0.02077481, 
    0.007483112, 0.3536391, 0.3212926, 0.2445854, 0.2078347, 0.2244244, 
    0.2129344, 0.2776971, 0.1677949, 0.08822817, 0.1937233, 0.3305392, 
    0.2392469, 0.2545877, 0.1069194, 0.1181627, 0.2014188, 0.2063789,
  0.2276053, 0.2321277, 0.2033669, 0.2534026, 0.2849262, 0.260983, 0.2147284, 
    0.2105076, 0.233339, 0.2423462, 0.2684079, 0.3059991, 0.2978179, 
    0.2870146, 0.1824167, 0.1715907, 0.1878818, 0.239635, 0.2050742, 
    0.2802361, 0.2701956, 0.2541667, 0.256862, 0.2541465, 0.2592013, 
    0.232125, 0.3253505, 0.2163759, 0.2525174,
  0.172587, 0.1527092, 0.1323835, 0.1611441, 0.1420658, 0.1092308, 
    0.08188558, 0.1207571, 0.1768102, 0.2368493, 0.1800908, 0.1966331, 
    0.1103608, 0.1192904, 0.09655333, 0.1120597, 0.1027126, 0.1210595, 
    0.1153679, 0.1175078, 0.1676354, 0.2086957, 0.2201247, 0.07438663, 
    0.09307821, 0.1628841, 0.130782, 0.1617031, 0.1682294,
  0.03812536, 0.01280078, 0.02436801, 0.1191909, 0.02564245, 0.1018925, 
    0.06727911, 0.07005493, 0.03331699, 0.009780012, 0.04859662, 0.0692206, 
    0.05449168, 0.007704246, 0.1514814, 0.1342764, 0.06057077, 0.07358596, 
    0.09817397, 0.1197784, 0.09866371, 0.04795498, 0.0001932836, 0.009163313, 
    0.04773019, 0.09134233, 0.06525755, 0.09470536, 0.04300252,
  -3.745358e-05, 8.124714e-06, 0.1252968, 0.01556999, 0.01681632, 0.1732566, 
    0.05634356, -0.000227484, -1.055519e-08, 0.001202937, 0.1398566, 
    0.04320026, 0.02001723, 0.03980958, 0.2243256, 0.01257208, 0.08427838, 
    0.1634236, 0.1079708, 0.03851493, 0.008386726, 0.0002189013, 
    -7.411807e-08, 0.0002621466, 0.01658698, 0.08188985, 0.02890849, 
    0.03991594, 0.001324467,
  4.106989e-05, 0.06022744, 0.04135392, 0.006327129, 0.2056311, 0.007727454, 
    0.001022384, 7.188235e-06, 6.642205e-06, 0.01112404, 0.1513053, 
    0.02490794, 0.001947572, 0.09566459, 0.2023945, 0.1103395, 0.1217602, 
    0.03764446, 0.004757137, 0.004892346, 5.940421e-07, 1.357023e-06, 
    1.015949e-07, 0.002760571, 0.07047089, 0.291906, 0.008321754, 
    0.0001023665, -3.455338e-06,
  0.007206009, 0.06315593, 0.2087698, 0.09542885, 0.01879029, 0.004895476, 
    0.009077111, 0.002424039, 0.001220965, 0.01120995, 0.03184869, 
    0.06611453, 0.1390864, 0.1181583, 0.2666351, 0.07114378, 0.01825692, 
    0.01318458, 0.003020902, 3.863209e-06, -9.406521e-08, -0.0001043011, 
    0.008745617, 0.1498378, 0.3406393, 0.2071095, 0.01338354, 0.0002705014, 
    0.002970272,
  0.1385132, 0.01791116, 0.02832594, 0.009151555, 0.122186, 0.09567922, 
    0.1358449, 0.1125475, 0.0839081, 0.03117629, 0.06460301, 0.01165705, 
    0.01203136, 0.05131203, 0.08103097, 0.004719607, 7.125416e-05, 
    1.392241e-05, 0.022939, 0.02329854, 0.01546688, 0.03491634, 0.07172934, 
    0.008659597, 0.03957001, 0.3423697, 0.01297148, 0.003585667, 0.05833245,
  4.191557e-05, 6.671032e-07, 1.69771e-06, 0.001380567, 0.03513927, 
    0.000630825, 4.644051e-05, -0.0003764374, 0.00136867, 0.04565802, 
    0.2015725, 0.04694227, 0.0759196, 0.04290409, 0.01462765, 0.02086034, 
    0.1023065, 0.1167545, 0.1139481, 0.1223909, 0.08114985, 0.002333268, 
    0.002446132, 0.001267144, 0.02118962, 9.842165e-05, -1.200161e-06, 
    0.00177304, 0.0004857246,
  2.916242e-06, 5.638315e-07, 1.332649e-07, 4.478125e-09, 1.113197e-06, 
    2.270726e-05, 9.654684e-05, 7.30579e-08, -7.776474e-10, 0.008328915, 
    0.1036105, 0.06398144, 9.935433e-06, 0.03139473, 0.0246961, 0.0002182252, 
    0.03083593, 0.07170022, 0.04112295, 0.01959343, 0.01833502, 0.009480921, 
    0.006952955, 0.0005964092, -9.560782e-07, 1.024139e-07, 0.0004082668, 
    0.01722951, 0.001793357,
  0.004815117, 0.0003511836, 0.0009134933, 0.01462188, 0.02403268, 
    0.04702487, 0.006371342, 0.001078072, 0.08503432, 0.2532564, 0.1452179, 
    0.05525981, 0.04121573, 0.0685083, 0.09055502, 0.07836776, 0.03093584, 
    0.07514013, 0.05815261, -1.096201e-05, 0.0135639, 0.06236171, 0.1244123, 
    0.03993949, 0.04073381, 0.03811421, 0.05607916, 0.08354881, 0.05113247,
  0.1641379, 0.07329653, 0.06010861, 0.1162142, 0.1360018, 0.1217028, 
    0.1417483, 0.1203369, 0.1189234, 0.09289151, 0.1435123, 0.09667751, 
    0.1113115, 0.170309, 0.1728064, 0.2744038, 0.2170094, 0.2268334, 
    0.06293238, 0.03806761, 0.08952041, 0.1190466, 0.1645469, 0.2532478, 
    0.2178051, 0.2122193, 0.1520628, 0.1317416, 0.1570105,
  0.124682, 0.1286502, 0.09385305, 0.09563324, 0.2321496, 0.1869586, 
    0.2028928, 0.06213431, 0.07387533, 0.03660427, 0.06301468, 0.04382922, 
    0.09308787, 0.2085022, 0.2552221, 0.1719488, 0.2487745, 0.3217036, 
    0.2795642, 0.2972575, 0.1857672, 0.1568717, 0.2047989, 0.158842, 
    0.2450795, 0.22466, 0.2744271, 0.1691901, 0.1455272,
  0.1942455, 0.2004974, 0.160008, 0.2630401, 0.2420084, 0.2177986, 0.2663439, 
    0.3411657, 0.2849356, 0.2166989, 0.213751, 0.06505714, 0.03143141, 
    0.1338753, 0.2975155, 0.3333297, 0.2529954, 0.3545942, 0.2113925, 
    0.2325274, 0.1064597, 0.1046999, 0.1460994, 0.1159879, 0.2573817, 
    0.3361236, 0.3076138, 0.2880318, 0.1920396,
  0.2221303, 0.2407493, 0.1644443, 0.1738788, 0.1492854, 0.09383532, 
    0.07997517, 0.1282587, 0.0965135, 0.1226903, 0.06444798, 0.0537736, 
    0.02069516, 0.05590913, 0.2386952, 0.2012093, 0.2815574, 0.2441398, 
    0.1681724, 0.1174229, 0.09219226, 0.0358217, 0.05247727, -0.008836762, 
    0.1557019, 0.07410114, 0.06032186, 0.313338, 0.2199055,
  0.1225379, 0.1385228, 0.1743746, 0.1921867, 0.1705882, 0.1250309, 
    0.1241536, 0.1631929, 0.1291586, 0.03506707, 0.01386493, 0.02811663, 
    0.04585449, 0.08149602, 0.1147231, 0.1103484, 0.08444511, 0.05914323, 
    0.09153675, 0.09496143, 0.06462776, 0.04975404, 0.03763875, -0.001541426, 
    0.0437723, 0.01753547, 0.04666733, 0.1473092, 0.2079387,
  0.00256033, 0.001952785, 0.00134524, 0.0007376951, 0.0001301503, 
    -0.0004773945, -0.001084939, -9.95753e-05, 0.0002460388, 0.0005916529, 
    0.000937267, 0.001282881, 0.001628495, 0.001974109, 0.009342709, 
    0.01048441, 0.0116261, 0.0127678, 0.0139095, 0.0150512, 0.0161929, 
    0.01787229, 0.01699253, 0.01611276, 0.01523299, 0.01435322, 0.01347346, 
    0.01259369, 0.003046365,
  0.09316878, 0.003576081, -0.0002209415, 0, -2.215946e-05, -0.0001789609, 0, 
    0, 0, 0, 0, 0, 0.004053868, 0.1989242, 0.1636462, 0.1992088, 0.2028638, 
    0.1638605, 0.08952257, 0.1422506, 0.1133433, 0.110351, 0.190852, 
    0.1281686, 0.1754295, 0.1698589, 0.3059222, 0.2500209, 0.1331942,
  0.3062257, 0.3613869, 0.3178314, 0.2713535, 0.2315172, 0.1235973, 
    0.01433133, 0.02605537, 0.04151473, 0.1309507, 0.08131336, 0.1393817, 
    0.3712608, 0.3022321, 0.2520263, 0.2153568, 0.2431164, 0.2187735, 
    0.2582299, 0.1658697, 0.1126748, 0.2185729, 0.3360848, 0.2871647, 
    0.2866308, 0.1038124, 0.1743124, 0.2042325, 0.2532209,
  0.2513246, 0.2481471, 0.2591307, 0.3127532, 0.3059868, 0.2938026, 
    0.2506773, 0.2268223, 0.2571459, 0.2561987, 0.2484949, 0.3296296, 
    0.326795, 0.2821954, 0.1871692, 0.1578857, 0.2118605, 0.2540996, 
    0.2206317, 0.2992629, 0.2948588, 0.2896917, 0.2519654, 0.2816017, 
    0.2872522, 0.2354817, 0.3151875, 0.2222341, 0.2571588,
  0.165391, 0.1451961, 0.1415517, 0.1674238, 0.1521216, 0.09402429, 
    0.07666861, 0.1147399, 0.1694515, 0.1980276, 0.1898222, 0.2079468, 
    0.1226122, 0.1185339, 0.09719581, 0.1014822, 0.09871407, 0.1157614, 
    0.1053601, 0.1295741, 0.1554907, 0.1875464, 0.1739011, 0.08174948, 
    0.1007159, 0.1686525, 0.1369314, 0.159251, 0.1968033,
  0.03857296, 0.01349621, 0.01761555, 0.1215971, 0.02723386, 0.1055624, 
    0.06555983, 0.07523023, 0.02764078, 0.01248211, 0.03859654, 0.06835796, 
    0.06262789, 0.01152195, 0.1310641, 0.1263573, 0.06547008, 0.06993847, 
    0.09280417, 0.105782, 0.09745316, 0.04725487, 0.0003553378, 0.007563941, 
    0.06339481, 0.09513523, 0.06103987, 0.09580102, 0.04146517,
  0.002719603, 6.662052e-07, 0.143165, 0.01943057, 0.01933306, 0.1574498, 
    0.04664971, 0.0005895746, 5.019745e-08, 0.008753022, 0.1149996, 
    0.1075314, 0.0259188, 0.04325655, 0.2374311, 0.01626843, 0.1093083, 
    0.1431675, 0.09792701, 0.04158625, 0.02240056, 0.0002213813, 
    -1.741408e-07, 0.00127083, 0.01638508, 0.08568466, 0.02990781, 0.0287252, 
    0.003255532,
  0.0001545524, 0.07779552, 0.05961872, 0.0103068, 0.233559, 0.01241424, 
    0.001324065, 2.484025e-05, -0.0001304507, 0.02008396, 0.1711674, 
    0.03777166, 0.004309847, 0.08351423, 0.2231681, 0.1186936, 0.1227478, 
    0.04187164, 0.004742988, 0.005596053, 8.505556e-07, 3.283365e-06, 
    -7.758655e-08, 0.001535481, 0.0808642, 0.2958066, 0.003880857, 
    0.0001324665, -1.75905e-05,
  0.005929887, 0.08506972, 0.2320887, 0.1126553, 0.02305104, 0.006744418, 
    0.01471381, 0.002881872, 0.001662089, 0.01312232, 0.05138843, 0.0784733, 
    0.1843046, 0.1658728, 0.2950276, 0.07364516, 0.01526855, 0.01315817, 
    0.00422306, 8.219979e-06, -9.638445e-08, 0.003798791, 0.00872934, 
    0.2052436, 0.3757803, 0.2365194, 0.01736663, 0.0002581175, 0.03261501,
  0.2117281, 0.04284234, 0.05222443, 0.01266849, 0.1177682, 0.1080673, 
    0.1501068, 0.1343807, 0.09555002, 0.03822934, 0.08444332, 0.02009621, 
    0.01710729, 0.05761556, 0.09200865, 0.009278026, 0.0001567692, 
    4.97041e-06, 0.007707091, 0.008246017, 0.035882, 0.06450363, 0.1114103, 
    0.02313809, 0.05195397, 0.3893507, 0.02161556, 0.005231485, 0.0468107,
  0.0002351456, 1.076885e-06, -6.176554e-06, 0.01047061, 0.01816543, 
    0.0008982122, 1.577659e-05, -7.570039e-05, 0.001376707, 0.04461751, 
    0.213932, 0.05099574, 0.0885044, 0.06878623, 0.01778337, 0.0222306, 
    0.1212529, 0.1441755, 0.1337857, 0.1192869, 0.09096693, 0.003741561, 
    0.003617895, 0.001470873, 0.009637558, 9.458086e-05, -7.204051e-08, 
    0.0009713, 7.258054e-06,
  5.108393e-06, 8.857153e-07, 8.504758e-08, 8.882775e-09, -1.061261e-05, 
    8.875296e-07, 2.489769e-06, 1.175678e-06, -1.259216e-08, 0.01612199, 
    0.09836788, 0.05165521, 1.427149e-06, 0.02160528, 0.03975321, 
    0.000739574, 0.03099924, 0.06713913, 0.02174214, 0.01684074, 0.007494588, 
    0.01521624, 0.01303647, 0.001119207, -3.798956e-06, 5.822512e-08, 
    0.0007785085, 0.01194466, 1.651144e-05,
  -3.677066e-05, 1.182901e-06, 0.006511711, 0.0181377, 0.03868129, 
    0.05843943, 0.00790792, 0.003757669, 0.1196869, 0.2877118, 0.1432246, 
    0.03769165, 0.03844018, 0.05626402, 0.0578954, 0.05769851, 0.03241641, 
    0.07943632, 0.04317927, -7.458546e-05, 0.01792924, 0.06330728, 0.1213543, 
    0.03526699, 0.04339764, 0.04653792, 0.04764636, 0.08521224, 0.06104689,
  0.1326067, 0.05775487, 0.05540211, 0.1005754, 0.1332496, 0.1285227, 
    0.2097572, 0.08060723, 0.1217972, 0.08563464, 0.1273023, 0.0889896, 
    0.10811, 0.1724576, 0.1769417, 0.2703669, 0.2046906, 0.2084156, 
    0.04578471, 0.03902664, 0.1234605, 0.1329643, 0.1654541, 0.243041, 
    0.2148727, 0.1879446, 0.148479, 0.1221172, 0.1398527,
  0.1215746, 0.1135117, 0.1025607, 0.1006474, 0.2229032, 0.1982043, 
    0.2140313, 0.1168772, 0.08417405, 0.03505829, 0.05073278, 0.03879109, 
    0.0878299, 0.2756686, 0.257809, 0.1524671, 0.2168438, 0.2822856, 
    0.274774, 0.3061644, 0.2280482, 0.1503378, 0.2102901, 0.1678493, 
    0.2566506, 0.2432526, 0.2759807, 0.1633243, 0.1304821,
  0.18423, 0.1899529, 0.1585699, 0.2774961, 0.2844732, 0.247682, 0.3502297, 
    0.4110307, 0.3013442, 0.2786723, 0.2249524, 0.07881668, 0.1756877, 
    0.1905896, 0.3113365, 0.3455195, 0.2786748, 0.3313666, 0.2870489, 
    0.2448442, 0.1005006, 0.1145443, 0.1887957, 0.1905368, 0.2801458, 
    0.3457824, 0.2873928, 0.2764474, 0.1732209,
  0.2139779, 0.2269359, 0.1895588, 0.1698148, 0.1398789, 0.1797866, 
    0.1424242, 0.2606935, 0.2305329, 0.2566413, 0.1364565, 0.1711304, 
    0.1938232, 0.2374738, 0.2714282, 0.2685562, 0.2994256, 0.2543822, 
    0.1587495, 0.1071414, 0.1092064, 0.05633517, 0.1306086, 0.03469109, 
    0.2110098, 0.1735787, 0.09369922, 0.314612, 0.2143025,
  0.1256185, 0.176698, 0.2247244, 0.2989759, 0.2430359, 0.1589846, 0.2020354, 
    0.2454416, 0.2257612, 0.1293673, 0.07932021, 0.122808, 0.2409103, 
    0.1991288, 0.1531589, 0.125615, 0.07710247, 0.08035605, 0.08301336, 
    0.08602889, 0.06431674, 0.04730817, 0.03979905, -0.002638107, 0.06308522, 
    0.03073268, 0.08287092, 0.1565644, 0.2096837,
  0.01556732, 0.01544515, 0.01532297, 0.0152008, 0.01507862, 0.01495645, 
    0.01483428, 0.03429533, 0.03673541, 0.0391755, 0.04161558, 0.04405566, 
    0.04649574, 0.04893582, 0.03728724, 0.03681803, 0.03634882, 0.03587961, 
    0.0354104, 0.03494119, 0.03447198, 0.02081973, 0.01897104, 0.01712234, 
    0.01527364, 0.01342495, 0.01157625, 0.009727555, 0.01566506,
  0.1029392, 0.0490526, 0.02798517, 0.01455064, -0.0001597832, 0.0001488154, 
    1.154597e-05, 0, 0, 0, 0, 0.002418791, 0.1187467, 0.1958351, 0.1557342, 
    0.1950129, 0.1910012, 0.1817476, 0.09514116, 0.1434841, 0.1516636, 
    0.1463031, 0.2207764, 0.1763938, 0.3119608, 0.2081845, 0.2988011, 
    0.1921826, 0.126386,
  0.3484827, 0.3638379, 0.3595975, 0.3259404, 0.2429154, 0.1150164, 
    0.0122811, 0.06393398, 0.08819477, 0.2243007, 0.1988897, 0.352208, 
    0.3471033, 0.299427, 0.2694977, 0.2109019, 0.2259343, 0.2460219, 
    0.2863319, 0.168782, 0.1483699, 0.2809724, 0.3541339, 0.3968143, 
    0.3199244, 0.1656941, 0.2535834, 0.2417463, 0.2633038,
  0.2186674, 0.257938, 0.3363217, 0.324062, 0.3134462, 0.3262954, 0.2642692, 
    0.2539364, 0.2199588, 0.277258, 0.2960482, 0.3839517, 0.3370176, 
    0.3075191, 0.2334198, 0.1905687, 0.2456963, 0.2649464, 0.262109, 
    0.3326901, 0.3133513, 0.2911539, 0.2704998, 0.2982895, 0.2884377, 
    0.2228167, 0.304558, 0.2240229, 0.2333656,
  0.2119507, 0.1715571, 0.1555116, 0.1603186, 0.1631843, 0.08304828, 
    0.09056295, 0.1173249, 0.1938814, 0.2230742, 0.2022499, 0.2073432, 
    0.1228151, 0.1062259, 0.09011839, 0.09619865, 0.09369451, 0.1108002, 
    0.09998401, 0.1537132, 0.1716822, 0.1894812, 0.1586219, 0.0794041, 
    0.1064583, 0.1723639, 0.1322048, 0.1608401, 0.1826128,
  0.03709417, 0.01570508, 0.01631256, 0.1303642, 0.02229576, 0.1124457, 
    0.0638778, 0.08638145, 0.02256683, 0.01321628, 0.03557909, 0.05359478, 
    0.06995077, 0.01876429, 0.1367404, 0.1286527, 0.06420006, 0.06996388, 
    0.1037653, 0.1081893, 0.1014935, 0.04825374, 0.001927255, 0.009932422, 
    0.06966746, 0.08347953, 0.08382388, 0.09330247, 0.04389027,
  0.0004827497, -3.260641e-05, 0.1427868, 0.02471102, 0.02833497, 0.1834802, 
    0.04405573, 0.002305588, 9.292195e-08, 0.009852624, 0.08527233, 
    0.09976341, 0.02811556, 0.0494222, 0.2646316, 0.01812332, 0.1292963, 
    0.1281057, 0.1028893, 0.04640523, 0.03782546, 0.00128925, 7.404518e-08, 
    0.003333028, 0.01706861, 0.1129331, 0.03614438, 0.02153911, 0.00235011,
  0.0004267496, 0.09486245, 0.08067781, 0.01060731, 0.2425013, 0.01916437, 
    0.003614627, 3.309342e-05, 0.0004387113, 0.03912928, 0.1794292, 
    0.04697156, 0.009080946, 0.08593816, 0.2535186, 0.1246084, 0.1350947, 
    0.04937221, 0.007602206, 0.009347217, -1.139346e-07, 2.177132e-06, 
    2.322055e-06, 0.0002254065, 0.09136516, 0.3221427, 0.003532241, 
    0.0001928061, 1.09102e-05,
  0.006180988, 0.09684011, 0.2919741, 0.1367122, 0.04215069, 0.009918374, 
    0.01307626, 0.002601775, 0.003652255, 0.02067466, 0.05967039, 0.08768863, 
    0.2240019, 0.1745866, 0.322745, 0.0790629, 0.01780191, 0.02006734, 
    0.01087354, 1.268573e-05, -4.030911e-07, 0.0244721, 0.00858256, 
    0.2534794, 0.4081791, 0.2808739, 0.01638119, 0.0008023452, 0.01126966,
  0.1716344, 0.05741544, 0.06686509, 0.02310728, 0.1237045, 0.1192937, 
    0.1676314, 0.1607137, 0.1200575, 0.06456309, 0.1042738, 0.02483351, 
    0.02198385, 0.07102569, 0.09776787, 0.01524665, 7.340219e-06, 
    -0.0001959948, 0.001606615, 0.01888169, 0.07495248, 0.05195078, 
    0.1328097, 0.04337467, 0.07708501, 0.403281, 0.02307652, 0.004595474, 
    0.02559857,
  7.102362e-06, 6.351356e-06, 0.0001320411, 0.03034708, 0.01641066, 
    0.001591653, 1.60569e-05, -1.091769e-05, 0.001486172, 0.04332983, 
    0.2305875, 0.0617429, 0.09821417, 0.08300745, 0.01495568, 0.01958766, 
    0.1114123, 0.1514534, 0.1477915, 0.1212409, 0.0997813, 0.003899148, 
    0.005759349, 0.002284261, 0.002752141, 0.0001825299, 9.147806e-08, 
    7.014948e-06, 5.974923e-05,
  4.315838e-06, 1.679058e-06, 2.936348e-08, 5.492853e-08, 0.0002799185, 
    3.901144e-07, 8.829676e-07, 0.0001440649, -9.648153e-08, 0.02040249, 
    0.08577874, 0.05400702, 1.568552e-06, 0.007329568, 0.03335411, 
    0.0007709841, 0.02682928, 0.0640022, 0.02133371, 0.05337754, 0.009613125, 
    0.02380568, 0.01497384, 0.001503578, -1.495396e-05, -4.575841e-07, 
    0.001598073, 6.798974e-05, -6.552458e-05,
  -2.541644e-06, 1.736351e-07, 0.004625341, 0.01939558, 0.05396337, 
    0.06267727, 0.009926789, 0.01294739, 0.1488969, 0.305977, 0.1438011, 
    0.03334394, 0.04106702, 0.04234663, 0.0506132, 0.06113312, 0.03352717, 
    0.08274601, 0.02445769, -3.997536e-05, 0.02306771, 0.05822195, 0.1147104, 
    0.03009597, 0.04700421, 0.04767419, 0.03453077, 0.05493931, 0.03833979,
  0.1166451, 0.05072584, 0.05025431, 0.0916549, 0.1223617, 0.1115554, 
    0.2263383, 0.04462335, 0.109074, 0.07709824, 0.1224476, 0.09102684, 
    0.1097965, 0.1724034, 0.1895165, 0.263724, 0.1921845, 0.1696997, 
    0.03685721, 0.04178936, 0.1553686, 0.158409, 0.1603536, 0.2384219, 
    0.190999, 0.1603359, 0.1692728, 0.1227263, 0.1401736,
  0.1139737, 0.1052497, 0.09883776, 0.1016961, 0.2106564, 0.1826245, 
    0.1858741, 0.121575, 0.07704058, 0.03151697, 0.04135968, 0.03222486, 
    0.09182522, 0.2623164, 0.2467859, 0.150306, 0.2036725, 0.2592162, 
    0.2572737, 0.3010523, 0.2353888, 0.1516147, 0.22196, 0.1674613, 
    0.2527203, 0.226097, 0.265045, 0.1752844, 0.1149986,
  0.1705312, 0.1871659, 0.1531367, 0.2760584, 0.2822817, 0.2353165, 
    0.3398531, 0.3637981, 0.3023928, 0.2624615, 0.2502938, 0.09922363, 
    0.2386987, 0.2231195, 0.2988647, 0.3449811, 0.2957801, 0.3120547, 
    0.2893798, 0.2422017, 0.109735, 0.1468498, 0.2118987, 0.2187815, 
    0.2723045, 0.3308707, 0.264401, 0.2573204, 0.188235,
  0.1958588, 0.216247, 0.2030266, 0.1704338, 0.1571486, 0.2312544, 0.144052, 
    0.326153, 0.3277446, 0.3578364, 0.1902234, 0.2862494, 0.2595056, 
    0.2129571, 0.2901748, 0.2540429, 0.2928572, 0.2469279, 0.1464832, 
    0.08997884, 0.1117502, 0.06817483, 0.1322624, 0.1052027, 0.1811941, 
    0.2491697, 0.1711787, 0.295487, 0.2098548,
  0.1212651, 0.1734356, 0.2241859, 0.3104326, 0.2325878, 0.1497211, 
    0.2116005, 0.2823451, 0.2525128, 0.1817422, 0.09852847, 0.2096781, 
    0.3128182, 0.2718441, 0.133687, 0.10339, 0.06967338, 0.07745539, 
    0.07500722, 0.0903824, 0.100029, 0.08017135, 0.04871071, 0.0135218, 
    0.059891, 0.04803326, 0.1153518, 0.1518333, 0.1958721,
  0.1294536, 0.1206586, 0.1118636, 0.1030686, 0.09427362, 0.08547864, 
    0.07668366, 0.0766302, 0.08159279, 0.08655537, 0.09151796, 0.09648054, 
    0.1014431, 0.1064057, 0.09275403, 0.09906659, 0.1053791, 0.1116917, 
    0.1180043, 0.1243168, 0.1306294, 0.1646213, 0.1621412, 0.159661, 
    0.1571809, 0.1547007, 0.1522205, 0.1497404, 0.1364895,
  0.1116929, 0.1003812, 0.07157033, 0.03715359, 0.02510357, 0.002680576, 0, 
    0, 0, 0, -0.00427977, 0.1481194, 0.2895257, 0.2107148, 0.165856, 
    0.1769595, 0.1893211, 0.1750403, 0.1124312, 0.1222151, 0.1625917, 
    0.1687317, 0.2450809, 0.1579088, 0.2697817, 0.2308732, 0.2575219, 
    0.1753239, 0.1083229,
  0.368625, 0.3896137, 0.3847209, 0.3867881, 0.2399429, 0.1046842, 
    0.02543358, 0.1055886, 0.1544977, 0.307203, 0.3090898, 0.3907622, 
    0.3209141, 0.2895963, 0.2710513, 0.2278012, 0.249191, 0.2258263, 
    0.2704743, 0.1634833, 0.2097493, 0.438999, 0.4731364, 0.3692366, 
    0.298324, 0.2220652, 0.2278562, 0.2820026, 0.306848,
  0.2970138, 0.2995096, 0.345392, 0.4026175, 0.3990913, 0.366847, 0.3404127, 
    0.317444, 0.3439054, 0.3050735, 0.329544, 0.3229758, 0.3426017, 
    0.2970819, 0.2408398, 0.2024804, 0.2371431, 0.286857, 0.248048, 
    0.3645943, 0.2970673, 0.2937591, 0.2702137, 0.3350401, 0.2873358, 
    0.2596965, 0.3357424, 0.2621808, 0.3192322,
  0.2254735, 0.1817468, 0.1832286, 0.1785718, 0.2010958, 0.08907477, 
    0.0913194, 0.1217079, 0.1849554, 0.2249852, 0.2350556, 0.2032143, 
    0.1244895, 0.09782164, 0.08333898, 0.09917756, 0.08997372, 0.1044927, 
    0.1247004, 0.1805587, 0.1758303, 0.1841004, 0.1491926, 0.08426322, 
    0.1090062, 0.1614073, 0.1349105, 0.1432908, 0.1911769,
  0.05872228, 0.02034175, 0.01347483, 0.1247719, 0.01892929, 0.1277036, 
    0.06989387, 0.09889898, 0.04582592, 0.01455233, 0.03459119, 0.04462383, 
    0.0773368, 0.01947226, 0.1432887, 0.1303297, 0.05633459, 0.07448685, 
    0.108078, 0.1131555, 0.1111846, 0.06330184, 0.002410041, 0.006067328, 
    0.06721801, 0.08312045, 0.1050721, 0.1074234, 0.05220683,
  -1.451713e-06, 5.535443e-07, 0.1462941, 0.01954699, 0.02898736, 0.188792, 
    0.0416526, 0.002729089, 8.909166e-08, 0.003377089, 0.04949839, 
    0.05527138, 0.05297429, 0.05630131, 0.2387635, 0.03059802, 0.156622, 
    0.1401818, 0.1174167, 0.0458747, 0.04525221, 0.004930143, 2.647944e-08, 
    0.002298699, 0.015418, 0.1370973, 0.04244447, 0.02235273, 0.004416357,
  0.0003181005, 0.09458288, 0.09848741, 0.009441137, 0.2203078, 0.0194077, 
    0.01392788, 4.408222e-05, 0.0003667478, 0.03038539, 0.1816946, 
    0.04808909, 0.01072625, 0.07994039, 0.1971659, 0.1259068, 0.1413016, 
    0.05622457, 0.00949748, 0.009535955, 1.105756e-05, 8.025772e-07, 
    1.294036e-06, 0.0001100374, 0.07372085, 0.372199, 0.004482314, 
    4.099534e-06, 3.024229e-07,
  0.0001554375, 0.0798251, 0.3568096, 0.1451169, 0.03680491, 0.01289559, 
    0.01320637, 0.005239504, 0.003467694, 0.02483979, 0.04726183, 0.05777658, 
    0.2140587, 0.1231844, 0.2482604, 0.06316988, 0.01970463, 0.03242813, 
    0.01517481, 0.0001041921, 1.597059e-07, 0.04106151, 0.0008787273, 
    0.2767309, 0.3782548, 0.3132314, 0.01453614, 0.0003104852, 0.000333491,
  0.07639918, 0.06911489, 0.09729745, 0.027478, 0.1128892, 0.1164682, 
    0.1729419, 0.1861183, 0.1548808, 0.07690557, 0.1034505, 0.02395071, 
    0.01638591, 0.04934253, 0.08360115, 0.028267, -7.867945e-06, 
    0.0002818725, 0.001347388, 0.007294375, 0.0457163, 0.02332201, 0.1758434, 
    0.05228169, 0.1196394, 0.4059981, 0.02916505, 0.007166838, 0.002498115,
  6.969748e-07, 3.413108e-06, 0.002114768, 0.1311498, 0.01157312, 
    0.007884747, 2.963389e-05, 0.001039919, 0.003025858, 0.03836904, 
    0.2349845, 0.06725197, 0.08225898, 0.07324961, 0.01275665, 0.02301742, 
    0.1088828, 0.1518585, 0.1662682, 0.1267401, 0.1113487, 0.004235435, 
    0.007034278, 0.004234249, 0.006834455, 0.0002302566, -3.268163e-07, 
    5.77183e-06, -0.0001277348,
  2.442885e-06, 7.799616e-07, 2.006063e-07, 2.43739e-07, 0.00492389, 
    -7.457345e-07, 2.872072e-07, 2.317954e-05, 1.435936e-06, 0.01625252, 
    0.08627644, 0.04807261, -9.427907e-06, 0.003780823, 0.02679996, 
    0.001138865, 0.02849449, 0.07101796, 0.02518012, 0.03874582, 0.006313402, 
    0.03888251, 0.01397076, 0.003310661, 0.0003307702, 1.419914e-05, 
    0.002716483, 1.458408e-06, 7.749243e-05,
  2.282777e-07, -4.193711e-09, 0.005792141, 0.0182819, 0.07257037, 
    0.06042137, 0.01280416, 0.02100695, 0.1507878, 0.3135662, 0.1523729, 
    0.0465367, 0.04740291, 0.04004726, 0.08124999, 0.07683748, 0.03389273, 
    0.09610728, 0.003954007, 0.001548854, 0.02553012, 0.05550674, 0.1105197, 
    0.02677182, 0.05699227, 0.04968093, 0.03763016, 0.03624254, 0.02018782,
  0.1073189, 0.04332069, 0.04731031, 0.09299657, 0.1105706, 0.09954061, 
    0.2245989, 0.0283589, 0.08209093, 0.08135758, 0.1111898, 0.08800686, 
    0.105799, 0.1808554, 0.1993753, 0.2545922, 0.178283, 0.1555761, 
    0.03434877, 0.04750267, 0.1834311, 0.1625795, 0.1670609, 0.2435735, 
    0.1652016, 0.1693217, 0.1829737, 0.1205582, 0.1442301,
  0.1012831, 0.08551441, 0.09363761, 0.1211318, 0.1930634, 0.1732293, 
    0.1483853, 0.1173561, 0.06640956, 0.03254014, 0.04088522, 0.03746725, 
    0.08754008, 0.2682461, 0.2555262, 0.1459148, 0.2002034, 0.2552025, 
    0.2496282, 0.2836245, 0.2508271, 0.1523114, 0.2437059, 0.1894901, 
    0.2652678, 0.221697, 0.2749743, 0.1652222, 0.1116117,
  0.1426326, 0.1908648, 0.1566708, 0.2590215, 0.2841194, 0.2236838, 
    0.3489928, 0.3679283, 0.2893465, 0.2634244, 0.2845753, 0.1125936, 
    0.2713965, 0.2342113, 0.2845728, 0.3355695, 0.2915881, 0.3210702, 
    0.2950492, 0.2380853, 0.1062659, 0.1902474, 0.2337976, 0.2572741, 
    0.2779623, 0.3097177, 0.2463768, 0.2499477, 0.1941159,
  0.1856313, 0.2176257, 0.2134757, 0.1940109, 0.1911012, 0.2122408, 
    0.1650207, 0.3647997, 0.3319373, 0.4354088, 0.2478489, 0.3120213, 
    0.1960036, 0.1783637, 0.3224125, 0.2704314, 0.2883296, 0.257967, 
    0.1487485, 0.07273419, 0.1099424, 0.07178554, 0.1416047, 0.129985, 
    0.1481918, 0.3087187, 0.2793064, 0.2939478, 0.1984052,
  0.1151084, 0.1692899, 0.2280996, 0.3287851, 0.2176038, 0.138804, 0.2074409, 
    0.3092482, 0.2956683, 0.2531392, 0.1845676, 0.2671657, 0.2714496, 
    0.2566777, 0.139874, 0.1015136, 0.06588838, 0.07248639, 0.1033046, 
    0.1665091, 0.1327742, 0.1265702, 0.07597548, 0.02877132, 0.06076474, 
    0.05859401, 0.1188072, 0.1359554, 0.1807548,
  0.2422447, 0.2411297, 0.2400147, 0.2388997, 0.2377847, 0.2366697, 
    0.2355547, 0.2220762, 0.2281189, 0.2341615, 0.2402042, 0.2462469, 
    0.2522895, 0.2583322, 0.269016, 0.26841, 0.2678039, 0.2671979, 0.2665918, 
    0.2659858, 0.2653798, 0.2642555, 0.2599339, 0.2556123, 0.2512906, 
    0.246969, 0.2426474, 0.2383258, 0.2431367,
  0.1337328, 0.1191146, 0.1626411, 0.04623549, 0.04380885, 0.01434937, 
    9.777895e-05, 0, 0, 0.0001016415, 0.07435144, 0.240513, 0.3479039, 
    0.2406854, 0.1429972, 0.1584449, 0.2161851, 0.1967986, 0.1447313, 
    0.1604692, 0.2222331, 0.2228237, 0.2858723, 0.2477538, 0.2778411, 
    0.2252254, 0.2150092, 0.1665857, 0.09041143,
  0.3864876, 0.358072, 0.3525341, 0.4284711, 0.2540665, 0.08965838, 
    0.08010203, 0.133454, 0.1789073, 0.312451, 0.3158166, 0.3818173, 
    0.2919859, 0.2907253, 0.2689704, 0.3061861, 0.2675573, 0.2985503, 
    0.3248907, 0.2559396, 0.2375662, 0.3700237, 0.4184048, 0.3972819, 
    0.2702606, 0.1512451, 0.1527688, 0.2289166, 0.38828,
  0.2711147, 0.3660074, 0.3349021, 0.3150021, 0.3216218, 0.3104268, 
    0.2899068, 0.2520894, 0.2732508, 0.334119, 0.3587359, 0.4230572, 
    0.3446418, 0.2938269, 0.2365461, 0.1988598, 0.2175366, 0.2750748, 
    0.2694302, 0.3041897, 0.2916401, 0.265184, 0.2810516, 0.3304369, 
    0.2929096, 0.2475339, 0.3386855, 0.2449808, 0.340652,
  0.2433965, 0.2010387, 0.1879584, 0.1706751, 0.1762576, 0.09884308, 
    0.09385124, 0.1300029, 0.2060578, 0.214973, 0.2272204, 0.2066309, 
    0.1392096, 0.09614889, 0.08361354, 0.08768782, 0.084548, 0.119632, 
    0.1385481, 0.1807887, 0.1768759, 0.1932012, 0.1707356, 0.09427133, 
    0.1033556, 0.1669883, 0.1243433, 0.1599438, 0.2378409,
  0.06119053, 0.03820808, 0.01743091, 0.1232195, 0.03558418, 0.1441334, 
    0.0825187, 0.09986869, 0.06406163, 0.01451976, 0.03533452, 0.02862511, 
    0.05495451, 0.01434795, 0.1659218, 0.1137533, 0.05904492, 0.07961754, 
    0.1149022, 0.1206103, 0.1058952, 0.05763283, 0.008577249, 0.003898669, 
    0.05200658, 0.08802087, 0.1428205, 0.1270203, 0.05742782,
  1.050163e-05, 3.963407e-06, 0.1686544, 0.02365868, 0.03527105, 0.1707783, 
    0.03438009, 0.001699954, 1.019425e-07, 0.001902978, 0.02774421, 
    0.02495313, 0.0730315, 0.05307072, 0.2087048, 0.05010691, 0.11937, 
    0.1420829, 0.08410782, 0.04513193, 0.05435752, 0.00736276, -1.882794e-06, 
    0.001091212, 0.0153161, 0.129284, 0.04320323, 0.0235023, 0.005434501,
  0.001408568, 0.06765041, 0.09933756, 0.00977798, 0.1711032, 0.02545763, 
    0.03151118, -7.857891e-06, -2.762479e-06, 0.003439293, 0.1542708, 
    0.04113198, 0.01351652, 0.0699525, 0.1484461, 0.1018413, 0.1158553, 
    0.04798663, 0.01478834, 0.02025799, 0.001296807, 3.34824e-07, 
    4.379215e-07, 0.0001514993, 0.06524137, 0.3860522, 0.0121033, 
    0.002004717, 3.134178e-05,
  0.0001737202, 0.03904967, 0.3991872, 0.1042241, 0.02427397, 0.015728, 
    0.02042264, 0.007401286, 0.00268682, 0.02150054, 0.03353409, 0.04117038, 
    0.1955285, 0.1010131, 0.2049312, 0.05379516, 0.01910495, 0.02701687, 
    0.01535434, 0.0003341837, -3.686208e-07, 0.01367047, 0.0004843473, 
    0.2139515, 0.2640478, 0.2493092, 0.01423023, 0.001273939, 1.00153e-05,
  0.03231301, 0.06054553, 0.06455418, 0.03977484, 0.0948372, 0.1125341, 
    0.1690034, 0.1883335, 0.1487639, 0.07507513, 0.0973219, 0.0205877, 
    0.01413735, 0.03505749, 0.0708695, 0.03558981, 1.682923e-05, 
    0.0008527893, 0.001042308, 0.01238449, 0.02047175, 0.01017971, 0.1811431, 
    0.06925387, 0.128469, 0.3839144, 0.03491048, 0.008373658, 0.0005755814,
  8.459041e-08, 1.022965e-06, 0.0002597276, 0.240599, 0.01330369, 0.01783906, 
    0.0001854072, 0.00166, 0.008454385, 0.04735815, 0.2474935, 0.07472987, 
    0.07026285, 0.06869164, 0.01462635, 0.02405259, 0.09208843, 0.1447996, 
    0.1467353, 0.1234738, 0.1203988, 0.003895918, 0.01048146, 0.009171924, 
    0.01159606, 0.0002562708, -6.085044e-06, 4.069761e-06, 2.781167e-05,
  1.32348e-06, 2.334752e-07, 6.849442e-08, 1.403664e-05, 0.001599397, 
    3.989933e-07, -1.217019e-07, 7.719346e-05, 7.211431e-05, 0.01916551, 
    0.1161369, 0.01817939, 1.727854e-05, 0.003401982, 0.03011438, 
    0.002452756, 0.03136871, 0.07111347, 0.01865463, 0.02057448, 0.001516626, 
    0.05995717, 0.01548179, 0.01404558, 0.002787813, 0.0008023293, 
    0.004444297, 1.159965e-06, 1.088392e-05,
  -2.351493e-08, 4.072323e-08, 0.007011923, 0.01812946, 0.08918795, 
    0.05930454, 0.01813346, 0.02188649, 0.1468812, 0.3237774, 0.129408, 
    0.05057773, 0.06331868, 0.04889589, 0.08928737, 0.08920933, 0.04945217, 
    0.1129892, 6.116895e-05, 0.00417234, 0.02734301, 0.05413954, 0.1147104, 
    0.04147982, 0.07703666, 0.05478071, 0.0480829, 0.02875992, 0.003400509,
  0.1122975, 0.03641949, 0.04215309, 0.1045902, 0.1115949, 0.08663035, 
    0.2190034, 0.01634778, 0.06292704, 0.1006431, 0.1109244, 0.0867257, 
    0.09804085, 0.2263944, 0.2025444, 0.2444775, 0.1655938, 0.1481082, 
    0.03407351, 0.05259328, 0.1962525, 0.1791727, 0.1958701, 0.2314325, 
    0.1444064, 0.1682793, 0.1964899, 0.1196767, 0.1429666,
  0.09842514, 0.07683089, 0.09581265, 0.1437921, 0.1908812, 0.2289438, 
    0.1330967, 0.1255899, 0.05985699, 0.03194328, 0.0408377, 0.04319058, 
    0.07582891, 0.2665258, 0.2901427, 0.1511943, 0.2026244, 0.2209812, 
    0.2420735, 0.2730794, 0.2479259, 0.1608476, 0.2578265, 0.1937795, 
    0.2812588, 0.2196046, 0.2619891, 0.1719027, 0.1051593,
  0.1402498, 0.187897, 0.1671238, 0.2593596, 0.3137538, 0.2359504, 0.3794689, 
    0.3854214, 0.2824691, 0.288845, 0.2994008, 0.1231677, 0.2908327, 
    0.246222, 0.2943231, 0.3554354, 0.3160205, 0.3294098, 0.2990806, 0.26047, 
    0.1305144, 0.2224259, 0.2491299, 0.2600934, 0.2708925, 0.3152809, 
    0.2331503, 0.2560026, 0.1785725,
  0.1934817, 0.2411496, 0.2272003, 0.2150712, 0.2155102, 0.2185531, 
    0.1927328, 0.3822727, 0.3451285, 0.4585012, 0.2566258, 0.2945612, 
    0.1777091, 0.1738949, 0.3325801, 0.2557398, 0.321466, 0.2709788, 
    0.1393609, 0.06863379, 0.1066474, 0.1166167, 0.1691014, 0.1382681, 
    0.1323917, 0.402701, 0.366805, 0.3206296, 0.2065547,
  0.1078101, 0.1818083, 0.2341674, 0.3622701, 0.2108815, 0.1505097, 
    0.2183984, 0.3051116, 0.3031907, 0.279525, 0.1712572, 0.2809479, 
    0.2579361, 0.2299525, 0.1588284, 0.1036424, 0.08225415, 0.0760424, 
    0.1085587, 0.1819036, 0.1432523, 0.1393196, 0.1324229, 0.04319767, 
    0.06528179, 0.06770805, 0.1207763, 0.125156, 0.1653686,
  0.256148, 0.2574337, 0.2587193, 0.2600049, 0.2612906, 0.2625762, 0.2638618, 
    0.2700847, 0.2802829, 0.290481, 0.3006792, 0.3108774, 0.3210755, 
    0.3312737, 0.3429289, 0.3360464, 0.3291639, 0.3222815, 0.315399, 
    0.3085165, 0.301634, 0.2741586, 0.2695573, 0.2649559, 0.2603546, 
    0.2557533, 0.2511519, 0.2465506, 0.2551195,
  0.1633203, 0.1435377, 0.216681, 0.1800629, 0.06700139, 0.02666355, 
    -0.000138139, -7.318689e-05, -2.831252e-07, 0.004039646, 0.2208219, 
    0.2932307, 0.3443769, 0.2912158, 0.1288623, 0.1341699, 0.1993051, 
    0.2099385, 0.1475243, 0.1434651, 0.2634954, 0.2651453, 0.2919984, 
    0.151091, 0.2036768, 0.1935126, 0.1802169, 0.1679832, 0.08786323,
  0.3692642, 0.411583, 0.4093236, 0.5484127, 0.2601216, 0.06913361, 
    0.1008773, 0.1938211, 0.1979289, 0.3140467, 0.3101827, 0.3428136, 
    0.2923513, 0.3211235, 0.2832143, 0.290823, 0.2717608, 0.2624958, 
    0.4009149, 0.3252754, 0.3764374, 0.3883367, 0.5378963, 0.4625233, 
    0.2175056, 0.1327975, 0.2209502, 0.3229378, 0.4406662,
  0.3058927, 0.3780274, 0.4075057, 0.3613275, 0.3986503, 0.3804947, 
    0.3335387, 0.3228316, 0.3140709, 0.3841664, 0.3632685, 0.4188908, 
    0.3591967, 0.2790289, 0.2542717, 0.2164947, 0.2355951, 0.3315617, 
    0.3016477, 0.3577499, 0.3654226, 0.2899643, 0.2894031, 0.3392855, 
    0.3125281, 0.2851797, 0.3230512, 0.3001533, 0.3508733,
  0.2352555, 0.1957083, 0.2095753, 0.1994893, 0.1724681, 0.09964297, 
    0.1140701, 0.1361464, 0.2093417, 0.2411431, 0.2772332, 0.213273, 
    0.1484338, 0.0970047, 0.08938672, 0.09312551, 0.08671539, 0.120518, 
    0.1642706, 0.1952043, 0.1852626, 0.2034751, 0.1728778, 0.1159493, 
    0.09150346, 0.1901158, 0.1059943, 0.1567055, 0.2341662,
  0.07153916, 0.03802678, 0.02902161, 0.1331348, 0.04499826, 0.1438044, 
    0.0849306, 0.1123105, 0.07487738, 0.03150913, 0.03611046, 0.01645585, 
    0.02358118, 0.009972936, 0.1962812, 0.1006485, 0.05524537, 0.07696922, 
    0.107948, 0.1163561, 0.1009742, 0.05795275, 0.01176935, 0.00127544, 
    0.04007201, 0.08229885, 0.1302357, 0.1244136, 0.04868401,
  0.0001511492, 2.423087e-06, 0.1517966, 0.03569221, 0.03822352, 0.1627183, 
    0.02561842, 0.001106951, 5.613698e-08, -0.0002686274, 0.02523047, 
    0.01587222, 0.06814461, 0.05333028, 0.2037525, 0.07007472, 0.1035215, 
    0.1128141, 0.0573982, 0.04354322, 0.06706435, 0.007396853, -1.240739e-05, 
    0.0006290162, 0.01138035, 0.1357226, 0.04183122, 0.02168521, 0.007918755,
  0.0003974688, 0.05249697, 0.08087073, 0.01493694, 0.1374462, 0.03597319, 
    0.03501023, 0.0001166902, 5.848096e-08, -6.985925e-05, 0.1348559, 
    0.03309025, 0.02070871, 0.05225431, 0.1274441, 0.08907994, 0.1003976, 
    0.03779115, 0.02352146, 0.04820877, 0.02006665, 9.112692e-06, 
    7.292768e-08, 8.299124e-05, 0.07625237, 0.3485199, 0.02745413, 
    0.01460352, 0.002037653,
  5.003937e-06, 0.01325447, 0.2962696, 0.08420848, 0.01890433, 0.01647253, 
    0.02929913, 0.01166086, 0.003762689, 0.0152311, 0.02214066, 0.03234593, 
    0.1489194, 0.08429679, 0.1875973, 0.06070159, 0.02543193, 0.01958534, 
    0.01751188, 0.004878475, 2.524093e-05, 0.003448563, 0.000407117, 
    0.2000419, 0.2134604, 0.2090093, 0.01728159, 0.003347459, 2.803346e-06,
  0.01161388, 0.03329688, 0.03129987, 0.05902313, 0.08972446, 0.1113798, 
    0.1578358, 0.1989963, 0.1767606, 0.09764949, 0.07835817, 0.01734041, 
    0.01436546, 0.03600285, 0.07664531, 0.06943731, -0.0001895794, 
    0.003461447, 0.003741043, 0.005070942, 0.002290851, 0.009224633, 
    0.1473622, 0.05852436, 0.133511, 0.3537526, 0.04953894, 0.0127248, 
    0.0007733072,
  9.004864e-08, 3.227543e-07, 1.073316e-05, 0.2918363, 0.01642862, 
    0.02170718, 0.0003144143, 0.002444924, 0.02568869, 0.06230665, 0.2573856, 
    0.08234345, 0.06252532, 0.06306759, 0.02261158, 0.03353671, 0.08271953, 
    0.1374631, 0.1378298, 0.1283026, 0.1169942, 0.003995185, 0.0219136, 
    0.01727455, 0.01654371, 0.0003439751, -2.036067e-05, 2.041414e-06, 
    -0.0004456738,
  1.432059e-06, 8.893868e-08, 4.765951e-08, 0.001079514, 0.01511868, 
    3.842653e-07, -6.705235e-06, 2.933045e-05, 0.00700059, 0.02719448, 
    0.1558474, 0.01087747, 0.000813516, 0.04592628, 0.02953223, 0.008270678, 
    0.03435055, 0.06242606, 0.01217225, 0.0147303, 0.0002633616, 0.07723728, 
    0.01288684, 0.02470661, 0.006573453, 0.001789506, 0.006204718, 
    4.463444e-07, 5.015408e-06,
  1.514568e-07, -2.099176e-06, 0.02380283, 0.02064781, 0.1107617, 0.0663131, 
    0.004309229, 0.01918341, 0.1386239, 0.3231232, 0.1511461, 0.05301902, 
    0.07038516, 0.06253839, 0.0990492, 0.1101987, 0.09944775, 0.1354426, 
    1.365675e-05, 0.008324945, 0.03674361, 0.0611688, 0.11319, 0.06300335, 
    0.07660384, 0.05293604, 0.05149281, 0.03075969, 0.0001524366,
  0.1180762, 0.02715773, 0.03989748, 0.1331373, 0.1276003, 0.07348739, 
    0.2196909, 0.006804198, 0.04382347, 0.1054017, 0.1138011, 0.09911158, 
    0.1021248, 0.2365173, 0.1919575, 0.2389968, 0.1469658, 0.140924, 
    0.04169475, 0.0603322, 0.1931501, 0.165536, 0.1883746, 0.1988823, 
    0.1388675, 0.1772237, 0.1990508, 0.1184552, 0.145014,
  0.09765759, 0.0645496, 0.1010049, 0.1744024, 0.2207069, 0.2971038, 
    0.1458992, 0.1224211, 0.04688507, 0.02674283, 0.04069325, 0.05310714, 
    0.07579117, 0.2912522, 0.3165492, 0.1819935, 0.2090466, 0.2328387, 
    0.2401725, 0.2635749, 0.2447277, 0.1596406, 0.2050342, 0.2133273, 
    0.2880269, 0.2318639, 0.2776281, 0.1633687, 0.09605896,
  0.1530765, 0.1749707, 0.1654882, 0.2875594, 0.3438364, 0.2750834, 
    0.3998525, 0.4364806, 0.2862793, 0.3143997, 0.3055554, 0.1227346, 
    0.2945593, 0.2778765, 0.293891, 0.3585096, 0.3086664, 0.3485449, 
    0.2873823, 0.2630056, 0.142078, 0.2285818, 0.2309794, 0.2621468, 
    0.259982, 0.3432099, 0.2377984, 0.2645631, 0.1727334,
  0.1911932, 0.2229277, 0.2336818, 0.2307162, 0.2333903, 0.2034473, 
    0.2274225, 0.4183881, 0.3583291, 0.454188, 0.2742127, 0.2854522, 
    0.1678951, 0.2091715, 0.3461229, 0.2745448, 0.3297185, 0.2450736, 
    0.134744, 0.08080929, 0.09780253, 0.1818836, 0.1676458, 0.112988, 
    0.1178278, 0.4886838, 0.3978683, 0.3303198, 0.2155178,
  0.1176431, 0.1956717, 0.2458392, 0.3864132, 0.2125657, 0.1678519, 
    0.2459152, 0.3379637, 0.3130616, 0.2983263, 0.2181487, 0.3149375, 
    0.259124, 0.2087814, 0.154809, 0.09695503, 0.09691907, 0.06793287, 
    0.09103432, 0.1780955, 0.1361221, 0.1402082, 0.1522019, 0.09571531, 
    0.08183371, 0.0663798, 0.1191668, 0.1395226, 0.1701845,
  0.2635781, 0.2676706, 0.2717631, 0.2758557, 0.2799482, 0.2840407, 
    0.2881332, 0.2916895, 0.3050501, 0.3184108, 0.3317714, 0.3451321, 
    0.3584927, 0.3718534, 0.3826526, 0.3712971, 0.3599416, 0.3485861, 
    0.3372306, 0.3258751, 0.3145196, 0.2942927, 0.288195, 0.2820974, 
    0.2759997, 0.269902, 0.2638044, 0.2577067, 0.2603041,
  0.1995254, 0.1901483, 0.2466969, 0.339144, 0.1199497, 0.04271504, 
    -0.004761435, -0.005938487, 0.001707348, 0.1933287, 0.2975616, 0.3131662, 
    0.3559496, 0.275305, 0.1929058, 0.1696932, 0.1486781, 0.1955005, 
    0.134621, 0.1382216, 0.2937438, 0.3075839, 0.2681619, 0.07108933, 
    0.1007649, 0.1626002, 0.1408821, 0.1697619, 0.1774857,
  0.3772948, 0.4381663, 0.4094429, 0.4915593, 0.2810471, 0.05582555, 
    0.08723737, 0.2604658, 0.2489447, 0.3698511, 0.3125952, 0.3211854, 
    0.2853532, 0.3168587, 0.3405583, 0.3122647, 0.294282, 0.3679165, 
    0.4243264, 0.2148518, 0.3255678, 0.3300267, 0.5565194, 0.4511425, 
    0.1708218, 0.1127966, 0.1928385, 0.2456065, 0.4173397,
  0.3227083, 0.3557429, 0.3879865, 0.3622577, 0.3371899, 0.3333962, 
    0.3093929, 0.2982997, 0.2954385, 0.3788229, 0.3224103, 0.3819014, 
    0.3350566, 0.304606, 0.2517923, 0.2208154, 0.2422757, 0.3210581, 
    0.3606454, 0.3471385, 0.3132337, 0.2689969, 0.30843, 0.3379169, 
    0.3839837, 0.288995, 0.3143363, 0.3278846, 0.3512551,
  0.257844, 0.2238617, 0.2275505, 0.2074082, 0.1804757, 0.1127547, 0.113539, 
    0.130417, 0.2213406, 0.2913501, 0.3035696, 0.2376629, 0.1650897, 
    0.08995815, 0.1028267, 0.09044896, 0.09394556, 0.1361889, 0.1893661, 
    0.2183303, 0.2158771, 0.2330574, 0.1850697, 0.1586266, 0.07761057, 
    0.1491391, 0.1093735, 0.1830019, 0.2514634,
  0.05862566, 0.04137019, 0.05041987, 0.1638868, 0.0408483, 0.1311418, 
    0.06207115, 0.1294798, 0.08088828, 0.03286374, 0.03214523, 0.007226864, 
    0.01335494, 0.01021797, 0.1919694, 0.09779967, 0.04173771, 0.07097687, 
    0.09754462, 0.1130829, 0.1130918, 0.05785289, 0.03203931, 3.74335e-05, 
    0.01975041, 0.07665783, 0.1250862, 0.09911025, 0.04740488,
  0.001702594, 2.402418e-07, 0.1334332, 0.04558735, 0.04552136, 0.1480292, 
    0.02974431, 0.008231259, -7.61629e-08, -9.587343e-06, 0.01785886, 
    0.01105784, 0.05792392, 0.04160825, 0.2245792, 0.08406656, 0.103258, 
    0.1180142, 0.05384582, 0.03980077, 0.0694965, 0.01411495, -6.08275e-05, 
    0.0003499429, 0.012213, 0.1346059, 0.03899623, 0.02461523, 0.01675907,
  0.000354146, 0.03963607, 0.1020828, 0.01826473, 0.129985, 0.03960235, 
    0.03686367, 0.007840415, 5.84846e-08, -1.623169e-05, 0.1189303, 
    0.03595135, 0.03609693, 0.0500329, 0.1086036, 0.07918844, 0.08740006, 
    0.02860954, 0.03143731, 0.0514542, 0.07953165, 0.002469083, 1.472496e-08, 
    2.38769e-05, 0.08586539, 0.3225917, 0.03376224, 0.03794384, 0.01636276,
  2.151119e-06, 0.004058518, 0.2512717, 0.07323992, 0.01880152, 0.01667594, 
    0.03396238, 0.01452111, 0.005953397, 0.01697015, 0.02511086, 0.02681909, 
    0.1256818, 0.07148595, 0.1771539, 0.06172397, 0.03477287, 0.02298658, 
    0.02437916, 0.01274078, 0.003968874, 0.0008707746, 0.0006048856, 
    0.1811724, 0.1801723, 0.1651704, 0.0200342, 0.002746492, -7.299117e-06,
  0.002266723, 0.01790943, 0.01640646, 0.0638425, 0.08974612, 0.1004377, 
    0.1467863, 0.1932763, 0.2088133, 0.1076487, 0.05896109, 0.01562459, 
    0.01473959, 0.03572278, 0.0763154, 0.07163244, 0.001236074, 0.001290895, 
    0.006171024, 0.007986737, 0.003000979, 0.01760473, 0.1101689, 0.04860596, 
    0.1375061, 0.3234939, 0.0498071, 0.01927623, 0.001173823,
  4.057101e-08, 1.032811e-07, 1.4488e-06, 0.1946819, 0.01455189, 0.02834028, 
    0.001455253, 0.002981717, 0.03309618, 0.06603931, 0.2631657, 0.08314428, 
    0.06083247, 0.06362504, 0.02558722, 0.04011652, 0.06871155, 0.1373693, 
    0.1297095, 0.1299779, 0.119898, 0.007726693, 0.03463503, 0.03972098, 
    0.03537013, 0.0007463064, -1.348127e-05, 7.28668e-07, -8.391927e-05,
  1.665614e-06, 3.905689e-08, 4.353534e-08, 0.00272368, 0.009995208, 
    2.8663e-07, -1.105787e-06, 2.70887e-05, 0.02983658, 0.02861701, 
    0.1715568, 0.0149034, 0.006571287, 0.04460507, 0.03945632, 0.01949021, 
    0.03386538, 0.05486786, 0.01066835, 0.02172035, 0.000319051, 0.09399573, 
    0.01715269, 0.02672406, 0.01040323, 0.004927137, 0.008380425, 
    1.555051e-07, 2.452856e-06,
  3.942949e-07, 0.0003103254, 0.05975225, 0.0440913, 0.1128736, 0.05968551, 
    -0.002010104, 0.01762508, 0.1198248, 0.3020951, 0.1706376, 0.05384184, 
    0.0957326, 0.1102989, 0.1211068, 0.1255354, 0.09720113, 0.1647699, 
    0.002662733, 0.009365987, 0.03591804, 0.08715791, 0.139018, 0.07291744, 
    0.07488147, 0.05688754, 0.05183152, 0.03571114, 0.0002841653,
  0.1255529, 0.02614963, 0.04727578, 0.1806662, 0.1219421, 0.07131059, 
    0.2257931, 0.007008856, 0.03032366, 0.09881406, 0.1076226, 0.125204, 
    0.1434315, 0.2462597, 0.1920243, 0.2324632, 0.1890513, 0.1438666, 
    0.05742903, 0.07294479, 0.1909002, 0.1416036, 0.1827149, 0.1598388, 
    0.163086, 0.1947, 0.2029684, 0.1281387, 0.1396353,
  0.1035962, 0.05640972, 0.1068043, 0.1979612, 0.2571859, 0.302618, 
    0.1612076, 0.1105442, 0.03445562, 0.01878708, 0.03789791, 0.04854891, 
    0.08638586, 0.3195778, 0.3203626, 0.1788025, 0.2096702, 0.2377287, 
    0.2421525, 0.2504413, 0.228782, 0.1499273, 0.2018227, 0.2420337, 
    0.2542412, 0.2628189, 0.2633229, 0.190929, 0.08687158,
  0.1497101, 0.1693181, 0.1638016, 0.3261586, 0.392551, 0.3316211, 0.4776873, 
    0.4869756, 0.2693966, 0.2995482, 0.2865044, 0.1158653, 0.2784, 0.2941002, 
    0.2818147, 0.3340645, 0.3195714, 0.3632815, 0.2817793, 0.2640453, 
    0.1225235, 0.1899049, 0.2218407, 0.2948786, 0.2342114, 0.3828973, 
    0.264022, 0.2704721, 0.189136,
  0.2266291, 0.2307931, 0.2576563, 0.2399049, 0.2601729, 0.2159137, 
    0.2542724, 0.4482722, 0.3580653, 0.4583482, 0.2953315, 0.2829625, 
    0.1663531, 0.2647383, 0.3794533, 0.2584521, 0.304251, 0.2553168, 
    0.09054685, 0.06198634, 0.102224, 0.1776529, 0.1429766, 0.06887478, 
    0.1177828, 0.4945846, 0.4329746, 0.3323755, 0.2390876,
  0.1482746, 0.2343214, 0.318087, 0.382388, 0.207017, 0.1930958, 0.3126732, 
    0.3970481, 0.3466352, 0.3057804, 0.2498931, 0.3209281, 0.2676179, 
    0.2172966, 0.1491106, 0.08452617, 0.08045333, 0.07259732, 0.09331255, 
    0.1716711, 0.1318138, 0.1252491, 0.1660544, 0.1014506, 0.07962037, 
    0.05582337, 0.1198826, 0.1663456, 0.1838489,
  0.2649513, 0.270602, 0.2762529, 0.2819037, 0.2875544, 0.2932053, 0.298856, 
    0.2982433, 0.3130539, 0.3278646, 0.3426752, 0.3574858, 0.3722965, 
    0.3871071, 0.3966208, 0.3841082, 0.3715955, 0.3590828, 0.3465701, 
    0.3340574, 0.3215447, 0.3065403, 0.2985916, 0.2906429, 0.2826941, 
    0.2747454, 0.2667966, 0.2588479, 0.2604306,
  0.2281703, 0.2253346, 0.2800858, 0.3794158, 0.1596916, 0.05809788, 
    0.02678952, 0.04442529, 0.1469372, 0.2578386, 0.3044807, 0.3172175, 
    0.3625285, 0.2120968, 0.1410394, 0.1453892, 0.1285764, 0.1474376, 
    0.09658906, 0.1538533, 0.3473227, 0.3586226, 0.2282297, 0.07091682, 
    0.115141, 0.134445, 0.1421858, 0.1675139, 0.1809298,
  0.3025595, 0.4502653, 0.3394493, 0.396933, 0.2413967, 0.03575946, 
    0.06137836, 0.3033751, 0.2846683, 0.3834302, 0.3402464, 0.3179787, 
    0.279211, 0.3025806, 0.2971436, 0.3159319, 0.2936946, 0.3300701, 
    0.291356, 0.2050311, 0.2011757, 0.3031933, 0.3656253, 0.4088037, 
    0.1463033, 0.1766861, 0.255833, 0.2442615, 0.2394032,
  0.3318994, 0.3565181, 0.3166838, 0.3523814, 0.3022388, 0.2958638, 0.301535, 
    0.228568, 0.2967268, 0.3379014, 0.3208017, 0.349132, 0.3217667, 
    0.3087288, 0.2847667, 0.240212, 0.2417169, 0.3135261, 0.3644655, 
    0.3331913, 0.2908188, 0.2704032, 0.2814144, 0.3665814, 0.3863657, 
    0.2616908, 0.3078389, 0.2959864, 0.3192133,
  0.23873, 0.2228007, 0.223923, 0.2037931, 0.1864496, 0.1051106, 0.1136069, 
    0.124582, 0.2033787, 0.3089752, 0.3238482, 0.2344937, 0.1684554, 
    0.09269681, 0.1145438, 0.1040673, 0.1117358, 0.1430179, 0.1992959, 
    0.2508844, 0.2247263, 0.2313599, 0.1901289, 0.1788184, 0.05954604, 
    0.1056272, 0.1266764, 0.1688136, 0.244781,
  0.06200351, 0.08089971, 0.05084904, 0.1651574, 0.04652356, 0.1295812, 
    0.07573855, 0.1507588, 0.07334569, 0.03341635, 0.04745502, 0.01003486, 
    0.01664635, 0.01552319, 0.1853877, 0.09897434, 0.02650661, 0.0759258, 
    0.112621, 0.1247892, 0.1409896, 0.06795894, 0.03061277, 0.001371661, 
    0.005396944, 0.07850619, 0.1227301, 0.09019238, 0.04741678,
  0.01103699, 0.0001037847, 0.131457, 0.04836778, 0.06622659, 0.126549, 
    0.03945304, 0.02226986, 4.75733e-05, -2.77132e-07, 0.0172125, 0.01036627, 
    0.04174994, 0.05020512, 0.2333048, 0.09105539, 0.1102515, 0.1238808, 
    0.04480389, 0.03335928, 0.06957211, 0.0275912, 0.0003197648, 
    0.0001435928, 0.01241288, 0.1255539, 0.03821897, 0.03217605, 0.04746731,
  0.005090227, 0.02982107, 0.1131625, 0.02233525, 0.1194656, 0.03323878, 
    0.03116055, 0.03849976, 5.670022e-05, 1.513947e-05, 0.1127764, 
    0.03724126, 0.03549425, 0.04062634, 0.08313642, 0.07233903, 0.07219626, 
    0.02213332, 0.02676105, 0.04845826, 0.1040099, 0.03271345, 2.919596e-05, 
    1.674297e-05, 0.09096014, 0.2922886, 0.03031462, 0.06075355, 0.03930495,
  -1.695568e-05, 0.007434944, 0.2122719, 0.06283269, 0.01819494, 0.01624174, 
    0.02683618, 0.01579286, 0.01233769, 0.02055358, 0.03056397, 0.02400864, 
    0.1028667, 0.0549242, 0.1422512, 0.05084581, 0.02680506, 0.02046847, 
    0.02424015, 0.01222118, 0.007153163, 0.0007078173, 9.32297e-05, 
    0.1552636, 0.159076, 0.1316941, 0.02322034, 0.00478992, 0.0003922535,
  0.001077052, 0.0103625, 0.009139528, 0.0496609, 0.08760259, 0.08723824, 
    0.1275484, 0.183985, 0.2104371, 0.1201061, 0.04334391, 0.01495417, 
    0.01578772, 0.03455626, 0.07253785, 0.06937409, 0.005397573, 0.002845717, 
    0.01630859, 0.01297385, 0.007931999, 0.02853223, 0.08190556, 0.04188391, 
    0.1413326, 0.2860778, 0.042182, 0.01842392, 0.002682364,
  8.39768e-09, 2.849695e-08, 1.907659e-07, 0.08663749, 0.01951683, 
    0.03702054, 0.001591582, 0.002350847, 0.0358158, 0.06705806, 0.2404846, 
    0.06896418, 0.05848523, 0.05572518, 0.0310673, 0.04456872, 0.06034451, 
    0.1418524, 0.1273427, 0.1265228, 0.1140814, 0.01008894, 0.04906888, 
    0.03171862, 0.03790015, 0.003798258, -1.359329e-05, 1.128766e-07, 
    -7.918576e-06,
  1.498843e-06, 2.019515e-08, 2.426673e-08, 0.01348626, 0.001246109, 
    4.368433e-05, -1.37852e-08, 0.002434275, 0.05928243, 0.04837244, 
    0.1962321, 0.02174198, 0.0217023, 0.03758353, 0.05632855, 0.02179702, 
    0.02813832, 0.06132478, 0.03062124, 0.03701586, 0.0004669822, 0.1199954, 
    0.01728658, 0.02314097, 0.02754172, 0.01769306, 0.01709694, 
    -2.879792e-06, 1.607801e-06,
  1.135915e-06, 0.01183705, 0.07047314, 0.04456392, 0.102251, 0.0473127, 
    -0.002233072, 0.008481675, 0.09321306, 0.2545512, 0.1842426, 0.09978001, 
    0.1240284, 0.1398695, 0.1312951, 0.1382767, 0.09546417, 0.1752647, 
    0.01818545, 0.01377921, 0.02983192, 0.1032833, 0.126368, 0.08339505, 
    0.07262044, 0.06366038, 0.05597318, 0.04018464, 9.376156e-05,
  0.1335895, 0.03448723, 0.04612996, 0.2179321, 0.1168689, 0.07419392, 
    0.230941, 0.006870292, 0.02682921, 0.1084564, 0.09579702, 0.1818309, 
    0.1900922, 0.2873725, 0.2183799, 0.2373846, 0.205705, 0.1417527, 
    0.06348332, 0.07314873, 0.185442, 0.1275755, 0.1806006, 0.1396706, 
    0.242279, 0.2395831, 0.2251333, 0.1325928, 0.141055,
  0.1100458, 0.06291009, 0.1128061, 0.170915, 0.2229616, 0.3006781, 
    0.1348432, 0.09124995, 0.0284469, 0.01007239, 0.02915119, 0.04197189, 
    0.1215188, 0.341157, 0.3228652, 0.1969547, 0.2051719, 0.2555721, 
    0.2358813, 0.2637497, 0.2273858, 0.1335253, 0.230373, 0.2514586, 
    0.2414411, 0.3166435, 0.2679294, 0.1976362, 0.1120873,
  0.1711055, 0.1618597, 0.1699216, 0.3173221, 0.4048159, 0.3321383, 
    0.5119593, 0.5268993, 0.2760055, 0.2990344, 0.2665295, 0.1077166, 
    0.251817, 0.2805765, 0.2731254, 0.2876699, 0.3351411, 0.3726223, 
    0.2867898, 0.2712023, 0.1053667, 0.1531482, 0.2011486, 0.2902606, 
    0.2222157, 0.4181893, 0.2987495, 0.302599, 0.2035078,
  0.26498, 0.2674078, 0.2596167, 0.2629522, 0.2799887, 0.1880458, 0.2429307, 
    0.4657097, 0.3334973, 0.4522649, 0.3203532, 0.282957, 0.1864753, 
    0.2759468, 0.3922568, 0.2598322, 0.3201555, 0.2418115, 0.08942024, 
    0.04790375, 0.09987899, 0.1637721, 0.1577467, 0.04283258, 0.08757307, 
    0.511751, 0.4282777, 0.3129585, 0.2503541,
  0.1300282, 0.2262765, 0.3345388, 0.3727517, 0.2054901, 0.2058319, 
    0.3414297, 0.398953, 0.3659245, 0.3075732, 0.2423469, 0.3164847, 
    0.2953573, 0.2227431, 0.1762786, 0.1516851, 0.1143867, 0.09742443, 
    0.1298449, 0.1735453, 0.135944, 0.1109447, 0.1641213, 0.1156539, 
    0.0695703, 0.05610776, 0.1154931, 0.1934897, 0.1844234,
  0.2521323, 0.2565313, 0.2609302, 0.2653291, 0.269728, 0.2741269, 0.2785259, 
    0.2826222, 0.3011923, 0.3197623, 0.3383323, 0.3569024, 0.3754724, 
    0.3940424, 0.401199, 0.3883169, 0.3754348, 0.3625528, 0.3496707, 
    0.3367887, 0.3239066, 0.3225138, 0.312427, 0.3023401, 0.2922532, 
    0.2821663, 0.2720794, 0.2619925, 0.2486132,
  0.2523987, 0.2356615, 0.3396672, 0.4186821, 0.1909771, 0.09955412, 
    0.1022737, 0.08547015, 0.1967745, 0.3262464, 0.3076435, 0.3187424, 
    0.3711815, 0.1399688, 0.1129364, 0.1729032, 0.1321802, 0.1025611, 
    0.03807912, 0.1082444, 0.3652908, 0.3270738, 0.1695515, 0.05698546, 
    0.09630418, 0.1521698, 0.09941707, 0.1429494, 0.2278028,
  0.2679989, 0.3409349, 0.3526255, 0.3898211, 0.2627919, 0.01831823, 
    0.1182048, 0.2349543, 0.3348101, 0.3711827, 0.3428018, 0.2798183, 
    0.2555197, 0.332282, 0.360609, 0.3804564, 0.3789177, 0.3276348, 
    0.2962905, 0.1701885, 0.22602, 0.3077366, 0.3994026, 0.3883478, 
    0.2143261, 0.2620994, 0.2532736, 0.3453235, 0.3574485,
  0.4066495, 0.3457684, 0.2966307, 0.3759262, 0.3091007, 0.3505912, 
    0.2960484, 0.2233762, 0.3024218, 0.3497446, 0.3851336, 0.4066412, 
    0.3611841, 0.3443543, 0.2882056, 0.2531856, 0.2765149, 0.3263586, 
    0.3681758, 0.3776643, 0.3189031, 0.275362, 0.2984341, 0.3727815, 
    0.3259314, 0.2893288, 0.3418576, 0.3502078, 0.3684171,
  0.2619156, 0.2613402, 0.2732832, 0.2217718, 0.1794043, 0.1337255, 
    0.1269897, 0.1645458, 0.263, 0.3409142, 0.3368123, 0.2766142, 0.1935446, 
    0.1221695, 0.1259409, 0.1234562, 0.1269283, 0.1794778, 0.2626802, 
    0.2957271, 0.2560138, 0.253335, 0.2340887, 0.1733532, 0.04836513, 
    0.09243041, 0.1281747, 0.1585609, 0.2536044,
  0.09445313, 0.1093053, 0.09295396, 0.181383, 0.08527857, 0.1530733, 
    0.09012732, 0.1609955, 0.132456, 0.0988964, 0.1218328, 0.03891272, 
    0.02748001, 0.04190949, 0.186887, 0.108411, 0.03561798, 0.08893729, 
    0.1383425, 0.1282231, 0.1511964, 0.09776966, 0.05893242, 0.003221597, 
    0.004796638, 0.08494711, 0.1304778, 0.1036997, 0.06999215,
  0.02474631, 0.002010376, 0.1270005, 0.06098485, 0.08171518, 0.1113439, 
    0.04498845, 0.04243608, 0.005417321, -4.554327e-06, 0.0294145, 
    0.009581983, 0.01742395, 0.1052819, 0.2361322, 0.1125453, 0.1163363, 
    0.1330692, 0.03659599, 0.02934074, 0.06025308, 0.04459403, 0.007951465, 
    9.770903e-05, 0.01338044, 0.1242713, 0.03614086, 0.03873155, 0.07425986,
  0.01439885, 0.02324966, 0.09912212, 0.02268685, 0.08915137, 0.02562412, 
    0.02936506, 0.04802368, 0.002691763, 0.00148235, 0.1112658, 0.03852075, 
    0.03420261, 0.0376568, 0.06376429, 0.06851778, 0.06130648, 0.01994921, 
    0.02367936, 0.03342817, 0.06896979, 0.1302167, 0.003967131, 5.662409e-06, 
    0.0955959, 0.2766421, 0.02858255, 0.04598917, 0.05614515,
  0.002992418, 0.004889582, 0.1824039, 0.06056581, 0.0185388, 0.01762269, 
    0.02570516, 0.02552094, 0.03185089, 0.02128947, 0.02891419, 0.02003134, 
    0.0861252, 0.04177593, 0.1111934, 0.04451935, 0.02126594, 0.02008862, 
    0.02387858, 0.02888763, 0.007257754, 0.005274377, 0.002229837, 0.1256995, 
    0.131753, 0.1050953, 0.02630601, 0.02591884, 0.01211527,
  0.001281029, 0.009215813, 0.00543943, 0.03922351, 0.08210325, 0.0709138, 
    0.09517642, 0.1600856, 0.1800658, 0.1424387, 0.03088559, 0.01681202, 
    0.01875455, 0.03309194, 0.06374565, 0.04976966, 0.01025825, 0.00969678, 
    0.02527972, 0.02414663, 0.02728512, 0.0340259, 0.06231213, 0.03811787, 
    0.1347891, 0.2282922, 0.03419392, 0.01768102, 0.001817116,
  3.021438e-09, 6.022335e-09, 2.731818e-08, 0.04155909, 0.05197007, 
    0.03821142, 0.002039523, 0.003959159, 0.0326149, 0.06858507, 0.2131645, 
    0.05774703, 0.05516184, 0.04658715, 0.03290984, 0.04226803, 0.05181602, 
    0.1372105, 0.1270146, 0.1127188, 0.08927459, 0.01095782, 0.06055474, 
    0.02595183, 0.02936058, 0.005902698, 0.0001004396, 2.18094e-08, 
    -1.905037e-06,
  8.790431e-07, 8.644771e-09, 1.820415e-08, 0.03029388, 9.791341e-05, 
    0.001065897, 9.056465e-10, 0.000988095, 0.02054403, 0.1191622, 0.2205189, 
    0.03430716, 0.0577318, 0.07319802, 0.08313656, 0.02447557, 0.02772588, 
    0.06628413, 0.04224896, 0.04746641, -3.005894e-05, 0.173249, 0.01456827, 
    0.01867042, 0.06807495, 0.05965408, 0.04110552, -1.011827e-05, 
    9.868538e-07,
  7.795921e-07, 0.06706014, 0.1350748, 0.05773382, 0.0998802, 0.03689077, 
    -0.001919334, 0.003278364, 0.07855311, 0.2209461, 0.1717143, 0.2060823, 
    0.1981149, 0.2115065, 0.1619044, 0.1539798, 0.1324491, 0.1788603, 
    0.06263842, 0.01721648, 0.04663508, 0.123476, 0.1533866, 0.108549, 
    0.0816325, 0.08445606, 0.0722437, 0.04546645, -3.408522e-06,
  0.1657054, 0.03392401, 0.05316941, 0.257565, 0.1251146, 0.09290735, 
    0.2308483, 0.003079718, 0.03016962, 0.1217493, 0.08863297, 0.2273462, 
    0.2548338, 0.2419868, 0.2681042, 0.2460077, 0.1931957, 0.186369, 
    0.1007273, 0.08511125, 0.1940713, 0.1099461, 0.1716316, 0.1420452, 
    0.3209447, 0.3073399, 0.2478187, 0.148143, 0.1662175,
  0.1069198, 0.08092932, 0.1209229, 0.2122665, 0.2256293, 0.3107896, 
    0.1268028, 0.08076336, 0.02207177, 0.009131077, 0.02509205, 0.03843004, 
    0.1601178, 0.3711242, 0.3278357, 0.2073204, 0.2329182, 0.2982076, 
    0.232301, 0.27025, 0.2165653, 0.1033182, 0.2770767, 0.2662672, 0.2474753, 
    0.375283, 0.2663077, 0.2051922, 0.1162498,
  0.2142702, 0.1489903, 0.1995514, 0.2482979, 0.4204883, 0.2957554, 
    0.5043837, 0.5812588, 0.3424985, 0.3222851, 0.2769104, 0.1033866, 
    0.2184613, 0.2853831, 0.3163905, 0.3026889, 0.3991634, 0.3838725, 
    0.3018275, 0.2730006, 0.08555239, 0.1342163, 0.2160359, 0.2978887, 
    0.2684569, 0.3985579, 0.2885207, 0.324026, 0.2908537,
  0.2878121, 0.2729532, 0.3208118, 0.2646142, 0.2422362, 0.1994287, 0.303403, 
    0.4947948, 0.3129688, 0.4606631, 0.3710621, 0.2981105, 0.2097237, 
    0.2695605, 0.3964536, 0.2237324, 0.2604508, 0.1745871, 0.07626222, 
    0.08711193, 0.122413, 0.1697192, 0.1589262, 0.02514514, 0.08393119, 
    0.5098748, 0.4348232, 0.3261114, 0.2997321,
  0.1235157, 0.2595346, 0.3440845, 0.3798048, 0.1764814, 0.2036422, 
    0.3515548, 0.3939045, 0.3916779, 0.3286772, 0.2761964, 0.3435112, 
    0.3274551, 0.2371792, 0.1786509, 0.1616499, 0.1747425, 0.1213108, 
    0.1479862, 0.1853461, 0.1495677, 0.1175821, 0.1705501, 0.1089721, 
    0.07579946, 0.05402843, 0.111891, 0.2135006, 0.1799646,
  0.2345039, 0.2399323, 0.2453607, 0.250789, 0.2562174, 0.2616458, 0.2670741, 
    0.2644005, 0.2851658, 0.3059312, 0.3266965, 0.3474618, 0.3682272, 
    0.3889925, 0.4050315, 0.3923219, 0.3796121, 0.3669025, 0.3541928, 
    0.3414831, 0.3287734, 0.3093756, 0.2958916, 0.2824076, 0.2689236, 
    0.2554396, 0.2419555, 0.2284715, 0.2301612,
  0.275351, 0.2403952, 0.3546252, 0.4591104, 0.1895719, 0.08913073, 
    0.1647563, 0.1879506, 0.2730716, 0.3857879, 0.3716697, 0.3735576, 
    0.3867072, 0.1091236, 0.1111318, 0.09984504, 0.1855656, 0.06482223, 
    0.02123357, 0.07911049, 0.3703596, 0.3394849, 0.1374745, 0.06884509, 
    0.04537233, 0.142735, 0.1111424, 0.1221529, 0.221373,
  0.3466717, 0.3999205, 0.3567941, 0.3897966, 0.2656278, 0.02330213, 
    0.1639265, 0.2072408, 0.3433965, 0.3622028, 0.3602348, 0.2271084, 
    0.2563413, 0.3011894, 0.3860074, 0.4538606, 0.4484913, 0.4404669, 
    0.3602581, 0.1954312, 0.2386528, 0.3997161, 0.4187092, 0.4155176, 
    0.3333392, 0.3817292, 0.3565941, 0.4750986, 0.5357282,
  0.461391, 0.398806, 0.3912829, 0.4012905, 0.3937734, 0.4575639, 0.3726374, 
    0.2826753, 0.322386, 0.3941547, 0.3736648, 0.4468741, 0.4291036, 
    0.4134375, 0.3504045, 0.3009553, 0.3560863, 0.3812652, 0.4223593, 
    0.3808044, 0.3729859, 0.3013629, 0.3404709, 0.4469406, 0.3212422, 
    0.3969672, 0.4407978, 0.4593763, 0.4348559,
  0.3785585, 0.3188383, 0.2920514, 0.2819181, 0.200055, 0.154576, 0.1418338, 
    0.2075771, 0.3077109, 0.3918186, 0.3619638, 0.3161544, 0.2583277, 
    0.1580263, 0.1637072, 0.1512481, 0.1727997, 0.2518533, 0.3265719, 
    0.2961653, 0.2808641, 0.2968982, 0.2374558, 0.1738735, 0.02775946, 
    0.1101635, 0.1469911, 0.1942459, 0.3119772,
  0.1860649, 0.1909009, 0.2204148, 0.1873895, 0.1094612, 0.2016633, 
    0.1243581, 0.2128757, 0.1894418, 0.2019652, 0.1831292, 0.08349593, 
    0.06285051, 0.0696518, 0.2153099, 0.1261411, 0.0633295, 0.1668262, 
    0.1746902, 0.1852523, 0.1671546, 0.149077, 0.1247794, 0.006327257, 
    0.007392642, 0.1037735, 0.1384083, 0.1352425, 0.1563397,
  0.07946367, 0.01692083, 0.1224162, 0.07825299, 0.07896563, 0.09735765, 
    0.04429901, 0.05753808, 0.05744095, 0.009850835, 0.02732426, 0.01200281, 
    0.004595865, 0.1330428, 0.2496137, 0.1202979, 0.1188749, 0.13998, 
    0.03354298, 0.04366662, 0.05103504, 0.06518393, 0.05964213, 0.0001583635, 
    0.01130955, 0.1504904, 0.03590421, 0.04358122, 0.09045223,
  0.07604458, 0.02225774, 0.07792734, 0.02725914, 0.0693514, 0.02702453, 
    0.04246328, 0.06909654, 0.04196832, 0.008075054, 0.1031648, 0.02695862, 
    0.04246139, 0.04128973, 0.03914496, 0.05818189, 0.05654632, 0.02271021, 
    0.02751945, 0.02983394, 0.05253992, 0.2137656, 0.02571052, -1.697278e-05, 
    0.08692097, 0.2780607, 0.03163374, 0.04744337, 0.07661963,
  0.01802406, 0.007269382, 0.1470029, 0.06762385, 0.02222201, 0.02278677, 
    0.02930987, 0.03664131, 0.05939346, 0.02557377, 0.02350461, 0.02037682, 
    0.07462071, 0.04043935, 0.0952865, 0.04283029, 0.02302252, 0.0235022, 
    0.02746722, 0.03209742, 0.02694404, 0.01771379, 0.03256745, 0.1036008, 
    0.1094304, 0.08723335, 0.0345005, 0.04719197, 0.05329077,
  0.003019127, 0.01027714, 0.00218733, 0.03157439, 0.07583717, 0.05903589, 
    0.08338501, 0.1274765, 0.1626263, 0.1475401, 0.02412946, 0.02179725, 
    0.02410144, 0.03378376, 0.06049712, 0.03533319, 0.008882089, 0.01274949, 
    0.01940172, 0.02318719, 0.03859859, 0.02957085, 0.05941099, 0.03635101, 
    0.1263674, 0.1623593, 0.0301477, 0.02320695, 0.002123638,
  1.327513e-09, 1.332704e-09, 6.919432e-09, 0.0166006, 0.07516789, 
    0.03984669, 0.00185527, 0.01286623, 0.01568318, 0.07547003, 0.1875285, 
    0.053245, 0.0523472, 0.04218335, 0.04270868, 0.04823651, 0.04771838, 
    0.123023, 0.1398701, 0.131503, 0.06671833, 0.01584434, 0.08241111, 
    0.02360957, 0.03446066, 0.02051431, 0.0005944714, 1.500068e-08, 
    -1.252649e-06,
  3.436981e-07, 2.980174e-09, -6.863463e-07, 0.00655228, 3.493533e-05, 
    0.01415218, 7.185895e-10, 0.0005040851, 0.004860761, 0.1214662, 
    0.2688081, 0.1091306, 0.07032828, 0.1365557, 0.1211241, 0.05247117, 
    0.04569726, 0.07907942, 0.07914124, 0.09026241, 0.01408935, 0.2225046, 
    0.02215295, 0.01335948, 0.08068117, 0.1250364, 0.08302685, -4.015623e-05, 
    4.596944e-07,
  -2.352629e-05, 0.08622339, 0.2182749, 0.05780563, 0.09913471, 0.026768, 
    -0.001867717, 0.001381121, 0.07149331, 0.1884343, 0.2434204, 0.2208131, 
    0.2001142, 0.2209722, 0.1513974, 0.2194344, 0.1498182, 0.1939977, 
    0.08406404, 0.0214952, 0.053286, 0.1590724, 0.142534, 0.142057, 
    0.1260946, 0.1607226, 0.09183418, 0.06162431, -9.227498e-05,
  0.1986829, 0.04920429, 0.08790161, 0.3093762, 0.1738559, 0.04595319, 
    0.2131439, 0.0005953843, 0.03565359, 0.123171, 0.07943451, 0.2466171, 
    0.3487221, 0.2262972, 0.2503336, 0.2426358, 0.2369385, 0.2429761, 
    0.1488673, 0.09296658, 0.1985989, 0.1037044, 0.1663483, 0.1719267, 
    0.4171055, 0.3281004, 0.2395908, 0.1756259, 0.1602742,
  0.1038529, 0.08233849, 0.1405992, 0.2553152, 0.3046585, 0.3617571, 
    0.1232819, 0.08045359, 0.01748162, 0.007815924, 0.03502615, 0.03842206, 
    0.2554614, 0.3581285, 0.278039, 0.2338655, 0.2349419, 0.3268525, 
    0.257547, 0.2696523, 0.1912956, 0.1052232, 0.2742209, 0.2747969, 
    0.3015759, 0.4141057, 0.244175, 0.2143386, 0.1472581,
  0.2436337, 0.1563157, 0.1705869, 0.2881347, 0.404844, 0.3224058, 0.5044754, 
    0.5657308, 0.4146661, 0.4238203, 0.3206593, 0.1035458, 0.172242, 
    0.3610649, 0.3357615, 0.3175278, 0.4224298, 0.4020047, 0.3379653, 
    0.1995593, 0.08867832, 0.1615878, 0.245942, 0.3016597, 0.4015622, 
    0.3587611, 0.2310607, 0.3248141, 0.305714,
  0.3899667, 0.2240417, 0.3320851, 0.32081, 0.2644115, 0.1982362, 0.3765815, 
    0.5126579, 0.3239951, 0.4849828, 0.4575119, 0.3217171, 0.2244048, 
    0.3276667, 0.3955232, 0.2176666, 0.2464842, 0.1613999, 0.07942921, 
    0.1381432, 0.1469329, 0.2130029, 0.1789276, 0.02959545, 0.06966773, 
    0.5074318, 0.4581316, 0.3327752, 0.3221068,
  0.1388243, 0.2707255, 0.381422, 0.3848498, 0.1446373, 0.2150835, 0.3676345, 
    0.4380898, 0.4335451, 0.3955586, 0.332688, 0.3702878, 0.3687583, 
    0.2924497, 0.1991005, 0.1882014, 0.1836472, 0.170436, 0.1853808, 
    0.2033902, 0.1685762, 0.135628, 0.1753877, 0.1184826, 0.07239052, 
    0.04535471, 0.1080528, 0.2011702, 0.1930323,
  0.230301, 0.235682, 0.241063, 0.246444, 0.2518249, 0.2572059, 0.2625869, 
    0.2785393, 0.3016201, 0.3247009, 0.3477817, 0.3708625, 0.3939433, 
    0.4170241, 0.4423902, 0.4298896, 0.417389, 0.4048884, 0.3923878, 
    0.3798872, 0.3673865, 0.3296242, 0.313663, 0.2977018, 0.2817406, 
    0.2657795, 0.2498183, 0.2338571, 0.2259962,
  0.3093794, 0.2580776, 0.3560147, 0.4746858, 0.1961635, 0.08612974, 
    0.2024786, 0.2411069, 0.3440909, 0.4198003, 0.4004832, 0.3923487, 
    0.4001745, 0.1190764, 0.07545539, 0.07887165, 0.118582, 0.09916868, 
    0.02914973, 0.06330005, 0.3386881, 0.307215, 0.1125996, 0.1306986, 
    0.05768783, 0.2430792, 0.1328254, 0.1712893, 0.3027215,
  0.34757, 0.3911003, 0.3666564, 0.3268484, 0.2571579, 0.02965131, 0.183892, 
    0.2232806, 0.3390239, 0.3771893, 0.3526069, 0.1939812, 0.246903, 
    0.2522976, 0.3861637, 0.4008945, 0.357204, 0.4103161, 0.4573822, 
    0.3642313, 0.3303354, 0.5137516, 0.4426762, 0.451725, 0.3748281, 
    0.4259379, 0.4792793, 0.4971377, 0.548781,
  0.4603663, 0.4255019, 0.4829684, 0.5013097, 0.5067661, 0.5061486, 
    0.4348188, 0.3665614, 0.3669604, 0.3671064, 0.3477128, 0.4703843, 
    0.504297, 0.4812202, 0.3927546, 0.3841272, 0.4467555, 0.4919127, 
    0.519546, 0.3547271, 0.3848967, 0.2949183, 0.3827246, 0.5030161, 
    0.4407312, 0.535729, 0.4460028, 0.5830718, 0.549078,
  0.4140382, 0.3316692, 0.3391183, 0.325156, 0.2765676, 0.2177674, 0.1966707, 
    0.3002979, 0.3196916, 0.3944634, 0.3018721, 0.3542958, 0.2884272, 
    0.3033038, 0.2539834, 0.2283707, 0.327601, 0.3158913, 0.2792622, 
    0.2978899, 0.2456325, 0.3194575, 0.3387749, 0.1720905, 0.01639082, 
    0.1353945, 0.19566, 0.293436, 0.4343463,
  0.2542576, 0.3006525, 0.2680289, 0.3037593, 0.2423707, 0.3318027, 
    0.2243404, 0.3505677, 0.2963017, 0.2786482, 0.1698413, 0.1558599, 
    0.06621185, 0.1472114, 0.2415195, 0.221628, 0.2070901, 0.353492, 
    0.2852945, 0.2200304, 0.1972013, 0.1752016, 0.1954704, 0.005973586, 
    0.05038653, 0.1354315, 0.1710587, 0.1914198, 0.240573,
  0.1317626, 0.07122124, 0.1270088, 0.1347696, 0.07652482, 0.09592248, 
    0.05907954, 0.1488335, 0.2186699, 0.001736445, 0.02732575, 0.01058154, 
    0.003763069, 0.1211139, 0.2887027, 0.1444527, 0.1169479, 0.1560091, 
    0.0370173, 0.0810623, 0.05428481, 0.1051355, 0.1973305, 0.0002418547, 
    0.0064667, 0.1572533, 0.05858662, 0.0649401, 0.1473596,
  0.1747932, 0.02373169, 0.05919905, 0.04786552, 0.06137799, 0.03893134, 
    0.06559501, 0.08550859, 0.1394738, 0.01306791, 0.08872107, 0.01937896, 
    0.0526449, 0.05708981, 0.03335215, 0.07241448, 0.06549688, 0.02835897, 
    0.04104966, 0.04071576, 0.05514555, 0.1675052, 0.3168733, -0.000177086, 
    0.0589397, 0.2808603, 0.07887835, 0.05115695, 0.09734219,
  0.06032987, 0.01589952, 0.1185733, 0.05938278, 0.02975224, 0.03314845, 
    0.03806801, 0.06716517, 0.08414954, 0.03205721, 0.02946233, 0.02511656, 
    0.06115501, 0.04684547, 0.07929889, 0.05191019, 0.03171822, 0.04171832, 
    0.04935044, 0.05385581, 0.0675005, 0.07898936, 0.1021752, 0.09277286, 
    0.08883407, 0.0617864, 0.04984106, 0.05782108, 0.1018267,
  0.003663375, 0.008744889, 0.001220853, 0.03073744, 0.07489888, 0.05427859, 
    0.07059509, 0.1060534, 0.1883896, 0.1397636, 0.03202803, 0.03088737, 
    0.0288908, 0.03922708, 0.06146659, 0.0371803, 0.009085702, 0.008190845, 
    0.018889, 0.02055255, 0.03159392, 0.03121474, 0.03863871, 0.0230645, 
    0.1106408, 0.1078191, 0.03241495, 0.037834, 0.004461303,
  6.858252e-10, 2.951505e-10, 1.356087e-09, 0.003547688, 0.07868443, 
    0.1220492, 0.001650369, 0.09281086, 0.008946273, 0.09098695, 0.1809273, 
    0.05131938, 0.07034206, 0.03891675, 0.04869445, 0.07082064, 0.05449049, 
    0.1273691, 0.140212, 0.1277564, 0.05659049, 0.02970959, 0.09050581, 
    0.02105841, 0.0491907, 0.1883694, 0.008862419, 4.901808e-09, -1.160473e-06,
  8.772252e-08, 1.53384e-09, -8.888085e-06, 0.001251883, -2.949745e-06, 
    0.01805962, 4.005407e-10, 0.0003779379, 0.001914158, 0.2079267, 
    0.3241558, 0.1418241, 0.1039786, 0.1367543, 0.1743166, 0.148596, 
    0.1044056, 0.087101, 0.1676925, 0.2445166, 0.002263136, 0.2669581, 
    0.03976387, 0.02216823, 0.06146337, 0.0982435, 0.1232731, -0.0001011308, 
    2.954706e-07,
  -7.373324e-06, 0.07022467, 0.1402931, 0.05900273, 0.09623262, 0.02061388, 
    -0.001701553, 0.0007476647, 0.06318184, 0.2149247, 0.2343136, 0.1573512, 
    0.140376, 0.1704519, 0.1659323, 0.1979474, 0.1726899, 0.2405546, 
    0.1857914, 0.02059532, 0.05538356, 0.2293932, 0.1508539, 0.1491169, 
    0.129732, 0.1957499, 0.1223488, 0.135653, -0.0003352854,
  0.2455768, 0.08526456, 0.1093159, 0.3539207, 0.1568056, 0.03590317, 
    0.1916885, -6.993463e-05, 0.04392616, 0.1148416, 0.08480853, 0.2475785, 
    0.2730056, 0.1669793, 0.1811569, 0.2352331, 0.2870669, 0.2899626, 
    0.1973139, 0.09304111, 0.2094556, 0.1167123, 0.1911537, 0.2070229, 
    0.3401652, 0.2694131, 0.2097526, 0.1965346, 0.1635012,
  0.1575262, 0.1194136, 0.1647356, 0.2798133, 0.3779614, 0.3670461, 
    0.1332092, 0.08146121, 0.01395918, 0.008759887, 0.0348059, 0.0425668, 
    0.3200609, 0.2504388, 0.2185525, 0.2083394, 0.314926, 0.3323112, 
    0.2280513, 0.2848457, 0.2040062, 0.1769239, 0.3079443, 0.3011467, 
    0.378356, 0.3478865, 0.206241, 0.2809084, 0.1699595,
  0.2745025, 0.141554, 0.1688663, 0.358944, 0.4542896, 0.3427795, 0.5022284, 
    0.5421427, 0.4462906, 0.4750244, 0.3747569, 0.12601, 0.1289682, 
    0.3419358, 0.4778328, 0.2747663, 0.4640497, 0.4112178, 0.3639902, 
    0.1518403, 0.1159191, 0.1882263, 0.2657855, 0.3448111, 0.6175634, 
    0.2930499, 0.1705034, 0.297033, 0.3077994,
  0.3538164, 0.2389627, 0.3079335, 0.3090862, 0.3174416, 0.2420262, 
    0.4007234, 0.5387552, 0.330883, 0.5214974, 0.5672894, 0.3730972, 
    0.2431876, 0.335797, 0.4131648, 0.2592505, 0.2424149, 0.1936809, 
    0.09455722, 0.1483296, 0.1374467, 0.2450887, 0.207089, 0.03512542, 
    0.0566569, 0.4698935, 0.476808, 0.3423799, 0.36766,
  0.1636756, 0.2966236, 0.3982019, 0.3782843, 0.2431686, 0.325802, 0.4396814, 
    0.4822147, 0.4981097, 0.4647757, 0.3993056, 0.3927571, 0.4107639, 
    0.3475308, 0.2455202, 0.2653745, 0.2148389, 0.220016, 0.2367919, 
    0.2419546, 0.189891, 0.1706168, 0.1946239, 0.1133591, 0.07732175, 
    0.03873824, 0.08996958, 0.1855167, 0.2298289,
  0.254095, 0.2581178, 0.2621406, 0.2661634, 0.2701863, 0.2742091, 0.2782319, 
    0.2864665, 0.3091934, 0.3319203, 0.3546472, 0.3773741, 0.4001009, 
    0.4228278, 0.4433235, 0.4298043, 0.416285, 0.4027658, 0.3892465, 
    0.3757273, 0.362208, 0.3359456, 0.3227151, 0.3094847, 0.2962542, 
    0.2830238, 0.2697933, 0.2565629, 0.2508768,
  0.4140086, 0.3246003, 0.3688025, 0.5145157, 0.2081046, 0.09048621, 
    0.2153872, 0.2931584, 0.3914036, 0.4584728, 0.4201387, 0.394087, 
    0.4121762, 0.09897739, 0.0757194, 0.1032707, 0.1613713, 0.138814, 
    0.05351537, 0.05263087, 0.3418684, 0.3466946, 0.1300058, 0.1581767, 
    0.07560217, 0.2402341, 0.08914563, 0.2071088, 0.3388495,
  0.3484689, 0.3693139, 0.336657, 0.2573736, 0.2459712, 0.03679253, 0.163555, 
    0.259643, 0.3930796, 0.4105173, 0.3591991, 0.1489691, 0.1998407, 
    0.2278369, 0.3056452, 0.3654387, 0.332441, 0.3821616, 0.4318691, 
    0.4009095, 0.3989268, 0.4820634, 0.51035, 0.472369, 0.2763019, 0.4563543, 
    0.3605464, 0.4148754, 0.4621173,
  0.4568111, 0.4183536, 0.489913, 0.5888364, 0.5525717, 0.5302916, 0.4513475, 
    0.3769682, 0.3649183, 0.2924559, 0.3575034, 0.499587, 0.5280266, 
    0.5353179, 0.4217254, 0.4547464, 0.4806765, 0.5504578, 0.4823028, 
    0.3146703, 0.3430251, 0.3083694, 0.463389, 0.4957792, 0.5275975, 
    0.4741333, 0.5097255, 0.5678632, 0.5177619,
  0.3919688, 0.3446676, 0.4090163, 0.3621845, 0.3596453, 0.3239468, 
    0.3479246, 0.3090053, 0.3243313, 0.3724262, 0.2872784, 0.4132791, 
    0.3246416, 0.3282227, 0.2971099, 0.4351376, 0.4167533, 0.3693357, 
    0.2481358, 0.2660103, 0.2463876, 0.3613569, 0.3489888, 0.1825006, 
    0.01359534, 0.1468497, 0.3431015, 0.4410771, 0.4613517,
  0.3606768, 0.2532984, 0.2038909, 0.3588455, 0.3517207, 0.3271519, 
    0.2925364, 0.3537275, 0.3990682, 0.314324, 0.2423004, 0.1642, 0.06809386, 
    0.2401086, 0.2580263, 0.3640022, 0.3194917, 0.3100933, 0.2827516, 
    0.268539, 0.2453149, 0.1592501, 0.3507749, 0.007800578, 0.02839836, 
    0.2149528, 0.217215, 0.2578227, 0.2989281,
  0.1241877, 0.1260396, 0.1095619, 0.1268044, 0.1106217, 0.09408194, 
    0.1091813, 0.1958845, 0.2418444, 0.007883427, 0.04398009, 0.01511379, 
    0.003386403, 0.0941088, 0.3081947, 0.1423807, 0.1221844, 0.2110951, 
    0.1188462, 0.06022499, 0.1642132, 0.1443384, 0.3040334, 0.0008980179, 
    0.002129414, 0.1696937, 0.04721079, 0.07777949, 0.1734466,
  0.27009, 0.03279832, 0.03519985, 0.1408362, 0.05821236, 0.0765924, 
    0.07152079, 0.07197112, 0.2366642, 0.05889845, 0.06747734, 0.01000236, 
    0.03543411, 0.06819022, 0.08210662, 0.08343007, 0.08403576, 0.06188913, 
    0.04136541, 0.04024213, 0.04167507, 0.08801458, 0.4386512, 0.0007656962, 
    0.03667606, 0.2769933, 0.05110701, 0.03386367, 0.07080858,
  0.1983892, 0.0953275, 0.07742319, 0.05673862, 0.07682328, 0.1073866, 
    0.1143238, 0.07026234, 0.167205, 0.05531608, 0.03699942, 0.03589821, 
    0.04718826, 0.05115408, 0.1129564, 0.08458994, 0.03614838, 0.05037307, 
    0.06167236, 0.06024972, 0.09413925, 0.1492315, 0.1745065, 0.05782371, 
    0.06616542, 0.04161571, 0.06265136, 0.09036272, 0.1891397,
  0.0596418, 0.005937821, 0.0005073372, 0.02258413, 0.06916677, 0.05496275, 
    0.1370712, 0.07627476, 0.1362178, 0.1170346, 0.04777069, 0.07617087, 
    0.1218262, 0.041844, 0.06716423, 0.06264833, 0.01781736, 0.008831151, 
    0.02495226, 0.02110335, 0.03388685, 0.03736006, 0.03093785, 0.009565186, 
    0.0665374, 0.1163339, 0.03975942, 0.08794789, 0.07895899,
  4.720849e-10, 1.091861e-10, 2.78372e-10, -0.001546519, 0.09536068, 
    0.1270757, 0.0005314762, 0.09457956, 0.006246936, 0.1081547, 0.1771999, 
    0.04526598, 0.03585386, 0.05028293, 0.07686803, 0.06915387, 0.1266914, 
    0.121081, 0.1450364, 0.1148217, 0.06436519, 0.07760146, 0.1523145, 
    0.03576636, 0.02108913, 0.06288547, 0.2918626, -2.640802e-06, 
    -1.053442e-06,
  2.65515e-08, 7.553596e-10, -5.027935e-06, 0.0004222326, -3.572735e-07, 
    0.01242629, 3.081866e-10, 0.0009689921, 0.001015307, 0.3478617, 
    0.2725324, 0.07965801, 0.09824938, 0.1167568, 0.1309306, 0.06394985, 
    0.05928679, 0.08093126, 0.08837435, 0.1940119, 0.01123729, 0.2750632, 
    0.07709092, 0.01808382, 0.0314044, 0.0648881, 0.1497411, 0.004914425, 
    2.380419e-07,
  -1.626647e-06, 0.07311729, 0.05900552, 0.06301476, 0.08770059, 0.01344679, 
    -0.001504377, 0.000459235, 0.04273286, 0.2074319, 0.1853077, 0.1081191, 
    0.1201482, 0.1306152, 0.1794991, 0.1811574, 0.2224841, 0.2776691, 
    0.1588394, 0.04282625, 0.06365348, 0.2478854, 0.1761189, 0.1441664, 
    0.2327171, 0.1619722, 0.06583425, 0.1486672, -0.0003533119,
  0.2241019, 0.04868951, 0.0936962, 0.3895977, 0.09950173, 0.02788975, 
    0.1763381, -0.0001718564, 0.03080753, 0.08837255, 0.1088263, 0.1520528, 
    0.1368153, 0.1384446, 0.1272751, 0.2179124, 0.3067999, 0.2827596, 
    0.1675147, 0.1046357, 0.215146, 0.1044396, 0.2340973, 0.232194, 
    0.2598952, 0.2340661, 0.2069718, 0.2101078, 0.1739631,
  0.2500759, 0.1481755, 0.2145531, 0.3139443, 0.4980449, 0.3583786, 
    0.1287159, 0.08481936, 0.01291267, 0.01253544, 0.02796749, 0.03861891, 
    0.3868011, 0.1464205, 0.1808879, 0.1871897, 0.2848807, 0.3466005, 
    0.2128413, 0.3180904, 0.1937106, 0.2671838, 0.2859792, 0.3396144, 
    0.4332663, 0.2309298, 0.178533, 0.2200876, 0.337483,
  0.3404315, 0.1455718, 0.195854, 0.4428053, 0.4936381, 0.3229996, 0.5326422, 
    0.5400578, 0.4273018, 0.4923462, 0.4052975, 0.1820965, 0.1160734, 
    0.2515391, 0.5636244, 0.2935624, 0.4766549, 0.4142682, 0.3484923, 
    0.1869218, 0.1768158, 0.2106195, 0.2869495, 0.3344067, 0.7397031, 
    0.209599, 0.1516391, 0.2858219, 0.2680706,
  0.2563853, 0.1894166, 0.3251152, 0.2609755, 0.3425753, 0.3106105, 
    0.4548398, 0.5485936, 0.3475819, 0.5620475, 0.6169849, 0.3815328, 
    0.2514887, 0.3656741, 0.4819729, 0.2839436, 0.2996488, 0.2089705, 
    0.09467722, 0.1723083, 0.1171096, 0.2752192, 0.2361321, 0.04181465, 
    0.05109954, 0.4216274, 0.49582, 0.3432833, 0.3449372,
  0.2428768, 0.3572987, 0.4054381, 0.3738754, 0.3163123, 0.3932588, 
    0.5277226, 0.5601346, 0.5960912, 0.5156776, 0.4650125, 0.3996422, 
    0.4572142, 0.4347047, 0.2857367, 0.3429678, 0.2867692, 0.2522779, 
    0.2736109, 0.3082433, 0.2576197, 0.2024469, 0.1931832, 0.1027509, 
    0.08392263, 0.0371975, 0.07844389, 0.1801654, 0.2709882,
  0.2995879, 0.3040421, 0.3084962, 0.3129504, 0.3174045, 0.3218587, 
    0.3263128, 0.3550571, 0.3767049, 0.3983527, 0.4200005, 0.4416482, 
    0.463296, 0.4849438, 0.4962378, 0.4801895, 0.4641411, 0.4480927, 
    0.4320444, 0.415996, 0.3999476, 0.3835415, 0.373488, 0.3634344, 
    0.3533809, 0.3433273, 0.3332737, 0.3232202, 0.2960246,
  0.4318767, 0.4084997, 0.4479497, 0.5724508, 0.2153327, 0.1015488, 
    0.2368651, 0.3438516, 0.4668736, 0.4784752, 0.4868489, 0.4338696, 
    0.4724007, 0.07988884, 0.07571665, 0.1751399, 0.2142976, 0.2055379, 
    0.1196021, 0.04991034, 0.4141198, 0.4015514, 0.1683446, 0.1754162, 
    0.2000363, 0.3239364, 0.05399354, 0.2082555, 0.2829373,
  0.3230177, 0.2838615, 0.3068804, 0.1957815, 0.1973367, 0.02698017, 
    0.1152371, 0.2360236, 0.3991003, 0.3918134, 0.3332161, 0.1356956, 
    0.1451007, 0.1863379, 0.2353215, 0.3243813, 0.2917512, 0.3458295, 
    0.4035098, 0.2949244, 0.4105923, 0.4295237, 0.5492354, 0.4130411, 
    0.2020532, 0.3426979, 0.3161246, 0.3027482, 0.3471563,
  0.4788278, 0.4625606, 0.4646475, 0.5972314, 0.5770901, 0.5707906, 
    0.5052502, 0.3459864, 0.2924032, 0.2052294, 0.336569, 0.4966929, 
    0.5111922, 0.5302869, 0.4244777, 0.4421483, 0.4910757, 0.544699, 
    0.3987803, 0.2701834, 0.3013954, 0.3284824, 0.4045626, 0.4748706, 
    0.5273308, 0.4353321, 0.5400689, 0.5019299, 0.47185,
  0.3912909, 0.3557621, 0.465978, 0.3973198, 0.3757676, 0.3783343, 0.3490308, 
    0.3637195, 0.3513886, 0.3519155, 0.2559997, 0.3562315, 0.2637413, 
    0.2926502, 0.3560853, 0.4324951, 0.3888249, 0.3099568, 0.2563628, 
    0.2144386, 0.2233077, 0.3768482, 0.3808252, 0.1836618, 0.01192938, 
    0.1667567, 0.3810976, 0.4100539, 0.4446953,
  0.2305669, 0.1942808, 0.1264697, 0.2985568, 0.2808496, 0.322199, 0.3099325, 
    0.3384024, 0.3946586, 0.2377117, 0.1689191, 0.09779387, 0.03699037, 
    0.1645926, 0.2876636, 0.2384185, 0.1701362, 0.3121907, 0.2602921, 
    0.1839323, 0.2537801, 0.2738232, 0.3613578, 0.007565084, 0.01136241, 
    0.2986892, 0.3130032, 0.2761828, 0.2475727,
  0.1018131, 0.0885704, 0.09523983, 0.09842239, 0.08777851, 0.08221731, 
    0.08150972, 0.1355477, 0.2265979, 0.007587658, 0.04001125, 0.01850091, 
    0.0043098, 0.04079939, 0.2870765, 0.1334021, 0.1095858, 0.1252407, 
    0.1012206, 0.01997588, 0.1649935, 0.03703556, 0.1537148, 0.005307129, 
    0.0006054484, 0.1371922, 0.03172534, 0.04215103, 0.09223216,
  0.1101303, 0.05199654, 0.0146739, 0.0274975, 0.06151843, 0.01998952, 
    0.0578823, 0.02507237, 0.1703258, 0.06723024, 0.05412209, 0.003763332, 
    0.008405012, 0.02845788, 0.04335178, 0.06556501, 0.08330484, 0.01616019, 
    0.007211626, 0.007280847, 0.008144636, 0.04164891, 0.2233317, 0.1601069, 
    0.02661438, 0.2741748, 0.03356733, 0.01897184, 0.0183447,
  0.2386498, 0.1176972, 0.05368677, 0.05851735, 0.1004535, 0.08520206, 
    0.02144195, 0.01883223, 0.05226653, 0.07676467, 0.03049455, 0.02388459, 
    0.03008962, 0.02896581, 0.08282924, 0.0246671, 0.01271269, 0.01363442, 
    0.01318514, 0.01658247, 0.02929387, 0.0580233, 0.1557745, 0.03069662, 
    0.05856787, 0.02761344, 0.02871232, 0.07506943, 0.1534564,
  0.0112005, 0.005697143, 0.0002537667, 0.01382922, 0.07627165, 0.05287553, 
    0.08060896, 0.07608154, 0.08539464, 0.09612645, 0.04574159, 0.03577083, 
    0.02757769, 0.03500982, 0.05368797, 0.02986243, 0.02667518, 0.0146079, 
    0.0325649, 0.02917692, 0.06643479, 0.1591451, 0.05511481, 0.002566259, 
    0.03758745, 0.1197893, 0.03089588, 0.01773041, 0.07314479,
  3.946848e-10, 7.956982e-11, 2.127394e-10, -0.003669755, 0.1065495, 
    0.03158816, -5.410553e-05, 0.02604086, 0.002701218, 0.1030715, 0.1542539, 
    0.02390393, 0.0131064, 0.02373616, 0.02254265, 0.02021068, 0.061235, 
    0.1212168, 0.1286694, 0.08647768, 0.04827467, 0.0514832, 0.3600969, 
    0.08360727, 0.003613355, 0.01833193, 0.1330671, -0.0001608605, 
    -8.562846e-07,
  1.562478e-08, 3.52317e-10, -4.718069e-06, 2.511757e-05, -1.046594e-07, 
    0.01112455, 2.799118e-10, 0.001883152, 0.0009780251, 0.3111982, 0.217218, 
    0.05536985, 0.02394373, 0.04933434, 0.07573385, 0.03232242, 0.02028847, 
    0.06717828, 0.02565093, 0.1163619, 0.01200326, 0.2462076, 0.02718237, 
    0.004046448, 0.004895201, 0.01023134, 0.07638842, 0.001031305, 
    2.110093e-07,
  -4.628318e-07, 0.0598767, 0.02082381, 0.05005033, 0.07757998, 0.0103959, 
    -0.001352983, 0.0002744918, 0.02651432, 0.2505586, 0.1536884, 0.06172618, 
    0.08395689, 0.1225406, 0.1394433, 0.1557461, 0.2046685, 0.1943842, 
    0.07375807, 0.01644806, 0.06145605, 0.2284219, 0.1792141, 0.2239129, 
    0.2607615, 0.1290377, 0.1332208, 0.1289677, -0.0002052795,
  0.178748, 0.0166783, 0.0731015, 0.4326276, 0.05279089, 0.03480764, 
    0.1705111, -0.000105453, 0.01578356, 0.09212039, 0.1169951, 0.1041689, 
    0.09321644, 0.1217489, 0.1015101, 0.1864089, 0.34054, 0.338535, 
    0.1567809, 0.1066333, 0.2128824, 0.110308, 0.2657314, 0.188577, 
    0.2215053, 0.202898, 0.2140578, 0.1325557, 0.173722,
  0.2726482, 0.1925616, 0.2586386, 0.2892914, 0.4622398, 0.2782089, 
    0.1030442, 0.09325252, 0.0123455, 0.02520767, 0.0168467, 0.03113616, 
    0.2748161, 0.08597235, 0.1612142, 0.1460665, 0.262177, 0.352486, 
    0.2182591, 0.350632, 0.1725271, 0.2544051, 0.2112154, 0.3796229, 
    0.3813421, 0.1484235, 0.1727505, 0.1930304, 0.2554977,
  0.3386983, 0.1657863, 0.2353296, 0.5003288, 0.5108001, 0.3188989, 
    0.5757405, 0.543285, 0.4061347, 0.4646118, 0.4161299, 0.2550829, 
    0.1254426, 0.1878045, 0.5659661, 0.285462, 0.4779848, 0.4059588, 
    0.3208476, 0.1850863, 0.2736988, 0.2612879, 0.2846275, 0.2748503, 
    0.762177, 0.1474997, 0.1268349, 0.2927827, 0.2345756,
  0.21426, 0.1580264, 0.2659548, 0.1804563, 0.4062016, 0.3264668, 0.5307113, 
    0.5637027, 0.3716289, 0.5761756, 0.650303, 0.3962373, 0.3089572, 
    0.3946764, 0.5337798, 0.3021748, 0.3504339, 0.2400337, 0.1215286, 
    0.2481063, 0.1329733, 0.3116378, 0.2321134, 0.04498259, 0.03810041, 
    0.376589, 0.5069547, 0.3262727, 0.2885262,
  0.2777242, 0.4910058, 0.4299213, 0.4031585, 0.3588076, 0.4658528, 
    0.6120657, 0.6242885, 0.6436254, 0.5790074, 0.546759, 0.4587899, 
    0.4872603, 0.4891547, 0.35999, 0.4207768, 0.3646025, 0.2808625, 
    0.3105688, 0.3845477, 0.3500826, 0.2208561, 0.1850476, 0.1158418, 
    0.1028074, 0.03973061, 0.05527047, 0.1897334, 0.3302908,
  0.358198, 0.3646259, 0.3710538, 0.3774818, 0.3839097, 0.3903376, 0.3967656, 
    0.4189372, 0.437162, 0.4553867, 0.4736115, 0.4918362, 0.510061, 
    0.5282858, 0.5220819, 0.5050768, 0.4880717, 0.4710665, 0.4540614, 
    0.4370563, 0.4200512, 0.41311, 0.4054624, 0.3978148, 0.3901672, 
    0.3825196, 0.374872, 0.3672245, 0.3530557,
  0.4401007, 0.4582294, 0.5569969, 0.6286439, 0.2226892, 0.1343998, 
    0.2533581, 0.4105389, 0.4988115, 0.5245231, 0.5667013, 0.4190443, 
    0.4892358, 0.04938579, 0.1829557, 0.2672449, 0.2550698, 0.1794269, 
    0.1058815, 0.05752437, 0.4348811, 0.4304759, 0.1636076, 0.1462844, 
    0.2012504, 0.2614504, 0.1026741, 0.1843696, 0.2342291,
  0.2508906, 0.2607607, 0.2847385, 0.1221638, 0.1080047, 0.01594561, 
    0.09180559, 0.1744778, 0.309704, 0.3175228, 0.2976894, 0.1378036, 
    0.09668361, 0.1447051, 0.1763451, 0.2893364, 0.2545389, 0.3452069, 
    0.3542156, 0.1951822, 0.3405189, 0.4463572, 0.6542112, 0.3543587, 
    0.2173356, 0.2602822, 0.2518075, 0.2120938, 0.2733696,
  0.4535708, 0.4741339, 0.4365765, 0.5281873, 0.6027136, 0.5849138, 
    0.5006621, 0.3101919, 0.2143523, 0.1615978, 0.2787654, 0.4531425, 
    0.497723, 0.4860561, 0.4115905, 0.4521548, 0.4829661, 0.5476077, 
    0.3346274, 0.2119925, 0.2718926, 0.319551, 0.3548045, 0.4691235, 
    0.5057457, 0.4596962, 0.5160492, 0.4599563, 0.4323939,
  0.3699456, 0.3697237, 0.4879924, 0.4073883, 0.4035669, 0.3539248, 
    0.3853303, 0.3788736, 0.3555755, 0.3241065, 0.2039401, 0.2783539, 
    0.2312045, 0.2675796, 0.3435845, 0.3073746, 0.293525, 0.2158433, 
    0.2005997, 0.1931713, 0.2135995, 0.3439256, 0.395899, 0.169136, 
    0.01462272, 0.2386643, 0.356185, 0.3713492, 0.4162124,
  0.1809797, 0.1273593, 0.07484022, 0.237892, 0.2261409, 0.2511143, 
    0.2623754, 0.34472, 0.3617357, 0.1365163, 0.08938266, 0.052221, 
    0.02903968, 0.09426446, 0.3288317, 0.1985529, 0.08582626, 0.2117855, 
    0.1951949, 0.1361432, 0.2759976, 0.2887304, 0.247932, 0.007818356, 
    0.02589924, 0.250158, 0.4043833, 0.2978349, 0.1938436,
  0.0933515, 0.04973548, 0.0977096, 0.02616834, 0.0544348, 0.04546332, 
    0.02219919, 0.06200007, 0.1547239, 0.001725838, 0.02328956, 0.009957116, 
    0.002591074, 0.01754867, 0.2275389, 0.09959482, 0.09982591, 0.0877686, 
    0.02048952, 0.004398962, 0.05214546, 0.009733799, 0.04182157, 0.06698263, 
    0.0001250169, 0.08710618, 0.01462738, 0.005884887, 0.05340351,
  0.03097833, 0.08649857, 0.01327617, 0.007923734, 0.02331356, 0.002634743, 
    0.0153265, 0.006505896, 0.05686423, 0.06697506, 0.04134881, 0.00115331, 
    0.001257317, 0.01257023, 0.01849084, 0.04235176, 0.03607996, 0.00254006, 
    0.0004434374, 0.0003295354, 0.0004230029, 0.0110467, 0.06358311, 
    0.1010674, 0.01880362, 0.2505699, 0.008067724, 0.007998543, 0.003197114,
  0.05889805, 0.03791016, 0.04606216, 0.04679716, 0.01626162, 0.01058243, 
    0.003171525, 0.001321856, 0.008866713, 0.009855816, 0.008736233, 
    0.003098493, 0.01307717, 0.006723793, 0.07704113, 0.009948803, 
    0.0006153189, 0.001656419, 0.001692759, 0.002013451, 0.005462092, 
    0.009915292, 0.03133148, 0.02029771, 0.04846616, 0.02163347, 0.002205033, 
    0.009666185, 0.0327259,
  0.001393807, 0.007146219, 0.0002848748, 0.008801228, 0.06316901, 
    0.02764403, 0.03139096, 0.0602147, 0.05022945, 0.0756768, 0.00740975, 
    0.003644813, 0.007180318, 0.009294337, 0.02341065, 0.0119903, 
    0.009264322, 0.01950317, 0.01631068, 0.02781747, 0.07207809, 0.2064927, 
    0.1423373, 0.0008280673, 0.02558402, 0.09199328, 0.005310114, 
    0.002117456, 0.01120997,
  3.630014e-10, 7.573296e-11, 2.055832e-10, -0.002420652, 0.08017755, 
    0.008794939, -0.0004896971, 0.00551442, 0.0008878359, 0.06652193, 
    0.1143513, 0.007644762, 0.003719121, 0.006919683, 0.002990899, 
    0.003256076, 0.0277506, 0.09185404, 0.08641303, 0.07655721, 0.02184991, 
    0.008230921, 0.4010298, 0.09382951, 0.000140356, 0.00655006, 0.05040024, 
    0.0001550278, -6.05174e-07,
  1.301152e-08, 1.684572e-10, -1.864527e-06, -3.420507e-05, -1.410619e-07, 
    0.002362686, 2.43446e-10, 0.0005838964, 0.0006698516, 0.2218676, 
    0.1565762, 0.02907202, 0.006331413, 0.02057441, 0.03701621, 0.007393644, 
    0.009953471, 0.03971933, 0.008650971, 0.05178288, 0.01567518, 0.2093656, 
    0.006458067, -0.0007109112, 0.000650371, 0.003607459, 0.02632825, 
    0.0003775017, 2.021193e-07,
  -1.505434e-07, 0.02151776, 0.01197599, 0.02719425, 0.06941453, 0.007920913, 
    -0.001145478, 0.0001635807, 0.0158063, 0.2725543, 0.1188661, 0.04424361, 
    0.06747863, 0.1017876, 0.09731085, 0.298752, 0.1455072, 0.1602022, 
    0.02293889, 0.005380108, 0.05203801, 0.2058212, 0.182372, 0.3425953, 
    0.14056, 0.07143667, 0.0669056, 0.06343449, -0.000128325,
  0.1294447, 0.006463026, 0.03417784, 0.4298553, 0.02667279, 0.06791251, 
    0.1636153, -7.454384e-05, 0.01333627, 0.08325329, 0.1202184, 0.08181472, 
    0.08078904, 0.1055071, 0.07480226, 0.1752, 0.3807769, 0.3237413, 
    0.1350694, 0.0980354, 0.2143092, 0.1063018, 0.2350152, 0.1444207, 
    0.1774375, 0.1605994, 0.1732827, 0.09106583, 0.1547646,
  0.2605032, 0.2190073, 0.3019969, 0.3131725, 0.3834269, 0.2579547, 
    0.09115479, 0.08913054, 0.009712552, 0.02370027, 0.007751235, 0.02160536, 
    0.1852609, 0.04737784, 0.1349797, 0.1262221, 0.2514399, 0.3620996, 
    0.232271, 0.3764342, 0.1485905, 0.1921042, 0.1621381, 0.433031, 
    0.3101099, 0.1066133, 0.1479585, 0.1597711, 0.2070943,
  0.2716337, 0.2000048, 0.2526699, 0.5760715, 0.4911786, 0.3132607, 
    0.5577124, 0.5159796, 0.4134766, 0.4367236, 0.4380316, 0.3303418, 
    0.1177864, 0.1598942, 0.4886919, 0.2953073, 0.470782, 0.3752481, 
    0.3117267, 0.1840729, 0.2908367, 0.3116977, 0.3078837, 0.2361513, 
    0.7179474, 0.1100177, 0.1195937, 0.2662124, 0.1950191,
  0.1890793, 0.1219296, 0.2321928, 0.1249004, 0.4485947, 0.4013948, 
    0.6079792, 0.577783, 0.3445481, 0.5883388, 0.6854289, 0.4918393, 
    0.3786573, 0.4548034, 0.5506861, 0.3965981, 0.4100649, 0.2331098, 
    0.1898957, 0.3167006, 0.1665572, 0.3536257, 0.1923673, 0.06971264, 
    0.04488521, 0.3405695, 0.5150814, 0.2957684, 0.2587971,
  0.3286465, 0.5042451, 0.4536609, 0.4409929, 0.3699639, 0.5223622, 
    0.6938642, 0.7026649, 0.7140833, 0.6763086, 0.5862454, 0.4953026, 
    0.5467826, 0.5647654, 0.4195353, 0.49226, 0.3895864, 0.3146806, 0.333713, 
    0.4594611, 0.4110053, 0.2383334, 0.1888479, 0.1603175, 0.1393353, 
    0.04715423, 0.05133107, 0.2056561, 0.4038661,
  0.4173191, 0.4248479, 0.4323767, 0.4399055, 0.4474342, 0.4549631, 
    0.4624918, 0.4544098, 0.4693805, 0.4843513, 0.499322, 0.5142927, 
    0.5292635, 0.5442342, 0.5208071, 0.5022901, 0.4837731, 0.4652561, 
    0.4467391, 0.4282221, 0.4097051, 0.4225257, 0.4185432, 0.4145607, 
    0.4105782, 0.4065956, 0.4026131, 0.3986306, 0.411296,
  0.4079661, 0.5115343, 0.6600119, 0.653678, 0.2463226, 0.1445636, 0.266823, 
    0.489029, 0.5772257, 0.5326946, 0.4650939, 0.3801453, 0.4967052, 
    0.02909042, 0.2207209, 0.2060569, 0.2480907, 0.1653684, 0.09226913, 
    0.09521756, 0.434834, 0.4513844, 0.1461308, 0.1486617, 0.1749403, 
    0.1828376, 0.1087774, 0.1459614, 0.1897272,
  0.1848499, 0.1731696, 0.216477, 0.07793817, 0.05697552, 0.007954068, 
    0.05606166, 0.1162963, 0.2236219, 0.2438332, 0.2594295, 0.1323285, 
    0.06779508, 0.1162997, 0.1283476, 0.2433781, 0.2376505, 0.266306, 
    0.3024325, 0.132284, 0.255735, 0.4024093, 0.6449634, 0.2945483, 
    0.1969276, 0.2170474, 0.2300286, 0.1764515, 0.2042171,
  0.3892669, 0.4061221, 0.3721152, 0.4675909, 0.5615498, 0.5555423, 0.463527, 
    0.2705588, 0.1577294, 0.1275588, 0.2425826, 0.4105212, 0.480132, 
    0.4629157, 0.3498443, 0.4120665, 0.4369364, 0.503709, 0.2980213, 
    0.1814471, 0.2254329, 0.2723625, 0.2984, 0.4142721, 0.4750885, 0.4539928, 
    0.4958802, 0.4195578, 0.3859563,
  0.3154453, 0.3233549, 0.4025172, 0.3446405, 0.3824294, 0.3833336, 
    0.4089437, 0.342774, 0.3271961, 0.2643726, 0.1537929, 0.2118739, 
    0.2140543, 0.2433585, 0.2931165, 0.2280803, 0.1909364, 0.150438, 
    0.1597835, 0.1583454, 0.1857729, 0.29957, 0.3436819, 0.1465481, 
    0.05428193, 0.2514916, 0.3100726, 0.3243996, 0.3691411,
  0.1461897, 0.07980874, 0.04688226, 0.197398, 0.1599968, 0.2075647, 
    0.2326415, 0.345333, 0.2671842, 0.06927389, 0.05335364, 0.02301404, 
    0.01923828, 0.06671582, 0.3410187, 0.1448247, 0.04178548, 0.1676375, 
    0.1403135, 0.1097516, 0.2321217, 0.2062389, 0.1466581, 0.01377416, 
    0.02691204, 0.2138282, 0.3920589, 0.2575533, 0.1426363,
  0.04029651, 0.02576978, 0.08798005, 0.00809642, 0.02443881, 0.02068901, 
    0.004948254, 0.02305382, 0.06113672, 0.0003983024, 0.01165712, 
    0.005589775, 0.001685701, 0.00805183, 0.1587344, 0.06733806, 0.0831975, 
    0.04627913, 0.006012593, 0.0007933326, 0.01814171, 0.003301891, 
    0.01400843, 0.1097222, -6.671649e-07, 0.04624718, 0.00467157, 
    0.001342161, 0.0233585,
  0.008825413, 0.0989375, 0.006003403, 0.001925326, 0.004740328, 
    0.0006096383, 0.005809409, 0.002085813, 0.01973319, 0.0539065, 0.0296445, 
    0.0002036478, 4.851365e-05, 0.004959073, 0.005216868, 0.02016483, 
    0.01954411, 0.0005200633, 2.911193e-05, 1.874228e-05, 0.0001032147, 
    0.003241983, 0.02074908, 0.03538501, 0.01367766, 0.2234793, 0.003135229, 
    0.0005009237, 0.0005212566,
  0.0208513, 0.008425881, 0.04113552, 0.03546896, 0.004675106, 0.003260946, 
    0.0008711542, 0.0003719981, 0.003057781, 0.001349003, 0.00258491, 
    0.0001566818, 0.002394836, 0.000675463, 0.04528103, 0.00526713, 
    3.856709e-05, 0.0005323709, 0.0003750133, 0.0001059282, 0.001547406, 
    0.00281834, 0.009958193, 0.02116494, 0.0439655, 0.01095873, -0.000530566, 
    0.002313459, 0.01188272,
  0.0004589304, 0.007470433, 0.0002586706, 0.00802234, 0.0357003, 0.01583863, 
    0.0308282, 0.03835855, 0.03247402, 0.04849983, 0.001774791, 0.0007599666, 
    0.00138093, 0.003143955, 0.01799287, 0.002860757, 0.0008901866, 
    0.003014983, 0.001063484, 0.007268639, 0.0189281, 0.04169434, 0.05959729, 
    0.0003203999, 0.01849306, 0.04846953, 0.0004664685, 0.0007814494, 
    0.003529962,
  3.480918e-10, 7.363336e-11, 1.945082e-10, -0.0007553999, 0.03954767, 
    0.002807257, -0.0009152625, 0.002334734, 7.408038e-05, 0.02539893, 
    0.06358176, 0.001705298, 0.00110737, 0.001076251, 0.0003181903, 
    0.000599712, 0.01131644, 0.03934452, 0.04301561, 0.02813201, 0.008571187, 
    0.002152722, 0.3022341, 0.07909445, -8.838681e-06, 0.003094029, 
    0.02324252, -2.007641e-05, -1.089771e-06,
  1.230119e-08, 1.098955e-10, -5.435753e-07, -5.908702e-06, -1.094891e-07, 
    0.001112894, 2.368185e-10, 5.525647e-05, 0.0004859403, 0.1661279, 
    0.09328608, 0.01162249, 0.002814155, 0.006706827, 0.01097568, 
    0.002906981, 0.004844959, 0.01737138, 0.004138367, 0.02798965, 
    0.02380784, 0.171265, 0.001630738, -0.001206615, 0.0003151647, 
    0.001807488, 0.01289859, 0.0001834286, 1.913978e-07,
  -1.632815e-08, 0.007308512, 0.006062288, 0.01295671, 0.06251727, 
    0.005367192, -0.0009608361, 9.060113e-05, 0.01030206, 0.2638902, 
    0.09664826, 0.03352892, 0.04149608, 0.08046937, 0.08037332, 0.2784463, 
    0.08138641, 0.1284104, 0.01106957, 0.002087333, 0.04251701, 0.1766843, 
    0.1454959, 0.2377986, 0.07196718, 0.0310446, 0.02412524, 0.02837006, 
    4.134255e-05,
  0.09850534, 0.002603037, 0.01651408, 0.408186, 0.0134977, 0.06329045, 
    0.1545327, -3.842395e-05, 0.01325204, 0.05731287, 0.1107188, 0.06818315, 
    0.07060297, 0.08972537, 0.05405305, 0.1503271, 0.3468568, 0.2772767, 
    0.09722462, 0.09359442, 0.2006426, 0.070349, 0.1819182, 0.1200181, 
    0.1428149, 0.110416, 0.1084095, 0.04808475, 0.1256632,
  0.1986497, 0.2153532, 0.2900803, 0.2998344, 0.3116174, 0.2289422, 
    0.06368435, 0.08105177, 0.005693228, 0.02419575, 0.003092, 0.02033065, 
    0.1323164, 0.02610681, 0.1098699, 0.1102617, 0.2092379, 0.3299977, 
    0.2093127, 0.3736793, 0.1231128, 0.1331035, 0.1254742, 0.4334273, 
    0.2552027, 0.08098935, 0.1173482, 0.1158223, 0.1495716,
  0.2005035, 0.2238495, 0.251124, 0.5831594, 0.4805084, 0.3217398, 0.4899337, 
    0.422696, 0.3778853, 0.3790422, 0.4078949, 0.3957009, 0.1140815, 
    0.1334682, 0.4161839, 0.302268, 0.4512898, 0.3495535, 0.31063, 0.1711041, 
    0.3235829, 0.292275, 0.3359117, 0.2109734, 0.6770776, 0.08289308, 
    0.1082903, 0.2095404, 0.1384369,
  0.1610303, 0.09284699, 0.2039475, 0.08623618, 0.4629528, 0.443301, 
    0.6862045, 0.5444641, 0.3503591, 0.6445851, 0.7492435, 0.5686015, 
    0.4556755, 0.5217823, 0.5354459, 0.5348007, 0.4263574, 0.2420178, 
    0.2318816, 0.3734562, 0.1825496, 0.3794785, 0.2150707, 0.1210795, 
    0.057019, 0.3000225, 0.5153053, 0.2517941, 0.2230299,
  0.4306765, 0.4995745, 0.4627345, 0.4326322, 0.3552786, 0.5605334, 
    0.6999528, 0.7296959, 0.8046473, 0.7281616, 0.665867, 0.6084763, 
    0.6335701, 0.655687, 0.6016153, 0.5882704, 0.4736308, 0.4216651, 
    0.4857277, 0.534336, 0.4835744, 0.2681614, 0.1928794, 0.2229994, 
    0.1598651, 0.06728608, 0.03054201, 0.2168762, 0.5035459,
  0.4153857, 0.4225698, 0.4297539, 0.436938, 0.4441221, 0.4513063, 0.4584903, 
    0.4220374, 0.4387548, 0.4554722, 0.4721896, 0.4889069, 0.5056244, 
    0.5223417, 0.5625827, 0.54353, 0.5244774, 0.5054247, 0.486372, 0.4673194, 
    0.4482667, 0.4450679, 0.4402191, 0.4353702, 0.4305214, 0.4256725, 
    0.4208237, 0.4159749, 0.4096384,
  0.3494994, 0.4846241, 0.5965579, 0.658792, 0.3129088, 0.1295786, 0.2642592, 
    0.515193, 0.401558, 0.3631147, 0.3594262, 0.3182997, 0.4283205, 
    0.01341037, 0.2329455, 0.214969, 0.2285122, 0.1933046, 0.07210254, 
    0.1273244, 0.4134165, 0.4581203, 0.1013714, 0.09864166, 0.146779, 
    0.1857174, 0.1238971, 0.1121768, 0.1465687,
  0.1215252, 0.1121813, 0.1411038, 0.04760361, 0.02611893, 0.002635277, 
    0.03775344, 0.07994143, 0.1511302, 0.1831379, 0.1910438, 0.1322262, 
    0.04394391, 0.09315415, 0.09180398, 0.2034325, 0.184584, 0.189541, 
    0.2284809, 0.08306892, 0.1773495, 0.3255208, 0.6084119, 0.2333878, 
    0.1769363, 0.189024, 0.191703, 0.141225, 0.1593441,
  0.2816689, 0.3066787, 0.291788, 0.4099408, 0.4574598, 0.4605158, 0.3638116, 
    0.2088101, 0.118408, 0.09965923, 0.2181702, 0.3624931, 0.4178383, 
    0.3936141, 0.2654047, 0.335042, 0.3663805, 0.4346541, 0.2519003, 
    0.1432633, 0.1714331, 0.2180378, 0.2314645, 0.3286652, 0.4247198, 
    0.4097249, 0.4360956, 0.3667027, 0.321309,
  0.2401338, 0.2385499, 0.2965422, 0.2600029, 0.315625, 0.3642095, 0.3691744, 
    0.2823124, 0.2565587, 0.1968614, 0.09748024, 0.1440437, 0.1637834, 
    0.2170738, 0.267863, 0.1778431, 0.1598987, 0.1007373, 0.107814, 
    0.1142154, 0.1345036, 0.2363258, 0.2603005, 0.1173963, 0.063719, 
    0.2326834, 0.2755232, 0.2708634, 0.2983049,
  0.102337, 0.04450796, 0.02737185, 0.1529062, 0.1097165, 0.1758588, 
    0.1756598, 0.3163605, 0.1854752, 0.04165206, 0.03200353, 0.01171548, 
    0.01446133, 0.04367328, 0.3008797, 0.1096797, 0.03057016, 0.1396025, 
    0.09969544, 0.07940212, 0.1712216, 0.115997, 0.09331635, 0.01925166, 
    0.0343319, 0.1695591, 0.3144737, 0.1880881, 0.09752651,
  0.01992812, 0.01500439, 0.07062496, 0.003463099, 0.006836071, 0.01540172, 
    0.002142376, 0.0105461, 0.02859285, 0.0001683179, 0.005226873, 
    0.002950476, 0.0003977662, 0.00313891, 0.1027552, 0.05353651, 0.07747742, 
    0.02524642, 0.002898614, 0.0003569039, 0.008863288, 0.00181807, 
    0.007083519, 0.08788865, -8.209083e-05, 0.02141112, 0.001433516, 
    0.0006138734, 0.00698108,
  0.004181285, 0.09654544, 0.002226551, 0.0008701692, 0.0004699139, 
    0.0003299518, 0.002613414, 0.0009853226, 0.009229676, 0.02634266, 
    0.02045823, 0.0001044653, 1.83483e-05, 0.001775663, 0.000686082, 
    0.00944226, 0.0108975, 0.0002450202, 9.195467e-06, 6.347349e-06, 
    4.865924e-05, 0.001328674, 0.009782302, 0.01956487, 0.009364407, 
    0.1889568, 0.001742849, 8.731816e-05, 0.0001953462,
  0.01098963, 0.002718032, 0.04079177, 0.0243125, 0.00204457, 0.001647049, 
    0.0004592791, 0.0002071227, 0.001680037, 0.0005810109, 0.0008946763, 
    6.40466e-05, 0.001052553, 0.0001072829, 0.0273105, 0.002482447, 
    1.304855e-05, 0.0003185382, 0.0001868165, 3.410435e-05, 0.0008718835, 
    0.001448706, 0.00509325, 0.02890357, 0.04754002, 0.006763322, 
    -0.0001503685, 0.001104967, 0.006395726,
  0.0002342909, 0.004279988, 0.0003314614, 0.009934776, 0.02066959, 
    0.01112231, 0.02536912, 0.02017106, 0.03282103, 0.03382922, 0.000877061, 
    0.0003538541, 0.0004813324, 0.002352997, 0.02011342, 0.000629345, 
    0.0003843962, 0.0002048002, 0.0002212729, 0.0009026428, 0.002901612, 
    0.01265064, 0.02025971, 0.0001549996, 0.01336211, 0.01890795, 
    0.0001468674, 0.0004415158, 0.001874702,
  3.4483e-10, 7.106551e-11, 1.959285e-10, 0.0006771224, 0.01931535, 
    0.001334864, -0.0009779397, 0.00142535, -6.300698e-07, 0.01110652, 
    0.02832857, 0.0003277559, 0.0003541122, 0.0002454808, 0.0002343839, 
    0.0002647261, 0.003176988, 0.02162266, 0.01767218, 0.01035663, 
    0.002873199, 0.001042444, 0.1938114, 0.05540112, -1.66514e-06, 
    0.001816208, 0.01299926, -3.346476e-05, -5.737038e-06,
  1.19989e-08, 9.700345e-11, -2.188425e-07, 3.767399e-06, -8.260799e-08, 
    0.0006959796, 2.750782e-10, 1.313611e-05, 0.0001707248, 0.1263457, 
    0.04746722, 0.004956103, 0.001655765, 0.002636202, 0.002561986, 
    0.001753155, 0.002579163, 0.006821759, 0.002503539, 0.01743176, 
    0.01173474, 0.146624, 0.0006755349, -0.0008516714, 0.0001941792, 
    0.001116161, 0.007876685, 0.0001085177, 1.857306e-07,
  3.455312e-08, 0.0037615, 0.003183001, 0.006705583, 0.05576153, 0.003962223, 
    -0.0008228131, 3.646093e-05, 0.009414435, 0.2188654, 0.07849151, 
    0.01555702, 0.02552769, 0.06133367, 0.06342585, 0.1509209, 0.04917651, 
    0.09222055, 0.006811192, 0.001217073, 0.03654128, 0.1415751, 0.1031041, 
    0.08947165, 0.04082216, 0.01657347, 0.01236357, 0.01267306, 1.025085e-05,
  0.07735668, 0.001526142, 0.009737791, 0.3753786, 0.008152057, 0.04627763, 
    0.1426419, -2.205703e-05, 0.01250657, 0.05108338, 0.1002745, 0.05511006, 
    0.05769958, 0.07366372, 0.03860808, 0.120152, 0.268012, 0.2183482, 
    0.06386711, 0.08044133, 0.1737832, 0.04778152, 0.1377369, 0.1021702, 
    0.110053, 0.07135645, 0.06622554, 0.02717226, 0.0968151,
  0.2035963, 0.2064628, 0.2406034, 0.269594, 0.2385925, 0.1892267, 
    0.03961309, 0.07337432, 0.004315337, 0.02863648, 0.001179391, 0.02067971, 
    0.0961588, 0.01490509, 0.0889093, 0.08980242, 0.1784993, 0.277966, 
    0.1614669, 0.3598204, 0.09243743, 0.08767179, 0.08746734, 0.3996454, 
    0.20507, 0.06168007, 0.09270665, 0.0743429, 0.1094076,
  0.1356912, 0.2342146, 0.2159633, 0.5403792, 0.4475788, 0.2938352, 
    0.3774464, 0.2921626, 0.3061734, 0.2935156, 0.3643956, 0.483733, 
    0.1070675, 0.1427855, 0.3713109, 0.2718979, 0.4480152, 0.3189505, 
    0.281599, 0.1861648, 0.364053, 0.2386385, 0.2867234, 0.1653384, 0.648438, 
    0.06094183, 0.09447093, 0.1466686, 0.08610567,
  0.1262612, 0.07225411, 0.2092126, 0.05873395, 0.4681278, 0.4208169, 
    0.7631572, 0.5794985, 0.3519521, 0.6463995, 0.7723231, 0.5394977, 
    0.6529745, 0.5040274, 0.5455718, 0.5847752, 0.4192571, 0.2414154, 
    0.2873465, 0.3627637, 0.2977449, 0.545593, 0.306963, 0.204671, 
    0.09786244, 0.2573621, 0.5142438, 0.2050626, 0.189461,
  0.5120667, 0.5087218, 0.5302676, 0.4737807, 0.4493077, 0.6631492, 0.726473, 
    0.7154371, 0.7421462, 0.7248898, 0.7281728, 0.6081035, 0.6162525, 
    0.6894701, 0.6525051, 0.7246175, 0.6572664, 0.6049152, 0.5488135, 
    0.5257771, 0.5601954, 0.2647463, 0.2229064, 0.2741514, 0.1418745, 
    0.1044239, 0.01937705, 0.2147129, 0.5448129,
  0.3278913, 0.3377218, 0.3475522, 0.3573826, 0.367213, 0.3770435, 0.3868739, 
    0.3759026, 0.3947988, 0.4136949, 0.4325911, 0.4514872, 0.4703833, 
    0.4892795, 0.6024239, 0.5785264, 0.5546288, 0.5307313, 0.5068338, 
    0.4829362, 0.4590387, 0.3801849, 0.3753558, 0.3705268, 0.3656977, 
    0.3608687, 0.3560396, 0.3512106, 0.320027,
  0.2879099, 0.3980478, 0.4689595, 0.5784779, 0.377424, 0.1063478, 0.2382001, 
    0.4142144, 0.2913897, 0.278329, 0.2391403, 0.235842, 0.3251642, 
    0.00836623, 0.2606661, 0.2398228, 0.1535779, 0.193307, 0.05396953, 
    0.1693558, 0.3599415, 0.440773, 0.07451001, 0.07044557, 0.1243229, 
    0.1689109, 0.1349046, 0.07837989, 0.1194581,
  0.07514335, 0.0827539, 0.09104179, 0.03076309, 0.01250583, 0.0009480263, 
    0.02727776, 0.05612962, 0.1202885, 0.1401498, 0.1452369, 0.1278107, 
    0.02671496, 0.06282493, 0.06386802, 0.1523678, 0.1249194, 0.131141, 
    0.1657572, 0.0554725, 0.1108357, 0.2560999, 0.5318149, 0.177715, 
    0.1705088, 0.1561179, 0.1544629, 0.09887411, 0.1119557,
  0.2002383, 0.2086724, 0.2258758, 0.3197483, 0.3452518, 0.336076, 0.2648375, 
    0.1580735, 0.07966699, 0.08371346, 0.1776293, 0.2853032, 0.317189, 
    0.2857448, 0.1969911, 0.253019, 0.2886693, 0.3547705, 0.1927692, 
    0.1045873, 0.1190592, 0.152794, 0.1542049, 0.2297008, 0.3442317, 0.35499, 
    0.361765, 0.2805166, 0.2323129,
  0.1710668, 0.1655233, 0.2208911, 0.1918398, 0.2522029, 0.2990333, 
    0.3044075, 0.2074012, 0.1878382, 0.130375, 0.05799007, 0.09049603, 
    0.1106896, 0.1720641, 0.2505622, 0.1316461, 0.1123262, 0.06479124, 
    0.07305343, 0.07546613, 0.08781204, 0.1654801, 0.176224, 0.09190789, 
    0.05995918, 0.1944516, 0.2366717, 0.2103024, 0.2271557,
  0.06525715, 0.02658814, 0.01615989, 0.1059969, 0.07672834, 0.1166313, 
    0.1322927, 0.2638217, 0.1271495, 0.02333239, 0.02017519, 0.006427453, 
    0.01048025, 0.02511013, 0.2523307, 0.07854439, 0.02409773, 0.1044319, 
    0.06142418, 0.04766763, 0.1233253, 0.06348733, 0.04303538, 0.02540044, 
    0.02524795, 0.1133426, 0.2445042, 0.1195686, 0.06386457,
  0.008033978, 0.007026821, 0.04710307, 0.001969506, 0.002375241, 
    0.009142954, 0.00150047, 0.006461997, 0.01781089, 9.640955e-05, 
    0.002723579, 0.001603501, 8.092268e-05, 0.001497562, 0.05460847, 
    0.03073102, 0.05768804, 0.0110465, 0.001824046, 0.0002316419, 
    0.005403657, 0.001236624, 0.004502122, 0.05424701, -8.391571e-05, 
    0.007579131, 0.0005798822, 0.0003801662, 0.00238662,
  0.002563147, 0.07926993, 0.0007466188, 0.000539405, -0.0005488073, 
    0.0002164277, 0.001584339, 0.0005902231, 0.005559681, 0.01479459, 
    0.01342422, -4.97121e-05, 1.055597e-05, 0.0005963783, 0.0002570793, 
    0.004824118, 0.005740833, 0.0001512394, 5.209616e-06, 3.499394e-06, 
    2.91617e-05, 0.0007106746, 0.005840095, 0.01336261, 0.005358549, 
    0.1415942, 0.0011526, 3.359489e-05, 0.0001077928,
  0.007101007, 0.001046657, 0.03988298, 0.01900703, 0.001202788, 0.001018614, 
    0.0002943946, 0.0001418544, 0.001114946, 0.0005048325, 0.0003906721, 
    5.822931e-05, 0.0003129879, 7.294414e-05, 0.01259101, 0.001160018, 
    8.162076e-06, 0.000220873, 0.0001340433, 1.638248e-05, 0.0005911662, 
    0.0009238691, 0.003244731, 0.02125551, 0.05098302, 0.006673616, 
    -2.911423e-05, 0.0006806553, 0.004166022,
  0.0001446473, 0.003152808, 0.00035488, 0.008743901, 0.009735323, 
    0.006159009, 0.01493743, 0.009157632, 0.03161018, 0.02897366, 
    0.0004878448, 0.0002236425, 0.0003032523, 0.001332389, 0.01258958, 
    0.0002934558, 0.0002495221, 6.851938e-05, 0.0001132189, 0.0003631022, 
    0.001237999, 0.006619262, 0.01003584, 0.0001316211, 0.007885941, 
    0.007348091, 5.143126e-05, 0.0002961715, 0.001216901,
  3.476316e-10, 6.956759e-11, 1.982325e-10, -0.0005965257, 0.0108486, 
    0.0008740434, -0.000808957, 0.001003268, -2.263096e-05, 0.004790578, 
    0.01261356, 0.0001283385, 0.000112933, 0.0001080567, 0.0001941857, 
    0.000162631, 0.00118203, 0.01114929, 0.006589598, 0.003827828, 
    0.0009791787, 0.000635393, 0.1525809, 0.03385134, -8.051628e-07, 
    0.001233325, 0.008520497, -2.303669e-05, -0.0001045762,
  1.197675e-08, 9.556281e-11, -1.270643e-07, 4.158691e-06, -8.312966e-08, 
    0.0004970296, 2.856213e-10, 6.492491e-06, 1.269354e-05, 0.07896496, 
    0.01968009, 0.001978475, 0.001138482, 0.001533969, 0.001008143, 
    0.001222885, 0.001305902, 0.002694838, 0.001743629, 0.01154813, 
    0.005678821, 0.1222838, 0.000376241, -0.0007478725, 0.0001372724, 
    0.0007847204, 0.005547305, 7.362295e-05, 1.802409e-07,
  3.532033e-08, 0.003517386, 0.002008667, 0.004833951, 0.0470937, 
    0.002269767, -0.0007300774, 3.742424e-06, 0.01003777, 0.1564693, 
    0.0658911, 0.008896548, 0.01499055, 0.04053883, 0.04213561, 0.08871823, 
    0.02913844, 0.06094741, 0.004807377, 0.0008361812, 0.03023354, 0.1094241, 
    0.07034813, 0.04746177, 0.0218557, 0.01041243, 0.008226814, 0.007278936, 
    5.942351e-06,
  0.05690828, 0.001042644, 0.008679023, 0.3493307, 0.005961565, 0.03410965, 
    0.1266611, -1.251593e-05, 0.01117892, 0.05676058, 0.0846503, 0.04496302, 
    0.04431613, 0.05763832, 0.02524151, 0.08800075, 0.1909411, 0.1477712, 
    0.0337538, 0.0701715, 0.1493116, 0.03692624, 0.1136848, 0.08342055, 
    0.08248848, 0.04513528, 0.03623408, 0.01545689, 0.06739392,
  0.177334, 0.1867983, 0.1987754, 0.2335984, 0.1667678, 0.1451496, 
    0.02382858, 0.07118037, 0.01615691, 0.03421703, 0.0005009657, 0.03267634, 
    0.07883414, 0.009715783, 0.07063559, 0.07077216, 0.1425641, 0.2075185, 
    0.1048843, 0.3418028, 0.07519829, 0.05945637, 0.06368315, 0.363807, 
    0.1698593, 0.04734597, 0.07073251, 0.04503454, 0.08416118,
  0.1009624, 0.2286805, 0.184727, 0.4942652, 0.3980902, 0.2326968, 0.2770501, 
    0.2326668, 0.2384349, 0.235683, 0.3005152, 0.534156, 0.149767, 0.1439109, 
    0.3353816, 0.2497889, 0.4266395, 0.2851265, 0.2513514, 0.2175668, 
    0.3912286, 0.2663341, 0.2252654, 0.1727066, 0.6274465, 0.04737111, 
    0.07813373, 0.1014689, 0.0525852,
  0.09717118, 0.05589648, 0.2165664, 0.04460963, 0.4334965, 0.3941196, 
    0.7674459, 0.5323163, 0.4145754, 0.6761693, 0.7800612, 0.5245686, 
    0.7871433, 0.3415722, 0.4828456, 0.5124009, 0.4200327, 0.229527, 
    0.3373345, 0.340987, 0.3271672, 0.6722066, 0.5333738, 0.3174122, 
    0.1370222, 0.2029182, 0.5156795, 0.1694012, 0.1468329,
  0.5554347, 0.5507134, 0.5508811, 0.4845088, 0.5291604, 0.6713941, 
    0.6868156, 0.6431353, 0.6606421, 0.5444815, 0.6407927, 0.5994784, 
    0.5493046, 0.5115314, 0.6203527, 0.6010383, 0.5994999, 0.5825809, 
    0.4963729, 0.4926341, 0.4701725, 0.2750737, 0.2784471, 0.3509804, 
    0.1155068, 0.09033512, 0.02160658, 0.1933777, 0.5037616,
  0.2220206, 0.2291644, 0.2363082, 0.2434521, 0.2505959, 0.2577398, 
    0.2648836, 0.2840192, 0.2998556, 0.3156919, 0.3315283, 0.3473647, 
    0.3632011, 0.3790375, 0.4729172, 0.4572284, 0.4415396, 0.4258508, 
    0.410162, 0.3944732, 0.3787844, 0.2635179, 0.2562265, 0.2489351, 
    0.2416437, 0.2343523, 0.2270609, 0.2197694, 0.2163055,
  0.2400485, 0.3074589, 0.3499801, 0.4445128, 0.3406, 0.1082597, 0.1742987, 
    0.3024546, 0.2293474, 0.167166, 0.1494373, 0.1841293, 0.2466507, 
    0.003131939, 0.2706915, 0.2368301, 0.1360325, 0.1543108, 0.03873401, 
    0.1828624, 0.2946025, 0.4203358, 0.06030199, 0.054184, 0.1077274, 
    0.1578856, 0.165846, 0.06319149, 0.109435,
  0.05565972, 0.05867954, 0.06890178, 0.0214869, 0.007226553, 0.0002724747, 
    0.02422995, 0.0427812, 0.09876613, 0.1196818, 0.1302048, 0.121534, 
    0.02108712, 0.04171675, 0.04934757, 0.1112184, 0.08635379, 0.09943639, 
    0.1305512, 0.04481724, 0.07707465, 0.1995343, 0.4390019, 0.1370053, 
    0.1471918, 0.1293329, 0.1255861, 0.07145875, 0.08370487,
  0.1597001, 0.1618508, 0.1783102, 0.2657557, 0.2748826, 0.2647652, 0.210794, 
    0.1240244, 0.05931356, 0.07457442, 0.1390923, 0.2222049, 0.2415768, 
    0.215114, 0.15183, 0.1949334, 0.2327746, 0.2962999, 0.1519769, 0.0845167, 
    0.08394903, 0.1050441, 0.1042185, 0.1545329, 0.2688569, 0.2797542, 
    0.3047795, 0.2225037, 0.179923,
  0.1314917, 0.1233412, 0.1779127, 0.1535753, 0.2025313, 0.2418167, 
    0.2386501, 0.1615329, 0.1433747, 0.09251256, 0.03784464, 0.05798938, 
    0.07568078, 0.1294379, 0.2155112, 0.09170124, 0.07264762, 0.0450261, 
    0.05287202, 0.05331159, 0.06014327, 0.1243348, 0.1298228, 0.0771112, 
    0.04853997, 0.1517166, 0.201339, 0.1715933, 0.1850466,
  0.04331226, 0.01821337, 0.01047608, 0.07033701, 0.0530876, 0.07319904, 
    0.09636031, 0.2059919, 0.0882588, 0.01449853, 0.0127387, 0.004518581, 
    0.008131127, 0.0166055, 0.2171011, 0.05735626, 0.01565297, 0.07596837, 
    0.04054336, 0.03044288, 0.07856777, 0.04041307, 0.02091385, 0.03471738, 
    0.01772968, 0.06799997, 0.1736414, 0.08077965, 0.04324419,
  0.004057655, 0.003457146, 0.02978613, 0.00138899, 0.001428515, 0.004731002, 
    0.001173682, 0.004709988, 0.0131263, 6.634897e-05, 0.001449945, 
    0.001045242, -1.485186e-05, 0.0009662606, 0.03001731, 0.01778312, 
    0.03859606, 0.004421409, 0.001351006, 0.0001756577, 0.003940997, 
    0.0009422271, 0.00329459, 0.04024542, 8.103142e-06, 0.003816482, 
    0.0003417481, 0.0002765737, 0.001445448,
  0.001843861, 0.0592191, 0.000374071, 0.0003933601, -0.0004490522, 
    0.0001607848, 0.001129234, 0.0004154481, 0.003923963, 0.00976677, 
    0.007587074, 2.12399e-05, 7.550071e-06, 0.0002906487, 0.0001730765, 
    0.00271751, 0.003210515, 0.0001071702, 3.747904e-06, 2.600702e-06, 
    2.050819e-05, 0.000459171, 0.00407734, 0.01025748, 0.003382326, 
    0.1019872, 0.0008555638, 1.82844e-05, 7.344879e-05,
  0.005220134, 0.0005663457, 0.04488946, 0.02876621, 0.0008620846, 
    0.000722326, 0.0002141136, 0.0001083298, 0.0008335687, 0.0003924257, 
    0.0002528928, 5.381193e-05, 0.0001179242, 5.026531e-05, 0.005633428, 
    0.0006419604, 5.873387e-06, 0.0001709872, 0.0001067463, 1.017874e-05, 
    0.0004506518, 0.0006771348, 0.002371307, 0.02226294, 0.04354924, 
    0.006585398, 1.88355e-05, 0.0004861456, 0.00307957,
  0.0001024837, 0.01235435, 0.0008654255, 0.009337923, 0.004441651, 
    0.00289169, 0.007708513, 0.004486803, 0.03403025, 0.03904253, 
    0.0003263847, 0.0001649713, 0.0002306309, 0.0006676902, 0.005842966, 
    0.0001673192, 0.0001853214, 3.836034e-05, 7.601448e-05, 0.0001706608, 
    0.0007801598, 0.004405783, 0.005925016, 0.001504091, 0.004353568, 
    0.003227339, 2.585958e-05, 0.0002227168, 0.0008980342,
  3.532122e-10, 6.751243e-11, 2.000771e-10, -0.0003524244, 0.007255807, 
    0.0006477432, -0.0005779523, 0.0007604523, -3.641357e-05, 0.002155656, 
    0.005606384, 7.420983e-05, 7.050232e-05, 5.942663e-05, 0.0001519372, 
    0.0001170801, 0.0006530847, 0.005742321, 0.002958156, 0.001797104, 
    0.0004133917, 0.0004498188, 0.1087246, 0.01883108, -6.179381e-07, 
    0.0009415878, 0.006314618, -1.725032e-05, -0.0001746314,
  1.221788e-08, 1.004989e-10, -8.866691e-08, 3.804348e-06, -6.860232e-08, 
    0.000391549, 2.947204e-10, 4.369155e-06, -6.0637e-05, 0.04944279, 
    0.01078639, 0.001050944, 0.0008656977, 0.001103871, 0.0006306978, 
    0.0009472722, 0.0006699265, 0.001450634, 0.001353436, 0.008498177, 
    0.003297703, 0.1040854, 0.0002684913, -0.000708771, 0.0001072556, 
    0.0006070219, 0.004316996, 5.6046e-05, 1.789921e-07,
  3.277788e-08, 0.003152983, 0.001517271, 0.003933711, 0.04069365, 
    0.0009628592, -0.0007129479, -6.537387e-05, 0.01287833, 0.1153836, 
    0.05195063, 0.004997149, 0.008765377, 0.02681437, 0.02820923, 0.04952363, 
    0.01776025, 0.03629524, 0.003758132, 0.0006431874, 0.02477885, 
    0.08714589, 0.05352844, 0.02824031, 0.01249654, 0.007360579, 0.006268725, 
    0.004978243, 6.587155e-06,
  0.04002609, 0.000606413, 0.007394423, 0.3247055, 0.004867936, 0.02924299, 
    0.1091693, -8.170285e-06, 0.007281734, 0.06402717, 0.07372957, 
    0.03997867, 0.03297813, 0.04547445, 0.01781903, 0.0642799, 0.1431886, 
    0.1032607, 0.01880035, 0.06134463, 0.1382138, 0.03149761, 0.09573419, 
    0.06974709, 0.06361137, 0.02953028, 0.02142645, 0.01046577, 0.04773475,
  0.1571906, 0.167902, 0.1749372, 0.2078826, 0.1369508, 0.1426506, 
    0.01727871, 0.08740927, 0.03266687, 0.03261752, 0.000698764, 0.04949988, 
    0.06904733, 0.007461476, 0.06034731, 0.05718468, 0.1146611, 0.1573066, 
    0.07740308, 0.3352422, 0.06866539, 0.0475852, 0.05282059, 0.3184673, 
    0.1511529, 0.03850644, 0.0550644, 0.03151152, 0.06805473,
  0.08340862, 0.2312703, 0.174934, 0.460394, 0.3587455, 0.1916905, 0.218987, 
    0.201605, 0.1887297, 0.1865577, 0.2527537, 0.6336944, 0.2426497, 
    0.154707, 0.309948, 0.2217395, 0.4201436, 0.2738098, 0.2617461, 0.233743, 
    0.379328, 0.301532, 0.1244369, 0.1554163, 0.6124517, 0.04140468, 
    0.06398533, 0.07577153, 0.03591802,
  0.07805458, 0.04460768, 0.2243452, 0.0358832, 0.4205545, 0.3012149, 
    0.6978616, 0.5396189, 0.5235912, 0.6698493, 0.7860794, 0.5264034, 
    0.7123756, 0.1924, 0.3402275, 0.3986978, 0.4532145, 0.2094885, 0.3411163, 
    0.2657793, 0.3400038, 0.5337639, 0.3485543, 0.3850197, 0.1518175, 
    0.1605002, 0.5469408, 0.1588467, 0.1213297,
  0.5430065, 0.5109746, 0.539454, 0.4176169, 0.4829469, 0.5436199, 0.5131895, 
    0.4345033, 0.5024615, 0.4009695, 0.446234, 0.4628523, 0.3284924, 
    0.2952184, 0.3954174, 0.4530898, 0.4413593, 0.4161125, 0.3100573, 
    0.302803, 0.350151, 0.3246369, 0.3089049, 0.4301963, 0.08954581, 
    0.06287985, 0.03022687, 0.1765304, 0.3957359,
  0.1362991, 0.1385082, 0.1407173, 0.1429263, 0.1451354, 0.1473444, 
    0.1495535, 0.14565, 0.1617251, 0.1778003, 0.1938754, 0.2099506, 
    0.2260257, 0.2421008, 0.3342765, 0.3243312, 0.3143859, 0.3044406, 
    0.2944952, 0.2845499, 0.2746046, 0.221341, 0.2130021, 0.2046632, 
    0.1963244, 0.1879855, 0.1796466, 0.1713078, 0.1345319,
  0.2256765, 0.2887464, 0.2803885, 0.3107904, 0.2605087, 0.0888455, 
    0.1224496, 0.209882, 0.1772457, 0.1162502, 0.1095533, 0.1505283, 
    0.195976, 0.002470352, 0.2942161, 0.2274349, 0.1260891, 0.1417742, 
    0.03518659, 0.1949931, 0.2579995, 0.4013121, 0.06147605, 0.05459906, 
    0.09568171, 0.1643264, 0.1744353, 0.06364714, 0.1039434,
  0.0458244, 0.04945482, 0.05734179, 0.01795254, 0.009453236, -2.682987e-05, 
    0.02208511, 0.03610712, 0.08872257, 0.1120885, 0.1188749, 0.1183302, 
    0.01794653, 0.03354004, 0.04262323, 0.09250962, 0.06977472, 0.08163482, 
    0.1083829, 0.03960589, 0.06309023, 0.1646921, 0.3830518, 0.1194289, 
    0.1334333, 0.1061943, 0.1064684, 0.05950529, 0.07050443,
  0.1349688, 0.1398031, 0.1496522, 0.236474, 0.2373998, 0.2281322, 0.1812017, 
    0.1038786, 0.04876169, 0.06108418, 0.1102057, 0.1819559, 0.2030723, 
    0.1723337, 0.126683, 0.1655915, 0.197989, 0.2487712, 0.123691, 
    0.07305072, 0.06567005, 0.08032023, 0.07927377, 0.1162788, 0.2066633, 
    0.2177253, 0.2632527, 0.1822287, 0.1548568,
  0.1107006, 0.1032364, 0.1470389, 0.128338, 0.1621483, 0.2010335, 0.1992113, 
    0.1357191, 0.1192122, 0.07478373, 0.02881067, 0.04132665, 0.05628759, 
    0.09756029, 0.1711652, 0.06951718, 0.05532895, 0.03380473, 0.04132429, 
    0.04166827, 0.04468841, 0.09873685, 0.1058365, 0.08089026, 0.03907652, 
    0.1208613, 0.1678104, 0.143881, 0.1576675,
  0.03215691, 0.0134785, 0.007703945, 0.04813287, 0.03872335, 0.05070072, 
    0.06893439, 0.156827, 0.06617318, 0.01064343, 0.009337368, 0.003721935, 
    0.006832214, 0.01306855, 0.2207166, 0.04191806, 0.01116349, 0.05585457, 
    0.02765595, 0.01881012, 0.05713337, 0.02866225, 0.01303158, 0.04136656, 
    0.01482164, 0.04666971, 0.1267674, 0.05844967, 0.03261893,
  0.002791753, 0.002366664, 0.02298284, 0.001136435, 0.00108975, 0.002991038, 
    0.0009868438, 0.003863871, 0.01083916, 5.570018e-05, 0.001054038, 
    0.0007811078, 0.0006255971, 0.0007685106, 0.01613867, 0.008430404, 
    0.02479315, 0.002768045, 0.001114616, 0.0001507725, 0.003178934, 
    0.0007897061, 0.002725546, 0.03332178, 0.007302403, 0.002609483, 
    0.0002574937, 0.0002247815, 0.001122961,
  0.001521233, 0.04589945, 0.006916927, 0.0003228401, -0.000474856, 
    0.0001335391, 0.0009168258, 0.000339782, 0.003192456, 0.007549281, 
    0.008394828, 0.0009807791, 6.353518e-06, 0.0002127506, 0.0001395627, 
    0.001862652, 0.002200968, 8.709254e-05, 3.167664e-06, 2.212508e-06, 
    1.681957e-05, 0.0003526423, 0.00329119, 0.008589911, 0.01339281, 
    0.121368, 0.000705576, 1.25356e-05, 5.702097e-05,
  0.004276001, 0.000261322, 0.08189362, 0.1512136, 0.0006975096, 
    0.0005755487, 0.0001739256, 9.13825e-05, 0.0006887913, 0.0003293923, 
    0.0002000288, 4.90147e-05, 6.19611e-05, 4.028618e-05, 0.003516123, 
    0.0004499139, 5.039029e-06, 0.0001455284, 9.345031e-05, 8.053028e-06, 
    0.0003817785, 0.000563252, 0.0019438, 0.1617787, 0.06750878, 0.0271809, 
    -4.61096e-05, 0.0003949672, 0.002534486,
  8.16185e-05, 0.05804646, 0.002783072, 0.0086112, 0.002564168, 0.001853568, 
    0.004757731, 0.002949372, 0.05496657, 0.1064318, 0.0002617252, 
    0.0001361527, 0.0001919266, 0.0004512503, 0.003308547, 0.0001249158, 
    0.0001542579, 2.807038e-05, 6.086059e-05, 0.0001098715, 0.0005964789, 
    0.00344962, 0.004347577, 0.02958811, 0.0114379, 0.002082874, 
    1.842444e-05, 0.0001857329, 0.0007383751,
  3.607283e-10, 6.50184e-11, 2.004623e-10, 0.0008501146, 0.0057385, 
    0.0005509286, -0.0003840637, 0.0006481168, -0.0005711622, 0.00126413, 
    0.003400091, 5.481098e-05, 5.946697e-05, 4.576722e-05, 0.0001280801, 
    9.740367e-05, 0.0004977097, 0.003578573, 0.001827267, 0.001259926, 
    0.0002673647, 0.0003674015, 0.1224718, 0.01555429, -5.30736e-07, 
    0.0008148754, 0.005272143, -1.417348e-05, -0.0002013637,
  1.233116e-08, 1.037166e-10, -6.610765e-08, 3.696223e-06, -5.29704e-08, 
    0.0003371194, 3.163208e-10, 3.503287e-06, -7.662617e-05, 0.02997365, 
    0.006718702, 0.0007365988, 0.0007371513, 0.000913094, 0.000497783, 
    0.0008103342, 0.0005042875, 0.001064886, 0.001174238, 0.006954202, 
    0.002344566, 0.09550078, 0.0002212737, -0.0009761992, 9.265601e-05, 
    0.0005128034, 0.003687114, 4.817304e-05, 1.810332e-07,
  5.027268e-08, 0.002500267, 0.001186171, 0.0034468, 0.0382693, 0.0005166769, 
    -0.0007449948, -0.0001031619, 0.0249494, 0.1071064, 0.03609718, 
    0.003617801, 0.005565541, 0.01877909, 0.02051209, 0.03116692, 0.01157583, 
    0.02515631, 0.003243088, 0.000552466, 0.02210145, 0.0753066, 0.05288186, 
    0.01862242, 0.009151695, 0.006036261, 0.005270183, 0.003998588, 
    3.287283e-06,
  0.03216423, 0.0003999506, 0.007117235, 0.3238128, 0.004248142, 0.02638696, 
    0.1114808, -6.843053e-06, 0.005886576, 0.06636941, 0.07563592, 
    0.03178992, 0.02750015, 0.03905548, 0.01451965, 0.04738072, 0.1154972, 
    0.0794825, 0.01290722, 0.06015355, 0.1377099, 0.02831161, 0.08768946, 
    0.06245565, 0.05366532, 0.02221856, 0.01528191, 0.00857574, 0.03981792,
  0.1439251, 0.1553911, 0.1663543, 0.2063911, 0.1219875, 0.1558245, 
    0.0192099, 0.1685215, 0.1495616, 0.04502644, 0.002613182, 0.1267577, 
    0.06620299, 0.00644646, 0.05142227, 0.04930031, 0.09303813, 0.1263339, 
    0.06219705, 0.3591062, 0.06774294, 0.04947646, 0.07123856, 0.3172657, 
    0.1467568, 0.03395741, 0.04697829, 0.0251764, 0.05901936,
  0.07540641, 0.2994518, 0.1999265, 0.4584744, 0.3613107, 0.2228228, 
    0.2131205, 0.20332, 0.2118095, 0.2056675, 0.2768272, 0.7186487, 
    0.3584505, 0.1527865, 0.2982863, 0.214499, 0.4283873, 0.273889, 
    0.3140199, 0.298161, 0.4375939, 0.350627, 0.09589578, 0.1649509, 
    0.6077451, 0.04248615, 0.05672207, 0.0636438, 0.02836452,
  0.06794868, 0.03845707, 0.2794136, 0.03008977, 0.4121671, 0.2470384, 
    0.6350015, 0.5282483, 0.5936229, 0.6485104, 0.7790262, 0.6273101, 
    0.5072613, 0.1357684, 0.2759511, 0.3359789, 0.5424435, 0.2293513, 
    0.3207549, 0.2226102, 0.3254522, 0.4078861, 0.2705632, 0.4781545, 
    0.1559142, 0.152879, 0.5960979, 0.1526325, 0.1092882,
  0.4999634, 0.4922405, 0.504155, 0.3645059, 0.3735993, 0.4539641, 0.4095363, 
    0.3315294, 0.4414512, 0.3264482, 0.3564098, 0.3311793, 0.2318083, 
    0.2097417, 0.2634673, 0.2865834, 0.2917119, 0.2934052, 0.2568665, 
    0.2399154, 0.2581529, 0.3337352, 0.3425704, 0.5817615, 0.09160598, 
    0.05088319, 0.04584905, 0.1656636, 0.3429095,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0006266061, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, -5.037389e-06, 0, 0, 0, 0, 0, 0, 0, 0, -7.164392e-06, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 5.474724e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0008570054, 0.0004400414, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 5.067427e-05, 0, 0, -2.568102e-05, 0, 0, -1.384702e-05, 
    -4.020165e-05, 0, 0, 0, 0, -3.202425e-05, 0, 0, -2.977926e-06, 0, 0, 0, 
    0, 0, -2.693896e-05, -2.266856e-05, -1.222761e-05, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0001918, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 4.647254e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, -5.792723e-05, 3.022687e-05, 0, 0, 0, 0, 0, 0, 0, 0.002675694, 
    0.003442427, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2.409464e-05, 0, 0, 0,
  0, 0, -1.094549e-05, 0, 0, -0.0001039485, -7.738102e-06, 0.001250624, 
    -6.314457e-05, 0.000238327, 0, 0, 0.000272508, -9.322511e-05, 
    0.0007619599, 0.003907819, 0, -2.578099e-05, 0, 0, 0, 0, 0, 
    -3.589016e-05, -4.029537e-05, -3.067263e-05, 0, 0, 0,
  0, 0, 0, 0, 0, -1.643171e-08, -3.628938e-05, 0, -2.82487e-06, 0.001905516, 
    0, 0, -7.60217e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0.0001169772, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2.085876e-07, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 3.341457e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -5.609647e-05, 
    -7.228069e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, -3.13268e-05, 0, -0.0001844949, 0.002521491, 0, 0, 0, 0, 0, 0, 0, 
    0.004579957, 0.008165371, 0, 0, -0.0001347558, 0, 0, 0, 0, 0, 0, 0, 0, 
    -4.015774e-05, 0, 0, 0,
  0, 0, 0.001620554, 0, 0, -0.0001732851, -7.738102e-06, 0.002754573, 
    -9.411781e-05, 0.001981063, 0, 0, 0.001066845, -0.000251738, 0.002603951, 
    0.006874156, 0, -5.67553e-05, 0, 0, 0, 0, 0, 0.0003441847, 6.103497e-05, 
    -6.46635e-05, 0, 0, 0,
  0, 0, -4.525715e-05, 0, 1.643069e-05, -1.10734e-07, -4.770867e-05, 0, 
    2.327928e-05, 0.00670847, 0.003784203, 0, 1.4156e-05, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, -1.484031e-05, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0.0002863905, 0, -1.599945e-10, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -7.10058e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -6.622054e-07, 0, 0, 0,
  0, 0, -4.121613e-06, 0, 0.0002761371, 0, -5.605217e-06, 0, 0, 0, 0, 0, 0, 
    0.000216825, 0, -9.518552e-05, 0.0002451807, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0,
  0, -0.0001075302, 0, 0.0002368531, 0.01037568, 0, 0.004211544, 0, 0, 0, 0, 
    0, 0.01150737, 0.01178095, 0.006654056, -5.175322e-05, -0.0002913501, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.001270729, 0, 0, 0,
  0, 0, 0.00390712, 0, 0, -0.0002439443, -2.429195e-05, 0.004372887, 
    -0.0001004231, 0.002501729, 0.0001608681, -2.100229e-05, 0.001765484, 
    5.873019e-05, 0.00323251, 0.008406972, -1.620797e-05, 3.998259e-05, 0, 0, 
    0, 0, 0, 0.0003436158, 0.0002662597, 0.0003438768, 0, 0, 0,
  0, 0, 0.001452206, 0, 0.001110874, 9.635869e-05, -2.248898e-05, 0, 
    0.0002165561, 0.01181494, 0.01266203, 0, 0.0009889697, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.0007114107, 0, -2.444704e-05, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 6.477443e-06, -1.037153e-05, 0.0003131937, 0, 
    -6.315476e-05, 0, 0, 0, 0.000433439, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -7.053904e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, -1.345329e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0002675324, 0, 0, 0, 0, 0, 0, 0.0007105349, 0.001215178, 0, 0, 0,
  0, 0, -9.689051e-05, 0, 0.001346247, 0, 0.00417548, 0, 0, 0, 0, 0, 0, 
    0.005869114, 0, 0.00164032, 0.002320308, 0, 0, 1.500883e-05, 0, 0, 0, 0, 
    -5.370782e-07, -1.973549e-05, 0.000769638, 0, 0,
  0, 0.001239044, -1.977371e-06, 0.0008456747, 0.01712689, -7.815392e-06, 
    0.007307013, -7.569825e-06, 0, 0, 0, -2.802701e-05, 0.02238886, 
    0.0200111, 0.01146066, 0.001624697, 0.001564666, 0, 0, 0, 0, 0, 0, 0, 
    5.031443e-05, 0.001677033, -2.837593e-05, 0, 0,
  0, -6.746718e-05, 0.004831275, -4.85933e-07, -1.032263e-05, -4.641463e-05, 
    -0.0001034599, 0.006893596, -0.0003360455, 0.003878554, 0.0001696364, 
    0.00229392, 0.00232916, 0.005406597, 0.004299934, 0.01806334, 
    -8.104288e-05, -2.188162e-05, -1.097985e-05, 0, 0, 0, 0, 0.004045213, 
    0.002531223, 0.001038566, 0.0009286992, 0, 0,
  0, 0, 0.005342192, 0, 0.003592822, 0.0002414694, 0.0001032701, 
    -5.577214e-06, 0.001916784, 0.0201235, 0.02197473, 0, 0.003640665, 0, 
    -2.34346e-07, 0, 0, 0, 0, -1.339643e-05, 0, 0, 0, 0.00105552, 0, 
    -0.0001934559, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 8.438948e-06, -5.198565e-05, 0.001154088, 
    -3.674372e-05, 0.001234002, 0, 0, 0, 0.005234224, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0004575093, -8.715991e-06, 0, 0, 0, 0, 
    0, 0.002694346, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0006538601, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 1.865951e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, -1.754822e-05, 0, -5.653981e-07,
  0, 0, 0, 0, 0.00044776, -0.000150096, 0, 4.262123e-06, 0, 0, 0, 
    0.0007172175, 0, -4.097224e-05, 0, 0, -3.080747e-05, 0.0120176, 
    -2.633954e-05, 0, 0, 0, 0, 0, 0.004573252, 0.004148772, 0.0002344725, 0, 0,
  0, 0, -4.028647e-05, -3.226415e-07, 0.01075116, 0.0007708275, 0.01943737, 
    0, 0, 0, 0, 0, 0, 0.01326839, -6.338738e-06, 0.006016058, 0.004227667, 
    -4.538547e-05, -4.774854e-05, 0.0003639823, -2.615046e-05, 0, 0, 0, 
    0.0001897634, -0.0001302886, 0.004463742, 0, 0,
  0, 0.002585485, -5.15952e-05, 0.002215665, 0.02970436, 0.0004995633, 
    0.01465826, 0.0003231976, 0, 0, 0, 0.0009873383, 0.03163616, 0.03068329, 
    0.01583976, 0.002402948, 0.003427746, 0, 0, 0, 0.0003854294, 0, 0, 0, 
    0.000254923, 0.005210597, 0.003571017, 0, 0,
  0, -0.00024263, 0.01096514, -1.848309e-05, -8.418929e-05, 0.001498948, 
    -0.0002604421, 0.01474218, -0.000596157, 0.006206994, 0.001170912, 
    0.007096378, 0.00551942, 0.01372566, 0.006659058, 0.03355681, 
    0.0008489012, -0.0002817751, -0.0001170166, 0, 0, 0, 0, 0.007360684, 
    0.006273042, 0.002278524, 0.004182487, 0, 0,
  0, 0, 0.009577524, 0, 0.006788272, 0.0009685931, 0.0005049578, 
    -5.577214e-06, 0.002093066, 0.03373022, 0.02620498, 0, 0.005700885, 
    0.000130913, -3.995456e-06, -2.535057e-05, 0, 0, 0, -5.014278e-05, 0, 0, 
    0, 0.002994971, -8.044531e-06, 0.001596692, 2.282856e-05, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, -1.489666e-05, -9.357416e-05, 0.005447414, 
    0.00066536, 0.00567447, 0, 0, 0, 0.01315848, 0, 0, 8.639221e-05, 0, 0, 0, 
    0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, -1.928936e-07, 0, 0, 0, 0.00409818, -0.0001698195, 0, 
    0, 0, 0, -3.271041e-05, 0.008480152, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.536296e-05, 0, 0, 0, 0.0003058283, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.00192533, -1.245668e-05, 0, 0, 0, 0, 
    -8.970721e-07, 0, 0, 0, 0, -6.540778e-07, -1.872599e-05, -2.624975e-05, 
    0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0.004747126, -7.752583e-07, -2.469668e-05, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, -2.063404e-05, -9.262325e-06, 0, 0, 0, 0, 0, 0.0001809545, 
    -6.638244e-06, 0.0005695337,
  0, 0, 0, -1.660237e-05, 0.006241412, 0.003148975, -3.982554e-07, 
    0.001412282, 0, 0, 2.951552e-06, 0.001646517, 0.001497073, -0.0002085862, 
    -3.074628e-06, -4.635827e-06, 0.002280472, 0.02340933, 0.001492358, 
    0.0005608495, -1.423673e-05, 0.0008758858, 0, 0, 0.009661114, 0.00874468, 
    0.009842492, -4.041404e-05, 0,
  0, 0, 0.0005297615, -7.214203e-05, 0.01682561, 0.007248395, 0.04488162, 0, 
    0, 0, -9.002408e-05, 0, 0, 0.03611481, 0.0005587231, 0.02209451, 
    0.006334904, 0.0003914964, 0.003091199, 0.005092898, -0.0001554798, 0, 0, 
    0, 0.005155679, 0.001240357, 0.01193629, 0, 0,
  0, 0.0105104, 0.0002741014, 0.01100943, 0.06429746, 0.001951495, 
    0.02068399, 0.001214039, 0, 0, -9.260352e-06, 0.006204152, 0.04435403, 
    0.04653182, 0.0220963, 0.01190764, 0.0126218, -1.896173e-06, 
    -1.283326e-05, 0, 0.002297169, 0, 0, 0, 0.001358334, 0.006924676, 
    0.009190115, 0, 0,
  0, -0.0002892104, 0.01907938, 0.0004483979, 6.443696e-05, 0.006950792, 
    0.0007500495, 0.02794486, -0.0009035025, 0.0079453, 0.002957257, 
    0.009389634, 0.01151209, 0.03995501, 0.02294025, 0.06509709, 0.01267395, 
    0.0003985121, 3.861167e-05, 0, 0, 0, 0, 0.01169988, 0.01715199, 
    0.00483174, 0.008609273, 0, 0,
  0, 7.609522e-06, 0.01110215, 0, 0.009973533, 0.007386826, 0.005781509, 
    -1.115443e-05, 0.003731846, 0.04513646, 0.02894578, -3.663702e-08, 
    0.01387206, 0.0001121191, 0.001245205, 1.988333e-05, 5.012179e-05, 0, 
    -9.678816e-07, -0.0001272614, 0, 0, 0, 0.005284936, 0.0005331761, 
    0.004375583, 2.895694e-05, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0001519367, 4.040876e-05, 0.01108994, 
    0.004635937, 0.0147404, 0.00017263, 0, 0.001198776, 0.02617167, 
    0.0004184901, 0, 0.0004414829, 0, 0, 0, 0, 0, 0, 0, -7.826714e-06,
  0, 0, 0, 0, 0, 0, 0, 0.003752204, 0, 0, 0, 0.009177823, 0.004327995, 
    -9.53856e-06, 6.721827e-05, 0, 0, 0.00447507, 0.01411765, 0, 0, 0, 
    3.535701e-05, 0, 0, 0, 0, 6.628027e-06, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0.002733723, 0.0001973327, 0.004913043, 
    8.230059e-06, 0.001429079, 0, 0, 0, 0.004110227, 0, 0, 0, 0, 0, 0, 0, 
    -6.9536e-07, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, -2.785174e-07, 0.003425441, 0.002260916, 
    0.001747865, -6.713988e-10, -2.488634e-05, -3.513569e-05, -3.264289e-05, 
    -5.480538e-06, 0, 0, 0, -0.0001148376, 0.002570911, 0.0007374746, 
    -5.690835e-06, -1.351347e-05, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, -1.322182e-06, 0, 0, 0, 9.889867e-05, 0, 0, 0, 0, 
    3.355364e-05, 0, 0, 0, 0, 0, 0, 0, 0, -2.689897e-06, 0, 0, 0, 0, 0,
  0.001537597, 0.0001643752, 0, 0.0005458347, 0.01170084, -6.387766e-06, 
    -0.0001115609, 0, 0, 0, 0, 0, 0, 0.0008101513, -1.119705e-14, 
    -8.91166e-05, 0.001181872, 0.003987235, 0.002196208, 0.0003612654, 
    0.001696652, 0.001356009, -3.188793e-05, 3.56465e-05, 0, 0.0002290407, 
    0.007643567, -6.37424e-05, 0.004602101,
  -1.148416e-05, -5.028086e-05, 0, -0.0001527233, 0.00842082, 0.01002249, 
    0.0006515838, 0.007287886, 0, 0, 0.005810634, 0.002729771, 0.01019835, 
    0.002034297, -0.0001170795, -1.746885e-05, 0.01627756, 0.04279695, 
    0.007597736, 0.01125056, 0.0005939719, 0.007268524, 0, 0, 0.01495364, 
    0.01486652, 0.02748245, -0.0001367557, 0.0003626839,
  0, 0, 0.004484474, 0.003103556, 0.02423496, 0.01308866, 0.09136747, 
    -5.871162e-08, 0, 3.658521e-05, -3.516993e-05, -3.640408e-05, 
    -4.304449e-05, 0.04669436, 0.01526121, 0.05615004, 0.01731163, 
    0.002445001, 0.02411393, 0.007137554, 0.001035345, 0, 0, 0, 0.01654623, 
    0.007282821, 0.02762969, 0, 0,
  0, 0.01980721, 0.002310574, 0.0274281, 0.1240255, 0.01127121, 0.02955921, 
    0.003280548, -3.555287e-09, -2.625217e-07, 0.001142955, 0.01132302, 
    0.05257921, 0.05880892, 0.03774901, 0.03404861, 0.04159894, 0.0008925631, 
    0.0004441027, 0, 0.009702796, 0, 0, 0.000111654, 0.004302442, 0.01277472, 
    0.02906302, 0, 0,
  0, 0.002423327, 0.03221904, 0.008630433, 0.007323212, 0.01442894, 
    0.003424755, 0.04070864, 0.01035706, 0.01268627, 0.006494356, 0.01325387, 
    0.02987844, 0.07524747, 0.07604634, 0.0985925, 0.01924539, 0.003753528, 
    0.0008176878, -2.138878e-06, 0, 0, -7.630796e-06, 0.03349467, 0.05582951, 
    0.01183706, 0.009920243, -5.707565e-08, 0,
  0, 0.001959075, 0.0144487, -2.718603e-05, 0.02349733, 0.02078615, 
    0.02002734, 0.0003430881, 0.01764979, 0.08184882, 0.03507784, 
    0.002739479, 0.03980967, 0.01890912, 0.01119089, 0.001118306, 
    0.001864761, 0, 8.005634e-05, 0.0004972601, -5.380889e-07, 0, 
    -9.160003e-12, 0.02525599, 0.002476014, 0.01982159, 5.350883e-05, 
    -6.880957e-06, -3.449154e-11,
  -5.305424e-10, 0, -5.626813e-06, 0, -2.88193e-07, -3.340187e-07, 0, 0, 
    -1.423557e-08, 0.0007788952, 0.001472174, 0.03664861, 0.01543744, 
    0.02394634, 6.685754e-05, -2.337873e-05, 0.005318071, 0.05053524, 
    0.002954619, 0.0002947523, 0.003432459, -8.437312e-05, 2.290147e-06, 
    -3.684564e-10, -1.311575e-06, -5.241443e-08, 0, 0, -2.766748e-05,
  0, 0, 0, 3.536471e-05, 0, 2.915382e-08, 1.182154e-05, 0.008326859, 
    -2.735295e-06, 0, 0, 0.01341909, 0.01101536, 0.0001403796, 0.0009400922, 
    -5.620918e-07, -1.213892e-06, 0.02587502, 0.03089394, -1.152646e-06, 
    3.491543e-06, 0.001050004, 0.002106902, 0, 0, -6.680214e-08, 
    4.468482e-05, 0.003706096, 0,
  0, 0, 0, 0, 0, 0, 0, -2.352205e-05, 0, 0.006871973, 0.004767708, 
    0.01714217, 0.0001444708, 0.004976702, -3.901711e-09, 0, 0, 0.008966741, 
    0, 0, 0, -5.58797e-05, 0, -2.130211e-05, 0, 0.0003855175, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, -4.050735e-05, 0.005554302, 0.008158647, 
    0.004935764, 0.002533582, 0.0004783454, 0.003295739, 0.005604611, 
    0.0008520135, 0, -2.956864e-05, 0, 0.0008358912, 0.01267206, 0.006736086, 
    0.001573157, 4.35646e-05, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -3.448733e-05, 0, 0, 0, -3.167379e-06, 5.953275e-05, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -3.174605e-05, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0.000126138, 0.005398463, -3.656146e-06, 0, 0, 0.002766648, 0, 
    0, -5.49944e-05, -1.198627e-10, 0.01063568, 0, 0.000326623, 
    -6.716255e-05, -5.918638e-05, -7.412689e-06, 3.008566e-05, 0, 
    -2.484724e-05, 0.001067596, 0, 0, 0, 0, 0,
  0.004173639, 0.001051937, 0.0008847503, 0.003632177, 0.02147037, 
    0.004657053, 0.001597739, -6.075512e-06, 0, 0, 0, 0, 0.001142868, 
    0.003476387, 0.003146702, 0.0004098977, 0.003873507, 0.01022311, 
    0.008700199, 0.008898402, 0.006625093, 0.01267192, 0.001522287, 
    0.002583348, 0, 0.008373321, 0.02410206, 0.01003629, 0.01019754,
  -0.0001787108, -9.847913e-05, 9.46667e-08, 0.002098847, 0.01233412, 
    0.02336715, 0.004546292, 0.01203429, -1.929378e-10, 1.100402e-05, 
    0.01322621, 0.01164254, 0.01384802, 0.01048586, 0.001429883, 0.00336256, 
    0.0270719, 0.07825848, 0.0282554, 0.03237586, 0.007189651, 0.01879352, 
    -5.150056e-05, 0, 0.01873546, 0.02767924, 0.05900613, 0.004374369, 
    0.005863916,
  0, 8.875673e-11, 0.008299073, 0.01440139, 0.02624059, 0.02566101, 
    0.1220518, 0.0004574121, 1.918165e-05, 0.000486782, 0.003661588, 
    0.0002521568, 0.001287147, 0.05857829, 0.0833216, 0.1140313, 0.0471945, 
    0.01894755, 0.03721801, 0.01216697, 0.007803243, -0.0001009643, 0, 
    7.524469e-08, 0.0309877, 0.02782382, 0.06737805, -4.164636e-06, 
    -4.691517e-08,
  -6.203394e-09, 0.0383111, 0.01307382, 0.1367488, 0.2344166, 0.07621676, 
    0.06273665, 0.01713393, 9.89724e-06, 0.001898153, 0.01214246, 0.02044165, 
    0.06699383, 0.08627114, 0.1655592, 0.0845193, 0.07500651, 0.004079811, 
    0.00246648, -3.592395e-07, 0.02013481, 0, 0, 0.0311143, 0.08413796, 
    0.02321175, 0.04766738, -2.290244e-07, 0,
  -3.006352e-06, 0.03362506, 0.1146477, 0.03848314, 0.05133939, 0.04548376, 
    0.03975087, 0.07683676, 0.06000527, 0.07058014, 0.01194861, 0.05042267, 
    0.1834281, 0.2875243, 0.3204065, 0.144425, 0.08454353, 0.01692358, 
    0.009800161, -3.073618e-06, 0.0008151152, 1.651917e-08, -1.80582e-05, 
    0.115789, 0.2672044, 0.05615764, 0.0168298, 3.225023e-05, 0,
  -3.050158e-10, 0.01416508, 0.05775666, 0.0002337123, 0.04977266, 
    0.04331654, 0.04982534, 0.01554507, 0.05335211, 0.1551024, 0.05224415, 
    0.04719889, 0.1289048, 0.1375106, 0.1898514, 0.07081091, 0.006008781, 
    0.0004591001, 0.0004614503, 0.0008685294, -5.722111e-06, -6.448656e-06, 
    2.034223e-06, 0.1034875, 0.09769477, 0.100711, 0.006160974, 0.00014742, 
    -1.08654e-05,
  -3.366793e-06, 0, 0.0008115217, 0, -2.123906e-06, -3.360303e-05, 
    4.271865e-05, 4.251829e-08, 0.001754769, 0.01875405, 0.01497054, 
    0.08492629, 0.07721981, 0.04694309, 0.01438748, 0.0077768, 0.01675935, 
    0.0741027, 0.007980385, 0.0008356125, 0.01153058, -7.293683e-05, 
    3.966684e-06, 9.502251e-07, -1.213186e-05, 0.0001817219, 0.0003372626, 
    1.430075e-06, -0.0001129134,
  -1.863204e-11, -8.096588e-08, -1.299648e-09, 4.050647e-05, 5.435783e-10, 
    0.0001699347, 0.003722163, 0.01123085, 0.001188864, 1.347861e-07, 
    8.899731e-07, 0.01666066, 0.02728992, 0.003645637, 0.0006134285, 
    0.0001355204, -0.0001051353, 0.05254005, 0.06239215, 0.0003125183, 
    0.001256632, 0.01051089, 0.007115499, 0, -7.022231e-14, 1.236114e-05, 
    0.0008477163, 0.008985998, -1.19532e-06,
  0, 0, 0, 0, 0, 0, -4.559105e-11, -0.0001205983, -7.108151e-05, 0.01983245, 
    0.01507785, 0.0277853, 0.001445332, 0.007452944, 1.025981e-05, 
    -1.273281e-05, -1.095904e-05, 0.01270081, 0.000420686, 0.0002262779, 
    -3.234896e-10, 0.002948197, 0.0006389841, 0.0002304938, 0.005905703, 
    0.001941812, 0.001054478, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 6.724422e-06, 0.01081434, 0.01185593, 
    0.00814664, 0.01158672, 0.01087983, 0.01073159, 0.008244918, 0.006889034, 
    0.0003205199, -7.809063e-05, 0, 0.001056918, 0.02744502, 0.02053295, 
    0.0124436, 0.00103091, 0, 0, 0,
  0, 0, 0, 0, 0, -2.09344e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.0001951246, 0.0001227108, 0, 9.216907e-06, -5.149557e-05, 
    0.002130544, 6.439961e-06,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.018195e-05, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, -2.45529e-05, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    7.686098e-05, -4.160489e-05, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0001771129, 
    3.224314e-05, 0.0002156762, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  -2.275403e-05, 0, 0, 0, 0.002421854, 0.01509997, 0.0003596647, 
    -5.180988e-06, 0, 0.003207865, 0, 0, 0.004703723, 0.0008425671, 
    0.01504723, -6.433188e-05, 0.003345065, 0.0001153133, 0.00377807, 
    0.0005142424, 0.003443812, 4.608942e-05, 0.002901355, 0.004308291, 
    0.003793189, -4.763115e-05, -6.661797e-05, -6.254666e-06, 0,
  0.008781186, 0.008365462, 0.004504669, 0.009046481, 0.03300568, 0.02020342, 
    0.005041678, 0.002999305, 0.0003485302, -2.672208e-05, -6.169564e-07, 
    -0.0003058662, 0.005356014, 0.005753828, 0.01667557, 0.007038052, 
    0.0128577, 0.01687329, 0.0333585, 0.03406419, 0.0154972, 0.02912431, 
    0.01515551, 0.005988962, 0.0007426809, 0.02669857, 0.03737425, 
    0.02553424, 0.01805774,
  0.01495926, 0.00534108, 0.0001688595, 0.01401888, 0.02626863, 0.03854052, 
    0.02396151, 0.02574753, -4.230387e-05, 0.0001477734, 0.01669464, 
    0.01934146, 0.0200798, 0.02955225, 0.0307277, 0.06359161, 0.05681922, 
    0.1723845, 0.1315648, 0.09059846, 0.05461873, 0.03406478, 0.003286246, 
    0.0002172547, 0.025568, 0.04510534, 0.1178486, 0.04921467, 0.0157847,
  0.001474882, 1.751155e-06, 0.01719055, 0.07215986, 0.08080444, 0.2059052, 
    0.2583361, 0.05952306, 0.04542245, 0.01832868, 0.05489311, 0.02842248, 
    0.008233744, 0.05918926, 0.1037682, 0.1878911, 0.1045161, 0.1662033, 
    0.1549956, 0.03754736, 0.01503825, 0.0002676825, -2.812678e-05, 
    0.0001968812, 0.05116848, 0.07342548, 0.2311153, 0.02753135, 0.0001077359,
  2.743343e-07, 0.0784412, 0.09350565, 0.1355266, 0.230975, 0.1177017, 
    0.08733548, 0.05775186, 0.009289091, 0.009708244, 0.07142369, 0.04010794, 
    0.06757466, 0.08283344, 0.1422666, 0.08329909, 0.1522052, 0.1066808, 
    0.09307928, 0.008436145, 0.03843441, 9.929058e-07, 0.03781448, 
    0.03193456, 0.09590689, 0.1707897, 0.1516542, 0.0835296, 1.141993e-06,
  2.182704e-05, 0.08212031, 0.499267, 0.1576918, 0.05022199, 0.08639161, 
    0.07577846, 0.165364, 0.0904856, 0.09579868, 0.01753731, 0.06980886, 
    0.1685751, 0.2372058, 0.271232, 0.1491909, 0.2365916, 0.08465663, 
    0.06817786, 0.07259195, 0.01045876, 1.870769e-06, 0.001470054, 0.3126027, 
    0.4015369, 0.2850446, 0.1260261, 0.02318176, 7.897307e-05,
  0.0008420497, 0.1589879, 0.4380562, 0.01106488, 0.1352849, 0.1242955, 
    0.1734409, 0.108419, 0.2130862, 0.3342548, 0.08139381, 0.1105718, 
    0.1337042, 0.1409468, 0.1635485, 0.1198256, 0.03260186, 0.0008792616, 
    0.002228444, 0.02053078, 0.01135218, 2.320563e-05, 0.00049983, 0.2498219, 
    0.3204664, 0.2624955, 0.1550938, 0.01199323, 0.0004214101,
  0.03129801, 2.139294e-07, 0.06068935, -5.327956e-10, 3.134198e-05, 
    0.002066313, 0.002562296, 0.01059394, 0.003826659, 0.0303197, 0.05008202, 
    0.1015204, 0.07295597, 0.05240016, 0.01688803, 0.01414207, 0.08182365, 
    0.1944002, 0.06924757, 0.08140725, 0.222931, 0.04859067, 0.01110919, 
    0.0004008854, -6.154943e-05, 0.0164361, 0.001539901, 0.0006685546, 
    0.0005762704,
  0.000473724, 0.0005472902, -5.372379e-05, 0.006650885, 3.198313e-07, 
    0.007947912, 0.02546847, 0.01440722, 0.007512062, 0.01792352, 0.01184836, 
    0.01364591, 0.04974911, 0.006041122, 0.01158185, 0.02285743, 0.00185412, 
    0.1111504, 0.2469753, 0.07389864, 0.09807052, 0.07916613, 0.01482316, 
    -2.195427e-06, 3.494689e-07, 0.001400609, 0.01343433, 0.05894887, 
    0.002523355,
  -1.062938e-09, -7.046367e-09, -4.757728e-06, 8.684761e-08, 1.047525e-07, 
    1.131154e-08, 3.82141e-05, 0.0001424301, 0.0009300793, 0.03998432, 
    0.03494134, 0.04874188, 0.02489535, 0.01388707, 0.007625678, 
    0.0002892338, 0.002701754, 0.01688577, 0.00396271, 0.001235182, 
    -0.0002056147, 0.03268073, 0.02325789, 0.02028587, 0.01651994, 
    0.005347978, 0.007968035, -1.840526e-07, 0,
  -1.492643e-06, 0, 0, 0, 0.0006228526, 0, 1.484066e-05, 0, -8.411657e-07, 
    0.003319826, 0.01418648, 0.02878974, 0.02322016, 0.03585163, 0.02913032, 
    0.02554189, 0.01453086, 0.02134572, 0.00369281, -0.0002163372, 0, 
    0.002049775, 0.03971788, 0.03275775, 0.03588266, 0.01079855, 
    -5.320235e-05, 0, 0,
  0, 0, 0, 0, 0, 0.000587597, 0, 0, 0, 0, 0, 0, 0, -8.218439e-08, 
    -9.644331e-06, -1.003311e-07, 0.0001701931, 0.001633336, 0.0004484009, 0, 
    0, 0, 0.001609673, 0.003564199, 0.0005500821, 0.006694431, 0.00482141, 
    0.003913766, 0.001254969,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.824786e-05, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.001553131, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0005968841, 0.0005284272, 
    3.957853e-06, 0, 0, 0, 0.000232666, 0.0003254468, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, -2.350246e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001304019, 
    0.00134628, 0.01577906, 0.02643472, 0.003880824, 0.005743146, 
    0.0002155858, 0.0009436703, 0.0001902878, 0, 0, -0.0001869895, 0,
  0.0001223808, 0.001203496, -2.077572e-06, 0, 0.004872529, 0.01708851, 
    0.006353167, 3.312185e-05, 0, 0.003354474, 0, 0, 0.01229409, 0.005343805, 
    0.01612443, 0.00189592, 0.007190356, 0.01703858, 0.02251764, 0.01366765, 
    0.01134443, 0.002979837, 0.01101613, 0.01461821, 0.01205939, 
    0.0006995118, 0.00313263, 0.009384151, -0.0001786967,
  0.05075736, 0.0259262, 0.01033239, 0.02164846, 0.07898588, 0.05922127, 
    0.04790099, 0.04748733, 0.005606139, 0.002175884, 3.485032e-07, 
    0.006280801, 0.006940995, 0.0100764, 0.03573698, 0.02887456, 0.03754627, 
    0.02693905, 0.05712524, 0.1170908, 0.09021894, 0.07338601, 0.06430279, 
    0.01833122, 0.01626655, 0.06427398, 0.08876041, 0.07867486, 0.09005659,
  0.0982837, 0.05518845, 0.02986023, 0.04461138, 0.06335426, 0.1425041, 
    0.08662978, 0.07815774, 0.06694344, 0.05786408, 0.06366654, 0.08117575, 
    0.06893859, 0.08145152, 0.04587935, 0.1044235, 0.07113688, 0.2300077, 
    0.1944149, 0.2048082, 0.1733195, 0.1743906, 0.03816636, 0.002104983, 
    0.03860507, 0.09886678, 0.1955774, 0.1603968, 0.06653121,
  0.000345536, 1.082507e-05, 0.04983255, 0.06969223, 0.08631352, 0.1966894, 
    0.2876378, 0.1392671, 0.1057833, 0.04793943, 0.09007481, 0.05826766, 
    0.03464628, 0.05949832, 0.06836154, 0.1908736, 0.09512957, 0.1516557, 
    0.1702629, 0.1027647, 0.111964, 0.02505262, 0.002621014, 1.335677e-06, 
    0.08860151, 0.1059457, 0.2891221, 0.1013105, 0.004739139,
  2.791603e-07, 0.05638983, 0.06716575, 0.1160315, 0.2104258, 0.09001627, 
    0.07868956, 0.04778188, 0.007049796, 0.00500096, 0.06289956, 0.03668048, 
    0.05141246, 0.07018454, 0.1215204, 0.06731587, 0.1342132, 0.08878546, 
    0.07335984, 0.02722004, 0.1524836, 0.01377444, 0.01912699, 0.02303124, 
    0.09248185, 0.1655404, 0.1408239, 0.09589019, 5.383361e-07,
  1.657784e-05, 0.04668173, 0.4705385, 0.136514, 0.02839265, 0.05626912, 
    0.04628758, 0.106206, 0.08102883, 0.07463242, 0.0125267, 0.0529053, 
    0.1316661, 0.2038952, 0.2297816, 0.1503035, 0.1887418, 0.05954589, 
    0.07594429, 0.04785499, 0.002130817, -1.926145e-06, 0.002092818, 
    0.298085, 0.3142474, 0.2453844, 0.08553711, 0.006867826, 1.000702e-05,
  0.0003969049, 0.09987436, 0.3062447, 0.008627218, 0.09805561, 0.0887769, 
    0.1138172, 0.07038039, 0.1696464, 0.2811983, 0.06296694, 0.06774195, 
    0.09493408, 0.09669097, 0.1115878, 0.09386032, 0.02357204, 9.16611e-06, 
    0.005407203, 0.007116305, 0.001308797, 4.751704e-05, 0.001043871, 
    0.1758593, 0.2310296, 0.1921847, 0.119192, 0.005094002, 0.0001304451,
  0.03229114, 2.003515e-06, 0.04152033, 2.628596e-05, -1.272689e-05, 
    0.004484207, 0.001811992, 0.007961384, 0.001907601, 0.0143325, 
    0.02631995, 0.07307158, 0.06045096, 0.06060875, 0.02062265, 0.01498979, 
    0.08169303, 0.1842814, 0.05251484, 0.05441836, 0.1442873, 0.02372023, 
    0.008279541, 0.0003350601, -1.045525e-05, 0.01778668, 0.0001316024, 
    0.003342176, 0.009953771,
  0.07898023, 0.0508234, 0.01919291, 0.001328998, -1.897692e-08, 0.01315197, 
    0.02209959, 0.0296453, 0.02718437, 0.02017572, 0.03158477, 0.02035014, 
    0.06261034, 0.01652867, 0.0383659, 0.0206871, 0.04781799, 0.1099665, 
    0.2566076, 0.05874473, 0.08024128, 0.09197531, 0.01368202, 6.155929e-05, 
    7.075126e-05, 0.01977952, 0.04222359, 0.1214852, 0.1213862,
  8.404233e-06, -1.717329e-06, 0.02556816, 0.0001073448, 0.0004216873, 
    -5.131046e-07, 0.002203152, 0.0003053882, 0.004013124, 0.1060921, 
    0.1571623, 0.1534915, 0.0775251, 0.06674258, 0.1067217, 0.03608521, 
    0.02512964, 0.04695887, 0.06008683, 0.0401439, 0.008104268, 0.1488852, 
    0.151491, 0.1507634, 0.1159877, 0.06251776, 0.02060494, 0.003255417, 
    -7.90367e-08,
  0.0003796369, 0.0002562332, 5.69035e-06, 0.0004087342, 0.007051763, 
    -1.896242e-08, 0.0001166622, -2.71607e-05, -2.955957e-06, 0.01046764, 
    0.02083967, 0.05071501, 0.06663225, 0.06730665, 0.06533397, 0.04570891, 
    0.0378035, 0.05873443, 0.02811137, 0.006408062, 0, 0.004228813, 
    0.05598365, 0.05931563, 0.1043352, 0.07851136, 0.005075575, 0.006192081, 
    0.001035309,
  4.010016e-05, -1.244754e-06, -9.081019e-06, 0.001084743, 0.0008860022, 
    0.001082462, 0, 0, 0, 0, 0, 0, 0.0001106033, 0.0009820829, 0.000151823, 
    0.001608258, 0.00345426, 0.007176626, 0.001390255, 0, 0, 0, 0.003466156, 
    0.00846759, 0.004631825, 0.03086469, 0.01235839, 0.004804441, 0.002801435,
  7.032458e-05, -4.01435e-05, 0, 0.0001036622, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 6.726507e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, -4.535753e-06, 0.004056257, 
    0.003554955, -5.334058e-05,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, -1.036609e-05, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0.0004519843, 0.002413883, 
    0.001807802, 3.232202e-05, -9.965851e-08, 0, 0, 0.001039372, 
    0.0006472924, -1.969111e-05, 0, 0, 0, 0,
  0, 0, 0, 0, 3.479819e-07, 0.0007797487, 0.0005982271, 0, 0, 0, 
    -1.597355e-06, -5.716739e-05, 0, 0, 2.158637e-05, -0.0004281447, 
    0.01692953, 0.02626158, 0.04786168, 0.08319525, 0.04664562, 0.04008379, 
    0.01518331, 0.01958399, 0.002708589, 1.727925e-06, 9.519945e-06, 
    0.0009176381, 0,
  0.01042454, 0.008712718, 0.001790475, 0.005672239, 0.03726545, 0.03778738, 
    0.04009696, 0.03515056, 0.002010974, 0.005768845, 0.005563378, 
    0.0001607271, 0.03029116, 0.02239702, 0.04060216, 0.03064438, 0.03740297, 
    0.04518067, 0.04222632, 0.03436475, 0.02418789, 0.008980868, 0.03435917, 
    0.03997611, 0.04166235, 0.02860661, 0.007033275, 0.01094505, 0.004098518,
  0.1335998, 0.1127964, 0.1132321, 0.1331845, 0.2082221, 0.1603898, 
    0.1257809, 0.1259313, 0.1134624, 0.04015474, 0.04273896, 0.08185605, 
    0.1059202, 0.06702331, 0.07668921, 0.08329059, 0.08932838, 0.05786768, 
    0.1075624, 0.1180864, 0.1592842, 0.1316409, 0.189992, 0.07123218, 
    0.06895735, 0.2048308, 0.1472637, 0.1151038, 0.1465471,
  0.07379045, 0.06990048, 0.03871818, 0.0376384, 0.05883263, 0.137169, 
    0.08633733, 0.09187797, 0.09735613, 0.1032917, 0.1183526, 0.09444814, 
    0.08281022, 0.1328575, 0.1147753, 0.1072419, 0.107934, 0.2415013, 
    0.196917, 0.1966635, 0.186787, 0.1718416, 0.03260886, 0.0136967, 
    0.08023157, 0.1261595, 0.2013901, 0.1645426, 0.06075986,
  1.429008e-05, 1.75664e-05, 0.06802538, 0.06298958, 0.0667822, 0.1622025, 
    0.265097, 0.09613506, 0.07167428, 0.04773981, 0.1074199, 0.05581937, 
    0.03440586, 0.05538768, 0.05053055, 0.1822382, 0.07133342, 0.1472254, 
    0.1458848, 0.1018662, 0.07370453, 0.04385803, 0.000283235, -0.0001316871, 
    0.07620573, 0.1153454, 0.2738095, 0.04695395, 0.001088727,
  -1.204075e-05, 0.047718, 0.05823129, 0.09711016, 0.2007965, 0.0870735, 
    0.06850464, 0.03135607, 0.003460373, 0.003788572, 0.04429859, 0.03626212, 
    0.04165094, 0.07315028, 0.1106213, 0.05083794, 0.1281409, 0.06212043, 
    0.06580096, 0.01594727, 0.1103987, 0.01314023, 0.0079227, 0.01657432, 
    0.08747272, 0.1629565, 0.11971, 0.05797128, 2.302794e-06,
  3.760928e-06, 0.016125, 0.4242306, 0.1242096, 0.02413666, 0.04962813, 
    0.04123292, 0.08975728, 0.07397621, 0.06276484, 0.01081468, 0.05164706, 
    0.1076733, 0.1830432, 0.2209182, 0.1644999, 0.1664025, 0.05861545, 
    0.06402101, 0.01427585, 0.001491208, -9.997713e-07, 0.00586607, 0.29125, 
    0.2827369, 0.2347615, 0.0690236, 0.002786203, 3.821724e-06,
  0.0007110388, 0.06906734, 0.2519535, 0.007601805, 0.07722539, 0.0731765, 
    0.09614871, 0.04437262, 0.1274597, 0.2637957, 0.06005643, 0.02650996, 
    0.09698478, 0.07872821, 0.1010598, 0.07569388, 0.02424333, -1.351737e-06, 
    0.004431314, 0.003831197, 0.001626628, 3.079162e-05, 0.0012675, 0.120918, 
    0.1756307, 0.1553784, 0.102216, 0.006621104, 0.0001836566,
  0.004307233, -1.727281e-06, 0.02986113, 1.353596e-05, -1.064903e-05, 
    0.006961619, 0.002180102, 0.003013347, 0.001804495, 0.01489668, 
    0.02018981, 0.05174302, 0.0517299, 0.05517237, 0.01315244, 0.02844631, 
    0.08184855, 0.173292, 0.02819811, 0.04084504, 0.1066554, 0.02140347, 
    8.186494e-05, 3.041667e-05, -1.533936e-06, 0.02066134, 0.00854447, 
    0.002789148, 0.01994691,
  0.1179492, 0.1395229, 0.01818418, 5.526864e-05, -0.0002254148, 0.02071284, 
    0.01266492, 0.03879423, 0.03386963, 0.03409312, 0.02232215, 0.02616723, 
    0.06472622, 0.03809708, 0.06599637, 0.01475295, 0.05095397, 0.08075028, 
    0.2432318, 0.03131009, 0.06592015, 0.09039445, 0.01578848, 6.487528e-05, 
    0.002412519, 0.03277667, 0.05827362, 0.1300647, 0.1195868,
  0.01001966, 0.005656615, 0.02935744, 0.03282824, 0.004149206, 
    -5.774416e-05, 0.02539864, 0.002573439, 0.01079948, 0.1887638, 0.219604, 
    0.1708113, 0.09664699, 0.09583148, 0.1277562, 0.08748005, 0.077248, 
    0.1264128, 0.06962126, 0.01651607, 0.02980677, 0.1208378, 0.1439674, 
    0.1556206, 0.1057835, 0.1343323, 0.08236145, 0.09629698, 0.03147792,
  0.009065758, 0.02985372, 0.006655619, 0.0006687696, 0.01053017, 
    -1.429089e-05, 0.0002353467, 0.0003407028, 0.002571751, 0.01418674, 
    0.04579586, 0.09511096, 0.1249806, 0.1180567, 0.1224713, 0.1223387, 
    0.09060825, 0.1648868, 0.1014171, 0.0171039, -0.0001051426, 0.006464439, 
    0.08195578, 0.0821633, 0.171532, 0.1552153, 0.1417966, 0.02615268, 
    0.007391644,
  0.004664507, 0.0008510203, -6.482621e-05, 0.004667331, 0.004210673, 
    0.004225371, 0, 0, 0, 0, 0, -8.095231e-06, 0.002584696, 0.003380372, 
    0.01205899, 0.01839128, 0.02743284, 0.06949422, 0.04376704, 
    -2.445821e-06, 6.78736e-05, -9.054518e-06, 0.008293985, 0.02003786, 
    0.02443105, 0.06933407, 0.09309821, 0.03458378, 0.01982205,
  0.004437142, 0.001801762, -3.666578e-06, 0.003159221, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.007100525, -0.0002544317, 0.001803615, -0.000104968, 
    -5.981027e-05, 0, 0, 0, 0, 0, -0.0001155511, 0.02413278, 0.009529327, 
    0.002942651,
  0, 2.471089e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0002406863, 
    0.0005854227, -6.628833e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.21899e-05, 
    -9.497831e-05,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.007670267, 0.01306558, 
    0.01426565, 0.01279175, 0.00478017, -0.0004398355, -7.615774e-05, 
    0.001896065, 0.004772015, -0.0001281789, 0, 0, 0, 0,
  0, 0, 0, 0.0002513029, -0.0001110027, 0.002402725, 0.02893438, 0, 0, 0, 
    -6.006167e-06, 0.0006419905, -0.0001819252, 0.0004396531, 0.003766289, 
    0.01874327, 0.03251527, 0.04009523, 0.1149505, 0.1095239, 0.07385083, 
    0.03981371, 0.009393402, 0.01699776, 0.02508198, 0.009674747, 
    0.004880472, 0.01418519, 0.006222638,
  0.02963847, 0.01810973, 0.01569834, 0.0379836, 0.1007308, 0.08326789, 
    0.09587544, 0.09584154, 0.06226662, 0.0469299, 0.02421538, 0.02278188, 
    0.1030796, 0.1090704, 0.09412796, 0.07058237, 0.06459238, 0.09330433, 
    0.09421545, 0.07226297, 0.04199284, 0.02787328, 0.05564487, 0.06917652, 
    0.1095852, 0.10742, 0.07386082, 0.06179897, 0.02570841,
  0.1577103, 0.1621529, 0.157434, 0.1725951, 0.2271051, 0.1778728, 0.1526295, 
    0.1734841, 0.1590146, 0.1327832, 0.1744816, 0.186985, 0.1616191, 
    0.1122973, 0.1103969, 0.1032155, 0.1226824, 0.111341, 0.1343057, 
    0.1127623, 0.1461616, 0.1288643, 0.2029089, 0.1113835, 0.1040184, 
    0.2418844, 0.1685092, 0.1346658, 0.1457856,
  0.0418021, 0.05464637, 0.03122535, 0.04142067, 0.04976866, 0.1170768, 
    0.08306831, 0.08247848, 0.0874946, 0.1014102, 0.1025556, 0.07176156, 
    0.06844739, 0.1325958, 0.1212862, 0.08044725, 0.09337515, 0.2467661, 
    0.1740059, 0.1721206, 0.1469327, 0.1571153, 0.02447962, 0.01657174, 
    0.0747968, 0.1277352, 0.1937907, 0.1565977, 0.04700467,
  1.702128e-06, 6.994005e-06, 0.06038158, 0.05547025, 0.08418503, 0.1329405, 
    0.2240241, 0.08113603, 0.04706252, 0.03544775, 0.1244326, 0.05761633, 
    0.03254, 0.05115595, 0.03243055, 0.1801216, 0.06080454, 0.1500966, 
    0.1205477, 0.09598857, 0.05531401, 0.03193847, 0.0006098493, 
    -0.000188091, 0.06542224, 0.1184894, 0.2355804, 0.02402587, 3.33348e-05,
  6.383509e-07, 0.03752141, 0.05629852, 0.07433116, 0.1947435, 0.07888724, 
    0.07641406, 0.03263089, 0.002312467, 0.003387479, 0.03175472, 0.03197928, 
    0.03730197, 0.08624188, 0.1171116, 0.04845215, 0.119802, 0.05101229, 
    0.05817696, 0.0105078, 0.05908418, 0.03531051, 0.008568791, 0.01182693, 
    0.07909504, 0.1714907, 0.0973305, 0.01375337, 6.922372e-07,
  -9.665694e-05, 0.00711753, 0.3589297, 0.09972067, 0.01750448, 0.03189857, 
    0.03631964, 0.07173928, 0.06034875, 0.04634725, 0.009246274, 0.05465677, 
    0.08712135, 0.1502681, 0.1994155, 0.1708404, 0.1241794, 0.04885371, 
    0.05145234, 0.001729526, 0.01026844, -2.139995e-06, 0.01659091, 
    0.2513776, 0.2434004, 0.1997538, 0.04958595, 0.0001467196, 4.141632e-07,
  0.0008368078, 0.04468415, 0.1929293, 0.004126287, 0.06287176, 0.05649836, 
    0.06726521, 0.02891015, 0.07659645, 0.207688, 0.05632057, 0.01941161, 
    0.07672437, 0.06087533, 0.08253769, 0.06317315, 0.02208329, 5.245601e-06, 
    0.003256341, 0.0008183743, 0.01344114, 1.216123e-05, 0.0005440313, 
    0.08196753, 0.1186131, 0.1257157, 0.06827215, 0.005190968, 0.0001962785,
  5.353376e-05, 3.842181e-07, 0.02575972, 3.066127e-05, 8.68054e-05, 
    0.005829625, 0.001592059, 0.001033455, 0.002575217, 0.01048198, 
    0.01297847, 0.04117287, 0.04844559, 0.0600285, 0.003584442, 0.02865675, 
    0.09118332, 0.1493264, 0.01037675, 0.03196815, 0.07010217, 0.01811738, 
    0.0001953121, 1.28956e-05, 5.876175e-05, 0.02362896, 0.01807297, 
    0.003636695, 0.02365911,
  0.08291436, 0.10134, 0.007536721, 0.001197315, 0.002424499, 0.01644426, 
    0.003874481, 0.02568721, 0.03113956, 0.04613962, 0.01219012, 0.02850621, 
    0.05831033, 0.05547733, 0.0490169, 0.008651045, 0.03395967, 0.04506419, 
    0.1833402, 0.02949718, 0.05840883, 0.08419538, 0.01729573, 0.0001187878, 
    0.00333124, 0.02541202, 0.02552902, 0.1013194, 0.1343033,
  0.02782127, 0.005198353, 0.02145942, 0.04616686, 0.005939193, 0.0001293828, 
    0.02698808, 0.007697923, 0.02601625, 0.1837291, 0.1924261, 0.1528755, 
    0.09987902, 0.1082825, 0.084476, 0.0675862, 0.07128309, 0.1114099, 
    0.03992914, 0.00379665, 0.03445143, 0.08140107, 0.1205755, 0.1323298, 
    0.0869306, 0.09704701, 0.08590528, 0.08701315, 0.0810957,
  0.07880206, 0.09513691, 0.03414296, 0.00414658, 0.02347181, 0.02054547, 
    0.002319879, 0.03907074, 0.07047465, 0.03844273, 0.05552125, 0.1255214, 
    0.1594381, 0.1219997, 0.1476093, 0.1424476, 0.1186465, 0.2256029, 
    0.1478716, 0.1046308, -6.362394e-06, 0.1011567, 0.1626513, 0.1076819, 
    0.1930223, 0.2185708, 0.153238, 0.02595634, 0.0745229,
  0.06214793, 0.02596144, 0.01112154, 0.04390342, 0.03442256, 0.0128775, 
    3.175174e-05, 0, 0, 0.009617321, 0.001872522, 0.003945426, 0.01316263, 
    0.0165839, 0.0668959, 0.0558131, 0.1439079, 0.1305082, 0.116979, 
    0.02390761, 0.01882139, 0.004992029, 0.03723014, 0.04531394, 0.05610105, 
    0.1528165, 0.2563892, 0.1475812, 0.09326022,
  0.06038246, 0.007394479, 0.001680782, 0.01645543, 7.510911e-05, 
    9.693487e-06, 0, 1.031276e-06, 0, 0, 0, 0, 0, 0, -5.119236e-05, 
    0.03646052, 0.02462939, 0.05201014, 0.001623109, 0.009907059, 
    8.483582e-05, 0, 0, 0, -1.108254e-05, 0.01101107, 0.06156132, 0.0810467, 
    0.05913297,
  -4.264451e-05, 4.824728e-05, 0.0009445921, -3.64776e-05, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.01150533, 0.03508097, 0.030629, 0.02121189, 0.01380277, 
    0, 0, 0, 0, 0, 0, -1.43774e-07, 0.006848007, 0.006113873,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.656277e-11, 0.009199974, 
    0.03726863, 0.03592094, 0.0335832, 0.02091487, 0.01620561, 0.0004089618, 
    -1.463274e-05, 0.004146178, 0.04863732, 0.03505419, -0.002915112, 
    0.0001458675, 0, 0,
  0.01061387, -9.058323e-05, -0.0003351111, 0.002670256, -0.0009311941, 
    0.004495618, 0.05438283, -0.0005636335, -3.547522e-05, -5.562695e-07, 
    -1.040546e-05, 0.0006636982, -0.002050076, 0.08687603, 0.06084236, 
    0.04311468, 0.05639393, 0.07307031, 0.1226598, 0.1040322, 0.0976065, 
    0.1015331, 0.04754686, 0.04240017, 0.08923252, 0.0448724, 0.03174798, 
    0.0139443, 0.02207169,
  0.0670559, 0.05380999, 0.06478283, 0.09204478, 0.1419367, 0.1124174, 
    0.1258305, 0.1201989, 0.1270761, 0.09632798, 0.05580522, 0.1196142, 
    0.1812615, 0.206567, 0.17389, 0.1492022, 0.1834269, 0.153794, 0.1626478, 
    0.1270725, 0.09876803, 0.09405673, 0.1399876, 0.1307628, 0.1852115, 
    0.2028129, 0.1298793, 0.09855402, 0.05937983,
  0.1515318, 0.1770968, 0.2012721, 0.1881566, 0.2167895, 0.1467623, 
    0.1366948, 0.2014685, 0.1807434, 0.1574939, 0.222024, 0.1887603, 0.17908, 
    0.1104228, 0.1130513, 0.09707498, 0.1208405, 0.1280323, 0.1357206, 
    0.1183997, 0.1380344, 0.1374754, 0.1978339, 0.1318624, 0.1008719, 
    0.2326497, 0.1659997, 0.1385775, 0.1337178,
  0.0447857, 0.05058793, 0.02749383, 0.04729066, 0.05009855, 0.09368218, 
    0.04737159, 0.06473719, 0.0591414, 0.07826068, 0.06253623, 0.05504159, 
    0.06686603, 0.1253536, 0.1099987, 0.0675887, 0.08587643, 0.2407184, 
    0.1635348, 0.1550215, 0.1021585, 0.1350988, 0.01857286, 0.0223539, 
    0.07687164, 0.1119535, 0.1743081, 0.1474981, 0.03920609,
  5.40688e-06, 6.066158e-06, 0.0519681, 0.03717494, 0.07632116, 0.1270615, 
    0.212384, 0.07388626, 0.02964232, 0.01752976, 0.1331225, 0.04541861, 
    0.03380344, 0.04765201, 0.0240267, 0.1675013, 0.05104308, 0.1395538, 
    0.1052855, 0.07766613, 0.04427725, 0.0141537, 0.0004994057, 0.0001584675, 
    0.05940864, 0.1155196, 0.2278436, 0.009656159, 7.276861e-06,
  1.548081e-05, 0.02816654, 0.06848983, 0.04797913, 0.1908261, 0.07298987, 
    0.07585797, 0.02148566, 0.002044315, 0.002833165, 0.01568953, 0.03650545, 
    0.03682607, 0.07705911, 0.1054248, 0.06083787, 0.1074814, 0.04206739, 
    0.04338796, 0.008824117, 0.02201385, 0.02668396, 0.01700244, 0.00741713, 
    0.06714652, 0.1775765, 0.09275479, 0.003901364, 3.754597e-09,
  -1.995371e-05, 0.006830727, 0.2961287, 0.08874143, 0.01200284, 0.02043612, 
    0.02745276, 0.06265447, 0.04083199, 0.03872108, 0.01231788, 0.05152423, 
    0.06670652, 0.1084887, 0.1855575, 0.1741108, 0.07743463, 0.04732024, 
    0.0244162, 0.000547345, 0.009125684, -2.571996e-06, 0.00164838, 
    0.1962742, 0.1927033, 0.1727196, 0.03986662, -4.167051e-06, 9.06605e-08,
  0.0009404813, 0.02762128, 0.1556882, 0.005307063, 0.05437743, 0.04458733, 
    0.04097583, 0.01853859, 0.05215088, 0.173985, 0.0563296, 0.01315391, 
    0.05951866, 0.03762708, 0.05549113, 0.03908433, 0.02076219, 7.029895e-06, 
    0.001707313, 0.000421744, 0.001072683, 1.715293e-06, 0.002909826, 
    0.05246713, 0.08056647, 0.0918093, 0.0382435, 0.004455047, 0.0002225933,
  0.0001469271, 5.252498e-07, 0.01679215, 0.001328761, 0.000967863, 
    0.006807552, 0.001578966, 0.0121458, 0.002564098, 0.007692339, 
    0.008101526, 0.03344567, 0.04157346, 0.07286666, 0.001440417, 
    0.006327786, 0.1038401, 0.1303545, 0.005084698, 0.02070873, 0.04725854, 
    0.01414976, 0.0002295574, 6.460859e-06, 0.0001641861, 0.02000082, 
    0.01477772, 0.006701945, 0.029547,
  0.04579576, 0.05333997, 0.003744086, 0.003704978, 0.006503773, 0.005355721, 
    0.003515171, 0.01909238, 0.01887463, 0.03382146, 0.007160195, 0.01749454, 
    0.06525309, 0.0753039, 0.03251605, 0.002575059, 0.02446046, 0.02955348, 
    0.1607196, 0.004034313, 0.05080254, 0.08803145, 0.02406118, 6.206724e-05, 
    0.002486131, 0.01237496, 0.01081222, 0.06754922, 0.08301681,
  0.01672935, 0.006421025, 0.01886997, 0.03053286, 0.004753387, 0.003022854, 
    0.05630618, 0.02059645, 0.05825358, 0.1503134, 0.1731987, 0.1202691, 
    0.1054338, 0.08085706, 0.05194576, 0.06073327, 0.06594279, 0.09060435, 
    0.01677993, 0.001810671, 0.02720877, 0.05128755, 0.1097279, 0.09959678, 
    0.06249549, 0.07762577, 0.06671089, 0.08663575, 0.06209682,
  0.07625898, 0.1061452, 0.04726595, 0.0202721, 0.06716547, 0.1080483, 
    0.007816416, 0.1656457, 0.0970206, 0.04889896, 0.07598998, 0.1606716, 
    0.1678938, 0.1376189, 0.1770548, 0.1496119, 0.1814739, 0.2461318, 
    0.1538349, 0.1207459, 0.02571406, 0.1475623, 0.2066044, 0.1441121, 
    0.2186617, 0.2023484, 0.1016879, 0.01390956, 0.0716682,
  0.06994967, 0.09732136, 0.1100882, 0.1480719, 0.1353446, 0.1010604, 
    0.02051103, 4.761716e-05, 0.003907405, 0.05400511, 0.02115043, 
    0.01733067, 0.03966239, 0.04858249, 0.09714091, 0.09198506, 0.1767853, 
    0.1918688, 0.2197947, 0.04322344, 0.06544192, 0.1026929, 0.09921688, 
    0.06662147, 0.08845159, 0.2078482, 0.3140498, 0.1502688, 0.09808762,
  0.1194777, 0.03281501, 0.03861877, 0.0780713, 0.01921897, 0.04258804, 
    0.02552631, 0.01111103, 0.01151291, -5.740822e-05, 0, 0, 0, 0.0001648397, 
    0.04733937, 0.08551206, 0.1175719, 0.09655629, 0.06598434, 0.07296476, 
    0.01810401, 0.01182278, 1.488624e-05, 0, -4.229464e-05, 0.03768357, 
    0.1076305, 0.1420819, 0.1156317,
  0.02106858, 0.01031476, 0.004777063, 0.001991975, 0.003464416, 0.009506063, 
    0.005715425, -5.522014e-08, -4.029527e-07, 0.0004155087, -3.818824e-07, 
    0, 0, 2.738716e-05, 0.04094997, 0.0456658, 0.05079416, 0.04166288, 
    0.0299579, 0.03351656, 0.0239704, -0.0002134038, 0, 0, 0, 0, 
    -7.562419e-05, 0.03138863, 0.03154277,
  -1.865569e-07, 0, 0, 0, 0, 0, -1.416751e-05, -7.003938e-05, -9.900605e-06, 
    0, 0, 0, 0, 0, 0, 0, -3.144821e-06, -2.05192e-05, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7.355041e-05, 0.04530444, 
    0.05175997, 0.06234319, 0.08989497, 0.03020035, 0.03661925, 0.02027997, 
    0.004310427, 0.03015018, 0.09991075, 0.1080988, 0.03573842, 0.00457408, 
    -0.0004213493, 0,
  0.02983602, 0.0318951, 0.06838485, 0.06477333, 0.008548085, 0.03132273, 
    0.08419307, -0.00220515, -0.001422297, -0.001431011, -4.107653e-05, 
    0.001465335, 0.03157051, 0.1610867, 0.1285693, 0.1098611, 0.1060159, 
    0.1504734, 0.1509744, 0.09648377, 0.1157155, 0.1895079, 0.1083136, 
    0.09397878, 0.1843073, 0.1120552, 0.05000173, 0.01788153, 0.0287804,
  0.1294279, 0.0952111, 0.104375, 0.1339534, 0.1904029, 0.179104, 0.1955051, 
    0.1709158, 0.1853852, 0.1463002, 0.09998049, 0.2017295, 0.2625203, 
    0.2448992, 0.210517, 0.1940422, 0.2337122, 0.2374027, 0.2454006, 
    0.1941574, 0.1991189, 0.1380721, 0.1807786, 0.1842607, 0.205134, 
    0.2332433, 0.1883207, 0.1597879, 0.1229972,
  0.145412, 0.1950564, 0.2145918, 0.1820882, 0.2032414, 0.1345326, 0.1335523, 
    0.2083047, 0.1585428, 0.1550231, 0.2337315, 0.1740604, 0.1719312, 
    0.09376094, 0.09386585, 0.09483946, 0.1272887, 0.1166585, 0.1421068, 
    0.1151769, 0.1267757, 0.1465756, 0.193394, 0.1320781, 0.1016739, 
    0.2482655, 0.1756103, 0.1277548, 0.1368523,
  0.05433502, 0.05237108, 0.03013593, 0.05675499, 0.04719861, 0.08215892, 
    0.03679303, 0.04488554, 0.03101085, 0.05640317, 0.04243889, 0.04493872, 
    0.06330288, 0.1277331, 0.09708057, 0.04862323, 0.07092207, 0.2102672, 
    0.1568327, 0.1507722, 0.08512332, 0.1145428, 0.02127855, 0.01928159, 
    0.04920691, 0.09890248, 0.1519316, 0.128836, 0.04463287,
  2.378756e-06, 4.571279e-06, 0.04624254, 0.03162813, 0.0606074, 0.1211148, 
    0.1739388, 0.04537631, 0.01049006, 0.00876032, 0.1105706, 0.04613191, 
    0.0416883, 0.04614193, 0.02186039, 0.1551112, 0.04254333, 0.1277957, 
    0.08701131, 0.07069308, 0.02972328, 0.009827643, 0.0009559594, 
    0.002877129, 0.060801, 0.09229145, 0.2012622, 0.004554895, 3.238069e-06,
  -1.544392e-06, 0.02784045, 0.07254981, 0.02921915, 0.1749823, 0.06831035, 
    0.07154615, 0.02268087, 0.001820009, 0.003971365, 0.007335119, 
    0.02846407, 0.03981429, 0.06783105, 0.1108588, 0.0838107, 0.09841222, 
    0.04021625, 0.02456187, 0.006131857, 0.001455037, 0.00216365, 
    0.006835161, 0.01116719, 0.05264555, 0.1672094, 0.0763517, 0.0004889425, 
    1.985022e-08,
  -6.140417e-05, 0.005759949, 0.224268, 0.05772875, 0.008129148, 0.01512202, 
    0.01978187, 0.05834758, 0.02887741, 0.03151102, 0.01610576, 0.05988655, 
    0.05806173, 0.08142774, 0.1854883, 0.1740018, 0.0483886, 0.04941379, 
    0.008041252, 0.0003182972, 0.003207057, -6.871442e-07, -2.771386e-05, 
    0.1693998, 0.1644592, 0.1462607, 0.03124565, 0.0001035552, -3.517478e-08,
  0.002427928, 0.02186105, 0.1263194, 0.008346885, 0.04104844, 0.03696148, 
    0.02460347, 0.01382969, 0.04808269, 0.1807658, 0.05684149, 0.01079225, 
    0.0504266, 0.02429253, 0.03761568, 0.02702861, 0.02661739, 7.028902e-06, 
    0.0007952236, 0.0005650181, 0.004264491, 2.242213e-05, 0.005463534, 
    0.03721629, 0.06369054, 0.08703303, 0.02113642, 0.003861929, 0.0004787428,
  0.0001481214, 2.854967e-07, 0.008030019, 0.002156792, 4.425232e-05, 
    0.001887493, 0.001385651, 0.004934607, 0.002124797, 0.00836337, 
    0.007984482, 0.03141567, 0.03658446, 0.08029807, 0.002448867, 
    0.0002152909, 0.07698337, 0.1194594, 0.00436877, 0.01008478, 0.03641262, 
    0.01100988, 0.0001555364, 1.685866e-05, 0.0002575443, 0.02524268, 
    0.01505889, 0.009247662, 0.02494955,
  0.01418229, 0.01841918, 0.003154001, 0.009099449, 0.009392413, 0.000238454, 
    0.006994397, 0.01563235, 0.0166897, 0.02092985, 0.003765413, 0.01615823, 
    0.06656959, 0.07702427, 0.01286234, 0.0008800131, 0.01720824, 0.02444059, 
    0.1181199, 0.001802528, 0.03427405, 0.08093958, 0.01833867, 4.997078e-05, 
    0.001500394, 0.009008872, 0.005961725, 0.03903908, 0.06728685,
  0.01485955, 0.0182647, 0.02047985, 0.01653412, 0.009181174, 0.01043197, 
    0.0669676, 0.03731983, 0.1370405, 0.1350224, 0.1648932, 0.1078152, 
    0.1007711, 0.0687722, 0.03321837, 0.06654454, 0.06037574, 0.06344304, 
    0.01003215, 3.0225e-06, 0.01278546, 0.03537076, 0.0824016, 0.06542219, 
    0.04337954, 0.06001884, 0.0442104, 0.098029, 0.03270793,
  0.05603263, 0.09413099, 0.07309342, 0.04335298, 0.09353165, 0.1241447, 
    0.03377195, 0.1996899, 0.110937, 0.04998488, 0.1206957, 0.1558467, 
    0.1948115, 0.1381167, 0.1656741, 0.1894071, 0.1685956, 0.230881, 
    0.1222098, 0.1421718, 0.08327182, 0.1634405, 0.1900576, 0.1406837, 
    0.2158402, 0.1702818, 0.07002971, 0.002784638, 0.05034102,
  0.07819186, 0.1189818, 0.1520347, 0.1930017, 0.2213523, 0.1837157, 
    0.1048295, 0.003638288, 0.05960869, 0.09524028, 0.06011117, 0.05159939, 
    0.0683408, 0.09336942, 0.1634524, 0.1231239, 0.2150412, 0.2139183, 
    0.2172437, 0.1282852, 0.131445, 0.1350871, 0.1475866, 0.1175507, 
    0.1283451, 0.2011109, 0.2823006, 0.1379538, 0.083005,
  0.1786056, 0.1073594, 0.1132161, 0.1846528, 0.1175544, 0.1117447, 
    0.1294768, 0.07150393, 0.02371434, 0.01753365, 0.01905031, -0.0003935389, 
    -0.0001162211, 0.08119686, 0.2268928, 0.1206499, 0.1625342, 0.1531964, 
    0.1279089, 0.1649628, 0.06308574, 0.03846538, 0.0056351, 3.174614e-08, 
    0.0002297115, 0.06563807, 0.1227096, 0.1768198, 0.1610435,
  0.06514321, 0.08131187, 0.04220581, 0.1103544, 0.1203695, 0.04996936, 
    0.0226418, 0.0171257, 0.01978992, 0.03026335, 0.002773199, 5.759972e-05, 
    0, 0.06123694, 0.1286215, 0.04826357, 0.06779729, 0.04305389, 0.05947109, 
    0.04109079, 0.04659227, 0.009877197, 0, 0, 0.005070387, 1.62812e-05, 
    -0.0003576816, 0.05989061, 0.05723183,
  0.01161436, 0.01129062, 0.008596478, 0.001893738, 0.03041643, 0.03383232, 
    0.03044127, 0.01329, 0.001480373, -0.0001189652, 0, 0, 0, -3.689946e-08, 
    -2.861702e-05, 3.687749e-05, 0.003308297, 0.005557833, 0.003912005, 
    -0.000133151, -9.213217e-06, 0, 0, 0, 0, 0, 0, -0.0001957312, 0.005507942,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.002644943, 0.06332865, 0.09379461, 
    0.1102968, 0.1518612, 0.1045298, 0.05259158, 0.04190214, 0.02196346, 
    0.06026297, 0.1554973, 0.1691074, 0.05023091, 0.02737527, -0.001109299, 0,
  0.1300866, 0.1543662, 0.1947255, 0.1697609, 0.03766404, 0.0589852, 
    0.1174781, 0.003986234, 0.008755236, -0.003130613, 9.887899e-05, 
    0.01064097, 0.09973918, 0.2364667, 0.1796712, 0.1967893, 0.1613205, 
    0.2724523, 0.2694719, 0.1528038, 0.2218158, 0.2421794, 0.2259916, 
    0.177671, 0.295564, 0.1999154, 0.1025015, 0.07632354, 0.1111077,
  0.1737788, 0.183967, 0.1576645, 0.2168864, 0.2242993, 0.2315486, 0.2556188, 
    0.2362577, 0.275566, 0.2861175, 0.1685818, 0.2393977, 0.2619276, 
    0.2497762, 0.2293063, 0.2406663, 0.2313257, 0.2499137, 0.2910997, 
    0.2344591, 0.2790223, 0.2120837, 0.2295803, 0.2396863, 0.2717865, 
    0.2580978, 0.2021932, 0.1636984, 0.1494006,
  0.1423731, 0.1922929, 0.2158778, 0.1834033, 0.2060207, 0.1483847, 
    0.1406024, 0.2140497, 0.1570179, 0.1766952, 0.2280964, 0.1855546, 
    0.1797445, 0.09752534, 0.08961853, 0.1065283, 0.1500514, 0.1221801, 
    0.144059, 0.1260876, 0.1170777, 0.1510967, 0.1722848, 0.1300935, 
    0.1053241, 0.2075439, 0.1626151, 0.1267768, 0.1251744,
  0.04410025, 0.04079305, 0.02919317, 0.06191097, 0.04690706, 0.06947915, 
    0.03253414, 0.03977884, 0.02227914, 0.03386012, 0.0391349, 0.04064625, 
    0.06353255, 0.1272035, 0.09380981, 0.04359981, 0.05136151, 0.1895939, 
    0.1364453, 0.1392312, 0.07398341, 0.09974267, 0.01988574, 0.01796944, 
    0.0381425, 0.08716127, 0.1437262, 0.1114244, 0.03345088,
  1.23371e-06, 1.411119e-07, 0.04514027, 0.03118364, 0.05883913, 0.1154105, 
    0.1410896, 0.04116825, 0.001963901, 0.001613451, 0.1046297, 0.03523212, 
    0.04369688, 0.04676588, 0.02138657, 0.1279841, 0.05015876, 0.1158506, 
    0.07519808, 0.0614626, 0.02206055, 0.01221773, 0.0002319992, 
    0.0004461446, 0.05985013, 0.07887684, 0.183915, 0.002698577, 9.748216e-06,
  -3.972358e-06, 0.02512207, 0.08001875, 0.02552707, 0.168001, 0.06154586, 
    0.07888918, 0.01410496, 0.001239448, 0.005711925, 0.005112372, 
    0.02267565, 0.04949306, 0.06568138, 0.1163304, 0.09601925, 0.1016794, 
    0.03209537, 0.01404137, 0.004954314, 0.0001504853, 1.379236e-05, 
    0.002288127, 0.01232292, 0.04157877, 0.1555972, 0.07166503, 8.013196e-05, 
    -9.03778e-10,
  0.0002522432, 0.006325188, 0.1723689, 0.04132872, 0.006607346, 0.01287903, 
    0.01546099, 0.04595336, 0.0268514, 0.03261133, 0.03416049, 0.07306801, 
    0.04756802, 0.06665537, 0.1937795, 0.1600999, 0.03139595, 0.06167815, 
    0.007254887, 0.0004113222, -8.877207e-05, 2.695892e-07, 0.00062655, 
    0.1368285, 0.1751753, 0.1321964, 0.03373236, 0.0002643406, 3.139831e-08,
  0.004531926, 0.02117402, 0.1150868, 0.01295826, 0.03307396, 0.03519981, 
    0.02122918, 0.01189133, 0.04293948, 0.2207021, 0.05716154, 0.01045791, 
    0.03690024, 0.0171847, 0.03487139, 0.02199321, 0.005428448, 1.055502e-05, 
    0.001609875, 0.000608116, 0.009674313, -6.415835e-07, 0.02556643, 
    0.03884639, 0.07166147, 0.0949254, 0.01406587, 0.005910066, 0.003527677,
  8.886214e-05, 1.096464e-07, 0.001999175, 0.004757514, 0.0001039921, 
    0.002010501, 0.00118527, 0.000726991, 0.001747105, 0.01026826, 
    0.009528744, 0.0342748, 0.03782503, 0.06444884, 0.002276855, 
    0.0005325997, 0.03828667, 0.1141095, 0.003467953, 0.007882329, 
    0.03069935, 0.009071579, 0.0002507569, 7.430758e-06, 0.001604939, 
    0.05190375, 0.01990836, 0.002540257, 0.02232349,
  0.008570044, 0.001986325, 6.454358e-05, 0.01744547, 0.009595661, 
    9.17979e-05, 0.00312018, 0.01424009, 0.01255496, 0.006011849, 
    0.002389489, 0.04000981, 0.05736728, 0.0397536, 0.008159497, 
    0.0001910196, 0.01320766, 0.0118451, 0.1043938, 4.039802e-05, 0.02359325, 
    0.07281081, 0.007147771, 0.0001100341, 0.00106786, 0.008417008, 
    0.0009366553, 0.03914704, 0.05314448,
  0.0123717, 0.02829142, 0.0175997, 0.003352959, 0.02305065, 0.01858268, 
    0.05769325, 0.06500016, 0.2229884, 0.1299418, 0.1569657, 0.08135559, 
    0.09817515, 0.05700171, 0.03597474, 0.0548247, 0.0588604, 0.05677476, 
    0.005528614, -0.0001041895, 0.006930102, 0.03251595, 0.07611187, 
    0.03874757, 0.03615426, 0.04602211, 0.03453419, 0.128844, 0.005718932,
  0.03756008, 0.09945847, 0.09188943, 0.07720698, 0.07750524, 0.1055397, 
    0.06573807, 0.1596237, 0.09599248, 0.06524961, 0.1336489, 0.1440549, 
    0.1978584, 0.1370796, 0.1822218, 0.196518, 0.1559789, 0.2172331, 
    0.100684, 0.1639797, 0.1612725, 0.1549441, 0.1835492, 0.139878, 
    0.2234636, 0.1597756, 0.05818289, 0.0008595224, 0.04108368,
  0.1067726, 0.1396985, 0.1617342, 0.1809016, 0.2292472, 0.2197954, 
    0.1616856, 0.1041117, 0.07308893, 0.1708713, 0.09204016, 0.1173899, 
    0.1518896, 0.2503288, 0.2370254, 0.1788233, 0.2332408, 0.1985524, 
    0.2055438, 0.1828888, 0.1843731, 0.1751733, 0.1703772, 0.1657961, 
    0.1549039, 0.187801, 0.2723285, 0.1553297, 0.1102118,
  0.2361164, 0.1395941, 0.158832, 0.2574562, 0.2746379, 0.2052968, 0.2237931, 
    0.1218817, 0.03105952, 0.02060426, 0.02941371, 0.01700256, -0.002148194, 
    0.1390889, 0.2594188, 0.15798, 0.1705828, 0.1751092, 0.2041294, 0.189527, 
    0.1346017, 0.08689075, 0.07313493, 0.001302542, 0.05024255, 0.1075614, 
    0.1600128, 0.1823878, 0.2321501,
  0.08220466, 0.1585702, 0.1184907, 0.2202539, 0.1991463, 0.1045538, 
    0.06625976, 0.07117369, 0.07166538, 0.0824388, 0.08250692, 0.01432331, 
    0.0385699, 0.1382563, 0.1997493, 0.06229123, 0.09290635, 0.04222187, 
    0.08629001, 0.1061077, 0.08926735, 0.02853841, 0.0007298913, 
    -1.27826e-06, 0.01104619, 0.001949157, -0.0002570215, 0.06711926, 
    0.08542652,
  0.04697203, 0.04390157, 0.05168572, 0.08927253, 0.08409809, 0.06709105, 
    0.05529229, 0.04856949, 0.03013648, 0.01038405, 0.01101178, 0.02068684, 
    0.01807157, 0.01166349, 0.006846324, 0.01809173, 0.02556378, 0.02240496, 
    0.01208595, 0.01275097, 0.001105584, -8.17447e-05, 0, -4.415507e-05, 
    0.0002894979, -3.627093e-06, 0, -0.004460354, 0.04080221,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.036665, 0.1275247, 0.1346545, 
    0.1836983, 0.2575113, 0.1833292, 0.1115979, 0.07387499, 0.04154757, 
    0.1081036, 0.1712369, 0.1686049, 0.07679649, 0.09847445, 0.00450589, 0,
  0.1734669, 0.264466, 0.3541409, 0.2922167, 0.07532494, 0.08795781, 
    0.1198944, 0.04433324, 0.03836789, 0.01791384, -0.0004166529, 0.02009086, 
    0.1352475, 0.3042909, 0.2700989, 0.2219078, 0.2007575, 0.3281195, 
    0.2997827, 0.1782165, 0.2493674, 0.2618868, 0.3359732, 0.249276, 
    0.3488041, 0.2692447, 0.1621193, 0.1239927, 0.228589,
  0.1884059, 0.2455671, 0.2680972, 0.2707251, 0.2143996, 0.2450624, 
    0.2542208, 0.2536168, 0.3028111, 0.3102657, 0.2316794, 0.257246, 
    0.2635263, 0.2458538, 0.2265798, 0.2515326, 0.2327615, 0.2268772, 
    0.319664, 0.2765352, 0.292952, 0.223887, 0.2654849, 0.2537405, 0.2643694, 
    0.2587357, 0.2147876, 0.1847764, 0.1591651,
  0.1557799, 0.2010511, 0.2054033, 0.178842, 0.2127661, 0.1504555, 0.1322414, 
    0.2025648, 0.1605899, 0.1740691, 0.2409497, 0.1687832, 0.1731787, 
    0.09538715, 0.08960807, 0.09802476, 0.1479326, 0.1241849, 0.131944, 
    0.1363419, 0.1320231, 0.1725443, 0.1784267, 0.1214193, 0.1118961, 
    0.2063187, 0.17138, 0.1163771, 0.128639,
  0.04530187, 0.04417529, 0.03182124, 0.05675783, 0.05010917, 0.06319495, 
    0.02757446, 0.0382334, 0.0158101, 0.06367494, 0.03892446, 0.04987426, 
    0.05960819, 0.1289428, 0.07294181, 0.03614934, 0.05030262, 0.179795, 
    0.1295395, 0.116039, 0.06654177, 0.1118251, 0.02137392, 0.01006664, 
    0.03284078, 0.08349334, 0.1336301, 0.09209363, 0.04102286,
  6.056682e-07, 2.117141e-06, 0.04911372, 0.02414056, 0.05885007, 0.1117007, 
    0.1143003, 0.03796095, 6.03074e-05, -0.0002212659, 0.1004119, 0.032878, 
    0.05059042, 0.04691691, 0.02597178, 0.1105925, 0.06778397, 0.1091933, 
    0.06907932, 0.05703885, 0.01781697, 0.009877396, 4.585967e-05, 
    0.0002829642, 0.0599541, 0.06203144, 0.1644105, 0.001914154, 1.885674e-05,
  -1.143784e-05, 0.03201945, 0.08559379, 0.02563159, 0.1610447, 0.05432909, 
    0.08078329, 0.01788573, 0.0007255035, 0.003514202, 0.003535365, 
    0.02561743, 0.06009786, 0.06764883, 0.1152141, 0.11376, 0.1037567, 
    0.02924336, 0.01060634, 0.004505333, 0.0001082311, 1.761949e-06, 
    8.288564e-05, 0.01072236, 0.04034335, 0.1510078, 0.06586688, 
    2.081453e-05, -5.937121e-10,
  0.0003197829, 0.03841013, 0.1434554, 0.0323521, 0.006287903, 0.0116525, 
    0.01223808, 0.04508437, 0.02339864, 0.04825088, 0.03942281, 0.07334235, 
    0.04992754, 0.05772714, 0.1768834, 0.1392046, 0.01996774, 0.06527077, 
    0.007031109, 0.0001758856, -5.400917e-05, -2.225994e-07, 0.002419754, 
    0.1074131, 0.1815436, 0.129695, 0.02622998, 0.000828093, 3.820894e-06,
  0.01922545, 0.02616506, 0.08631436, 0.01468321, 0.03260472, 0.02964236, 
    0.02799077, 0.01056915, 0.05399217, 0.2274674, 0.03991204, 0.01008327, 
    0.03115773, 0.01415439, 0.03654291, 0.01853078, 0.001270532, 
    0.0001438256, 0.002556329, 0.001473165, 0.0007414221, -6.441386e-05, 
    0.06146009, 0.04481991, 0.07685933, 0.1111774, 0.01227642, 0.00914517, 
    0.005544964,
  0.0004103681, 6.586987e-07, 0.004233405, 0.001935961, 0.0005908781, 
    0.003223016, 0.001234691, 0.0002379239, 0.001585224, 0.01114299, 
    0.007669493, 0.03602475, 0.04268574, 0.06993953, 0.001568746, 
    0.0006669094, 0.01912722, 0.1032896, 0.003367742, 0.00869635, 0.01906886, 
    0.008853276, 0.0003997787, 3.741748e-05, 0.003146219, 0.01853616, 
    0.001732116, 0.0003824612, 0.01343416,
  0.01084714, -1.593481e-05, 4.015345e-06, 0.01390711, 0.01990181, 
    0.002233285, 0.0001748763, 0.01472782, 0.01150424, 0.002085753, 
    0.003798828, 0.03882813, 0.04552557, 0.02593577, 0.003554325, 
    0.0001818479, 0.01186103, 0.003326445, 0.09278765, 4.647819e-05, 
    0.02388963, 0.0638893, 0.001200383, 0.0002605416, 0.001246545, 
    0.01059251, 0.0004965222, 0.02782149, 0.03475986,
  0.01422753, 0.02766117, 0.009467476, 0.000150355, 0.0352219, 0.02233657, 
    0.06344891, 0.1014603, 0.2515408, 0.1414086, 0.1402084, 0.06360284, 
    0.1065798, 0.06100611, 0.03644786, 0.04714854, 0.05032283, 0.05473142, 
    0.005197207, 0.0005623556, 0.002861412, 0.042543, 0.07293665, 0.03098472, 
    0.02235545, 0.0336891, 0.02364103, 0.1194494, -2.57045e-05,
  0.02719831, 0.08825023, 0.1007722, 0.1014443, 0.06990261, 0.08275431, 
    0.147467, 0.1272526, 0.07737269, 0.06522292, 0.1412068, 0.1452316, 
    0.1956315, 0.1414574, 0.1794129, 0.1787636, 0.1463761, 0.1959258, 
    0.08639058, 0.1655377, 0.2104446, 0.1720346, 0.177484, 0.1392322, 
    0.235175, 0.1222898, 0.0432627, 0.002952242, 0.02381098,
  0.09621881, 0.138184, 0.1479321, 0.1608815, 0.2170725, 0.2174471, 
    0.1819083, 0.1662988, 0.1124739, 0.2055794, 0.1528749, 0.1750505, 
    0.1795643, 0.2776089, 0.2686803, 0.1805839, 0.2698589, 0.2098687, 
    0.1916982, 0.2052195, 0.1765154, 0.1657439, 0.1970866, 0.1932122, 
    0.1657817, 0.185277, 0.2563437, 0.1785409, 0.1114603,
  0.2536356, 0.1534601, 0.162746, 0.3097981, 0.3200271, 0.2601801, 0.2902749, 
    0.2080991, 0.1322796, 0.04895574, 0.04188659, 0.03112504, 0.08039618, 
    0.2442447, 0.3029521, 0.1920135, 0.176996, 0.2067561, 0.2240985, 
    0.2119658, 0.1567264, 0.1521112, 0.1603916, 0.02318353, 0.1122935, 
    0.1894915, 0.1984548, 0.2100293, 0.2337499,
  0.1448557, 0.2382276, 0.2886485, 0.2686689, 0.3145678, 0.1952588, 
    0.1304156, 0.1307087, 0.1114147, 0.09313718, 0.1045584, 0.09492341, 
    0.1044413, 0.1478747, 0.1817295, 0.0826473, 0.1192098, 0.07982312, 
    0.1277403, 0.2068514, 0.1296408, 0.07299709, 0.1039678, -0.003072961, 
    0.05403405, 0.007813197, 0.00193833, 0.07789946, 0.1325693,
  0.1332255, 0.1454534, 0.1193699, 0.1332187, 0.08029281, 0.06262692, 
    0.06653277, 0.07349246, 0.08089966, 0.08958438, 0.08653676, 0.08019611, 
    0.08226851, 0.08775471, 0.1102352, 0.1010937, 0.09131766, 0.0655045, 
    0.0412668, 0.03029164, 0.01167613, 0.0006061494, 0.0001239099, 
    -0.0002221652, -0.00181842, -6.905691e-05, -0.004382314, 0.03737045, 
    0.1154717,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -0.0006035925, -0.0006035925, -0.0006035925, -0.0006035925, 
    -0.0006035925, -0.0006035925, -0.0006035925, 0,
  -4.678266e-06, 0, 0, 0, 0, -0.0003685764, 0, 0, 0, 0, 0, -5.963342e-05, 
    0.0001606615, 0.08457266, 0.1762862, 0.1587288, 0.2369577, 0.3295046, 
    0.2613517, 0.2158643, 0.1514649, 0.0817484, 0.1844418, 0.1598191, 
    0.1468477, 0.1030617, 0.1412887, 0.03203667, 0.001400164,
  0.2672195, 0.3448693, 0.3849893, 0.3952406, 0.1512702, 0.1230415, 
    0.1263067, 0.1012727, 0.07850026, 0.02608073, 0.008242684, 0.07893975, 
    0.1364672, 0.3132712, 0.2705694, 0.2359821, 0.2307721, 0.3476012, 
    0.3291751, 0.2199611, 0.2503574, 0.26283, 0.3246196, 0.2903496, 0.368426, 
    0.2759824, 0.181837, 0.1633422, 0.2951438,
  0.20037, 0.265359, 0.322096, 0.2816501, 0.2390435, 0.2800786, 0.2999554, 
    0.316935, 0.347566, 0.3263969, 0.2311983, 0.2633269, 0.2685538, 
    0.2389353, 0.2088387, 0.2428542, 0.247676, 0.2594842, 0.3116285, 
    0.2708765, 0.3072611, 0.2434619, 0.2626502, 0.2884936, 0.2724645, 
    0.2648349, 0.1952659, 0.1709866, 0.1627797,
  0.1559775, 0.1998626, 0.2094056, 0.1714834, 0.1890548, 0.1477959, 
    0.1502457, 0.1971296, 0.1793021, 0.1697481, 0.2329583, 0.1980757, 
    0.157438, 0.0893034, 0.08880926, 0.08859554, 0.1517844, 0.1105627, 
    0.1269789, 0.1290885, 0.1368936, 0.1596927, 0.186015, 0.116785, 
    0.1101922, 0.1964396, 0.1429857, 0.1302455, 0.1168775,
  0.04684158, 0.04866017, 0.02357933, 0.06882943, 0.05676813, 0.06307316, 
    0.02210358, 0.04816183, 0.005282784, 0.03489405, 0.03170557, 0.04026494, 
    0.05358214, 0.1260616, 0.07788533, 0.03489868, 0.06647689, 0.1934736, 
    0.1307315, 0.1194127, 0.06516191, 0.09839722, 0.0224541, 0.007848221, 
    0.03170886, 0.08120647, 0.1200732, 0.08284109, 0.05219581,
  4.581371e-07, 1.763032e-07, 0.0566732, 0.01836799, 0.05079104, 0.1169253, 
    0.08552597, 0.02400523, -3.077248e-05, -6.243778e-05, 0.09920292, 
    0.03142316, 0.04174894, 0.04317678, 0.02329526, 0.09119265, 0.07593514, 
    0.08864128, 0.064031, 0.0546115, 0.01753237, 0.01555362, 1.609745e-05, 
    0.0009703182, 0.06260089, 0.04873745, 0.1506262, 0.00129687, 1.230463e-05,
  -1.029829e-06, 0.02340605, 0.09027037, 0.03101262, 0.1683512, 0.0512443, 
    0.0864721, 0.01023984, 0.0004297392, 0.001775962, 0.002901604, 
    0.03057339, 0.06678446, 0.07842357, 0.1433411, 0.1395701, 0.1175321, 
    0.03036926, 0.009693664, 0.004925286, 0.0001873258, 4.366089e-07, 
    4.249983e-06, 0.01429066, 0.04679069, 0.1424995, 0.05527912, 
    1.216955e-05, -1.647153e-09,
  0.005484565, 0.07488919, 0.1288774, 0.04001864, 0.006782318, 0.01211615, 
    0.01097072, 0.04303983, 0.0237317, 0.06273032, 0.04527827, 0.07325983, 
    0.06481348, 0.06126842, 0.1790472, 0.1134891, 0.01642115, 0.06481656, 
    0.0116898, 9.037981e-05, 5.172804e-05, 0.0006620842, 0.008778154, 
    0.1042118, 0.2079165, 0.1311729, 0.02589907, 0.0008260423, 4.648103e-07,
  0.07872206, 0.05602457, 0.07485972, 0.01573085, 0.02800974, 0.02744836, 
    0.02642064, 0.009183566, 0.05441509, 0.2250259, 0.03402237, 0.007607561, 
    0.02985166, 0.01357405, 0.03192692, 0.01868912, 0.002935805, 
    0.0004323359, 0.003146083, 0.01013191, 0.01053594, 0.00151036, 0.1087404, 
    0.05983878, 0.1298667, 0.1157817, 0.01310557, 0.01102459, 0.007344239,
  0.0006001503, 0.001112352, 0.02027128, 0.004149035, 0.0001521328, 
    0.005843513, 0.001443101, 0.0004358911, 0.002287495, 0.01122825, 
    0.01207968, 0.03495489, 0.05576503, 0.08139534, 0.001176201, 
    0.0009850824, 0.005808258, 0.1063075, 0.007923928, 0.01036135, 
    0.01304839, 0.009490164, 0.001101246, 0.001217034, 0.004081904, 
    0.0006058135, 0.0001304257, 1.050845e-05, 0.01390219,
  0.008217392, 7.392872e-06, 1.249616e-05, 0.01020954, 0.01861494, 
    8.370798e-05, 6.936999e-06, 0.01473785, 0.01189471, 0.00512154, 
    0.01312132, 0.03602957, 0.03713964, 0.01480658, 0.002100509, 
    0.0002673244, 0.01319558, 0.006142627, 0.07498113, 8.530715e-06, 
    0.02447111, 0.05960457, 0.0009030343, 0.001878554, 0.001638319, 
    0.01452831, 7.550024e-05, 0.01736846, 0.02302231,
  0.02263771, 0.01350539, -4.439824e-05, 0.0001999972, 0.0418341, 0.02313863, 
    0.08589263, 0.1480844, 0.2588147, 0.1667272, 0.148201, 0.0922294, 
    0.1210217, 0.05704103, 0.02739696, 0.03259274, 0.05525688, 0.05100632, 
    0.01141017, 0.001915764, 0.0004919716, 0.05891778, 0.06830796, 
    0.02828332, 0.01432945, 0.0324741, 0.01931417, 0.07750308, 0.0002844802,
  0.0191162, 0.08252143, 0.09790161, 0.1186388, 0.06704286, 0.06732628, 
    0.2028033, 0.08913098, 0.06893519, 0.05977746, 0.1529282, 0.1455442, 
    0.1695279, 0.1458589, 0.1734601, 0.2001278, 0.1512638, 0.171845, 
    0.06597272, 0.1430576, 0.2024181, 0.1964173, 0.1763117, 0.1492806, 
    0.2475979, 0.1369638, 0.03715983, 0.006341254, 0.01604525,
  0.08798613, 0.1306379, 0.1493927, 0.1571029, 0.2211254, 0.2232419, 
    0.1686207, 0.2388815, 0.1437472, 0.2436815, 0.1714742, 0.1984922, 
    0.1859854, 0.2699268, 0.2826514, 0.2043276, 0.2758052, 0.2259033, 
    0.1770096, 0.1768138, 0.1628962, 0.1615617, 0.2325915, 0.2075294, 
    0.1897606, 0.203348, 0.2724567, 0.1805557, 0.1092248,
  0.2479515, 0.1501492, 0.1668256, 0.3289593, 0.32863, 0.2662187, 0.3005388, 
    0.2732795, 0.2139511, 0.1522317, 0.08038999, 0.0710887, 0.1062293, 
    0.3059792, 0.3059441, 0.1559637, 0.1832251, 0.2132515, 0.2333038, 
    0.2259252, 0.1473702, 0.1833048, 0.2100524, 0.1288081, 0.1910126, 
    0.2476267, 0.2130082, 0.2412909, 0.2422257,
  0.2748796, 0.2997418, 0.3386524, 0.253799, 0.3138565, 0.2387184, 0.2128229, 
    0.1951374, 0.1896347, 0.1464791, 0.1616919, 0.1336582, 0.1339991, 
    0.1224917, 0.1595192, 0.1014149, 0.1504627, 0.1034472, 0.1259129, 
    0.2041744, 0.2061329, 0.07358641, 0.1770793, 0.02820558, 0.09118226, 
    0.01999854, 0.01363616, 0.1208139, 0.2353124,
  0.1848284, 0.1679939, 0.1334184, 0.1352092, 0.06932236, 0.05724258, 
    0.1195239, 0.1177493, 0.1126771, 0.1213358, 0.1311196, 0.1586116, 
    0.1785261, 0.1791684, 0.2044776, 0.2037217, 0.1807989, 0.1436896, 
    0.1411022, 0.1341522, 0.09121242, 0.08042628, 0.02340945, -0.004079978, 
    0.03719165, 0.004974834, 0.003955011, 0.08715986, 0.2901953,
  0.01948665, 0.01714497, 0.01480328, 0.0124616, 0.01011991, 0.007778226, 
    0.005436542, 0.003259401, 0.003207441, 0.003155481, 0.003103521, 
    0.003051561, 0.002999601, 0.002947641, 0.005238319, 0.00703079, 
    0.008823262, 0.01061573, 0.0124082, 0.01420067, 0.01599314, 0.01148495, 
    0.01208612, 0.0126873, 0.01328847, 0.01388965, 0.01449082, 0.01509199, 
    0.02136,
  -0.001379295, -1.435289e-05, 0, 0, -2.573e-06, -0.002710296, -0.0002486106, 
    0, 0, 0, 0, 0.001078875, 0.003975067, 0.132015, 0.1705277, 0.1676577, 
    0.2727205, 0.3320634, 0.2860756, 0.2542961, 0.2518023, 0.2113813, 
    0.240025, 0.1580018, 0.1200572, 0.0807965, 0.1280739, 0.07541315, 
    0.01214056,
  0.3356517, 0.3510031, 0.3619073, 0.4046612, 0.2590648, 0.1724031, 
    0.1297365, 0.1527679, 0.1337747, 0.05241074, 0.05764928, 0.1360606, 
    0.1423797, 0.3260415, 0.2925039, 0.2373425, 0.2490145, 0.344049, 
    0.3066299, 0.2411234, 0.2468995, 0.2709257, 0.3542119, 0.2847058, 
    0.3935161, 0.2535154, 0.2523874, 0.1759061, 0.3238939,
  0.2284022, 0.306738, 0.3329646, 0.2854575, 0.227602, 0.2606517, 0.3145653, 
    0.3482304, 0.3558491, 0.3096683, 0.2484355, 0.2731637, 0.279711, 
    0.2449638, 0.213376, 0.2469919, 0.2427515, 0.2395489, 0.2911166, 
    0.2822412, 0.3049709, 0.2706495, 0.2339509, 0.2568908, 0.281623, 
    0.2600082, 0.192487, 0.1982143, 0.1890986,
  0.1465956, 0.1834828, 0.2148768, 0.185389, 0.1873583, 0.1427009, 0.1466687, 
    0.1688242, 0.1610136, 0.18466, 0.2563695, 0.1873068, 0.165468, 
    0.08434596, 0.08074319, 0.08990005, 0.1661478, 0.1289414, 0.1290306, 
    0.1201404, 0.1137843, 0.1468606, 0.1864603, 0.1233657, 0.1120173, 
    0.1715443, 0.1318061, 0.1335639, 0.1176556,
  0.04608178, 0.04404337, 0.01880552, 0.08854892, 0.0524849, 0.06879587, 
    0.02440755, 0.04399067, 0.01716596, 0.02546871, 0.03406004, 0.03995199, 
    0.04900206, 0.1219336, 0.08182217, 0.04330547, 0.06735167, 0.1952079, 
    0.1195531, 0.09436963, 0.07219771, 0.09035984, 0.02039123, 0.007440849, 
    0.04310447, 0.08095173, 0.117228, 0.07944573, 0.0433363,
  1.766519e-06, -9.780173e-07, 0.0645564, 0.01373295, 0.05000138, 0.1347205, 
    0.07064738, 0.01957623, 6.829962e-07, 0.0004399065, 0.09603727, 
    0.03080312, 0.04907011, 0.04572184, 0.02244339, 0.08217946, 0.08074534, 
    0.07843115, 0.06401673, 0.0456163, 0.0195662, 0.01654747, -1.007013e-05, 
    0.001340062, 0.06001123, 0.04459042, 0.1405596, 0.003001194, 4.437479e-06,
  1.326734e-06, 0.02642961, 0.1056239, 0.04560121, 0.1845132, 0.04649675, 
    0.1018344, 0.006735086, 0.0005580838, 0.002281703, 0.003231235, 
    0.03825986, 0.0691645, 0.07642408, 0.1729731, 0.1483342, 0.1222113, 
    0.03666598, 0.01405079, 0.00543625, 0.0003332622, 7.230553e-07, 
    3.913058e-06, 0.006768648, 0.08495831, 0.1435799, 0.04910637, 
    2.42142e-05, 3.556267e-09,
  0.000129223, 0.0651937, 0.1404803, 0.04849594, 0.01043776, 0.0143357, 
    0.01349023, 0.05401262, 0.0353244, 0.08309347, 0.0427508, 0.06451438, 
    0.09051441, 0.08306675, 0.195923, 0.09747768, 0.01900584, 0.06873255, 
    0.0211086, 0.0006509775, 0.0006153945, 0.0131616, 0.003666352, 0.1316017, 
    0.2545403, 0.1564901, 0.02578355, 0.0009124282, 1.635445e-05,
  0.1007705, 0.1243409, 0.08586972, 0.01766589, 0.03124899, 0.03425094, 
    0.03116911, 0.01270081, 0.073675, 0.2459888, 0.03905933, 0.008738184, 
    0.03874951, 0.01814848, 0.04051035, 0.02669355, 0.00476715, 0.0005969371, 
    0.004911963, 0.01214296, 0.007647627, 0.01087591, 0.1111728, 0.1015097, 
    0.1115435, 0.1386744, 0.01425236, 0.01039822, 0.007667528,
  0.004274002, 0.001423237, 0.04422896, 0.04540727, 9.661577e-06, 
    0.005521544, 0.001851181, 0.0009368818, 0.004199251, 0.01293824, 
    0.02316938, 0.03710371, 0.06824151, 0.08850273, 0.002476716, 0.001744144, 
    0.003787341, 0.09206448, 0.008479683, 0.01408202, 0.0138631, 0.01255013, 
    0.001517754, 0.004001685, 0.005098272, 0.001107164, 0.0001253, 
    0.0001882877, 0.01626499,
  0.002039626, 2.183841e-06, 0.003245476, 0.01418217, 0.01151417, 
    1.359074e-05, 4.735067e-05, 0.01045485, 0.01187156, 0.04103229, 
    0.009214338, 0.03433771, 0.02776717, 0.01216474, 0.0002173577, 
    0.0004966278, 0.02263632, 0.03384195, 0.06135517, 1.290286e-05, 
    0.02756809, 0.07115795, 0.001693143, 0.004404404, 0.002353976, 0.01647, 
    -9.63108e-05, 0.007215168, 0.02324106,
  0.01281702, 0.00300832, 0.001286162, 0.001113221, 0.04862086, 0.02346758, 
    0.1050219, 0.1588217, 0.2533932, 0.1858718, 0.1402626, 0.1019337, 
    0.1325179, 0.05392374, 0.0280259, 0.03100582, 0.05906206, 0.05073849, 
    0.01899297, 0.002639952, 0.004047724, 0.07063047, 0.06373932, 0.02255797, 
    0.01093873, 0.03534289, 0.01806054, 0.0468683, 0.005626745,
  0.01656432, 0.07027236, 0.09936953, 0.1255751, 0.06304094, 0.0550563, 
    0.2030652, 0.05536591, 0.05899817, 0.05678993, 0.1514294, 0.1411005, 
    0.1511178, 0.1405514, 0.1716423, 0.181233, 0.1648735, 0.1616993, 
    0.05419102, 0.120451, 0.2009835, 0.1937905, 0.1621573, 0.1477246, 
    0.2264664, 0.1234292, 0.03073831, 0.0105767, 0.005974145,
  0.07775966, 0.1301078, 0.1525129, 0.1608765, 0.2177957, 0.2342655, 
    0.1621213, 0.2750345, 0.1907681, 0.2448159, 0.178964, 0.2213173, 
    0.1941174, 0.2862703, 0.3113513, 0.2013799, 0.2579662, 0.2409621, 
    0.1574837, 0.1647627, 0.1582801, 0.1601886, 0.2419339, 0.2181834, 
    0.2151912, 0.206584, 0.2648112, 0.178116, 0.09758329,
  0.2664907, 0.139779, 0.1722995, 0.3089553, 0.3156646, 0.2838511, 0.2913834, 
    0.2722377, 0.2237632, 0.1862212, 0.1021132, 0.09292979, 0.1543432, 
    0.3607014, 0.3382458, 0.146124, 0.1858593, 0.2289907, 0.2189809, 
    0.2268722, 0.1405054, 0.1753343, 0.2352528, 0.1418368, 0.2633258, 
    0.2640203, 0.2025012, 0.2250457, 0.2582627,
  0.279584, 0.2867008, 0.3510736, 0.2505629, 0.3026915, 0.2419142, 0.242186, 
    0.2145442, 0.2532277, 0.1891692, 0.1538082, 0.1304813, 0.1351735, 
    0.1285664, 0.1454423, 0.1063022, 0.1464032, 0.1297686, 0.1223077, 
    0.1954051, 0.226438, 0.09139359, 0.2201696, 0.03341474, 0.1609132, 
    0.04557244, 0.02586534, 0.1956016, 0.2182199,
  0.1814853, 0.1517566, 0.114079, 0.1344275, 0.0850976, 0.06270064, 
    0.1367177, 0.1812431, 0.1795036, 0.1776087, 0.1682525, 0.2105689, 
    0.1828641, 0.1992593, 0.2232009, 0.2065459, 0.238179, 0.2243109, 
    0.2049421, 0.226225, 0.1782361, 0.2012865, 0.1507641, 0.04197351, 
    0.09058751, 0.02670691, 0.02514045, 0.2549092, 0.3029723,
  0.07102598, 0.06937036, 0.06771474, 0.06605913, 0.06440351, 0.0627479, 
    0.06109228, 0.0575835, 0.056624, 0.0556645, 0.054705, 0.0537455, 
    0.052786, 0.0518265, 0.03744094, 0.04303411, 0.04862728, 0.05422044, 
    0.05981361, 0.06540678, 0.07099994, 0.08724054, 0.08426248, 0.08128443, 
    0.07830638, 0.07532834, 0.07235029, 0.06937224, 0.07235046,
  0.014405, -0.0001785445, -1.040956e-06, -6.170875e-11, -0.0008826389, 
    0.01111808, 0.006090676, -0.0005593578, 1.908405e-06, 3.573486e-05, 
    -0.001204282, 0.01620335, 0.03879087, 0.15777, 0.1254223, 0.1639969, 
    0.3079684, 0.3492506, 0.2938813, 0.3181429, 0.3466936, 0.3021307, 
    0.2128753, 0.1607942, 0.1403933, 0.1291173, 0.1374376, 0.07954632, 
    0.02605088,
  0.322928, 0.3518443, 0.343824, 0.4222583, 0.3444307, 0.2147987, 0.1398751, 
    0.1849504, 0.160597, 0.1344336, 0.1437234, 0.1688395, 0.1461641, 
    0.3426636, 0.2942844, 0.2293577, 0.3010396, 0.3525595, 0.3384372, 
    0.2583393, 0.2914182, 0.3049082, 0.3676427, 0.32643, 0.4062608, 
    0.2531167, 0.2794345, 0.1554289, 0.3612172,
  0.245636, 0.3489891, 0.3406116, 0.3112971, 0.25779, 0.2608228, 0.3463234, 
    0.3036984, 0.3382367, 0.3406446, 0.2623098, 0.2858507, 0.2612995, 
    0.2503137, 0.2171033, 0.2551063, 0.2767613, 0.2538005, 0.3149216, 
    0.2744411, 0.3053042, 0.2540473, 0.2384721, 0.2674165, 0.2845812, 
    0.2485704, 0.1824038, 0.1984926, 0.2101349,
  0.1473145, 0.1820267, 0.1993339, 0.2088821, 0.1882649, 0.1386517, 
    0.1204449, 0.1662892, 0.1788805, 0.2069332, 0.2704222, 0.2046202, 
    0.1690779, 0.1125128, 0.086336, 0.09441798, 0.1682351, 0.1261395, 
    0.1152411, 0.1248517, 0.1174463, 0.1388697, 0.1926845, 0.1282138, 
    0.1027288, 0.165546, 0.1316722, 0.1329429, 0.1227013,
  0.04579607, 0.04795029, 0.01664152, 0.07202654, 0.04268872, 0.05735242, 
    0.0265073, 0.04041531, 0.01630701, 0.02045941, 0.04619092, 0.04475322, 
    0.04959844, 0.1208856, 0.08051284, 0.05170184, 0.07314632, 0.184597, 
    0.1163987, 0.0892607, 0.08364352, 0.0917673, 0.01925057, 0.009050804, 
    0.06059295, 0.08492634, 0.112557, 0.08156838, 0.04757336,
  3.808338e-05, -1.613819e-06, 0.06680282, 0.0168884, 0.05502475, 0.1579584, 
    0.07266601, 0.02286202, 1.059193e-06, 0.002987354, 0.1052417, 0.02998453, 
    0.07115302, 0.05066508, 0.03787755, 0.08548071, 0.07788749, 0.06945229, 
    0.0798635, 0.04379419, 0.02512978, 0.02187543, 1.513804e-05, 
    0.0002782189, 0.06484241, 0.04475094, 0.153617, 0.00843794, 6.619674e-05,
  6.43973e-05, 0.03906269, 0.113261, 0.05272287, 0.1982471, 0.05429894, 
    0.117893, 0.009555421, 0.001597218, 0.003475222, 0.006154009, 0.04629613, 
    0.07217479, 0.06994475, 0.1684316, 0.1600309, 0.1279494, 0.04581109, 
    0.01514378, 0.006198122, 0.0008203516, 4.713453e-07, 3.72936e-06, 
    0.002912594, 0.0941631, 0.1483681, 0.05390172, 5.864148e-05, 1.555568e-08,
  2.958455e-05, 0.04363593, 0.1746145, 0.06453137, 0.01318472, 0.01598843, 
    0.01694947, 0.0597046, 0.0446837, 0.09552716, 0.04061574, 0.06765709, 
    0.1282157, 0.1053941, 0.2094544, 0.121074, 0.02504924, 0.07499168, 
    0.01759064, 0.001876675, 0.0001716215, 0.01965537, 0.02427551, 0.1627736, 
    0.2891323, 0.1821318, 0.02639534, 0.0005913008, 9.563901e-05,
  0.1098015, 0.1902575, 0.1307245, 0.02920976, 0.02984873, 0.04011406, 
    0.03577637, 0.01622719, 0.07704625, 0.27957, 0.05540093, 0.007446158, 
    0.0478493, 0.02370686, 0.0546135, 0.03275517, 0.004183729, 0.0004405034, 
    0.005016755, 0.01264588, 0.00799151, 0.002998827, 0.1201347, 0.1607089, 
    0.1252297, 0.137653, 0.01369828, 0.009273945, 0.007888043,
  0.01979003, 0.008030726, 0.02903967, 0.1434046, 1.915589e-05, 0.004654353, 
    0.001976444, 0.00122608, 0.00325707, 0.01386715, 0.03019625, 0.03886832, 
    0.07852252, 0.0931559, 0.007650519, 0.001369113, 0.007306859, 0.108055, 
    0.008157866, 0.02081576, 0.015855, 0.01021882, 0.004833033, 0.004756919, 
    0.004688535, 0.001952892, 2.763672e-06, 0.00213817, 0.03766965,
  3.820692e-05, 3.017033e-06, 0.02761145, 0.03041835, 0.003263536, 
    4.437056e-07, 0.001756824, 0.007804618, 0.01983168, 0.03336923, 
    0.002879499, 0.02894842, 0.03509263, 0.01048752, 0.0001698618, 
    0.001643298, 0.02733566, 0.02292963, 0.04986826, 2.1886e-05, 0.04969157, 
    0.07204102, 0.002027281, 0.00329216, 0.006121506, 0.02051174, 
    0.0007339962, 0.00124793, 0.0004323873,
  0.005752136, 0.0007188896, 0.002404841, 0.0002407834, 0.04573727, 
    0.02047163, 0.09658197, 0.1637228, 0.2261069, 0.2104336, 0.1353357, 
    0.1074853, 0.1321785, 0.06374634, 0.03463386, 0.04615675, 0.05265768, 
    0.05568196, 0.02484129, 0.003356864, 0.009263038, 0.06377966, 0.05815578, 
    0.02094032, 0.01758722, 0.04777528, 0.01826612, 0.04558286, 0.005568319,
  0.01762912, 0.05801468, 0.09027512, 0.1361208, 0.06161015, 0.04344933, 
    0.1945902, 0.03642407, 0.04049578, 0.05834547, 0.1487567, 0.1347438, 
    0.149307, 0.1304096, 0.1822355, 0.1776787, 0.1782812, 0.1549404, 
    0.04936317, 0.1125604, 0.2106465, 0.1880368, 0.1819457, 0.1506644, 
    0.2301672, 0.1194576, 0.03370199, 0.008353302, 0.005384053,
  0.0893289, 0.147525, 0.1520523, 0.1976127, 0.2256526, 0.2357648, 0.1682557, 
    0.2968233, 0.1900962, 0.235696, 0.170132, 0.2230312, 0.1758197, 
    0.3086813, 0.3122938, 0.2140336, 0.2632021, 0.2384517, 0.1430678, 
    0.1493476, 0.1425539, 0.1643568, 0.232219, 0.2297285, 0.2213692, 
    0.2133752, 0.2587782, 0.1862428, 0.1060888,
  0.2831594, 0.1431357, 0.1792601, 0.305283, 0.3427425, 0.3053662, 0.305387, 
    0.2939566, 0.2140926, 0.2044811, 0.08994966, 0.1120548, 0.2190007, 
    0.3662958, 0.3502049, 0.1841827, 0.1820478, 0.2353174, 0.2016945, 
    0.224294, 0.1338919, 0.1832885, 0.2418856, 0.1554023, 0.2917702, 
    0.2716815, 0.2046457, 0.2158993, 0.2766585,
  0.267866, 0.2720161, 0.3646649, 0.2589813, 0.3017775, 0.2879507, 0.2406994, 
    0.2248825, 0.2849582, 0.2309162, 0.1586908, 0.1484474, 0.1708905, 
    0.1178798, 0.1313785, 0.1024643, 0.1375272, 0.1366123, 0.115602, 
    0.1961879, 0.2342778, 0.1454001, 0.2165146, 0.0608603, 0.147402, 
    0.09876633, 0.05339198, 0.1724494, 0.2083871,
  0.1643929, 0.1394447, 0.1113905, 0.1356202, 0.1060129, 0.08186631, 
    0.1464344, 0.1821424, 0.2227095, 0.2094531, 0.1982706, 0.2699854, 
    0.1891219, 0.1869554, 0.2064287, 0.2318644, 0.2756473, 0.2237403, 
    0.2167212, 0.2315011, 0.1883228, 0.2145391, 0.2176719, 0.05180254, 
    0.1106468, 0.08594695, 0.07474024, 0.2588258, 0.2905994,
  0.08739972, 0.08723405, 0.08706837, 0.0869027, 0.08673703, 0.08657135, 
    0.08640568, 0.1003769, 0.1051038, 0.1098308, 0.1145578, 0.1192847, 
    0.1240117, 0.1287386, 0.1391175, 0.141325, 0.1435325, 0.14574, 0.1479474, 
    0.1501549, 0.1523624, 0.1213316, 0.1145628, 0.1077941, 0.1010253, 
    0.09425657, 0.08748782, 0.08071906, 0.08753226,
  0.01928135, 0.007921161, 0.0006761605, 5.530166e-05, 0.0006484587, 
    0.03121893, 0.03112524, 0.01302169, 0.0001791837, 0.001311956, 
    0.01989499, 0.0368504, 0.06788551, 0.1622291, 0.1218623, 0.2101938, 
    0.3846735, 0.4088983, 0.3001823, 0.3657868, 0.4037401, 0.3738627, 
    0.204587, 0.1653385, 0.1352791, 0.1356046, 0.1086792, 0.09477473, 
    0.05126037,
  0.3381766, 0.3848143, 0.3761386, 0.4536473, 0.4409175, 0.2518722, 
    0.1668107, 0.2126284, 0.175244, 0.1757868, 0.2008726, 0.1769646, 
    0.1501475, 0.3152294, 0.291419, 0.2642312, 0.3579032, 0.3465962, 
    0.3001299, 0.2511463, 0.2747571, 0.314292, 0.3246555, 0.3673706, 
    0.4462016, 0.28085, 0.2512123, 0.126575, 0.3943286,
  0.2739986, 0.3473046, 0.3771371, 0.3424028, 0.2909767, 0.2997693, 
    0.3673111, 0.3577348, 0.3981322, 0.326111, 0.3167433, 0.3132696, 
    0.2611209, 0.2277995, 0.224277, 0.2503053, 0.2638942, 0.27321, 0.3113831, 
    0.2727761, 0.3294822, 0.2488547, 0.2461203, 0.2837508, 0.3179309, 
    0.2911663, 0.1908633, 0.2128371, 0.2126035,
  0.1632122, 0.2039184, 0.2092524, 0.1989876, 0.1780548, 0.1380074, 0.122277, 
    0.1607712, 0.1751046, 0.1896916, 0.2549363, 0.1980902, 0.1764892, 
    0.09270915, 0.07496581, 0.1071484, 0.1726521, 0.1315097, 0.1176336, 
    0.1312875, 0.1307433, 0.1404638, 0.1857445, 0.1252563, 0.09929939, 
    0.1492383, 0.1250684, 0.1280388, 0.1283543,
  0.05403826, 0.05476234, 0.02102612, 0.07189408, 0.04194511, 0.04838828, 
    0.02981247, 0.03660034, 0.02552531, 0.01921386, 0.05165222, 0.04752597, 
    0.05247775, 0.1235316, 0.09332569, 0.06961229, 0.1004924, 0.1785738, 
    0.1186081, 0.09229647, 0.09478117, 0.08793924, 0.02036848, 0.0111523, 
    0.05037693, 0.08755437, 0.1090819, 0.08161227, 0.05829783,
  0.002526004, -3.024616e-05, 0.07399083, 0.01154083, 0.06586896, 0.1774106, 
    0.08235558, 0.02560924, 2.097966e-06, 0.001909345, 0.106293, 0.044621, 
    0.1252394, 0.07583849, 0.06402934, 0.08026632, 0.07288361, 0.0680713, 
    0.0913662, 0.05344402, 0.03206745, 0.01801069, 5.027543e-05, 
    -2.866556e-05, 0.07069179, 0.05533297, 0.1665431, 0.01753551, 0.000326964,
  0.0004152627, 0.04109625, 0.1245422, 0.03517085, 0.1617617, 0.05052412, 
    0.1279145, 0.01740371, 0.0009821323, 0.003757347, 0.009400936, 
    0.05028431, 0.08064458, 0.06303626, 0.1617808, 0.1428734, 0.1320593, 
    0.03632078, 0.01265663, 0.00540079, 0.001187888, 2.248468e-07, 
    2.036403e-06, 0.0009046855, 0.0770072, 0.1806567, 0.05164187, 
    0.0002515713, 7.629595e-06,
  0.000144821, 0.01340325, 0.2244174, 0.06420686, 0.01284476, 0.01528124, 
    0.01729613, 0.05933596, 0.04429483, 0.08775305, 0.039095, 0.06122849, 
    0.1135952, 0.07355013, 0.1427485, 0.09480805, 0.02403269, 0.06104988, 
    0.0111685, 0.001698095, 4.070863e-05, 0.01726317, 0.01152715, 0.1727646, 
    0.2538786, 0.2133028, 0.02728398, 0.002177171, 4.89806e-05,
  0.03862369, 0.1907088, 0.1584264, 0.03357474, 0.02798698, 0.04243504, 
    0.03038572, 0.01995453, 0.06591672, 0.3013757, 0.07468572, 0.007909435, 
    0.03932296, 0.0187217, 0.04087936, 0.0232055, 0.001965878, 0.0008016928, 
    0.00412667, 0.01395391, 0.02682052, 0.005087132, 0.1216434, 0.1882445, 
    0.1295416, 0.1223354, 0.01320449, 0.01237335, 0.01030742,
  0.01551526, 0.002676362, 0.014817, 0.2081819, 1.522155e-05, 0.002285134, 
    0.00360698, 0.001555444, 0.004668474, 0.0114609, 0.03862949, 0.03505961, 
    0.07336761, 0.08606959, 0.0127269, 0.002331729, 0.01513066, 0.1052127, 
    0.0120537, 0.02479375, 0.01637599, 0.009930904, 0.01005477, 0.007199986, 
    0.005230322, 0.0001878201, 0.0003139343, 0.002757142, 0.0576287,
  7.805167e-06, 2.098578e-06, 0.002548101, 0.04722833, 0.0001137944, 
    1.686755e-07, 0.002944785, 0.009850373, 0.0180393, 0.01789667, 
    0.001295395, 0.02185933, 0.02238695, 0.00361848, 0.0001494875, 
    0.005339644, 0.03053583, 0.01299576, 0.05626492, 2.021939e-05, 
    0.05575654, 0.06943398, 0.002508738, 0.002850151, 0.008468585, 
    0.02883269, 0.001777834, 0.001780386, 1.261612e-05,
  0.002714794, 0.001985953, 0.003316575, 0.0007669898, 0.03006673, 
    0.01858884, 0.06579617, 0.1600527, 0.2040087, 0.2245883, 0.1349321, 
    0.1106054, 0.1199455, 0.05399305, 0.0526012, 0.04970512, 0.06298599, 
    0.06079938, 0.03029118, 0.00417661, 0.01906238, 0.05473624, 0.04889372, 
    0.04101719, 0.02985801, 0.06725989, 0.02330416, 0.02975888, 0.0001693228,
  0.02335648, 0.04439463, 0.08759373, 0.141562, 0.06732697, 0.03112795, 
    0.195715, 0.02038874, 0.02661672, 0.05924355, 0.1395674, 0.1256108, 
    0.1465783, 0.1266045, 0.1740215, 0.1730854, 0.1746505, 0.1470511, 
    0.05813047, 0.1190657, 0.2186652, 0.1778329, 0.1756898, 0.1502215, 
    0.2226212, 0.1320346, 0.03477724, 0.0116105, 0.007975564,
  0.07362696, 0.1410516, 0.1381313, 0.2024864, 0.1971909, 0.2008922, 
    0.1804373, 0.2986576, 0.1712284, 0.2298193, 0.170794, 0.217838, 
    0.1396748, 0.3011697, 0.3330967, 0.23097, 0.2392652, 0.2516246, 
    0.1624795, 0.1457268, 0.1285773, 0.1637759, 0.2244497, 0.2303728, 
    0.2105184, 0.2092935, 0.2634513, 0.1864801, 0.09448636,
  0.2627452, 0.1444439, 0.2338705, 0.3028397, 0.3413727, 0.3013426, 
    0.2624665, 0.3060856, 0.2181172, 0.209752, 0.09972143, 0.09630627, 
    0.2453188, 0.3764147, 0.3638135, 0.1741304, 0.1683266, 0.2634189, 
    0.1948916, 0.2381827, 0.1199535, 0.1874535, 0.2393525, 0.2068659, 
    0.3024645, 0.2848974, 0.2196182, 0.2547907, 0.2968822,
  0.264466, 0.3020601, 0.3660414, 0.2416767, 0.325863, 0.3007253, 0.2561615, 
    0.2642579, 0.2999652, 0.2460771, 0.1846561, 0.1716855, 0.1596511, 
    0.1203332, 0.1193024, 0.1064778, 0.1317303, 0.1426793, 0.1161242, 
    0.1933733, 0.2425645, 0.1492553, 0.2195432, 0.09187273, 0.152556, 
    0.1363167, 0.08312159, 0.150019, 0.1926779,
  0.1351027, 0.1303991, 0.1317272, 0.1491913, 0.1397941, 0.1274326, 
    0.1547703, 0.1753679, 0.2412461, 0.2234948, 0.2595942, 0.2941465, 
    0.2026572, 0.1801559, 0.1922718, 0.2219221, 0.2554769, 0.2242337, 
    0.2143669, 0.2259167, 0.1799356, 0.2163942, 0.1939217, 0.06857981, 
    0.09885146, 0.1023048, 0.1438795, 0.2517839, 0.2914654,
  0.1346407, 0.1336931, 0.1327455, 0.1317979, 0.1308503, 0.1299027, 
    0.1289551, 0.137109, 0.1479435, 0.158778, 0.1696125, 0.180447, 0.1912816, 
    0.2021161, 0.2108168, 0.2094486, 0.2080805, 0.2067123, 0.2053442, 
    0.203976, 0.2026079, 0.1894844, 0.1809656, 0.1724469, 0.1639281, 
    0.1554093, 0.1468906, 0.1383718, 0.1353988,
  0.05033576, 0.02380863, 0.01413197, 0.01344429, 0.0224495, 0.07340929, 
    0.05303349, 0.03571824, 0.01719528, 0.05565667, 0.08329163, 0.1167149, 
    0.1777577, 0.1942721, 0.1293574, 0.3501563, 0.4174471, 0.4304549, 
    0.3076677, 0.371184, 0.4536269, 0.4081814, 0.1916395, 0.1776708, 
    0.1783741, 0.1466539, 0.1283049, 0.1017932, 0.05456242,
  0.4035444, 0.4280886, 0.416326, 0.4901493, 0.4568181, 0.2511479, 0.2047869, 
    0.2336359, 0.1882326, 0.196819, 0.229379, 0.1803986, 0.1573332, 0.320516, 
    0.2790907, 0.2743026, 0.3007553, 0.2838971, 0.2751238, 0.4234205, 
    0.4275753, 0.3242937, 0.3592655, 0.323413, 0.4613332, 0.3102499, 
    0.2708603, 0.1544108, 0.4050705,
  0.3265608, 0.3875609, 0.3658777, 0.3571118, 0.3372106, 0.3099118, 
    0.3444099, 0.3913032, 0.3761084, 0.3577967, 0.3040175, 0.3088568, 
    0.2804565, 0.2619517, 0.2428867, 0.2586006, 0.2925598, 0.2696101, 
    0.3204783, 0.2910548, 0.3291626, 0.2717093, 0.2507046, 0.2897379, 
    0.2937967, 0.2382326, 0.1969721, 0.2424073, 0.2197794,
  0.1697291, 0.2280168, 0.2042927, 0.2289678, 0.1848823, 0.1567931, 
    0.1291489, 0.1699659, 0.1673688, 0.2000038, 0.2606681, 0.2171101, 
    0.1741384, 0.09995869, 0.06807626, 0.1161638, 0.1703214, 0.1411727, 
    0.120237, 0.1392302, 0.1231282, 0.1545461, 0.1831258, 0.1181368, 
    0.08766908, 0.1371692, 0.1429792, 0.1449378, 0.132254,
  0.08135372, 0.06737319, 0.02621822, 0.07944623, 0.05679026, 0.05305578, 
    0.03419754, 0.04004872, 0.03824255, 0.02537788, 0.06157485, 0.0602356, 
    0.06382631, 0.1333909, 0.1073502, 0.08069752, 0.1063404, 0.1818458, 
    0.1278126, 0.100549, 0.103601, 0.08854205, 0.03048941, 0.01390789, 
    0.03889113, 0.08967144, 0.1085371, 0.09027914, 0.06177209,
  0.006773916, 5.368028e-05, 0.07803632, 0.01810741, 0.07415067, 0.1562635, 
    0.1133873, 0.02635703, 3.731489e-05, 0.000199549, 0.0713037, 0.02461988, 
    0.1373377, 0.05267342, 0.0613966, 0.08559005, 0.07617234, 0.06019742, 
    0.07726409, 0.0609558, 0.04293417, 0.02257451, 2.186689e-06, 
    -1.233723e-05, 0.07149146, 0.05066673, 0.1603657, 0.02286995, 0.002742938,
  0.0001462337, 0.03233512, 0.1205952, 0.02368038, 0.1286926, 0.04789059, 
    0.1118694, 0.02550755, 0.001169034, 0.003047615, 0.009101946, 0.06827684, 
    0.08538528, 0.04964281, 0.1590628, 0.1201264, 0.1158322, 0.02593325, 
    0.01200635, 0.008790632, 0.003062939, 2.176391e-07, 4.231564e-07, 
    3.443663e-05, 0.05388564, 0.2089157, 0.03118416, 0.001697407, 0.0003006899,
  2.441397e-06, 0.00398599, 0.2590744, 0.03266887, 0.01108768, 0.01501842, 
    0.01864333, 0.05919318, 0.04107928, 0.0869722, 0.03715396, 0.05790399, 
    0.1090909, 0.05476196, 0.100131, 0.05500148, 0.0240642, 0.04088502, 
    0.009607873, 0.0008437754, 0.003914828, 0.0132329, 0.008551665, 
    0.1184309, 0.1767195, 0.1743137, 0.02817112, 0.005140433, 6.642012e-06,
  0.009563434, 0.1256401, 0.08733553, 0.04026386, 0.02739499, 0.04215515, 
    0.02893787, 0.01963919, 0.05860639, 0.2743214, 0.08617389, 0.008311839, 
    0.03591371, 0.01798322, 0.03375067, 0.01808806, 0.002276463, 0.002738031, 
    0.004682713, 0.01630221, 0.02715175, 0.004128003, 0.08817334, 0.159946, 
    0.08201858, 0.1122056, 0.01837424, 0.01428967, 0.004485246,
  0.002574377, 5.203908e-05, 0.0008941867, 0.2588295, 1.358499e-06, 
    0.001243705, 0.005010899, 0.00159226, 0.005731512, 0.01156993, 
    0.05016121, 0.03565948, 0.06843642, 0.07222595, 0.01186217, 0.005145988, 
    0.01745553, 0.08113049, 0.02124367, 0.02783777, 0.0163698, 0.01100855, 
    0.02350427, 0.01284786, 0.007467736, 0.0002911246, 8.013481e-05, 
    0.0003997143, 0.0298669,
  3.398562e-06, 7.60758e-07, 4.180826e-05, 0.0403757, 0.0001053308, 
    9.310993e-08, 0.0006348731, 0.01129163, 0.01494142, 0.005421034, 
    0.001971527, 0.01910049, 0.01955218, 0.001457403, 0.0002990406, 
    0.007785527, 0.02906419, 0.003978471, 0.03940707, 2.063521e-05, 
    0.01782027, 0.06886244, 0.005192722, 0.006121519, 0.01705044, 0.03139952, 
    0.002391193, 5.761537e-05, 6.247442e-06,
  0.001221171, 0.003014074, 0.008177633, 0.001955378, 0.01798015, 0.01164759, 
    0.03875763, 0.1498613, 0.1843119, 0.2160675, 0.1407304, 0.1206587, 
    0.1193663, 0.04936721, 0.07582566, 0.05613496, 0.06706919, 0.06943238, 
    0.04473538, 0.004863613, 0.02578687, 0.05436476, 0.06434671, 0.06523567, 
    0.03672723, 0.07189139, 0.01877517, 0.01405537, -0.0001852223,
  0.02628227, 0.03071991, 0.08309532, 0.1481707, 0.0654707, 0.0198081, 
    0.1876256, 0.009037322, 0.01814401, 0.06576353, 0.1328767, 0.1204817, 
    0.1534863, 0.1346743, 0.1730665, 0.1808934, 0.1587567, 0.1455196, 
    0.07884198, 0.1384926, 0.2225018, 0.1670818, 0.1747551, 0.1471851, 
    0.2137536, 0.1479812, 0.04632489, 0.01693977, 0.01812376,
  0.07945047, 0.13931, 0.1396486, 0.1986678, 0.1959771, 0.2179616, 0.1712837, 
    0.2648264, 0.1669498, 0.2160328, 0.1494653, 0.2092931, 0.1079353, 
    0.2976893, 0.3272716, 0.23837, 0.2276623, 0.2441439, 0.1709035, 
    0.1518809, 0.1215208, 0.1845219, 0.227389, 0.2129472, 0.194734, 
    0.2024482, 0.2669257, 0.1776654, 0.09454095,
  0.2589271, 0.1421412, 0.1943199, 0.3184284, 0.404154, 0.3173648, 0.3508576, 
    0.335861, 0.2214483, 0.2022767, 0.09426653, 0.08878601, 0.252571, 
    0.3765323, 0.3733722, 0.1735325, 0.1716676, 0.2636647, 0.202899, 
    0.2547469, 0.1088027, 0.2037286, 0.2357539, 0.2195212, 0.2946601, 
    0.3056328, 0.2547438, 0.2598557, 0.3102696,
  0.2756352, 0.3060315, 0.3852304, 0.2570496, 0.3561287, 0.3981453, 
    0.2806528, 0.2833371, 0.3676778, 0.2858995, 0.1864873, 0.1710469, 
    0.1466741, 0.1356277, 0.1190092, 0.1106696, 0.1258835, 0.1418584, 
    0.1192049, 0.2025361, 0.251046, 0.1414013, 0.2113166, 0.07608046, 
    0.1552099, 0.1709449, 0.1169962, 0.1425059, 0.18982,
  0.1364347, 0.1313327, 0.1167493, 0.1629442, 0.1581921, 0.1341433, 
    0.1533412, 0.181307, 0.2497858, 0.2477485, 0.2446528, 0.2692513, 
    0.2065266, 0.1959895, 0.1821521, 0.2518674, 0.2653487, 0.2266328, 
    0.2226485, 0.2129034, 0.1802334, 0.1978159, 0.1677195, 0.05014256, 
    0.08244164, 0.1234155, 0.1718815, 0.2541935, 0.3043617,
  0.1739201, 0.1771531, 0.1803861, 0.183619, 0.186852, 0.190085, 0.193318, 
    0.2194771, 0.2323422, 0.2452073, 0.2580723, 0.2709374, 0.2838024, 
    0.2966675, 0.312312, 0.3080706, 0.3038293, 0.2995878, 0.2953465, 
    0.2911051, 0.2868637, 0.2290854, 0.2172288, 0.2053721, 0.1935154, 
    0.1816588, 0.1698022, 0.1579455, 0.1713337,
  0.05990031, 0.06550848, 0.02706266, 0.04140416, 0.07705063, 0.1074122, 
    0.07488029, 0.0377974, 0.04190833, 0.1058544, 0.1085652, 0.1700867, 
    0.2012106, 0.233398, 0.1113357, 0.300089, 0.4373837, 0.4512299, 
    0.3003052, 0.3515874, 0.4445608, 0.4104406, 0.1892513, 0.2036981, 
    0.1641894, 0.1208497, 0.1306255, 0.1058803, 0.06253227,
  0.4181376, 0.3936252, 0.4540975, 0.5438553, 0.4586293, 0.2373431, 
    0.1948642, 0.2430255, 0.2146899, 0.2012774, 0.2719058, 0.1882322, 
    0.1656147, 0.3322732, 0.2520154, 0.2950969, 0.316691, 0.3222173, 
    0.3142608, 0.3731956, 0.3949187, 0.3091073, 0.325051, 0.339648, 
    0.4039017, 0.3235136, 0.3509595, 0.2082136, 0.3654772,
  0.3591509, 0.4138447, 0.3937138, 0.3580646, 0.3419238, 0.3871276, 
    0.3397682, 0.3815525, 0.4014086, 0.34801, 0.3494166, 0.377457, 0.2823241, 
    0.2574978, 0.2518597, 0.2733897, 0.2824192, 0.2701041, 0.3080186, 
    0.3360268, 0.3202459, 0.2848344, 0.2627019, 0.2981817, 0.3233998, 
    0.2424355, 0.2119345, 0.2487351, 0.2433053,
  0.2088036, 0.2323734, 0.2194446, 0.2183109, 0.180149, 0.153407, 0.1474777, 
    0.1832045, 0.1862831, 0.2134701, 0.271284, 0.2351084, 0.20468, 0.1338721, 
    0.08114766, 0.1399801, 0.1880195, 0.148128, 0.1335559, 0.1652802, 
    0.1374514, 0.14675, 0.2093817, 0.1290742, 0.084853, 0.1213709, 0.1545118, 
    0.1454844, 0.1393625,
  0.08324447, 0.07466479, 0.03644519, 0.09310521, 0.06430088, 0.05099405, 
    0.03689591, 0.0539729, 0.04631741, 0.04108711, 0.1046928, 0.06339629, 
    0.06975077, 0.1401083, 0.1137907, 0.08996113, 0.1066688, 0.1898592, 
    0.1177705, 0.0836853, 0.1112058, 0.09525725, 0.04274387, 0.01794212, 
    0.02369034, 0.09794981, 0.1227839, 0.08583556, 0.06482276,
  0.01039206, 0.0006040944, 0.08954454, 0.02140371, 0.07640166, 0.1520263, 
    0.1193521, 0.02977901, 0.00190417, 0.00114119, 0.03948487, 0.007844299, 
    0.1406469, 0.04042562, 0.05835955, 0.08423996, 0.08562372, 0.06762602, 
    0.07286167, 0.05988673, 0.04772437, 0.02598429, 1.812399e-05, 
    2.89427e-06, 0.07711811, 0.04494653, 0.1249254, 0.02600642, 0.004826528,
  8.741977e-05, 0.02117384, 0.1031746, 0.02329089, 0.1056419, 0.046344, 
    0.09698471, 0.03720254, 0.0006685474, 0.002575447, 0.01156444, 
    0.06702007, 0.08152913, 0.0427732, 0.1481266, 0.08802252, 0.09184807, 
    0.03002786, 0.01672024, 0.02209924, 0.01629324, 1.19705e-05, 
    1.805373e-07, -4.881119e-05, 0.04432625, 0.1951259, 0.0326342, 
    0.01580015, -1.445877e-05,
  1.72069e-06, 0.003871757, 0.1619751, 0.02337125, 0.01043116, 0.01712298, 
    0.02085497, 0.0619146, 0.03774009, 0.08660415, 0.03755046, 0.05611622, 
    0.1099456, 0.04505152, 0.07236248, 0.04649367, 0.02552493, 0.03421745, 
    0.01600713, 0.001764816, 0.0001058314, 0.00772885, 0.00154004, 0.1059092, 
    0.1522877, 0.1462554, 0.03547818, 0.006723943, 3.915005e-06,
  0.003456004, 0.0597938, 0.04427633, 0.05819695, 0.02616825, 0.04259285, 
    0.03358957, 0.02073754, 0.05805278, 0.2492734, 0.08587082, 0.007795829, 
    0.03894009, 0.02036369, 0.03055423, 0.01940213, 0.003400155, 0.0048043, 
    0.008479863, 0.02482385, 0.01456188, 0.003771399, 0.06639719, 0.1346046, 
    0.06335803, 0.1025205, 0.02567215, 0.01398153, 0.003556399,
  0.0004364897, 9.683205e-06, -0.0001088835, 0.235743, -9.250971e-05, 
    0.001477447, 0.006066756, 0.002678992, 0.005011075, 0.01275569, 
    0.05736852, 0.04530297, 0.0697643, 0.06892774, 0.01081725, 0.00571485, 
    0.02132369, 0.06851436, 0.02832192, 0.03529653, 0.02064571, 0.01492697, 
    0.03445717, 0.01980517, 0.01302838, 0.0006339545, 4.524363e-06, 
    4.776032e-05, 0.01093905,
  2.801338e-06, 2.61837e-07, 1.950291e-06, 0.02053369, 1.105424e-05, 
    -1.797993e-08, 2.884878e-05, 0.00618347, 0.01589326, 0.003626671, 
    0.002772517, 0.0188658, 0.02082903, 0.001659565, 0.002267065, 0.01189986, 
    0.02695395, 0.002308988, 0.008800005, 1.894801e-05, 0.0008590386, 
    0.07011972, 0.01101261, 0.01009399, 0.02184976, 0.03149534, 0.002587465, 
    8.962682e-06, 2.30922e-06,
  0.002290493, 0.001856817, 0.04049259, 0.004704393, 0.01045627, 0.008869902, 
    0.01911003, 0.1382338, 0.1673806, 0.2105431, 0.1320923, 0.1215273, 
    0.1241397, 0.04735804, 0.1030331, 0.06717473, 0.07836699, 0.09190758, 
    0.04706503, 0.006219238, 0.03505492, 0.06340977, 0.07521754, 0.08659387, 
    0.05997672, 0.07717673, 0.02324986, 0.01132246, -0.0003938922,
  0.02469099, 0.03171413, 0.08144371, 0.1639123, 0.05581001, 0.02803079, 
    0.1805224, 0.004138531, 0.01074133, 0.06899752, 0.1273392, 0.1225619, 
    0.1618061, 0.1500191, 0.1901365, 0.1855398, 0.167405, 0.183612, 0.086927, 
    0.1361182, 0.2443151, 0.1439122, 0.1811045, 0.1322345, 0.2079603, 
    0.164849, 0.06198911, 0.01932511, 0.02177701,
  0.09920692, 0.1365607, 0.1430447, 0.1828952, 0.1908355, 0.2720661, 
    0.2099166, 0.2394259, 0.1686208, 0.1944438, 0.1454664, 0.1955274, 
    0.09248653, 0.3248737, 0.35774, 0.2289004, 0.2566847, 0.2561362, 
    0.1805874, 0.1750254, 0.1183137, 0.187991, 0.2294397, 0.1900404, 
    0.1870598, 0.2181973, 0.2827952, 0.1754879, 0.09525471,
  0.2331126, 0.1660752, 0.1967687, 0.3145493, 0.4036412, 0.3236039, 
    0.3517851, 0.3002483, 0.2185478, 0.1945395, 0.1264596, 0.07850482, 
    0.2738098, 0.3657267, 0.3636733, 0.1675182, 0.1688543, 0.254993, 
    0.218638, 0.2637712, 0.08508062, 0.1961171, 0.2095573, 0.2176057, 
    0.27296, 0.3187104, 0.2832912, 0.2633999, 0.3007469,
  0.2902573, 0.3118671, 0.3778969, 0.2717355, 0.376866, 0.3520074, 0.3495362, 
    0.324053, 0.4000964, 0.2716761, 0.1862618, 0.1718529, 0.1498694, 
    0.1448512, 0.1182472, 0.1166901, 0.1251436, 0.143695, 0.121401, 
    0.2057399, 0.26385, 0.1363636, 0.2153511, 0.06215889, 0.151911, 
    0.2310529, 0.1543269, 0.1347429, 0.1960021,
  0.194901, 0.1637224, 0.1924253, 0.1780596, 0.147287, 0.1804757, 0.186228, 
    0.1969224, 0.2574318, 0.2391477, 0.2330103, 0.2411142, 0.187219, 
    0.1979607, 0.1879389, 0.2395955, 0.2397062, 0.2007539, 0.220273, 
    0.2063269, 0.1800708, 0.1901621, 0.1550037, 0.03541097, 0.06478375, 
    0.1639526, 0.1717275, 0.2572328, 0.3051236,
  0.1799833, 0.1854659, 0.1909486, 0.1964313, 0.2019139, 0.2073966, 
    0.2128793, 0.2349581, 0.2495499, 0.2641416, 0.2787333, 0.2933251, 
    0.3079168, 0.3225085, 0.3414608, 0.334382, 0.3273031, 0.3202243, 
    0.3131455, 0.3060668, 0.2989879, 0.2455676, 0.232572, 0.2195765, 
    0.2065809, 0.1935853, 0.1805897, 0.1675941, 0.1755972,
  0.0734354, 0.1228403, 0.07242585, 0.0575456, 0.1384725, 0.1437455, 
    0.0866485, 0.05473849, 0.09580711, 0.09499243, 0.2234072, 0.2411996, 
    0.2372611, 0.2283512, 0.1086705, 0.1722656, 0.3262783, 0.3741047, 
    0.3110988, 0.3102012, 0.4579088, 0.388532, 0.2076716, 0.1804907, 
    0.1173803, 0.1051237, 0.1270447, 0.1210633, 0.07409711,
  0.4137875, 0.3322375, 0.3636829, 0.4901541, 0.4513918, 0.2334218, 
    0.1649371, 0.2608394, 0.2389197, 0.2061869, 0.2978175, 0.1891167, 
    0.2089727, 0.2922063, 0.2113346, 0.3245985, 0.3341443, 0.3303966, 
    0.3010588, 0.2831677, 0.285249, 0.2393108, 0.3040794, 0.3855681, 
    0.3775699, 0.2983142, 0.3032783, 0.1629384, 0.3376801,
  0.3685911, 0.4086977, 0.3714003, 0.3791965, 0.3243265, 0.3234703, 
    0.3581394, 0.4152265, 0.4056278, 0.3166949, 0.3514712, 0.3218679, 
    0.2870921, 0.2818593, 0.2512428, 0.2712038, 0.3045957, 0.3124976, 
    0.3225881, 0.3588905, 0.3205247, 0.2931069, 0.2731964, 0.2993182, 
    0.3496645, 0.2406786, 0.2041346, 0.2473379, 0.2461523,
  0.2340802, 0.2324682, 0.2277336, 0.2368074, 0.181326, 0.1550415, 0.1578429, 
    0.1905019, 0.2108588, 0.2176069, 0.306461, 0.2495766, 0.22605, 0.1608609, 
    0.107242, 0.1555767, 0.2404253, 0.1624331, 0.1484815, 0.1992081, 
    0.1553511, 0.1716613, 0.2168813, 0.1347557, 0.09739842, 0.1060895, 
    0.1643315, 0.1660549, 0.1549322,
  0.08090873, 0.09116872, 0.04913744, 0.1101913, 0.07236475, 0.0494586, 
    0.03937085, 0.06666604, 0.06782203, 0.06593113, 0.1131568, 0.0899899, 
    0.05705646, 0.1249817, 0.1177728, 0.09346964, 0.122273, 0.1881018, 
    0.1139628, 0.08130468, 0.1191126, 0.1145628, 0.05125164, 0.02130502, 
    0.009361858, 0.108197, 0.1230686, 0.07976015, 0.05374795,
  0.01853672, 0.001534084, 0.09077621, 0.03194753, 0.07311019, 0.1309984, 
    0.08422821, 0.03713464, 0.006593406, 0.001671923, 0.01753918, 
    0.002886252, 0.1062325, 0.0583524, 0.06927174, 0.08341594, 0.09365159, 
    0.07732912, 0.06736108, 0.06209329, 0.0550859, 0.02893311, 0.001004425, 
    8.029188e-06, 0.07564809, 0.05821471, 0.1031628, 0.03230851, 0.008270847,
  1.821303e-05, 0.01417842, 0.1014748, 0.02706574, 0.09983241, 0.04172892, 
    0.07859799, 0.05099576, 0.000820459, 0.003599779, 0.01211119, 0.06452341, 
    0.09221434, 0.0468432, 0.1316763, 0.06570608, 0.07559781, 0.03283412, 
    0.02917353, 0.03415466, 0.06411546, 0.003146196, 5.224948e-08, 
    -6.614273e-05, 0.04297002, 0.1845979, 0.05421458, 0.06567921, 0.007450783,
  3.248748e-06, 0.002608938, 0.1415161, 0.02117682, 0.01270264, 0.02000647, 
    0.02276462, 0.0643371, 0.03236723, 0.08980966, 0.0471762, 0.05540448, 
    0.1059034, 0.03741865, 0.05705824, 0.0388009, 0.02702819, 0.03253387, 
    0.02802993, 0.009272523, -0.0004452236, 0.003942625, 0.004009342, 
    0.09654984, 0.133147, 0.1332034, 0.04614, 0.00751029, 0.0003333794,
  0.002435679, 0.02794775, 0.04136178, 0.05144883, 0.02861326, 0.03991106, 
    0.03891169, 0.02405628, 0.06523082, 0.2605746, 0.08765992, 0.008139181, 
    0.03699557, 0.02182208, 0.03178118, 0.02391077, 0.007214117, 0.007409262, 
    0.01937531, 0.0280586, 0.01794248, 0.008333595, 0.05631154, 0.1134393, 
    0.05862556, 0.09527642, 0.03189971, 0.01650988, 0.003173331,
  0.0001089207, 2.115948e-06, -9.387878e-05, 0.1581114, 0.0001082979, 
    0.004902985, 0.00919204, 0.003022397, 0.005089477, 0.01372462, 
    0.06302671, 0.05206696, 0.07093979, 0.07451547, 0.01415135, 0.006563824, 
    0.02644557, 0.06475485, 0.03814534, 0.04461683, 0.0258475, 0.018262, 
    0.05255811, 0.02030124, 0.0179295, 0.0005086565, 1.718408e-06, 
    3.709858e-06, 0.003303082,
  2.061196e-06, 8.688978e-08, 3.336874e-07, 0.005958835, 1.308398e-05, 
    -9.886309e-08, -1.626502e-07, 0.002602066, 0.01575981, 0.001070797, 
    0.005134697, 0.01887468, 0.03417588, 0.008944469, 0.009858792, 
    0.01895552, 0.0257091, 0.003582216, 0.001198161, 9.128407e-06, 
    0.0003252086, 0.08329128, 0.01552888, 0.01280618, 0.02336796, 0.03389131, 
    0.006645998, -1.758342e-05, 1.799097e-06,
  0.01119338, 0.004418329, 0.05670774, 0.007303603, 0.008626414, 0.003121864, 
    0.005122694, 0.1225251, 0.1491406, 0.2038857, 0.133553, 0.1171316, 
    0.1320961, 0.04952773, 0.1208582, 0.07725976, 0.07629211, 0.1101562, 
    0.04911584, 0.008635575, 0.05441589, 0.082602, 0.08005474, 0.09099654, 
    0.06500138, 0.0692802, 0.04379085, 0.003579071, -9.837772e-05,
  0.02080612, 0.03365432, 0.08260283, 0.18121, 0.04342593, 0.01361923, 
    0.17314, 0.003950777, 0.0125329, 0.07123521, 0.1271907, 0.1216815, 
    0.1614656, 0.1761294, 0.204608, 0.2007712, 0.1993008, 0.234153, 
    0.1159136, 0.1401655, 0.2058495, 0.1424252, 0.192697, 0.1142322, 
    0.2251974, 0.1960706, 0.08509742, 0.04507055, 0.02184728,
  0.1069924, 0.1489557, 0.156214, 0.1939727, 0.1568062, 0.2106707, 0.2084293, 
    0.2111298, 0.1524784, 0.1671909, 0.143544, 0.174052, 0.0872557, 
    0.3781399, 0.3256794, 0.215793, 0.2271013, 0.2533949, 0.1890624, 
    0.1810855, 0.1228079, 0.1777458, 0.1984345, 0.1763506, 0.208456, 
    0.2591451, 0.2967293, 0.172969, 0.1034986,
  0.2310819, 0.158671, 0.1720492, 0.3358344, 0.414051, 0.3438891, 0.2841333, 
    0.2669641, 0.2115594, 0.2024443, 0.1578913, 0.07320564, 0.3003715, 
    0.3440288, 0.344611, 0.1821444, 0.1899485, 0.2642733, 0.2349852, 
    0.2486529, 0.08650742, 0.1812168, 0.2035543, 0.2120548, 0.2754748, 
    0.3543522, 0.2977475, 0.2692721, 0.2972974,
  0.3151858, 0.3061277, 0.3452789, 0.2601401, 0.3324042, 0.3066001, 
    0.2977315, 0.3511316, 0.4287685, 0.3048368, 0.1963083, 0.1837044, 
    0.1801692, 0.1546432, 0.1178885, 0.1162123, 0.1257142, 0.1378435, 
    0.1252348, 0.2003646, 0.2881024, 0.1297062, 0.1975126, 0.06516114, 
    0.1556263, 0.3094177, 0.1853264, 0.1490462, 0.1851968,
  0.2270209, 0.198865, 0.1757459, 0.1748275, 0.2234611, 0.1855828, 0.1577188, 
    0.2103918, 0.2735125, 0.2377543, 0.2531295, 0.2552096, 0.2115855, 
    0.2124921, 0.1910127, 0.2074638, 0.2286932, 0.1947793, 0.2031989, 
    0.2091326, 0.1939045, 0.204478, 0.1540234, 0.02599318, 0.05634103, 
    0.1509309, 0.1586162, 0.2412829, 0.2961952,
  0.1714773, 0.1784899, 0.1855025, 0.1925152, 0.1995278, 0.2065404, 0.213553, 
    0.2352182, 0.250325, 0.2654317, 0.2805384, 0.2956452, 0.3107519, 
    0.3258587, 0.3511084, 0.3422759, 0.3334435, 0.324611, 0.3157786, 
    0.3069461, 0.2981137, 0.2323419, 0.219055, 0.2057681, 0.1924812, 
    0.1791943, 0.1659074, 0.1526204, 0.1658672,
  0.08743396, 0.1434198, 0.1094014, 0.07717911, 0.1593049, 0.174862, 
    0.0992462, 0.08444827, 0.1270301, 0.2050267, 0.301465, 0.2838867, 
    0.2884894, 0.1818548, 0.1874319, 0.1809561, 0.2796945, 0.3329774, 
    0.2630107, 0.3045259, 0.4795322, 0.3959395, 0.2286344, 0.1704905, 
    0.1038078, 0.08399617, 0.1260615, 0.1642013, 0.1231087,
  0.3815252, 0.3078581, 0.2729048, 0.4900723, 0.4533081, 0.2287139, 0.183379, 
    0.2948196, 0.2477664, 0.2048663, 0.2917859, 0.1872887, 0.2383265, 
    0.3378621, 0.2265355, 0.3175286, 0.3073938, 0.2911368, 0.3083364, 
    0.2667795, 0.3078948, 0.2110155, 0.2471847, 0.3598927, 0.3609077, 
    0.2519342, 0.2339448, 0.164047, 0.3069352,
  0.3377321, 0.369042, 0.3365916, 0.4011871, 0.2942402, 0.3048551, 0.3713805, 
    0.4123112, 0.387899, 0.3246301, 0.31519, 0.3012804, 0.3017898, 0.2923605, 
    0.2796443, 0.2943294, 0.3165903, 0.3039344, 0.335912, 0.3431507, 
    0.3317783, 0.3157212, 0.2737492, 0.308565, 0.2918947, 0.2387302, 
    0.2135744, 0.2426605, 0.3119965,
  0.2263432, 0.2850532, 0.2145645, 0.2391278, 0.1847131, 0.1619125, 
    0.1639307, 0.1954882, 0.2256029, 0.2416708, 0.3231735, 0.2674266, 
    0.2278197, 0.1427836, 0.114989, 0.1883038, 0.2530834, 0.1944312, 
    0.1763815, 0.1929341, 0.1698644, 0.2057368, 0.2362799, 0.1453013, 
    0.09526315, 0.1029766, 0.1660418, 0.201668, 0.1843134,
  0.08446227, 0.1028791, 0.07034367, 0.121982, 0.09770773, 0.06976489, 
    0.04915536, 0.06914721, 0.09129205, 0.1069265, 0.1203524, 0.1002086, 
    0.06044402, 0.1219844, 0.1171406, 0.08738797, 0.1339747, 0.2065971, 
    0.1201565, 0.07915209, 0.1100102, 0.1392021, 0.06885339, 0.02415081, 
    0.004961127, 0.105426, 0.1279278, 0.07192189, 0.06251422,
  0.02751534, 0.003215634, 0.09121405, 0.0357858, 0.06550433, 0.1117534, 
    0.09065294, 0.03324343, 0.009485859, 0.002520525, 0.007989984, 
    0.001197904, 0.06571863, 0.09248101, 0.0851443, 0.09512305, 0.1062083, 
    0.06894007, 0.06868427, 0.06825425, 0.0571449, 0.03954701, 0.001783561, 
    1.809854e-06, 0.07136276, 0.06544985, 0.09315061, 0.04673347, 0.01998696,
  0.0008649562, 0.008915436, 0.108181, 0.03579181, 0.0911628, 0.0344585, 
    0.06884105, 0.05331581, 0.001177058, 0.006343, 0.009755038, 0.06012872, 
    0.09475058, 0.04651623, 0.1125262, 0.05031961, 0.0717812, 0.0299909, 
    0.02704119, 0.03795318, 0.09846788, 0.03656575, 8.766739e-06, 
    -3.367276e-05, 0.05920196, 0.1910627, 0.03605468, 0.06943202, 0.0286283,
  5.737129e-06, 0.0008032004, 0.1357979, 0.0226809, 0.01358033, 0.01977618, 
    0.02649973, 0.06244542, 0.02654166, 0.08564009, 0.05934266, 0.05641384, 
    0.1064105, 0.03207648, 0.04739846, 0.03108095, 0.02383085, 0.03158714, 
    0.02864981, 0.01886501, 0.006177539, 0.005949461, 0.005112897, 
    0.09076367, 0.1212886, 0.1245628, 0.0557623, 0.01106192, 0.004028699,
  0.002033749, 0.02045946, 0.04233164, 0.03954748, 0.03305899, 0.03912213, 
    0.03900147, 0.02313604, 0.07854518, 0.2561806, 0.07567374, 0.01057597, 
    0.03486188, 0.02143028, 0.0303977, 0.02516676, 0.01122153, 0.01105849, 
    0.02143887, 0.02861611, 0.0245715, 0.01632058, 0.04212672, 0.09718182, 
    0.05855738, 0.08339261, 0.02944488, 0.01762441, 0.003954871,
  5.787273e-05, 7.446693e-07, -3.418591e-05, 0.08965292, 0.0001019368, 
    0.005156929, 0.007131041, 0.002674033, 0.00411462, 0.01434087, 
    0.06302311, 0.04737596, 0.05825197, 0.06383704, 0.01885928, 0.01004854, 
    0.03052338, 0.06484335, 0.05025218, 0.0484628, 0.02617637, 0.01739201, 
    0.05310662, 0.01978402, 0.01971364, 0.001075871, 5.006309e-07, 
    1.311343e-06, 0.001139511,
  1.322134e-06, 3.80578e-08, 4.058782e-08, 0.0003025693, 5.073199e-06, 
    -1.946469e-07, -6.776903e-08, 0.003387, 0.0161988, 0.005350428, 
    0.007670143, 0.02893753, 0.04546897, 0.01793245, 0.02117731, 0.02657634, 
    0.02618875, 0.006808421, 0.0008380314, 4.663209e-06, 3.184929e-05, 
    0.1049664, 0.02107381, 0.01466891, 0.02862941, 0.04069925, 0.01439931, 
    -2.453696e-05, 1.60065e-06,
  0.005032373, 0.00742646, 0.05224999, 0.01376877, 0.009373353, 0.0004490181, 
    -0.0009691889, 0.1030956, 0.1306532, 0.1904726, 0.1344757, 0.1214385, 
    0.1336478, 0.06469354, 0.1388822, 0.0965113, 0.09002958, 0.1084428, 
    0.05946964, 0.01527538, 0.04587751, 0.09107751, 0.0873571, 0.1139936, 
    0.05470084, 0.07307244, 0.0506313, 0.001714135, 0.0002096733,
  0.0142174, 0.03184373, 0.08171575, 0.1945094, 0.03850635, 0.001935151, 
    0.1655577, 0.001158674, 0.01715641, 0.0670554, 0.127422, 0.1398864, 
    0.1920403, 0.2299858, 0.2185184, 0.2262021, 0.2140401, 0.2551362, 
    0.1283776, 0.1522264, 0.1936856, 0.1508168, 0.1738144, 0.1014947, 
    0.2724162, 0.2116934, 0.09579427, 0.05275552, 0.02676869,
  0.1348207, 0.1516409, 0.169021, 0.2033894, 0.1543311, 0.1752036, 0.1694458, 
    0.1915993, 0.1493898, 0.1407898, 0.1102061, 0.1434624, 0.09866159, 
    0.4217322, 0.2980899, 0.2076879, 0.222149, 0.2480601, 0.2069534, 
    0.1823147, 0.1165138, 0.1535666, 0.1890855, 0.1885513, 0.1961345, 
    0.2995324, 0.3436841, 0.1766962, 0.1548792,
  0.2589211, 0.1499417, 0.1732318, 0.2919756, 0.3541381, 0.3066221, 
    0.2721959, 0.2623614, 0.1974275, 0.2094197, 0.1582127, 0.07330973, 
    0.3206444, 0.3377334, 0.3874345, 0.1733357, 0.1721178, 0.2878276, 
    0.2458565, 0.256245, 0.08452473, 0.2213256, 0.2039132, 0.2160383, 
    0.2929299, 0.3398378, 0.3053645, 0.2894183, 0.3135619,
  0.3217429, 0.3124852, 0.3600325, 0.3208663, 0.3268186, 0.2963299, 
    0.2720721, 0.3843796, 0.4172061, 0.3935734, 0.242017, 0.2027384, 
    0.2473319, 0.1911677, 0.1265625, 0.1731026, 0.1304384, 0.1097647, 
    0.09941532, 0.2115481, 0.2962557, 0.1501631, 0.1812064, 0.08557444, 
    0.1526769, 0.3390111, 0.2025331, 0.1505112, 0.2224133,
  0.2347441, 0.144768, 0.1924341, 0.1691294, 0.1953243, 0.1372266, 0.1792354, 
    0.23287, 0.2696805, 0.2568818, 0.2664266, 0.2363464, 0.2029718, 
    0.2274922, 0.1742719, 0.2073952, 0.2179412, 0.1856894, 0.2081942, 
    0.2263742, 0.1972955, 0.2032892, 0.1507606, 0.02114762, 0.0517397, 
    0.1279442, 0.1548746, 0.2248984, 0.2905323,
  0.1606044, 0.1686554, 0.1767063, 0.1847573, 0.1928082, 0.2008592, 
    0.2089102, 0.2257226, 0.2397977, 0.2538728, 0.2679479, 0.282023, 
    0.2960981, 0.3101732, 0.3299114, 0.3197563, 0.3096013, 0.2994463, 
    0.2892913, 0.2791362, 0.2689812, 0.209187, 0.197216, 0.1852449, 
    0.1732739, 0.1613028, 0.1493318, 0.1373608, 0.1541636,
  0.1164846, 0.1950328, 0.1315019, 0.1404974, 0.1848352, 0.174541, 
    0.08834389, 0.09490263, 0.1971764, 0.2494487, 0.3363, 0.2945904, 
    0.3216528, 0.1391199, 0.1976646, 0.2118287, 0.2478868, 0.2873744, 
    0.2138632, 0.3197641, 0.4655925, 0.3805585, 0.2445265, 0.1750982, 
    0.1149449, 0.08129126, 0.1319165, 0.2220497, 0.1597033,
  0.392369, 0.3856653, 0.3207203, 0.4876859, 0.4457282, 0.2269801, 0.1861273, 
    0.3260602, 0.2511992, 0.1908019, 0.2618321, 0.1837765, 0.2421937, 
    0.3801359, 0.3501402, 0.3739987, 0.3221889, 0.3445085, 0.4834165, 
    0.3312178, 0.3358358, 0.2409243, 0.2727738, 0.3580142, 0.3770325, 
    0.2979874, 0.24576, 0.2059918, 0.3861422,
  0.3586434, 0.3449761, 0.3167211, 0.3532323, 0.2959185, 0.3228227, 
    0.3899482, 0.467968, 0.4535907, 0.3511876, 0.3196467, 0.3058305, 
    0.3448281, 0.3463242, 0.3528005, 0.3565872, 0.352914, 0.3305879, 
    0.3952961, 0.3842406, 0.3411135, 0.3384435, 0.2865765, 0.3326321, 
    0.3279869, 0.2486449, 0.2838152, 0.2809659, 0.3382294,
  0.2847348, 0.2803648, 0.2099134, 0.247393, 0.2262967, 0.1829445, 0.1741362, 
    0.2585715, 0.2526022, 0.271517, 0.3529885, 0.30824, 0.2330286, 0.1844534, 
    0.1164403, 0.2376879, 0.2834105, 0.240309, 0.241374, 0.2197791, 
    0.1907342, 0.2311573, 0.2670375, 0.1561525, 0.07350901, 0.1190343, 
    0.2023229, 0.2220392, 0.209526,
  0.1279751, 0.1180528, 0.1475034, 0.1263662, 0.1264367, 0.1058573, 
    0.06382774, 0.1048241, 0.1348782, 0.1455968, 0.1566698, 0.08775061, 
    0.05305865, 0.1167361, 0.1246702, 0.1113192, 0.1720516, 0.2357601, 
    0.129181, 0.1039798, 0.1530464, 0.176823, 0.09707531, 0.02735233, 
    0.0344489, 0.1156705, 0.139153, 0.0877462, 0.09002222,
  0.04783136, 0.01322926, 0.08041774, 0.04877834, 0.06278109, 0.09792279, 
    0.1060878, 0.07358167, 0.0275758, 0.004246266, 0.006622516, 0.0003739517, 
    0.0497571, 0.09550683, 0.09211965, 0.1168592, 0.1229648, 0.07550897, 
    0.0715881, 0.08070558, 0.05901752, 0.07393387, 0.008530464, 1.242908e-05, 
    0.06337096, 0.05944101, 0.08500995, 0.045077, 0.08807994,
  0.01553993, 0.001755423, 0.1401023, 0.03407188, 0.08546131, 0.0290918, 
    0.06737515, 0.05405191, 0.004520874, 0.010775, 0.005030506, 0.05270684, 
    0.09235115, 0.03531668, 0.08144017, 0.04178563, 0.0686805, 0.02523408, 
    0.02653194, 0.03085675, 0.06980587, 0.1365274, 0.00511987, 8.502469e-05, 
    0.08392444, 0.1878446, 0.02877959, 0.04735902, 0.07431055,
  0.00115378, 0.004459219, 0.1220269, 0.02708851, 0.01462192, 0.01918073, 
    0.02782608, 0.05701414, 0.02080422, 0.0756641, 0.06429492, 0.04989964, 
    0.08192691, 0.02586657, 0.03519642, 0.02608071, 0.02051378, 0.02902537, 
    0.02927388, 0.01888615, 0.03054749, 0.01553397, 0.02518644, 0.07358548, 
    0.1215835, 0.1185187, 0.05569917, 0.02357936, 0.01471112,
  0.002633233, 0.02042262, 0.04057498, 0.02377882, 0.03358329, 0.04034395, 
    0.03151941, 0.02189725, 0.0938601, 0.2693592, 0.0631581, 0.01155941, 
    0.03255604, 0.02021222, 0.02671421, 0.02708726, 0.01309483, 0.01296229, 
    0.02421595, 0.02471899, 0.02023, 0.02135726, 0.03664041, 0.08375881, 
    0.06702849, 0.07096528, 0.0259833, 0.01731866, 0.005584579,
  1.437385e-05, 2.164905e-07, -1.232073e-05, 0.03710862, 0.0008530646, 
    0.005391751, 0.006812296, 0.003421458, 0.00698405, 0.02214267, 
    0.05875913, 0.03730669, 0.0448203, 0.05623687, 0.02016498, 0.0166232, 
    0.03620774, 0.06868761, 0.08133501, 0.04862862, 0.02332327, 0.01560319, 
    0.05502351, 0.01685483, 0.02429552, 0.004031612, 1.225162e-05, 
    1.970625e-07, 0.0004493383,
  6.350776e-07, 2.46014e-08, 1.651833e-08, 0.006229963, 1.39461e-06, 
    -4.388232e-06, -2.640035e-07, 0.001903107, 0.01706735, 0.02143551, 
    0.02444683, 0.03850112, 0.04961853, 0.02437888, 0.04397887, 0.05529968, 
    0.04073738, 0.03930528, 0.006841015, 1.066025e-05, 1.485669e-05, 
    0.1304009, 0.02492238, 0.01508145, 0.02488908, 0.03972718, 0.01435507, 
    -1.500362e-05, 1.432403e-06,
  0.00024707, 0.006658404, 0.03318982, 0.009133453, 0.008190013, 
    -0.0001424399, -0.00335206, 0.07987759, 0.1245924, 0.1623799, 0.1686157, 
    0.1328633, 0.1440147, 0.09442938, 0.1803115, 0.1531172, 0.1205349, 
    0.1036626, 0.08796043, 0.04439444, 0.04598921, 0.1208476, 0.09657065, 
    0.1014326, 0.07727587, 0.1021396, 0.06189394, 0.06424711, -9.457999e-05,
  0.005290123, 0.02947004, 0.06324016, 0.192957, 0.03943197, 0.005408139, 
    0.155543, 2.144638e-05, 0.01810732, 0.07543465, 0.1288517, 0.1930561, 
    0.2553108, 0.2743939, 0.2297756, 0.253038, 0.2494828, 0.2662976, 
    0.1695886, 0.1461635, 0.1641964, 0.1501616, 0.1434654, 0.1010646, 
    0.3691319, 0.2218181, 0.1011275, 0.08491122, 0.03804182,
  0.1187573, 0.1899664, 0.1979207, 0.2239258, 0.1646573, 0.1667162, 
    0.1614697, 0.199809, 0.143123, 0.1401837, 0.06181818, 0.1381379, 
    0.1444103, 0.4506409, 0.3138047, 0.2324701, 0.2666923, 0.2953012, 
    0.2098124, 0.1726266, 0.1102199, 0.1540845, 0.1843589, 0.1967653, 
    0.2423308, 0.3613174, 0.3697383, 0.1966651, 0.1924254,
  0.2948481, 0.1373443, 0.1878251, 0.3319326, 0.3923331, 0.3083954, 
    0.2180494, 0.2801813, 0.1768427, 0.1833718, 0.1682503, 0.06969725, 
    0.3303427, 0.3423117, 0.4429936, 0.1951186, 0.1654339, 0.2956887, 
    0.2700173, 0.2373836, 0.09418435, 0.2013475, 0.2348264, 0.2065796, 
    0.3079767, 0.312301, 0.3019772, 0.2749792, 0.3511945,
  0.3654168, 0.3838397, 0.3900863, 0.3609119, 0.3780859, 0.3436826, 
    0.3235576, 0.3717975, 0.3487675, 0.3347644, 0.2551739, 0.2262504, 
    0.2595121, 0.234764, 0.1669675, 0.1749096, 0.1517533, 0.1090447, 
    0.09388019, 0.2370308, 0.3023126, 0.148591, 0.1880713, 0.09100065, 
    0.1560908, 0.3316183, 0.2306415, 0.1516076, 0.2768817,
  0.2657399, 0.1445685, 0.1998421, 0.1966606, 0.2084828, 0.2579475, 
    0.2300537, 0.3325832, 0.3160512, 0.3138666, 0.2703764, 0.2483673, 
    0.2229986, 0.2317314, 0.1727986, 0.2126223, 0.2151843, 0.1681651, 
    0.2007168, 0.2468196, 0.2112998, 0.1992494, 0.1573083, 0.02364715, 
    0.05602525, 0.09930205, 0.1578809, 0.213241, 0.3446299,
  0.1634839, 0.1715128, 0.1795418, 0.1875707, 0.1955996, 0.2036285, 
    0.2116574, 0.2176277, 0.2301683, 0.242709, 0.2552497, 0.2677903, 
    0.280331, 0.2928717, 0.3143338, 0.3043292, 0.2943246, 0.28432, 0.2743154, 
    0.2643108, 0.2543062, 0.2038807, 0.1933157, 0.1827507, 0.1721857, 
    0.1616207, 0.1510558, 0.1404908, 0.1570608,
  0.1344189, 0.2055568, 0.2028284, 0.1556105, 0.2030965, 0.1878994, 
    0.1157287, 0.1192944, 0.2469695, 0.2509892, 0.345935, 0.3153513, 
    0.3495013, 0.1172395, 0.1398268, 0.190025, 0.2647454, 0.2734956, 
    0.2013435, 0.2911037, 0.457324, 0.3905912, 0.2369363, 0.1689979, 
    0.1126256, 0.095552, 0.2230642, 0.2247522, 0.1645953,
  0.4051106, 0.3632733, 0.3850558, 0.452179, 0.4316011, 0.2223532, 0.197503, 
    0.3541442, 0.2443027, 0.2156146, 0.2273149, 0.1823751, 0.2283856, 
    0.3628745, 0.5563048, 0.4343022, 0.4197389, 0.4666467, 0.4898018, 
    0.3918302, 0.3657109, 0.2771758, 0.3139578, 0.3341352, 0.3855922, 
    0.3928164, 0.3156137, 0.3855434, 0.4713327,
  0.4237568, 0.3532238, 0.3549979, 0.3166423, 0.3439282, 0.3431811, 
    0.4270696, 0.5116969, 0.5408486, 0.3648965, 0.346123, 0.3168354, 
    0.3839624, 0.3615456, 0.3580157, 0.4047519, 0.4317817, 0.4522702, 
    0.4780665, 0.3930452, 0.3309336, 0.3530957, 0.3212394, 0.3394954, 
    0.3864888, 0.3188787, 0.3636259, 0.3553035, 0.3528588,
  0.3499296, 0.2938083, 0.2584552, 0.3049549, 0.253747, 0.2102069, 0.1780488, 
    0.3256249, 0.3038466, 0.3054236, 0.3893397, 0.3239893, 0.3213134, 
    0.2245017, 0.1550377, 0.2813757, 0.3288992, 0.2793998, 0.2625074, 
    0.2598645, 0.2626227, 0.2404243, 0.2914478, 0.1683564, 0.07173791, 
    0.1560405, 0.236487, 0.2580356, 0.2628645,
  0.1965326, 0.1719232, 0.2314287, 0.1629617, 0.1873686, 0.1574485, 
    0.08104057, 0.1873257, 0.1982076, 0.2006834, 0.2333606, 0.06976448, 
    0.04705875, 0.1385673, 0.1459853, 0.1649678, 0.2443102, 0.3185001, 
    0.1886566, 0.1702497, 0.1815264, 0.2188898, 0.1763732, 0.03178778, 
    0.03226979, 0.1584668, 0.1550486, 0.1210447, 0.1151624,
  0.1130922, 0.02868686, 0.07805405, 0.06868065, 0.06620792, 0.08735577, 
    0.1033035, 0.1029335, 0.08926562, 0.02327533, 0.005780669, 0.001096904, 
    0.03128659, 0.09254006, 0.09945437, 0.1500273, 0.1402559, 0.08818794, 
    0.08850106, 0.08428957, 0.09380552, 0.1013552, 0.05352122, 4.713077e-05, 
    0.06259733, 0.06811763, 0.0758169, 0.04435163, 0.1056461,
  0.08737265, -0.0004338528, 0.140011, 0.03646066, 0.07635847, 0.0296712, 
    0.06482068, 0.05843495, 0.02595913, 0.008633792, 0.003642052, 0.04682139, 
    0.09187985, 0.03141444, 0.06628572, 0.04421864, 0.07977103, 0.02524764, 
    0.03380425, 0.03003383, 0.0528915, 0.1603296, 0.05875122, 0.0003369885, 
    0.1206168, 0.1964832, 0.03299694, 0.03996206, 0.1036323,
  0.02106661, 0.0155065, 0.1093735, 0.03241603, 0.01845394, 0.02112405, 
    0.03074462, 0.05288426, 0.0231208, 0.06371088, 0.05635725, 0.0434945, 
    0.06176765, 0.02299026, 0.02775586, 0.02506012, 0.01936003, 0.02800333, 
    0.03062275, 0.02201533, 0.02253137, 0.02886877, 0.04531489, 0.06502663, 
    0.1229513, 0.1117045, 0.06010256, 0.0340619, 0.05828531,
  0.005132275, 0.02316123, 0.03829138, 0.01284513, 0.03736436, 0.04090727, 
    0.02848288, 0.02559691, 0.1135023, 0.2547647, 0.05171085, 0.01608098, 
    0.02977111, 0.02315902, 0.02479992, 0.02894769, 0.01571072, 0.01585522, 
    0.02679937, 0.02127603, 0.01543427, 0.0240185, 0.03470071, 0.06744158, 
    0.07766, 0.05979436, 0.02409187, 0.01983867, 0.01788997,
  2.532602e-06, 7.096943e-08, -3.861664e-06, 0.01617974, 0.01451758, 
    0.0144327, 0.007442664, 0.005008997, 0.007145683, 0.02693785, 0.05901669, 
    0.03515959, 0.03880702, 0.05019362, 0.03291419, 0.03670711, 0.04052434, 
    0.07725739, 0.1111944, 0.04799245, 0.02308011, 0.01745958, 0.05374007, 
    0.0140329, 0.04095063, 0.02130497, 0.001155293, 1.864343e-07, 0.0002011693,
  2.323134e-07, 1.85083e-08, 8.636537e-09, 0.0008791076, 1.175424e-07, 
    0.0003749601, -1.290141e-05, 0.002016786, 0.0199, 0.03299299, 0.08266465, 
    0.06686247, 0.0555044, 0.03197917, 0.09445822, 0.1146714, 0.0742005, 
    0.06076484, 0.04118489, 0.00162936, 5.145476e-06, 0.1741813, 0.02479823, 
    0.01996921, 0.0495901, 0.05308257, 0.06857202, 1.133471e-05, 9.346963e-07,
  1.114845e-05, 0.0102652, 0.01249988, 0.008162889, 0.003391078, 
    -7.980874e-05, -0.00398644, 0.05765679, 0.1132921, 0.1455666, 0.185006, 
    0.173832, 0.2268338, 0.1530305, 0.2872842, 0.2240498, 0.171088, 
    0.1817586, 0.1740729, 0.04244751, 0.05666053, 0.1466542, 0.140376, 
    0.1382058, 0.1866033, 0.1345889, 0.06717906, 0.1485866, -0.0002649888,
  0.001219643, 0.01632064, 0.04603986, 0.1788689, 0.04257359, 0.001546784, 
    0.1526628, -7.139458e-05, 0.01562126, 0.05946205, 0.1299925, 0.185002, 
    0.3185129, 0.2723022, 0.2259129, 0.3094499, 0.3475829, 0.2898705, 
    0.2326518, 0.1516434, 0.1445134, 0.1481793, 0.1473739, 0.1175597, 
    0.4494943, 0.2551537, 0.1400844, 0.1091175, 0.04974532,
  0.1566696, 0.2266911, 0.2085388, 0.192904, 0.1024598, 0.1749967, 0.1706159, 
    0.2233658, 0.1457853, 0.1401037, 0.0571643, 0.1259753, 0.2505706, 
    0.427634, 0.4359882, 0.241767, 0.3737986, 0.3551782, 0.3095863, 
    0.1625963, 0.09437809, 0.1161667, 0.181896, 0.1888462, 0.3033406, 
    0.4357795, 0.3439571, 0.2437259, 0.1769707,
  0.3049844, 0.1395618, 0.2322743, 0.4158429, 0.4699092, 0.2714827, 0.247104, 
    0.3027097, 0.1941737, 0.1699927, 0.2075723, 0.07176478, 0.3372056, 
    0.3185601, 0.4898654, 0.2264877, 0.1775954, 0.3098891, 0.2778276, 
    0.2047882, 0.1330184, 0.2149183, 0.2582351, 0.1981874, 0.3973938, 
    0.2704624, 0.2425987, 0.2255077, 0.3246405,
  0.4043868, 0.3607283, 0.3934066, 0.4756958, 0.3410744, 0.3424156, 
    0.3776082, 0.2942043, 0.3058534, 0.2700018, 0.2902387, 0.2707633, 
    0.2425463, 0.22836, 0.1923837, 0.1481389, 0.1595772, 0.1058224, 
    0.08708754, 0.269272, 0.3120727, 0.1623371, 0.2124125, 0.09207258, 
    0.1440722, 0.3335482, 0.2423894, 0.1371187, 0.397114,
  0.2827143, 0.1441021, 0.2102337, 0.1866145, 0.1925017, 0.2315702, 
    0.2376661, 0.3209552, 0.2948909, 0.3033462, 0.3205489, 0.3031729, 
    0.2439272, 0.232381, 0.1960078, 0.195271, 0.202463, 0.1678239, 0.2392953, 
    0.304781, 0.2359958, 0.2092473, 0.1626733, 0.02963037, 0.0633835, 
    0.08342434, 0.1560425, 0.205612, 0.3346841,
  0.1690997, 0.1775773, 0.1860548, 0.1945324, 0.2030099, 0.2114875, 
    0.2199651, 0.2138364, 0.2247443, 0.2356522, 0.2465602, 0.2574681, 
    0.2683761, 0.279284, 0.301517, 0.2917796, 0.2820422, 0.2723049, 
    0.2625675, 0.2528302, 0.2430928, 0.1935263, 0.1838782, 0.17423, 
    0.1645819, 0.1549337, 0.1452856, 0.1356374, 0.1623176,
  0.1294883, 0.2164367, 0.2615474, 0.1897082, 0.2297818, 0.2199363, 
    0.1181614, 0.1384058, 0.2496293, 0.25747, 0.3590625, 0.3259205, 
    0.3866586, 0.1063634, 0.1203149, 0.2038346, 0.2447649, 0.2662207, 
    0.190596, 0.2534352, 0.4745774, 0.4367371, 0.2388977, 0.1417361, 
    0.1143342, 0.138539, 0.2544613, 0.1779713, 0.1835758,
  0.384138, 0.3474442, 0.3997301, 0.4271476, 0.4106201, 0.2324136, 0.15728, 
    0.3610205, 0.22705, 0.2366991, 0.2288913, 0.1961744, 0.2168902, 
    0.3505454, 0.412224, 0.4569111, 0.5117498, 0.5400615, 0.3849154, 
    0.4028856, 0.3864711, 0.3179419, 0.3660705, 0.3576306, 0.3882575, 
    0.4376881, 0.4450487, 0.4340586, 0.4177157,
  0.4498649, 0.4001218, 0.3464913, 0.3475256, 0.3457317, 0.4352384, 
    0.4825838, 0.4992547, 0.5248508, 0.3816946, 0.3519132, 0.3365341, 
    0.4178867, 0.3915679, 0.3595572, 0.4120318, 0.4907748, 0.502996, 
    0.502627, 0.3995007, 0.3588665, 0.4091621, 0.3561817, 0.368325, 0.48005, 
    0.4686807, 0.4151025, 0.4131739, 0.3630319,
  0.3814555, 0.3259396, 0.3018637, 0.2917495, 0.2784753, 0.2517479, 
    0.2199357, 0.3874192, 0.3531836, 0.325812, 0.3579717, 0.2940015, 
    0.3862786, 0.3172521, 0.2245828, 0.2700757, 0.3222519, 0.2729434, 
    0.2571737, 0.2547335, 0.2779207, 0.2434722, 0.3054092, 0.1697328, 
    0.08902704, 0.2261107, 0.3079215, 0.3582115, 0.3352466,
  0.2374275, 0.3271341, 0.2505994, 0.2314615, 0.2655923, 0.2496134, 0.152994, 
    0.2957147, 0.3375356, 0.2856922, 0.2079546, 0.1108558, 0.07089121, 
    0.2436687, 0.2024236, 0.2126253, 0.2644374, 0.3128859, 0.222252, 
    0.2273997, 0.2051881, 0.3315268, 0.2328825, 0.04369061, 0.01305352, 
    0.1775549, 0.2545204, 0.1653034, 0.173455,
  0.1997026, 0.0535408, 0.08121072, 0.1302617, 0.1106086, 0.09465314, 
    0.1081397, 0.119494, 0.1917007, 0.02070049, 0.004551751, 0.0002950274, 
    0.01331927, 0.09010557, 0.09772935, 0.1943897, 0.1541052, 0.1033492, 
    0.1081586, 0.08804404, 0.07472994, 0.1092723, 0.1977532, 7.769056e-05, 
    0.05978031, 0.1047488, 0.0736185, 0.05896837, 0.1046269,
  0.223033, -0.0006626485, 0.1327587, 0.05232971, 0.08336635, 0.04005121, 
    0.07123805, 0.0785462, 0.09213983, 0.007798005, 0.001326634, 0.03674458, 
    0.09132184, 0.06429528, 0.06705422, 0.05713064, 0.06965446, 0.03114561, 
    0.0403611, 0.03843687, 0.06165586, 0.1377599, 0.1953847, -6.2126e-05, 
    0.09379773, 0.1912214, 0.04713854, 0.04887711, 0.119695,
  0.0824477, 0.03483663, 0.0847699, 0.03311756, 0.0278421, 0.0291733, 
    0.03848355, 0.05613883, 0.03257447, 0.05365494, 0.06638006, 0.04788635, 
    0.06205138, 0.02413147, 0.03254907, 0.03211123, 0.02187696, 0.03184391, 
    0.06402984, 0.04586346, 0.04804403, 0.0545021, 0.06863507, 0.0411939, 
    0.09658538, 0.09325655, 0.07667415, 0.05161769, 0.07915346,
  0.01078468, 0.02203349, 0.03362737, 0.008435396, 0.05487045, 0.08916103, 
    0.0342875, 0.0325847, 0.1235119, 0.205509, 0.04653495, 0.02360341, 
    0.0332664, 0.03778937, 0.02646057, 0.03994881, 0.02133892, 0.01614852, 
    0.03296992, 0.02349971, 0.01580539, 0.02544562, 0.01790193, 0.05080143, 
    0.07133907, 0.05575404, 0.02836495, 0.02677108, 0.02109765,
  -9.489667e-07, 4.013606e-08, -2.557095e-06, 0.00621386, 0.0186961, 
    0.1091065, 0.006949069, 0.01156635, 0.009211786, 0.03593056, 0.07393871, 
    0.04926581, 0.04943132, 0.05029267, 0.08072881, 0.05219665, 0.04480651, 
    0.08666693, 0.1250508, 0.05063074, 0.02798636, 0.02595862, 0.07044009, 
    0.01934167, 0.05865302, 0.1243655, 0.02319673, 2.03304e-07, 0.0001522648,
  5.190284e-08, 1.381023e-08, 4.471816e-09, 0.0001745699, 1.423104e-08, 
    0.002319277, -1.160514e-05, 0.006730969, 0.02510657, 0.07280663, 
    0.122355, 0.08513165, 0.06702304, 0.06680876, 0.1013973, 0.1640782, 
    0.1741363, 0.06359155, 0.223277, 0.05475721, -1.824231e-05, 0.201249, 
    0.05326031, 0.03588085, 0.09921247, 0.0774519, 0.1556081, 0.003349872, 
    3.970294e-07,
  -1.72053e-05, 0.0130123, 0.008161074, 0.009151332, 0.003366058, 
    -2.749284e-05, -0.004058535, 0.03999698, 0.1097917, 0.1553295, 0.2097598, 
    0.2027973, 0.2512158, 0.2341935, 0.3520924, 0.2763626, 0.2432251, 
    0.2705991, 0.3032881, 0.05867963, 0.04922397, 0.176573, 0.1497049, 
    0.254689, 0.1979243, 0.1583066, 0.116502, 0.07503755, -0.0006652791,
  -7.429475e-05, 0.02306757, 0.03535669, 0.1649918, 0.04543563, 0.001062114, 
    0.1463853, -3.23515e-06, 0.01229885, 0.05325231, 0.1352994, 0.1972302, 
    0.2388138, 0.1897089, 0.1678234, 0.3042822, 0.3769899, 0.3322538, 
    0.3017007, 0.1350875, 0.1284023, 0.1731127, 0.162922, 0.1391967, 
    0.3548412, 0.254056, 0.1089922, 0.202846, 0.0739955,
  0.1470517, 0.2784775, 0.2103859, 0.1696623, 0.1382372, 0.1599965, 
    0.1854424, 0.2154402, 0.1346711, 0.1198672, 0.03167075, 0.1236221, 
    0.4009611, 0.3931733, 0.3547609, 0.3085665, 0.3999507, 0.4076862, 
    0.4305514, 0.1513398, 0.09424297, 0.09985997, 0.1794692, 0.1719668, 
    0.311334, 0.3769387, 0.3101803, 0.2860795, 0.1698511,
  0.2657248, 0.1351656, 0.2917954, 0.4940894, 0.489865, 0.2732576, 0.2599481, 
    0.2838245, 0.1750019, 0.1686889, 0.1936089, 0.07192723, 0.3125134, 
    0.2969797, 0.4830689, 0.2736136, 0.2494428, 0.3072608, 0.276425, 
    0.1761292, 0.139077, 0.2382766, 0.2729613, 0.1946993, 0.5518513, 0.21932, 
    0.1506462, 0.1806626, 0.2746725,
  0.3334621, 0.294784, 0.4180678, 0.4518265, 0.3249259, 0.277117, 0.3452467, 
    0.3118186, 0.3126196, 0.2733789, 0.3306323, 0.3180539, 0.252001, 
    0.2069586, 0.239771, 0.216478, 0.1329882, 0.1006127, 0.09775432, 
    0.3041869, 0.3153512, 0.1703805, 0.2282671, 0.09784134, 0.1324325, 
    0.3385874, 0.2442814, 0.1304041, 0.4599069,
  0.2865714, 0.1419283, 0.2344638, 0.207999, 0.2503022, 0.2388174, 0.3011032, 
    0.3442022, 0.3161708, 0.2978217, 0.3525273, 0.3315454, 0.3014703, 
    0.2940793, 0.2452738, 0.2136668, 0.2229361, 0.2029858, 0.27759, 
    0.3754787, 0.2653022, 0.2260258, 0.1695764, 0.04175144, 0.08077934, 
    0.08914452, 0.1465879, 0.2056229, 0.3043352,
  0.1861326, 0.1933555, 0.2005784, 0.2078013, 0.2150241, 0.222247, 0.2294699, 
    0.2124569, 0.2218668, 0.2312768, 0.2406868, 0.2500969, 0.2595069, 
    0.2689168, 0.2952984, 0.2846831, 0.2740678, 0.2634525, 0.2528372, 
    0.2422218, 0.2316065, 0.1946883, 0.1886708, 0.1826532, 0.1766357, 
    0.1706181, 0.1646006, 0.158583, 0.1803543,
  0.1323456, 0.2038834, 0.2980749, 0.229886, 0.2642602, 0.2126348, 0.1235807, 
    0.1729297, 0.2536393, 0.2506295, 0.3679906, 0.3342183, 0.4033398, 
    0.07450639, 0.1116787, 0.204302, 0.2207816, 0.2557714, 0.1700819, 
    0.2650611, 0.4698378, 0.4676238, 0.2423662, 0.09480856, 0.1143736, 
    0.1482617, 0.2355065, 0.1247813, 0.1932695,
  0.3575963, 0.2949791, 0.3456054, 0.3630293, 0.3948502, 0.234131, 0.1202562, 
    0.3754677, 0.2258673, 0.2497613, 0.2220631, 0.2178615, 0.2184887, 
    0.290567, 0.3269926, 0.4719315, 0.4828663, 0.5354037, 0.3519608, 
    0.3932007, 0.4657368, 0.3707288, 0.3977841, 0.3747248, 0.3698896, 
    0.5475363, 0.5316264, 0.3285716, 0.3238468,
  0.3611057, 0.3736447, 0.3079026, 0.3604771, 0.3445367, 0.453495, 0.5318509, 
    0.4863081, 0.468771, 0.3048762, 0.2981465, 0.3674217, 0.5246449, 
    0.4293466, 0.3362955, 0.3751892, 0.5065985, 0.5124959, 0.4735612, 
    0.3709126, 0.370772, 0.4377274, 0.4576004, 0.4251869, 0.5428788, 
    0.4779394, 0.4219189, 0.4178239, 0.3773264,
  0.3935591, 0.3651948, 0.2945486, 0.3059764, 0.277057, 0.3070314, 0.3002824, 
    0.4215327, 0.3670194, 0.3206956, 0.3381028, 0.3159349, 0.3408373, 
    0.3177566, 0.2552717, 0.2815001, 0.2969805, 0.2514492, 0.2371684, 
    0.2440549, 0.2128764, 0.2577707, 0.2928029, 0.1936824, 0.06152797, 
    0.1936415, 0.3495787, 0.4083108, 0.3447961,
  0.2558984, 0.326591, 0.1794402, 0.2443168, 0.2579152, 0.2880018, 0.252442, 
    0.2647463, 0.3753929, 0.2329984, 0.2134043, 0.1604694, 0.1402434, 
    0.2384878, 0.2456828, 0.2426276, 0.2329329, 0.2647053, 0.2074049, 
    0.1883139, 0.2329091, 0.3923908, 0.267074, 0.06130573, 0.006728269, 
    0.2053764, 0.2318502, 0.2099788, 0.2367202,
  0.2078296, 0.1581122, 0.08979392, 0.2310721, 0.1128055, 0.07551992, 
    0.1288981, 0.1138504, 0.2653316, 0.0667159, 0.006416691, -1.967803e-06, 
    0.01127139, 0.08260068, 0.09845804, 0.1601005, 0.1688838, 0.1103916, 
    0.07475214, 0.07685765, 0.06682267, 0.09850992, 0.3614444, 0.0003198934, 
    0.05523317, 0.09333563, 0.0994491, 0.08423429, 0.108872,
  0.2971945, 0.002469068, 0.1096653, 0.08782449, 0.1007031, 0.08634143, 
    0.08922029, 0.04851971, 0.1340184, 0.02513924, 0.0003776062, 0.0243214, 
    0.08002479, 0.05635365, 0.07215317, 0.1068279, 0.06338754, 0.04828417, 
    0.04692107, 0.04115778, 0.08749304, 0.06412153, 0.4909337, -0.002159636, 
    0.07256597, 0.1894329, 0.04634367, 0.03508615, 0.08762553,
  0.2561896, 0.06215145, 0.05456462, 0.02305519, 0.1158177, 0.05859479, 
    0.04467421, 0.1069865, 0.06504345, 0.1136687, 0.05555628, 0.1542097, 
    0.06320192, 0.0317648, 0.04273171, 0.09266641, 0.0261583, 0.07705722, 
    0.07856962, 0.07953058, 0.1611817, 0.1357241, 0.1492203, 0.02507455, 
    0.0620736, 0.06747966, 0.09252268, 0.07889283, 0.1378395,
  0.06098807, 0.01501323, 0.02817191, 0.006773489, 0.0620483, 0.1013043, 
    0.1214427, 0.1063408, 0.07570666, 0.1669354, 0.07626956, 0.08330554, 
    0.1274643, 0.04654235, 0.03268699, 0.05164037, 0.03441202, 0.01589377, 
    0.06719527, 0.03277533, 0.02909927, 0.03327191, 0.01409511, 0.03671344, 
    0.04038224, 0.06387664, 0.03740687, 0.05105978, 0.0432157,
  -1.096085e-06, 3.069224e-08, -5.796049e-07, 0.003130369, 0.01975828, 
    0.2573545, 0.04083619, 0.08666517, 0.02902201, 0.09610552, 0.07691341, 
    0.06943358, 0.04937791, 0.04537375, 0.04447614, 0.05536205, 0.05178932, 
    0.1000771, 0.1344637, 0.07603538, 0.05648312, 0.03502681, 0.1359107, 
    0.03041616, 0.0504698, 0.1081367, 0.132922, -6.594781e-07, 0.0001679175,
  2.61192e-08, 1.18446e-08, 2.564604e-09, 4.304987e-05, 4.514594e-09, 
    0.02857705, -1.784287e-05, 0.01345727, 0.02491446, 0.1154865, 0.1122535, 
    0.1140284, 0.1187129, 0.09657723, 0.06061624, 0.106487, 0.09336171, 
    0.07433965, 0.2204038, 0.1496959, -0.0004761143, 0.246634, 0.05815705, 
    0.02329048, 0.03775863, 0.0376051, 0.07984374, 0.04312219, 1.191639e-07,
  1.717134e-06, 0.02061816, 0.005896231, 0.012158, 0.0006414109, 
    -7.594643e-06, -0.003735452, 0.02856913, 0.1025553, 0.181145, 0.1959798, 
    0.1507441, 0.2189875, 0.2009008, 0.253647, 0.2523388, 0.1680204, 
    0.1973819, 0.2806191, 0.07086766, 0.04331671, 0.2108036, 0.1288244, 
    0.200485, 0.1843996, 0.1780563, 0.1295409, 0.1302122, 0.0008578894,
  -0.0009426957, 0.019734, 0.02804379, 0.1794391, 0.03933786, -6.169004e-06, 
    0.1417172, 8.285376e-07, 0.01426894, 0.06056661, 0.135931, 0.147084, 
    0.1802511, 0.1508559, 0.1408022, 0.2457154, 0.3486469, 0.3269525, 
    0.2792746, 0.119289, 0.1210173, 0.2356997, 0.1548593, 0.1249014, 
    0.2558142, 0.2337465, 0.1273616, 0.3324995, 0.09988485,
  0.2030123, 0.2822688, 0.1966707, 0.1342205, 0.1158647, 0.187475, 0.178892, 
    0.2140386, 0.1139835, 0.110341, 0.02206209, 0.1246609, 0.4272683, 
    0.329965, 0.2916224, 0.2543492, 0.369684, 0.4628646, 0.4446837, 
    0.1639667, 0.1266789, 0.0911713, 0.161516, 0.1613795, 0.2879441, 
    0.296118, 0.3025414, 0.2304256, 0.2447024,
  0.2542431, 0.141641, 0.2818789, 0.4525289, 0.4667316, 0.2889805, 0.3253775, 
    0.2745164, 0.1631231, 0.154347, 0.2054219, 0.06335956, 0.2379376, 
    0.2787456, 0.5154179, 0.241983, 0.2882613, 0.2840849, 0.2999063, 
    0.1510369, 0.1519444, 0.2027584, 0.2742642, 0.178589, 0.5840173, 
    0.136928, 0.112902, 0.1665695, 0.2502309,
  0.2142913, 0.2164523, 0.4381155, 0.3935556, 0.3448161, 0.2786653, 
    0.3038334, 0.3307631, 0.310046, 0.3679312, 0.3638862, 0.378177, 
    0.2868026, 0.2256196, 0.2534792, 0.1814797, 0.1280834, 0.1294534, 
    0.1043444, 0.3166586, 0.3207003, 0.1871034, 0.2358617, 0.09861212, 
    0.1291871, 0.3571493, 0.2558866, 0.1207482, 0.3915621,
  0.2546635, 0.186682, 0.2542659, 0.2929873, 0.2789888, 0.3169407, 0.3228983, 
    0.3619622, 0.3957443, 0.326753, 0.4144069, 0.4092787, 0.3508429, 
    0.3429478, 0.2605981, 0.2312341, 0.2679602, 0.3011685, 0.3371041, 
    0.4010107, 0.279122, 0.2270376, 0.1664076, 0.05900431, 0.1018931, 
    0.1088913, 0.1311889, 0.2006841, 0.2779624,
  0.2259647, 0.2321153, 0.238266, 0.2444167, 0.2505673, 0.256718, 0.2628687, 
    0.2344878, 0.2421779, 0.249868, 0.2575581, 0.2652482, 0.2729383, 
    0.2806285, 0.29553, 0.2842042, 0.2728785, 0.2615528, 0.250227, 0.2389012, 
    0.2275755, 0.1927697, 0.1902547, 0.1877396, 0.1852246, 0.1827096, 
    0.1801946, 0.1776795, 0.2210442,
  0.1449854, 0.2216627, 0.301686, 0.2636899, 0.3046098, 0.2054196, 0.1427531, 
    0.1979288, 0.2769846, 0.2815218, 0.339057, 0.3735398, 0.4179584, 
    0.04308817, 0.07121713, 0.2173395, 0.2592382, 0.2440526, 0.1460946, 
    0.2808705, 0.5386129, 0.4820924, 0.251193, 0.08604547, 0.1082347, 
    0.1741807, 0.1199055, 0.0894817, 0.1849965,
  0.2819679, 0.2435909, 0.3052622, 0.2907229, 0.3600875, 0.2227383, 
    0.09622756, 0.3848754, 0.2304042, 0.2561392, 0.2048533, 0.2426376, 
    0.2164428, 0.1843724, 0.2165726, 0.3616631, 0.4598109, 0.4434027, 
    0.35901, 0.4340672, 0.5103495, 0.4424129, 0.4138015, 0.4357745, 
    0.3499183, 0.5598383, 0.3561601, 0.1983733, 0.2466662,
  0.3021663, 0.3302997, 0.2815652, 0.3364441, 0.3681956, 0.3888549, 
    0.4643595, 0.4334787, 0.4328184, 0.2491751, 0.2639886, 0.3534818, 
    0.495852, 0.4398447, 0.3198074, 0.3717224, 0.4353693, 0.4687413, 
    0.4355899, 0.3337079, 0.3344372, 0.3661383, 0.4404365, 0.4467072, 
    0.5144733, 0.4613684, 0.4452229, 0.388085, 0.3756024,
  0.3912941, 0.3534759, 0.2980404, 0.2947529, 0.274774, 0.3013213, 0.3818544, 
    0.3867227, 0.3459067, 0.3059754, 0.3125804, 0.328524, 0.3343243, 
    0.2669248, 0.2338057, 0.2953755, 0.274516, 0.2454795, 0.2013723, 
    0.2372544, 0.1776692, 0.2241623, 0.2709458, 0.1859225, 0.034791, 
    0.1777305, 0.3586741, 0.3948419, 0.3775608,
  0.2987841, 0.2494518, 0.1368317, 0.2630909, 0.3015381, 0.2709584, 
    0.3136929, 0.1829701, 0.2379359, 0.1352978, 0.1882254, 0.1246397, 
    0.07553705, 0.2965546, 0.2691114, 0.1872852, 0.1774254, 0.2208994, 
    0.1982999, 0.1952384, 0.239131, 0.3844902, 0.243925, 0.08315842, 
    0.009057501, 0.1878229, 0.1949616, 0.2278154, 0.2271842,
  0.08466557, 0.1899845, 0.07772145, 0.08412728, 0.0856458, 0.05744642, 
    0.05435742, 0.02550272, 0.1445809, 0.02032726, 0.01409932, -3.030533e-05, 
    0.00850272, 0.05703398, 0.1085915, 0.1081208, 0.1089947, 0.1259318, 
    0.09364657, 0.03596736, 0.04177717, 0.03591937, 0.1375044, 0.00395449, 
    0.05511761, 0.06988189, 0.06748391, 0.01743315, 0.04928959,
  0.09855562, 0.01021781, 0.08588671, 0.07260747, 0.08087292, 0.08742995, 
    0.06148801, 0.01468018, 0.08038566, 0.04733511, 0.0001406242, 0.01844144, 
    0.07697924, 0.02247827, 0.04595243, 0.05089892, 0.04426642, 0.04217005, 
    0.01842531, 0.01114461, 0.02313955, 0.01412182, 0.2387348, 0.1110727, 
    0.05465467, 0.1907655, 0.01101006, 0.006418016, 0.02056013,
  0.2195976, 0.1501147, 0.03412134, 0.02299388, 0.04974448, 0.0514013, 
    0.027972, 0.09267313, 0.122011, 0.04833022, 0.02285982, 0.05994412, 
    0.0303613, 0.01878032, 0.03516372, 0.02757596, 0.01749192, 0.02883739, 
    0.01810591, 0.05202443, 0.07090354, 0.1207918, 0.1748903, 0.01479649, 
    0.03763585, 0.04719432, 0.03892587, 0.01990951, 0.05649289,
  0.11932, 0.007327276, 0.01609486, 0.006204389, 0.08269184, 0.03678364, 
    0.02844978, 0.02258139, 0.04186425, 0.1454633, 0.04562773, 0.1756373, 
    0.03368428, 0.03186215, 0.02691363, 0.03793581, 0.06609118, 0.03280133, 
    0.0676467, 0.1148822, 0.1615752, 0.176041, 0.03489591, 0.02365175, 
    0.01136519, 0.04199826, 0.04577326, 0.08973008, 0.1242293,
  -4.01421e-07, 2.787783e-08, -2.628728e-07, 0.001283168, 0.01812776, 
    0.06559721, 0.009678751, 0.06329785, 0.01754088, 0.06358363, 0.05992559, 
    0.07293266, 0.01991459, 0.02269501, 0.01187249, 0.01281482, 0.03521195, 
    0.08478166, 0.0861312, 0.06177754, 0.025732, 0.02029628, 0.2647103, 
    0.08629575, 0.007399048, 0.02494253, 0.04971546, -0.0001507236, 
    7.518449e-05,
  2.050925e-08, 1.112685e-08, 1.599369e-09, 0.0002796791, 2.611203e-09, 
    0.01183118, -1.911322e-05, 0.005182201, 0.0169043, 0.1549976, 0.12144, 
    0.06501113, 0.0647992, 0.05617965, 0.01396505, 0.03958181, 0.04077708, 
    0.07515544, 0.1455362, 0.1437704, -0.0001027512, 0.2334493, 0.01256877, 
    0.002399372, 0.009414016, 0.01205617, 0.04300186, 0.01189958, 7.581735e-08,
  -6.190564e-06, 0.01261244, 0.003446979, 0.01437088, 0.0006971718, 
    -4.348195e-06, -0.003340519, 0.02340386, 0.08938165, 0.1800908, 
    0.1759262, 0.1311963, 0.1657313, 0.1338251, 0.2085318, 0.1857816, 
    0.08536914, 0.1252356, 0.232035, 0.05129123, 0.03918102, 0.2378446, 
    0.12131, 0.139194, 0.1626575, 0.1558074, 0.09697897, 0.07439958, 0.002279,
  -0.001605692, 0.009560208, 0.02343307, 0.1697755, 0.02501331, 
    -0.0002532214, 0.1294535, 7.793446e-06, 0.01410537, 0.06480695, 
    0.1309599, 0.1256903, 0.1525676, 0.1201582, 0.1184751, 0.2062902, 
    0.3050508, 0.307355, 0.2674789, 0.1105071, 0.1199619, 0.2306762, 
    0.1327813, 0.1154663, 0.2111485, 0.2348233, 0.1306146, 0.2414352, 
    0.09453537,
  0.1894291, 0.2684779, 0.1497597, 0.0952695, 0.1052851, 0.1943084, 
    0.1448916, 0.1942137, 0.09477136, 0.09140848, 0.01777092, 0.1361483, 
    0.3114456, 0.2740831, 0.2506787, 0.2093995, 0.3818418, 0.4232449, 
    0.3708267, 0.1766373, 0.1158358, 0.08318719, 0.1269787, 0.1511018, 
    0.2243087, 0.2247437, 0.2818712, 0.199518, 0.256727,
  0.2550741, 0.1791378, 0.2704859, 0.409605, 0.4832058, 0.2916881, 0.3990448, 
    0.2327824, 0.119042, 0.1168291, 0.1761356, 0.06496809, 0.2127989, 
    0.2409035, 0.5780436, 0.202089, 0.2511588, 0.2666524, 0.3324899, 
    0.1733722, 0.1201523, 0.1519484, 0.2586234, 0.1407502, 0.4824989, 
    0.09142787, 0.08676517, 0.1695029, 0.2327842,
  0.1450722, 0.1484958, 0.3657368, 0.3047646, 0.3677697, 0.318388, 0.2977796, 
    0.3427232, 0.283752, 0.3761866, 0.4529384, 0.4267704, 0.3390246, 
    0.2574649, 0.2672554, 0.1733061, 0.1729915, 0.1416348, 0.1472625, 
    0.3428762, 0.3380832, 0.2307164, 0.2587112, 0.08720266, 0.1415943, 
    0.3661848, 0.2535377, 0.09578889, 0.2611014,
  0.2022688, 0.1847987, 0.3145785, 0.3719897, 0.3524875, 0.4564292, 
    0.4303274, 0.3969753, 0.4103175, 0.3566379, 0.4270538, 0.435332, 
    0.4029618, 0.3741229, 0.2864059, 0.2914065, 0.3203711, 0.3631078, 
    0.3895719, 0.461292, 0.3157219, 0.2300728, 0.1575195, 0.06435009, 
    0.1337519, 0.1402712, 0.1235792, 0.1865099, 0.2930182,
  0.2810682, 0.2852596, 0.289451, 0.2936424, 0.2978338, 0.3020251, 0.3062165, 
    0.2465499, 0.2524093, 0.2582686, 0.264128, 0.2699873, 0.2758467, 
    0.2817061, 0.286898, 0.275481, 0.264064, 0.252647, 0.2412301, 0.2298131, 
    0.2183962, 0.2012858, 0.202652, 0.2040183, 0.2053845, 0.2067507, 
    0.2081169, 0.2094831, 0.2777151,
  0.1853099, 0.2378492, 0.3103171, 0.3051883, 0.351772, 0.193737, 0.1721935, 
    0.2276445, 0.2691123, 0.2616282, 0.3016213, 0.4177616, 0.4124625, 
    0.01940116, 0.04907485, 0.260351, 0.277759, 0.2550918, 0.124749, 
    0.2658063, 0.5542116, 0.5110623, 0.2405335, 0.08481105, 0.09441794, 
    0.2086943, 0.06723721, 0.0424853, 0.1893694,
  0.2111264, 0.183447, 0.2789675, 0.210993, 0.303524, 0.2137714, 0.07615529, 
    0.3546182, 0.232485, 0.2367696, 0.1829136, 0.2699426, 0.1927199, 
    0.1240346, 0.1597434, 0.2833536, 0.4041296, 0.3532624, 0.3082039, 
    0.3549927, 0.4574835, 0.4397316, 0.4876918, 0.4739999, 0.3194128, 
    0.4399053, 0.2516366, 0.148961, 0.1827448,
  0.27213, 0.2850121, 0.2385064, 0.2802902, 0.3550478, 0.3528214, 0.4089161, 
    0.3895411, 0.3888977, 0.1866024, 0.2432515, 0.3217834, 0.4269666, 
    0.4091326, 0.3038554, 0.3636231, 0.4056968, 0.472924, 0.4296195, 
    0.3240173, 0.2799442, 0.3163729, 0.3492014, 0.4379435, 0.4943071, 
    0.4293747, 0.39499, 0.3622322, 0.3219197,
  0.3668423, 0.3185776, 0.3060063, 0.3153197, 0.3438336, 0.3433571, 
    0.3953376, 0.3413321, 0.3166898, 0.2657971, 0.2730751, 0.3074805, 
    0.3068084, 0.2582624, 0.2446848, 0.2584162, 0.2445387, 0.2263591, 
    0.178879, 0.2075016, 0.1687804, 0.1731699, 0.2390921, 0.16888, 0.0365228, 
    0.1815476, 0.3862514, 0.3518778, 0.3675286,
  0.2852303, 0.1572602, 0.1056198, 0.2476464, 0.2506303, 0.2059172, 
    0.1840899, 0.1631743, 0.1528619, 0.09670115, 0.1499448, 0.0870204, 
    0.04535884, 0.2136055, 0.2892087, 0.1062394, 0.1421871, 0.1850068, 
    0.161677, 0.2017471, 0.2229625, 0.3433748, 0.1798787, 0.104099, 
    0.02022537, 0.1953663, 0.2451629, 0.262839, 0.2328249,
  0.04194866, 0.06688886, 0.06112754, 0.04049655, 0.04928869, 0.04560062, 
    0.0226125, 0.00731806, 0.04986259, 0.00697355, 0.01924583, -2.169209e-05, 
    0.005003834, 0.02546482, 0.07205684, 0.07762131, 0.07579619, 0.1152231, 
    0.08532692, 0.01431177, 0.01822258, 0.006973463, 0.04236443, 0.0223756, 
    0.05545679, 0.02577413, 0.03671565, 0.003428367, 0.01158034,
  0.03269272, 0.03821478, 0.07068177, 0.01093675, 0.04391513, 0.02024999, 
    0.02684907, 0.003290075, 0.02893327, 0.007822964, 7.621171e-05, 
    0.0142859, 0.02769651, 0.005845988, 0.01943862, 0.01826483, 0.01950207, 
    0.0115758, 0.001287683, 0.0005689249, 0.002920442, 0.002154584, 
    0.07614143, 0.231446, 0.03810141, 0.19315, 0.002320434, 0.0005631691, 
    0.003146969,
  0.06123189, 0.03831594, 0.0279713, 0.01208794, 0.007085315, 0.00877491, 
    0.004590962, 0.02587378, 0.01464846, 0.01674434, 0.01245908, 0.02739577, 
    0.02118441, 0.003073631, 0.01130472, 0.01094405, 0.004005612, 0.01013291, 
    0.002891675, 0.008878618, 0.01619519, 0.0263046, 0.03399915, 0.01113726, 
    0.02007604, 0.04180555, 0.00887199, 0.001661086, 0.01200897,
  0.01487737, 0.003307343, 0.0126556, 0.006686231, 0.03941948, 0.01366157, 
    0.008014099, 0.002905062, 0.024885, 0.1136329, 0.01867764, 0.02941429, 
    0.009385559, 0.005229182, 0.01156532, 0.007757476, 0.01695397, 
    0.04127718, 0.01153419, 0.06732225, 0.1927014, 0.1996884, 0.2140206, 
    0.01133655, 0.003185346, 0.01832809, 0.00499728, 0.009406403, 0.01671227,
  -3.453999e-08, 2.689536e-08, 8.19968e-08, 0.0009256871, 0.01296372, 
    0.01845996, 0.003765514, 0.009812158, 0.001938054, 0.01286331, 0.0257731, 
    0.01878358, 0.00525571, 0.007624181, 0.001632118, 0.00169619, 
    0.006773845, 0.050183, 0.03939809, 0.02261655, 0.004750675, 0.002020002, 
    0.3704305, 0.0843287, 0.0005304778, 0.006344274, 0.01830419, 0.003137991, 
    3.198446e-05,
  1.872743e-08, 1.076569e-08, 1.1149e-09, 6.47393e-05, 2.139186e-09, 
    0.003293018, -3.414165e-05, 0.0007692775, 0.01147879, 0.23042, 
    0.04789515, 0.04995601, 0.02443128, 0.01065374, 0.003327493, 0.01007473, 
    0.01468394, 0.01668385, 0.05389655, 0.06082226, 2.870092e-05, 0.2027597, 
    0.002582399, -0.001715886, 0.002523082, 0.002596814, 0.01507353, 
    0.003910162, 6.589397e-08,
  -2.089486e-05, 0.005338737, 0.0008474235, 0.004608729, 0.001234938, 
    -1.598381e-05, -0.002966566, 0.01786061, 0.06844407, 0.1759904, 
    0.1719924, 0.1060956, 0.1405447, 0.09285513, 0.1776181, 0.1412268, 
    0.05979294, 0.1045888, 0.1468485, 0.02442287, 0.03402426, 0.2150871, 
    0.1091482, 0.09507043, 0.09890842, 0.1132368, 0.03843958, 0.0370019, 
    0.003802068,
  -0.002201297, 0.0149985, 0.01930167, 0.1638175, 0.01319577, 0.001868212, 
    0.1092416, 6.933644e-06, 0.01052214, 0.05168815, 0.1296742, 0.1057445, 
    0.1281046, 0.09657399, 0.09795599, 0.1681907, 0.2526745, 0.2540778, 
    0.2216489, 0.1094075, 0.094868, 0.2155362, 0.1172628, 0.09540533, 
    0.1749477, 0.2078015, 0.0989905, 0.1372845, 0.07867622,
  0.1560919, 0.2147432, 0.1088098, 0.07382613, 0.1191553, 0.1813177, 
    0.1011351, 0.1744908, 0.0774002, 0.07675261, 0.01860694, 0.1489881, 
    0.2057454, 0.2274137, 0.2145069, 0.184987, 0.4012076, 0.3762188, 
    0.2949564, 0.1850777, 0.09533595, 0.06635335, 0.09887767, 0.1615153, 
    0.1570806, 0.1835151, 0.2500874, 0.1814564, 0.2416596,
  0.2249401, 0.2125039, 0.2521718, 0.3803083, 0.4456222, 0.286915, 0.3402044, 
    0.2038716, 0.06529716, 0.09117162, 0.1439442, 0.08334625, 0.1852141, 
    0.2124196, 0.563817, 0.1932729, 0.246381, 0.247896, 0.3076128, 0.2121066, 
    0.1057115, 0.09580455, 0.2518699, 0.09677055, 0.383261, 0.06099411, 
    0.07034379, 0.1567226, 0.2184914,
  0.09297599, 0.1017141, 0.3034202, 0.2072815, 0.36286, 0.2977709, 0.351937, 
    0.3265377, 0.2598398, 0.359376, 0.529355, 0.4189844, 0.3855559, 
    0.2816228, 0.2748781, 0.2252786, 0.2603791, 0.1700804, 0.1714209, 
    0.3711373, 0.3297926, 0.3032694, 0.2738334, 0.08360881, 0.1323835, 
    0.3631229, 0.2527603, 0.07411323, 0.1752397,
  0.1921238, 0.1795577, 0.3665092, 0.4478653, 0.4455309, 0.523879, 0.4979955, 
    0.4362856, 0.4322597, 0.3730072, 0.414214, 0.4701846, 0.4668438, 
    0.4463271, 0.3440421, 0.4056879, 0.3744356, 0.4218075, 0.4658699, 
    0.5053468, 0.4055146, 0.2397071, 0.1536997, 0.08452635, 0.1648008, 
    0.1641731, 0.1230452, 0.2140193, 0.3532311,
  0.2707836, 0.2743719, 0.2779601, 0.2815483, 0.2851366, 0.2887248, 
    0.2923131, 0.2786284, 0.283732, 0.2888356, 0.2939392, 0.2990428, 
    0.3041464, 0.30925, 0.3056944, 0.2941234, 0.2825523, 0.2709813, 
    0.2594103, 0.2478392, 0.2362682, 0.2379149, 0.2407941, 0.2436733, 
    0.2465525, 0.2494317, 0.2523109, 0.2551901, 0.267913,
  0.2587493, 0.2474534, 0.3020123, 0.2972609, 0.3929994, 0.1908039, 
    0.1836174, 0.237002, 0.2427234, 0.2089725, 0.2564432, 0.3916791, 
    0.4254141, 0.01276962, 0.08870939, 0.2860687, 0.3328548, 0.2859488, 
    0.1441375, 0.2485164, 0.5470692, 0.5644061, 0.2141634, 0.0838576, 
    0.08928686, 0.2237344, 0.06304306, 0.03254515, 0.1829346,
  0.1406454, 0.1268599, 0.236935, 0.146067, 0.2275464, 0.199001, 0.05991264, 
    0.3109366, 0.2070269, 0.2089767, 0.1510887, 0.2698386, 0.1326621, 
    0.07255954, 0.1221529, 0.2124998, 0.350619, 0.2977725, 0.2612734, 
    0.2511634, 0.3419575, 0.4195707, 0.4777603, 0.4805533, 0.3262683, 
    0.3369633, 0.1801351, 0.1138427, 0.1499488,
  0.2433622, 0.2364848, 0.1931465, 0.2262733, 0.3088889, 0.328059, 0.3647448, 
    0.3267919, 0.3242947, 0.1329683, 0.2058243, 0.2734324, 0.3846443, 
    0.3557841, 0.2709012, 0.3395046, 0.3843004, 0.443569, 0.4005129, 
    0.2992665, 0.248611, 0.2713563, 0.2883483, 0.3660815, 0.4585309, 
    0.402768, 0.3397029, 0.312383, 0.2637061,
  0.3120133, 0.2593333, 0.275857, 0.3033715, 0.3662329, 0.368689, 0.3556772, 
    0.2987315, 0.28187, 0.2138106, 0.2301193, 0.2604391, 0.2516031, 
    0.2267488, 0.2033785, 0.1989593, 0.2090764, 0.1843114, 0.147442, 
    0.1774763, 0.1422326, 0.1469436, 0.1937702, 0.1490774, 0.08641561, 
    0.2045158, 0.3404647, 0.2969008, 0.3206868,
  0.2249904, 0.08443485, 0.08080452, 0.1998618, 0.1785916, 0.1697099, 
    0.1102611, 0.1829127, 0.1138122, 0.07027025, 0.118839, 0.04857359, 
    0.02797578, 0.1522104, 0.2684727, 0.05071861, 0.1151953, 0.1582721, 
    0.147728, 0.2051459, 0.1697098, 0.2821556, 0.1038343, 0.09628541, 
    0.02183537, 0.1457012, 0.2224488, 0.2180192, 0.1649961,
  0.01225852, 0.0267536, 0.05284608, 0.01985519, 0.02707902, 0.03321192, 
    0.01238625, 0.002788663, 0.02175554, 0.002644927, 0.02043837, 
    3.84363e-06, 0.004134773, 0.01498157, 0.03631347, 0.05396769, 0.05796056, 
    0.06787517, 0.03429163, 0.003439301, 0.006957332, 0.00244861, 0.01584814, 
    0.01338222, 0.04720431, 0.007652297, 0.0179741, 0.001136804, 0.003378039,
  0.01238273, 0.04375103, 0.05037362, 0.002241746, 0.01396099, 0.005988249, 
    0.01060025, 0.0005160628, 0.009330653, 0.002070247, 5.060457e-05, 
    0.008949252, 0.01327515, 0.001791815, 0.008841472, 0.005750046, 
    0.01341495, 0.0009412924, 0.0001073997, 7.553109e-05, 0.001073426, 
    0.0007399382, 0.02612726, 0.09299509, 0.02683739, 0.1771193, 
    0.0005348647, 0.0001025381, 0.001169215,
  0.02284619, 0.009762183, 0.0187679, 0.006065232, 0.002354685, 0.002147529, 
    0.0001194137, 0.01325853, 0.002882161, 0.004242486, 0.007957611, 
    0.01784005, 0.006692695, 0.0003583203, 0.002472924, 0.005129464, 
    0.0003880276, 0.003428603, 0.0006115125, 0.003376818, 0.005914109, 
    0.009270796, 0.01073734, 0.01342219, 0.01385967, 0.04574443, 0.001038009, 
    0.0004473853, 0.003405993,
  0.003771221, 0.001227039, 0.008995559, 0.006664562, 0.01385535, 0.01033569, 
    0.001588149, 0.0008501898, 0.01938386, 0.09778028, 0.007724067, 
    0.008325073, 0.005418812, 0.0006459292, 0.002182375, 0.001239478, 
    0.002082784, 0.004342517, 0.001004891, 0.00910832, 0.05148267, 
    0.03255382, 0.1446241, 0.008165788, 0.001209083, 0.01030121, 
    0.0002199726, 0.002065139, 0.004626377,
  -7.928522e-08, 2.651907e-08, 1.811748e-07, 0.002620878, 0.005624226, 
    0.007985621, 0.0002768891, 0.003531497, 0.0003241609, 0.002884972, 
    0.006372768, 0.008118747, 0.000819061, 0.002519501, 0.0004884807, 
    0.0002123396, 0.0005703706, 0.02273786, 0.01128115, 0.004094453, 
    0.0005944793, 8.972169e-05, 0.2977275, 0.0642869, 0.0002148193, 
    0.00291644, 0.007455228, 0.001186362, -8.910772e-06,
  1.827567e-08, 1.040982e-08, 9.173028e-10, 5.124985e-05, 1.983222e-09, 
    0.001142978, -1.114348e-05, 0.0002928454, 0.008128338, 0.1703931, 
    0.01719646, 0.02517107, 0.004179548, 0.003954399, 0.001569431, 
    0.002916769, 0.007782461, 0.002914479, 0.02398705, 0.02701461, 
    -2.65718e-05, 0.1631472, 0.0009777492, -0.001189368, 0.00131822, 
    0.001058701, 0.007750571, 0.001948557, 6.38451e-08,
  -4.253272e-06, 0.00470514, 0.0002334681, 0.001509315, 0.001048889, 
    -1.852691e-05, -0.002715116, 0.01312087, 0.05347437, 0.1594464, 0.174656, 
    0.07647766, 0.1185006, 0.05852962, 0.1462456, 0.0907241, 0.03849658, 
    0.08236884, 0.08909348, 0.01217664, 0.03046061, 0.1917074, 0.09442783, 
    0.07067322, 0.05681064, 0.06748211, 0.01557742, 0.01376481, 0.007291199,
  -0.001867169, 0.01349272, 0.01305418, 0.1536253, 0.007694263, 0.0005260044, 
    0.09152777, 7.656178e-06, 0.007828779, 0.03979849, 0.1291576, 0.09330083, 
    0.1088074, 0.08235235, 0.07396369, 0.1350462, 0.2046268, 0.2292398, 
    0.1818964, 0.1085146, 0.07265425, 0.1916251, 0.1046245, 0.0755222, 
    0.1380645, 0.1279747, 0.05345958, 0.08268945, 0.06158964,
  0.1109339, 0.1523692, 0.0771254, 0.06272948, 0.1039487, 0.1826542, 
    0.06900696, 0.1461215, 0.06423654, 0.07141295, 0.01999929, 0.1483882, 
    0.1517597, 0.181892, 0.1908894, 0.1671875, 0.3935613, 0.3532935, 
    0.2542921, 0.1698477, 0.08078945, 0.05260143, 0.07779348, 0.1808142, 
    0.1178621, 0.148097, 0.2069986, 0.1231079, 0.1979283,
  0.1656311, 0.225865, 0.2313862, 0.3555818, 0.3906563, 0.2330761, 0.258037, 
    0.1764024, 0.04625938, 0.06903609, 0.1279257, 0.1118072, 0.1624798, 
    0.1756784, 0.4914261, 0.1959619, 0.2277533, 0.2284251, 0.2614015, 
    0.2091213, 0.1066701, 0.07091736, 0.242793, 0.1054766, 0.3186979, 
    0.03996553, 0.05798716, 0.1322087, 0.1946221,
  0.0548795, 0.07725664, 0.270739, 0.1244322, 0.3276906, 0.2543816, 
    0.3539221, 0.2790271, 0.2359942, 0.3619266, 0.5322554, 0.4175507, 
    0.4560314, 0.3354238, 0.25588, 0.3165281, 0.2902534, 0.195838, 0.1755072, 
    0.3922047, 0.3031942, 0.3848727, 0.2882121, 0.08793522, 0.1264728, 
    0.3286646, 0.2662808, 0.05666686, 0.1197729,
  0.2110156, 0.1738014, 0.4675841, 0.4906239, 0.4552997, 0.5304193, 
    0.5327755, 0.5202435, 0.4930971, 0.4007508, 0.4470048, 0.5069188, 
    0.5249823, 0.4999783, 0.4017006, 0.4894863, 0.4452917, 0.5138996, 
    0.5735401, 0.5369578, 0.4534944, 0.2273964, 0.171119, 0.1457233, 
    0.1578803, 0.1727703, 0.1106261, 0.2395407, 0.4033494,
  0.3068349, 0.3060478, 0.3052606, 0.3044734, 0.3036863, 0.3028991, 
    0.3021119, 0.2476685, 0.2574751, 0.2672817, 0.2770883, 0.2868949, 
    0.2967014, 0.306508, 0.3797838, 0.3723371, 0.3648905, 0.3574438, 
    0.3499972, 0.3425505, 0.3351039, 0.3530459, 0.3514731, 0.3499003, 
    0.3483276, 0.3467548, 0.3451821, 0.3436093, 0.3074647,
  0.2940012, 0.2136553, 0.2605517, 0.2450943, 0.3730365, 0.1715431, 
    0.1738717, 0.2491561, 0.1562306, 0.1560695, 0.1957127, 0.3413951, 
    0.4237588, 0.006961151, 0.1395396, 0.3692552, 0.4568566, 0.380483, 
    0.1640221, 0.2635519, 0.5063616, 0.6240342, 0.1822486, 0.07412196, 
    0.09835909, 0.2934759, 0.06763744, 0.01880582, 0.1824495,
  0.09446543, 0.09022247, 0.1757598, 0.09472921, 0.165436, 0.1855497, 
    0.0466978, 0.2496488, 0.1740441, 0.1729049, 0.1195294, 0.2605527, 
    0.07871068, 0.03935043, 0.09354124, 0.1492298, 0.3064167, 0.2419579, 
    0.2120197, 0.1844606, 0.2685697, 0.3759289, 0.4461799, 0.4486187, 
    0.3086364, 0.2489185, 0.1323676, 0.08950792, 0.1096891,
  0.2032185, 0.1746472, 0.1461534, 0.1772042, 0.2627895, 0.280422, 0.3045111, 
    0.266839, 0.2520528, 0.1031599, 0.1655855, 0.2209313, 0.3390889, 
    0.2906267, 0.2160463, 0.298519, 0.3332243, 0.3922311, 0.35074, 0.2570804, 
    0.2006218, 0.2008902, 0.2201066, 0.2825633, 0.396433, 0.3480662, 
    0.2967322, 0.249649, 0.2018616,
  0.2414863, 0.2004124, 0.2045747, 0.2569002, 0.3188054, 0.3444511, 
    0.3050935, 0.2508753, 0.217529, 0.1567676, 0.1711859, 0.1998787, 
    0.1837829, 0.1662065, 0.1499396, 0.1663183, 0.1667687, 0.1420095, 
    0.1064995, 0.1355031, 0.1045767, 0.1176223, 0.1521467, 0.1172128, 
    0.1116632, 0.1916665, 0.2959957, 0.2662095, 0.2722343,
  0.1467166, 0.04299862, 0.06443081, 0.1517523, 0.1253853, 0.1361479, 
    0.07036559, 0.1663306, 0.08649966, 0.04452987, 0.08078194, 0.02176439, 
    0.01995504, 0.1098373, 0.236261, 0.02930704, 0.09267533, 0.1348771, 
    0.1516081, 0.1735474, 0.1311896, 0.1938709, 0.05828716, 0.09270136, 
    0.01340371, 0.1048051, 0.136888, 0.1360246, 0.09378341,
  0.003975013, 0.01387879, 0.0464534, 0.008128368, 0.01426081, 0.02141184, 
    0.006610576, 0.001447796, 0.01289501, 0.001317321, 0.01166387, 
    4.249819e-06, 0.002021846, 0.009532076, 0.01829795, 0.0317889, 
    0.03858646, 0.03176693, 0.015007, 0.001559542, 0.002235201, 0.0009709249, 
    0.008393649, 0.007352728, 0.03841839, 0.002573964, 0.01022407, 
    0.0006048781, 0.001694043,
  0.006408229, 0.03357261, 0.02630809, 0.0007187478, 0.003790206, 
    0.003105811, 0.003092552, 0.0002622013, 0.004187324, 0.001027956, 
    3.130077e-05, 0.004321597, 0.005989468, 0.0006088262, 0.00292192, 
    0.002202847, 0.007976047, -0.000212025, 4.21787e-05, 3.547869e-05, 
    0.0006347845, 0.0003564378, 0.01208466, 0.04813527, 0.01833647, 
    0.1508615, 0.0001348709, 5.364135e-05, 0.0006234253,
  0.01227998, 0.001969857, 0.0156827, 0.002185093, 0.001324947, 0.001020421, 
    1.98236e-05, 0.00793423, 0.001373004, 0.0006594859, 0.003529273, 
    0.010979, 0.002266878, 9.519872e-05, 0.0007137142, 0.002200969, 
    4.658047e-05, 0.001760678, 0.0002488552, 0.001875331, 0.003069493, 
    0.004901745, 0.005401282, 0.01542387, 0.01110028, 0.05175756, 
    -0.0008266324, 0.0002314106, 0.001824526,
  0.001856956, 0.0005969937, 0.01452521, 0.005312996, 0.006501263, 
    0.004779655, 0.0003876382, 0.0004606131, 0.02175752, 0.1142768, 
    0.004404458, 0.004066365, 0.004436044, 0.0002564919, 0.0004993957, 
    0.0002672456, 0.0008139738, 0.0005915253, 0.0002909692, 0.0022178, 
    0.01586678, 0.01250441, 0.03784123, 0.006641121, 0.0003230448, 
    0.004119183, 4.937072e-05, 0.001084769, 0.002293081,
  5.04696e-09, 2.633476e-08, 2.424732e-07, 0.002031328, 0.002361957, 
    0.004518203, -0.0004692138, 0.00198973, 0.0001412086, 0.001318652, 
    0.001177969, 0.003620659, 0.0001580581, 0.0005892347, 0.0002920659, 
    0.0001094675, 0.000161316, 0.008671895, 0.002382708, 0.0005659666, 
    0.0002441196, 3.418465e-05, 0.2034291, 0.04795776, 0.0001234594, 
    0.001686085, 0.003977267, 0.0003578915, -5.765307e-05,
  1.813364e-08, 1.015931e-08, 8.30825e-10, 2.571116e-06, 1.925593e-09, 
    0.0005732934, -2.640785e-05, 0.0001229197, 0.006043062, 0.05441156, 
    0.01130781, 0.01460046, 0.001068461, 0.002363928, 0.0009778297, 
    0.001113711, 0.004526369, 0.001278356, 0.01284653, 0.01628098, 
    -1.848147e-05, 0.1167087, 0.0005882239, -0.001013175, 0.0008430308, 
    0.0005229625, 0.004769491, 0.001227163, 6.394117e-08,
  2.540198e-07, 0.003378917, 0.0001363038, 0.0004514719, 0.001565241, 
    -1.002698e-05, -0.002618158, 0.009587274, 0.03944398, 0.1204793, 
    0.1432891, 0.05553392, 0.08740035, 0.04011877, 0.1088357, 0.05928515, 
    0.02617225, 0.06101634, 0.05597933, 0.007256194, 0.02413338, 0.1668225, 
    0.07518875, 0.04994299, 0.0310125, 0.03853488, 0.00833822, 0.007124758, 
    0.00809102,
  -0.001422044, 0.004197141, 0.01006301, 0.1409228, 0.004534268, 
    0.0001782268, 0.07931069, 7.657861e-06, 0.005162884, 0.03152076, 
    0.1154186, 0.07355621, 0.09258513, 0.06633846, 0.05117526, 0.1040516, 
    0.1560477, 0.219062, 0.1443605, 0.1046701, 0.06667221, 0.164546, 
    0.09187984, 0.05932869, 0.1077386, 0.07299984, 0.0276011, 0.06316454, 
    0.04598227,
  0.07190864, 0.101627, 0.04996694, 0.04515812, 0.1045654, 0.1462692, 
    0.04953497, 0.1221427, 0.05393461, 0.06733254, 0.02568529, 0.1284468, 
    0.1165016, 0.11892, 0.1657097, 0.1471968, 0.3515563, 0.2839088, 
    0.2125347, 0.147238, 0.06712482, 0.03662747, 0.05268966, 0.1667846, 
    0.08827636, 0.1146862, 0.1579645, 0.07273498, 0.1500231,
  0.1131809, 0.2200386, 0.1987529, 0.3138669, 0.3257295, 0.1876569, 
    0.1740185, 0.1331982, 0.03983547, 0.05813058, 0.1021873, 0.118081, 
    0.1602671, 0.1465746, 0.3840427, 0.1764982, 0.2501327, 0.2071657, 
    0.2175456, 0.1801686, 0.0990733, 0.05880213, 0.2276971, 0.1105727, 
    0.2754123, 0.0278681, 0.0461801, 0.1080745, 0.1382599,
  0.03077492, 0.05761674, 0.2528839, 0.07875426, 0.3064893, 0.2597609, 
    0.2902082, 0.2714429, 0.2042549, 0.371573, 0.5292196, 0.4026969, 
    0.5361802, 0.3843162, 0.259953, 0.3831441, 0.2829077, 0.2225223, 
    0.1842173, 0.4162148, 0.2716868, 0.5191607, 0.3772263, 0.1221592, 
    0.1023314, 0.2755376, 0.2689093, 0.03671073, 0.08204778,
  0.3485936, 0.2312172, 0.5424467, 0.4904614, 0.4787991, 0.5067372, 0.575842, 
    0.5277284, 0.5233356, 0.4363179, 0.5203174, 0.5025309, 0.4647878, 
    0.5026272, 0.4834679, 0.5244991, 0.4993073, 0.5054047, 0.5949978, 
    0.618084, 0.5809292, 0.2209169, 0.2010031, 0.2558131, 0.1231327, 
    0.1555591, 0.09301212, 0.2049567, 0.3874481,
  0.164152, 0.1618822, 0.1596123, 0.1573425, 0.1550727, 0.1528029, 0.1505331, 
    0.1085854, 0.1239563, 0.1393272, 0.154698, 0.1700689, 0.1854398, 
    0.2008106, 0.2958373, 0.2936177, 0.2913981, 0.2891785, 0.2869589, 
    0.2847393, 0.2825197, 0.2974204, 0.2865389, 0.2756575, 0.264776, 
    0.2538946, 0.2430131, 0.2321317, 0.1659678,
  0.2767366, 0.214793, 0.2282357, 0.1978236, 0.2467069, 0.1663571, 0.1352503, 
    0.09267824, 0.04262957, 0.08729021, 0.1735962, 0.2580064, 0.3671132, 
    0.006670859, 0.2146627, 0.4590739, 0.4488543, 0.4655587, 0.1367073, 
    0.3025497, 0.5023884, 0.6872541, 0.1559887, 0.06376255, 0.1628162, 
    0.3512397, 0.104766, 0.009479562, 0.1927451,
  0.06000226, 0.06209974, 0.1250492, 0.06897198, 0.1150228, 0.1651732, 
    0.04112238, 0.2062137, 0.1408435, 0.1301863, 0.09246376, 0.2632573, 
    0.04961511, 0.0205565, 0.06375972, 0.1016398, 0.2446924, 0.1823625, 
    0.1677035, 0.1358822, 0.2104705, 0.3080912, 0.3775827, 0.3866128, 
    0.2769836, 0.1882703, 0.09459049, 0.06561602, 0.07583083,
  0.1549779, 0.1172224, 0.111081, 0.1396189, 0.2026448, 0.2174762, 0.2327747, 
    0.19718, 0.1781909, 0.0767578, 0.1248956, 0.1664602, 0.2786586, 
    0.2309773, 0.1546779, 0.2295048, 0.2586672, 0.3365922, 0.2901983, 
    0.2106944, 0.1675868, 0.1304656, 0.1505368, 0.2073941, 0.3087026, 
    0.2802839, 0.2345604, 0.1914301, 0.1494723,
  0.1794793, 0.1426694, 0.1479603, 0.1979014, 0.2640421, 0.2786041, 
    0.2508862, 0.2051454, 0.1558161, 0.1048526, 0.1124456, 0.1306072, 
    0.1212413, 0.111472, 0.1216625, 0.1344829, 0.1195557, 0.09947319, 
    0.06908285, 0.09087278, 0.07299035, 0.07989202, 0.1051216, 0.09151763, 
    0.1064216, 0.1513885, 0.2382126, 0.2243149, 0.209719,
  0.08810169, 0.02355766, 0.04663825, 0.1058031, 0.07538188, 0.09803544, 
    0.04338169, 0.1172954, 0.05250152, 0.02192076, 0.04850477, 0.01195107, 
    0.01261977, 0.06717551, 0.2067952, 0.01731475, 0.06869406, 0.09900969, 
    0.1156186, 0.1235241, 0.08900569, 0.1222333, 0.03690972, 0.08406433, 
    0.006496633, 0.07098576, 0.09816778, 0.08020733, 0.05245068,
  0.002247144, 0.008872569, 0.03652854, 0.003857081, 0.006053775, 
    0.009622326, 0.002877541, 0.0008717794, 0.00892595, 0.0008729004, 
    0.005835738, -5.09825e-07, 0.002126899, 0.003297358, 0.008307637, 
    0.01490644, 0.01809277, 0.0123714, 0.005316869, 0.0007177047, 
    0.0009425251, 0.0005976366, 0.005382085, 0.004362458, 0.03029195, 
    0.0009447684, 0.004532421, 0.0003920495, 0.00110545,
  0.004048014, 0.02611789, 0.01104864, 0.0004376332, 0.0003384583, 
    0.00197698, 0.001136094, 0.0001654667, 0.002255794, 0.0006685374, 
    2.144567e-05, 0.00158043, 0.002641707, 0.0003741691, 0.001044632, 
    0.001120677, 0.003819233, -8.104651e-05, 2.41924e-05, 2.248241e-05, 
    0.0004405195, 0.0002176783, 0.00710159, 0.03077361, 0.01125446, 
    0.1167048, 6.485068e-05, 3.459812e-05, 0.0003986947,
  0.008010394, 0.0002304551, 0.01283796, 0.002341754, 0.0008672804, 
    0.0006263654, 2.475337e-05, 0.003628112, 0.001006292, -0.0004259727, 
    0.001724785, 0.005261709, 0.0008537216, 4.039861e-05, 0.0002348495, 
    0.001008603, 1.76817e-05, 0.0009108754, 0.0001849445, 0.001267248, 
    0.001922981, 0.003164397, 0.003389845, 0.01466351, 0.01612908, 
    0.04856057, -0.0008580574, 0.0001494978, 0.001180285,
  0.001146078, 0.0001818522, 0.0100321, 0.003693798, 0.002943228, 
    0.002200458, 0.0002344859, 0.0002992288, 0.02452349, 0.117043, 
    0.002180638, 0.002532547, 0.002306624, 0.0001570335, 0.0001645906, 
    0.0001229868, 0.0004886704, 0.0002798679, 0.0001549129, 0.001098117, 
    0.008276087, 0.007060126, 0.0184845, 0.005669089, -1.99982e-05, 
    0.001554337, 2.358145e-05, 0.0007219694, 0.001432874,
  9.654373e-09, 2.626886e-08, 2.303042e-07, 0.001630389, 0.0009592902, 
    0.002997021, -0.0005941462, 0.001429317, 7.874552e-05, 0.000864994, 
    0.000516715, 0.001479522, 5.724065e-05, 0.0001823228, 0.0002024479, 
    7.113266e-05, 4.642578e-05, 0.002857049, 0.0008772264, 0.0002547439, 
    0.0001529428, 1.900877e-05, 0.1511969, 0.03048722, 8.034736e-05, 
    0.00113126, 0.002566906, 0.0001979527, -0.0002057883,
  1.821497e-08, 9.990027e-09, 7.986979e-10, -1.590414e-06, 1.89113e-09, 
    0.0003540739, -6.407079e-05, 7.724926e-05, 0.004433237, 0.01515557, 
    0.008156309, 0.005739785, 0.0005456874, 0.001631457, 0.0006967956, 
    0.0006653937, 0.002863413, 0.0007991158, 0.008123951, 0.01143274, 
    -1.141002e-05, 0.09056963, 0.0004390664, -0.000946375, 0.0006079963, 
    0.0003585501, 0.003345251, 0.000878062, 6.433309e-08,
  -4.522142e-06, 0.002145439, 7.015563e-05, 0.0002315875, 0.001594324, 
    -4.195903e-06, -0.002443838, 0.01006002, 0.03205553, 0.07599287, 
    0.1197868, 0.03403668, 0.05418991, 0.02901077, 0.0754451, 0.03928652, 
    0.01950248, 0.04453833, 0.03624268, 0.005031788, 0.01867216, 0.1331306, 
    0.05137754, 0.03122827, 0.01787554, 0.02222892, 0.005424001, 0.004662494, 
    0.007146767,
  -0.001226419, 0.001908943, 0.007639902, 0.1299554, 0.002711394, 
    4.124301e-05, 0.0670734, 6.248915e-06, 0.003740749, 0.02480786, 
    0.09658322, 0.05579969, 0.07474034, 0.04739668, 0.03245229, 0.07387133, 
    0.1092865, 0.1708581, 0.1029105, 0.09641962, 0.06004796, 0.1305413, 
    0.08235118, 0.04678067, 0.08160102, 0.04243127, 0.01502887, 0.04427211, 
    0.03157764,
  0.04296122, 0.07069113, 0.03089296, 0.03128817, 0.08830201, 0.1478138, 
    0.03773984, 0.1061362, 0.05081677, 0.0638114, 0.02438432, 0.1046254, 
    0.09231403, 0.08329193, 0.1414344, 0.1124105, 0.2760383, 0.2150699, 
    0.1475771, 0.1322744, 0.05716582, 0.01674072, 0.03642874, 0.13395, 
    0.06873292, 0.09232299, 0.1162857, 0.04200291, 0.1002711,
  0.07443871, 0.1992119, 0.1567153, 0.258375, 0.2725247, 0.1563404, 
    0.1359978, 0.1001852, 0.04337918, 0.05369284, 0.07957609, 0.1233905, 
    0.1733114, 0.1251773, 0.3199364, 0.1584157, 0.2646008, 0.1843936, 
    0.170067, 0.1527081, 0.08614492, 0.05998995, 0.179583, 0.1447709, 
    0.2457226, 0.0216753, 0.03654703, 0.07929, 0.09130752,
  0.02081629, 0.04235681, 0.2362496, 0.05212883, 0.2877561, 0.2871343, 
    0.3147323, 0.2639755, 0.1790175, 0.3655142, 0.4883686, 0.3410083, 
    0.5653451, 0.3705739, 0.2525048, 0.401608, 0.2540186, 0.191054, 
    0.1962659, 0.3605266, 0.2157433, 0.5971173, 0.3416207, 0.2099038, 
    0.08849447, 0.183457, 0.2752193, 0.02389136, 0.05709291,
  0.4044425, 0.2370979, 0.5394688, 0.4673513, 0.4971722, 0.479369, 0.5085163, 
    0.4603063, 0.4607689, 0.4804412, 0.5312172, 0.4513823, 0.4190042, 
    0.4638894, 0.4566303, 0.3891575, 0.3967497, 0.4394919, 0.5399687, 
    0.5501336, 0.5442064, 0.211674, 0.241069, 0.3860603, 0.1142065, 
    0.08851494, 0.09504931, 0.2320069, 0.3415759,
  0.08443969, 0.08230194, 0.08016419, 0.07802643, 0.07588867, 0.07375091, 
    0.07161316, 0.0679916, 0.0776552, 0.08731882, 0.09698242, 0.106646, 
    0.1163096, 0.1259732, 0.1519034, 0.1539089, 0.1559144, 0.1579199, 
    0.1599254, 0.1619309, 0.1639364, 0.1987, 0.1891687, 0.1796373, 0.1701059, 
    0.1605746, 0.1510432, 0.1415119, 0.0861499,
  0.2978669, 0.2364064, 0.1597067, 0.04414133, 0.08969007, 0.1426584, 
    0.08972612, 0.03364779, 0.01594756, 0.0370524, 0.1112743, 0.2627877, 
    0.3104573, 0.006324554, 0.3048322, 0.5414567, 0.3718613, 0.459754, 
    0.1025645, 0.3079869, 0.4832693, 0.7016703, 0.1446165, 0.05843614, 
    0.2114241, 0.4021363, 0.1309277, 0.00760132, 0.1929209,
  0.04189728, 0.04859331, 0.09991778, 0.0546023, 0.08978738, 0.1358089, 
    0.03734702, 0.1865681, 0.1291121, 0.1143709, 0.07644081, 0.2453142, 
    0.03313877, 0.01621291, 0.04577562, 0.07699709, 0.1826915, 0.1390667, 
    0.1311461, 0.1077086, 0.1690712, 0.2517253, 0.3089728, 0.338584, 
    0.2358269, 0.1497813, 0.07265663, 0.05053148, 0.05813925,
  0.1268059, 0.09090538, 0.0875717, 0.1166311, 0.1601678, 0.1725312, 
    0.187102, 0.1536482, 0.1353775, 0.06239418, 0.1024271, 0.1364302, 
    0.2273581, 0.1824759, 0.1121883, 0.178851, 0.2015565, 0.2945093, 
    0.2346995, 0.1675185, 0.1179672, 0.09339712, 0.103831, 0.1543643, 
    0.2347409, 0.2210918, 0.188103, 0.1534781, 0.1220283,
  0.1407431, 0.1098756, 0.1129777, 0.1622034, 0.2113563, 0.2295552, 
    0.2116901, 0.1696954, 0.1237793, 0.07886475, 0.07981318, 0.08834057, 
    0.07947511, 0.07637285, 0.08828012, 0.1058696, 0.08622579, 0.06684382, 
    0.04927746, 0.06203472, 0.05381277, 0.06168848, 0.07850422, 0.07708424, 
    0.09127159, 0.1173657, 0.1929328, 0.180776, 0.1692331,
  0.05732019, 0.01526467, 0.03322675, 0.0661926, 0.04243811, 0.06585709, 
    0.02586862, 0.08388629, 0.0331133, 0.01146604, 0.04004222, 0.008256258, 
    0.008164953, 0.04090482, 0.1850507, 0.0111688, 0.04641251, 0.07285582, 
    0.07840571, 0.07373603, 0.05135098, 0.07428244, 0.02466201, 0.07657705, 
    0.004388661, 0.05374369, 0.05808419, 0.04772121, 0.03247374,
  0.001620926, 0.006458747, 0.03004117, 0.002409701, 0.002400112, 0.00372537, 
    0.001460631, 0.0006468006, 0.006896318, 0.0006576033, 0.003289119, 
    -8.382485e-07, 0.002032098, 0.001410689, 0.004547242, 0.007383166, 
    0.009760198, 0.006470799, 0.002686468, 0.0004485698, 0.0005140632, 
    0.0004378278, 0.003949173, 0.003239635, 0.01980826, 0.0004803907, 
    0.002125931, 0.0002905287, 0.0008279823,
  0.002949199, 0.02091291, 0.006609923, 0.0003267171, -0.0007132509, 
    0.001371697, 0.000556241, 0.0001215349, 0.001545454, 0.0004967656, 
    9.56902e-06, 0.0007281448, 0.001851826, 0.000281398, 0.0004753792, 
    0.0007400448, 0.002026399, 5.841256e-06, 1.689429e-05, 1.64254e-05, 
    0.0003405051, 0.000143641, 0.004946158, 0.02286285, 0.007441771, 
    0.09421495, 4.625809e-05, 2.55603e-05, 0.0002915386,
  0.005938478, -0.0002635006, 0.01336695, 0.00980811, 0.0006455574, 
    0.0004440372, 2.782518e-05, 0.001736056, 0.0008053986, -0.0003078834, 
    0.001087381, 0.002567694, 0.0003525279, 3.029215e-05, 0.0001430486, 
    0.0006081953, 1.097319e-05, 0.0004791533, 0.0001529074, 0.0009587992, 
    0.00138042, 0.002322968, 0.002454059, 0.01192326, 0.01314966, 0.03697754, 
    -0.0009233023, 0.0001105296, 0.0008766634,
  0.0008156968, 0.005627551, 0.006682286, 0.002366748, 0.001411941, 
    0.001079022, 0.00017009, 0.0002185151, 0.02488447, 0.1220774, 
    0.001043569, 0.001806422, 0.001253158, 0.0001180118, 8.364986e-05, 
    8.014074e-05, 0.0003453658, 0.0001763344, 0.0001074843, 0.0007001581, 
    0.00555456, 0.004887643, 0.01171329, 0.005904843, 0.0005149783, 
    0.0006985327, 1.507826e-05, 0.0005415177, 0.001030111,
  8.270838e-09, 2.631042e-08, 2.35795e-07, 0.0007518437, 0.0006083775, 
    0.002236086, -0.0004385836, 0.001093136, 1.211299e-05, 0.0005817582, 
    0.0003438185, 0.0007157547, 3.470004e-05, 0.0001088992, 0.0001557032, 
    5.322659e-05, 2.832947e-05, 0.001311718, 0.0005450385, 0.0001672028, 
    0.0001116548, 1.229761e-05, 0.100817, 0.01571039, 5.977522e-05, 
    0.0008529918, 0.001883607, 0.0001340817, -0.0004790954,
  1.831692e-08, 9.845041e-09, 7.66899e-10, -3.748573e-06, 1.880282e-09, 
    0.0002534215, -3.477692e-05, 5.796496e-05, 0.003285805, 0.008462298, 
    0.005339321, 0.002395749, 0.0003704799, 0.001257867, 0.0005474155, 
    0.0004834786, 0.001821343, 0.0005746272, 0.005997107, 0.008923245, 
    -9.177345e-06, 0.07398392, 0.0003506249, -0.0009064641, 0.0004807849, 
    0.0002789485, 0.002592469, 0.0006898809, 6.522372e-08,
  -5.428113e-06, 0.001804705, 2.058684e-05, 0.0001492132, 0.001425388, 
    -2.263142e-06, -0.002325249, 0.0105712, 0.03169838, 0.05614909, 
    0.1015736, 0.0197117, 0.03236794, 0.01886986, 0.05074877, 0.02355266, 
    0.01736796, 0.02624176, 0.02331864, 0.003943845, 0.01639993, 0.1052679, 
    0.03769543, 0.01942006, 0.01280959, 0.01521968, 0.004138318, 0.003494206, 
    0.005450298,
  -0.0011277, 0.001079443, 0.006535457, 0.1219182, 0.001981738, 
    -4.170533e-05, 0.05467403, 5.760782e-06, 0.003025077, 0.01987917, 
    0.08344505, 0.03972517, 0.06042762, 0.03510646, 0.02289797, 0.05271594, 
    0.07231374, 0.1223782, 0.06873245, 0.08671872, 0.05700898, 0.1108265, 
    0.07407547, 0.03974266, 0.06115192, 0.02731043, 0.009127022, 0.03347623, 
    0.02208764,
  0.03063656, 0.05217656, 0.02323441, 0.02984751, 0.08100685, 0.1434982, 
    0.03012331, 0.1035901, 0.05773707, 0.05894474, 0.02255285, 0.08942506, 
    0.0780886, 0.06425622, 0.123094, 0.08930149, 0.2047658, 0.164208, 
    0.1026071, 0.1243213, 0.04780857, 0.01591638, 0.02600098, 0.1033032, 
    0.05861105, 0.07733683, 0.08658946, 0.02829381, 0.06688541,
  0.05350897, 0.2099262, 0.1343403, 0.2311987, 0.2441006, 0.1356781, 
    0.1283102, 0.08795947, 0.04794509, 0.05583702, 0.06774047, 0.1878395, 
    0.2031032, 0.1162779, 0.2836319, 0.1475209, 0.265942, 0.1683002, 
    0.1526298, 0.135463, 0.08059849, 0.07886188, 0.1451858, 0.1807308, 
    0.2280139, 0.01829972, 0.02935921, 0.05933315, 0.06862251,
  0.01662909, 0.03324139, 0.2413545, 0.0401453, 0.2730085, 0.258288, 
    0.3257676, 0.2770384, 0.2252301, 0.4052883, 0.4732426, 0.3103858, 
    0.5729985, 0.3153943, 0.241303, 0.344806, 0.2545747, 0.1642756, 0.187067, 
    0.2723375, 0.1684249, 0.5566428, 0.3648019, 0.2212924, 0.101732, 
    0.1292214, 0.2799112, 0.02274647, 0.0446053,
  0.4254069, 0.290191, 0.4791551, 0.4098929, 0.4207113, 0.3820923, 0.3790518, 
    0.3362329, 0.3569509, 0.4084167, 0.3505739, 0.2695455, 0.2925145, 
    0.3044598, 0.3189493, 0.2453347, 0.2191715, 0.2386025, 0.2913729, 
    0.340854, 0.3481097, 0.2069642, 0.2727171, 0.5280143, 0.1053681, 
    0.03350636, 0.1028995, 0.2302092, 0.3076649,
  0.08015239, 0.07858247, 0.07701255, 0.07544263, 0.0738727, 0.07230278, 
    0.07073286, 0.05804318, 0.06595751, 0.07387184, 0.08178618, 0.08970051, 
    0.09761484, 0.1055292, 0.1338054, 0.1347969, 0.1357885, 0.13678, 
    0.1377715, 0.1387631, 0.1397546, 0.1505055, 0.1431696, 0.1358337, 
    0.1284977, 0.1211618, 0.1138258, 0.1064899, 0.08140833,
  0.2703884, 0.2191936, 0.08607888, 0.006991617, 0.03135999, 0.1043368, 
    0.06037698, 0.009359424, 0.01097459, 0.02209021, 0.0739506, 0.2487794, 
    0.2916582, 0.007503903, 0.3521692, 0.4914738, 0.320632, 0.4199767, 
    0.09327874, 0.3174949, 0.4600945, 0.6949031, 0.1581068, 0.05709052, 
    0.2360958, 0.441218, 0.1591323, 0.01371285, 0.1784165,
  0.03432482, 0.04203754, 0.08734035, 0.04770301, 0.07639213, 0.1143669, 
    0.04096604, 0.1697029, 0.1276224, 0.1038451, 0.06926267, 0.2439419, 
    0.02565665, 0.01387922, 0.03749271, 0.06578098, 0.1479978, 0.1176323, 
    0.110276, 0.08971764, 0.1469584, 0.2193385, 0.2635361, 0.3092672, 
    0.2174066, 0.130666, 0.06207789, 0.04287227, 0.04831973,
  0.1087662, 0.07725848, 0.07537425, 0.1028084, 0.1364965, 0.1476213, 
    0.1621915, 0.1268634, 0.1126241, 0.05199298, 0.08572023, 0.1178105, 
    0.1969137, 0.144404, 0.09122533, 0.1446512, 0.1656482, 0.2505792, 
    0.1948821, 0.1398787, 0.09141043, 0.07673905, 0.07994615, 0.1225914, 
    0.1896471, 0.1803901, 0.1611441, 0.1310697, 0.1055787,
  0.1206577, 0.09301095, 0.09339613, 0.1333881, 0.1810605, 0.1894134, 
    0.1829717, 0.1433821, 0.1063036, 0.06749157, 0.06270318, 0.0660315, 
    0.06132182, 0.05735726, 0.07041349, 0.08283629, 0.0658728, 0.04976023, 
    0.03852768, 0.04965208, 0.04286194, 0.05045858, 0.06353985, 0.08213264, 
    0.08006789, 0.09877916, 0.1579167, 0.1430025, 0.1413395,
  0.04131824, 0.01191786, 0.02414757, 0.04261949, 0.02663226, 0.04057651, 
    0.01789228, 0.05922873, 0.02239126, 0.007809453, 0.02764316, 0.006475323, 
    0.005795455, 0.02737813, 0.1868931, 0.008202258, 0.02976744, 0.05198736, 
    0.05608182, 0.05161369, 0.03603724, 0.04953391, 0.01715121, 0.07708811, 
    0.003454339, 0.04347293, 0.03733144, 0.0348954, 0.02333356,
  0.001330646, 0.005327936, 0.03574323, 0.001926705, 0.0013592, 0.001984868, 
    0.0009828872, 0.0005421399, 0.005884741, 0.0005580988, 0.00224384, 
    -7.312686e-07, 0.006307924, 0.001015287, 0.003192473, 0.004567401, 
    0.006544466, 0.004200184, 0.002052413, 0.0003488924, 0.0003796215, 
    0.0003611603, 0.003275577, 0.002592172, 0.04824961, 0.0003749634, 
    0.001385398, 0.0002428993, 0.0006922788,
  0.002465455, 0.0173973, 0.02533993, 0.0002582269, -0.001180908, 
    0.001112801, 0.0003930388, 0.0001029212, 0.001255072, 0.0004090285, 
    -3.066222e-05, 0.001268564, 0.001484123, 0.0002386199, 0.0003459422, 
    0.0005836721, 0.001385079, 2.560994e-05, 1.365832e-05, 1.342873e-05, 
    0.0002877606, 0.0001142131, 0.003992031, 0.01883739, 0.01907955, 
    0.1383326, 3.85747e-05, 2.151046e-05, 0.0002435127,
  0.004899989, -0.0006374699, 0.03651537, 0.08075745, 0.0004855675, 
    0.0003542499, 2.520582e-05, 0.001124321, 0.0006404468, -0.0002874067, 
    0.0008383488, 0.001656605, 0.0002175616, 2.421469e-05, 0.000110295, 
    0.0004655218, 8.464247e-06, 0.0003539987, 0.0001201836, 0.0007982156, 
    0.001132308, 0.001914684, 0.00199994, 0.05708574, 0.04881796, 0.06423792, 
    -0.0007422072, 9.264364e-05, 0.0007304978,
  0.0006536298, 0.1041057, 0.01002447, 0.001477024, 0.0009274636, 
    0.000728749, 0.0001383322, 0.0001781894, 0.03315398, 0.1384017, 
    0.0006722094, 0.001443657, 0.0008329798, 8.32925e-05, 5.938219e-05, 
    6.260119e-05, 0.0002782807, 0.0001437886, 8.800038e-05, 0.0005277706, 
    0.004265846, 0.003680327, 0.008864595, 0.03296178, 0.0312006, 
    0.0004371787, 1.214405e-05, 0.0004494515, 0.0008318104,
  -1.279609e-07, 2.636618e-08, 2.3576e-07, 0.001034359, 0.000268891, 
    0.001857673, -0.000397349, 0.0008265359, -7.921972e-05, 0.0004701825, 
    0.00027206, 0.0005002783, 2.798756e-05, 8.145429e-05, 0.0001359938, 
    4.582967e-05, 2.259683e-05, 0.0008450468, 0.0004249341, 0.0001352841, 
    9.256709e-05, 1.170295e-05, 0.1156796, 0.01343175, 5.043099e-05, 
    0.0007101728, 0.001557889, 0.0001057953, -0.001272571,
  1.840037e-08, 9.777056e-09, 7.586295e-10, -1.670094e-06, 1.875216e-09, 
    0.000205542, -2.546698e-05, 4.893739e-05, 0.01005674, 0.005931227, 
    0.003719791, 0.001604079, 0.000299112, 0.001025499, 0.0004738189, 
    0.00040737, 0.001372574, 0.0004724653, 0.00503033, 0.007640912, 
    -8.058675e-06, 0.06737334, 0.000304963, -0.001078653, 0.00041632, 
    0.0002387633, 0.002215251, 0.0005901219, 6.585103e-08,
  -4.767492e-06, 0.001308759, -5.368889e-05, 0.0001146201, 0.00132114, 
    -1.5201e-06, -0.002330509, 0.01811955, 0.04117473, 0.04888322, 
    0.07391479, 0.01291979, 0.02193551, 0.01170822, 0.03514995, 0.01489376, 
    0.00868772, 0.01289362, 0.01653863, 0.003388842, 0.01561541, 0.09273213, 
    0.04099472, 0.01305609, 0.007602413, 0.01127153, 0.003521822, 
    0.002924946, 0.004476623,
  -0.001009064, 0.0005564761, 0.006676799, 0.126101, 0.001580565, 
    -5.922422e-05, 0.05388568, 5.760926e-06, 0.002655638, 0.01666517, 
    0.08227753, 0.03101552, 0.05427581, 0.02915682, 0.01877123, 0.04090902, 
    0.0529104, 0.0935166, 0.05021959, 0.08229217, 0.06880145, 0.0968971, 
    0.0723917, 0.03477336, 0.04676482, 0.02072388, 0.006796096, 0.0243844, 
    0.01764208,
  0.02579206, 0.04238246, 0.02025882, 0.04783825, 0.09027007, 0.1575215, 
    0.02705211, 0.1379586, 0.09043465, 0.06340084, 0.02133024, 0.1003462, 
    0.07350179, 0.0550692, 0.1079328, 0.07211276, 0.1612837, 0.1291804, 
    0.07562058, 0.1305462, 0.04735264, 0.02503252, 0.0284834, 0.1062028, 
    0.05523032, 0.06907563, 0.07132906, 0.02208601, 0.05085897,
  0.04313881, 0.280559, 0.1441479, 0.2410622, 0.2559252, 0.1600253, 
    0.1468443, 0.1194123, 0.09780625, 0.1155356, 0.08556161, 0.3477122, 
    0.2647689, 0.1395641, 0.2655635, 0.1461111, 0.3121435, 0.1606356, 
    0.2048043, 0.131885, 0.1059514, 0.1528299, 0.114948, 0.2628096, 0.222353, 
    0.01763351, 0.0253228, 0.0492407, 0.0540595,
  0.01452609, 0.02886584, 0.288559, 0.03445327, 0.2572058, 0.2354974, 
    0.3834161, 0.3386992, 0.3472875, 0.4687094, 0.5259359, 0.3776151, 
    0.5372962, 0.325377, 0.2514066, 0.3006887, 0.3125418, 0.1802136, 
    0.1813791, 0.2325556, 0.1659609, 0.4634471, 0.3463341, 0.2763201, 
    0.08673499, 0.1203519, 0.2775029, 0.02691832, 0.04006677,
  0.4340492, 0.2299523, 0.4205144, 0.3330821, 0.3680149, 0.3097147, 
    0.3185539, 0.2628451, 0.2745905, 0.300802, 0.2500039, 0.2014058, 
    0.2240935, 0.2217972, 0.2418074, 0.1892049, 0.1793842, 0.1742767, 
    0.2134344, 0.2536407, 0.260989, 0.2157911, 0.3267428, 0.5245196, 
    0.1187265, 0.02057488, 0.1019644, 0.2545147, 0.279977,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -4.982908e-05, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.588639e-06, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.751537e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -3.394659e-05, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, -4.549313e-06, 0, -2.036557e-05, 0, 0, 0, 0.0002922295, 0, 
    4.35563e-05, -1.140437e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0005471823, 8.221478e-06, 
    -1.051745e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2.192507e-05, 0, 0, 
    -6.376654e-06, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 3.327438e-05, 0, -0.0002321914, 0, 0, 
    -9.17946e-07, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.113346e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0.001988176, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, -2.831459e-06, 0, 0, 0, 0, 0, 0, 0.0004110957, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, -5.864289e-06, -5.737459e-06, -5.029911e-05, -1.803457e-05, 0, 
    7.226855e-06, 0.0005012339, 0.001339714, 0, 0.0009596986, 0.002177034, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  -1.282235e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0.001085297, 0, 0, 0.001572357, 
    2.054957e-05, -6.980482e-06, 0, -1.09953e-05, 0, 0, 0, 0, 0, 0, 
    -1.664893e-05, -2.270639e-05, 0, -1.672077e-05, -1.529415e-05, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001979887, -5.380756e-05, -0.0003275873, 0, 
    -6.493764e-06, -8.720487e-06, 0, 0, 0, 0, 0, -1.410651e-05, 
    -7.552046e-06, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -4.931072e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0.005210693, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, -2.346175e-05, 0, 0, -3.069837e-05, 0, 0, 0, 0, 0, 0, 
    0.002183353, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, -4.990961e-05, 0, 0, -2.571323e-05, 0.0001440903, -0.0002043074, 
    0.0003909917, 0.0008157503, 7.226855e-06, 0.000290422, 0.001673114, 
    0.002016978, 0.001298395, 0.003515424, -6.009629e-06, 0, 0, 0, 0, 0, 0, 
    0, 0, -3.111212e-05, 0, 0, 0, 0,
  0.001031353, 0.002918942, 0, 0, -1.258949e-05, 0, 0, 0, 0, 0.001364971, 0, 
    0, 0.00507798, 1.232882e-05, -2.747804e-05, 0, -3.848357e-05, 0, 0, 0, 0, 
    0, 0, -0.000103633, 0.0007779457, 0, -8.39569e-05, 2.427104e-05, 
    -1.222183e-05,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0.006435046, -0.0001200141, 0.0004857879, 
    -3.215584e-05, 0.003646648, -1.009741e-05, -3.83336e-06, 0, 
    -3.009452e-06, 0, 0, 3.301667e-05, -2.214742e-05, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001071686, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0.0001166661, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.416201e-05, 
    0, 0, 0, 0, 0, 0, 0, -3.182071e-05, 0, 0, 0, 0,
  0, 0, 0, 0, 0.009324664, 0, -3.702887e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, -5.289266e-05, 0, 0, -9.300836e-05, 0, 0, 0, 0, 0, 0, 
    0.004408256, -2.524221e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, -4.993596e-05, 0, 0, 3.85595e-05, 0.0009725309, 0.0008010789, 
    0.0003690304, 0.003743603, 7.226855e-06, 0.006781443, 0.002286253, 
    0.005787685, 0.003232117, 0.007891246, 0.0005779298, 0, 0, 0, 0, 0, 0, 0, 
    -1.689933e-05, 8.40684e-05, 0, 0, 0, 0,
  0.001568581, 0.003357824, 0, 0, -2.636506e-05, 0, 0, 0, 0, 0.005062279, 0, 
    0, 0.009493031, -9.113965e-06, 0.006417122, 0, 2.445071e-07, 0, 
    -4.485226e-05, 0, 0, 0, 0, 0.0007095763, 0.002638463, -1.148966e-05, 
    0.0001905084, 8.516332e-06, -4.190482e-05,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01415502, -0.0001841759, 0.0009809866, 
    -5.175433e-05, 0.01091324, -4.279814e-05, 0.001648023, 0, -1.504726e-05, 
    0, 0, 0.0003237904, -8.730748e-05, 0, 0, -2.264747e-05, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.00778585, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 6.407183e-08, 0, 0, 0, 0, 0.0002350171, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0.0003753766, -2.664609e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0008581914, 0, 0, 0, 0, -4.762856e-05, 0, 0, -7.682097e-05, 
    0.0007835334, 0, 0.000345455, 0,
  0, 0, 0, 0, 0.01373675, 0, 0.001949758, 0, 0, 0, 0, 0, 0, 0, 0, 
    -0.0001112873, 0, 0, 0, 6.402638e-05, 0, 0, 0, 0, 0, 0.0003884704, 0, 0, 0,
  0, 0, 0, 0, 0.0006976846, 0, 0, -0.0001009488, 0, 0, 0, 0, 0, 0, 
    0.01411102, -0.0001310068, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, -5.808238e-05, 0, -5.254239e-06, -2.506715e-07, 0.00323106, 0.002365879, 
    0.000553872, 0.00624895, 1.7755e-05, 0.01481116, 0.004245217, 
    0.008288412, 0.00451867, 0.01807321, 0.002551986, 0, 0, 0, 0, 0, 0, 0, 
    -6.124311e-05, -2.522253e-05, 0, 0, 0, 0,
  0.005575981, 0.007856162, 0, 0, -5.582e-05, 0, 0, 0, -5.506668e-06, 
    0.0092134, 0, 0, 0.01549367, 0.001657553, 0.006338397, -5.26488e-06, 
    0.0004536364, 0, -4.221982e-05, -2.828489e-06, 0, 0, 0, 0.00361709, 
    0.006531043, -2.683687e-05, 0.005036314, 0.001079596, 0.0004132146,
  0, 0, 0, -6.466195e-07, 0, 0, 0, 0, 0, 0.02330115, -2.487402e-05, 
    0.009837273, 0.001698191, 0.01901486, -0.0001692335, 0.002645934, 
    0.0001965236, -9.756765e-05, 0, -1.301727e-05, 0.0003162728, 
    -0.0001806971, 0, -2.152322e-06, -4.999885e-05, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.02053204, -2.062076e-05, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, -1.515242e-05, 0.0002380376, 0, 0, 0, 0, 0.00576581, 
    -5.954401e-05, 0, -2.731707e-05, -6.945463e-06, 0, 0, 0, 0, 0, 0, 0, 
    -0.000176945, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -9.997801e-06, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  -1.565651e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0.002312988, 0.0009096214, 0, -2.98903e-05, 0.001326647, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.003165649, 0, -5.766179e-05, -8.045085e-06, 0.002018158, 
    0.001891381, 0, 0, 0.0003589709, 0.00188274, 0.0003979768, 0.003418199, 0,
  0, 0, -8.032872e-06, 2.270813e-05, 0.0190688, 0, 0.005614171, 0, 0, 0, 0, 
    0, 0, 0, -0.0001251815, 9.755229e-05, 0, 0, -4.108694e-07, 0.001166473, 
    0, 0, 0, 0, -5.717887e-07, 0.002813481, -1.06845e-05, 0, 0,
  0, 0, 0, -6.619791e-06, 0.003239863, 0, 0, -0.0001541325, 0, 0, 0, 0, 0, 0, 
    0.03077478, 6.817542e-05, 0, 0, 0.001696173, 0, 0, 0, 0, 0, 
    -4.322786e-06, 0, 0, 0, 0,
  0, 0.002456032, -8.834115e-06, 9.837589e-05, -5.895288e-05, 0.005318365, 
    0.007201771, 0.003662288, 0.009661874, -2.073634e-05, 0.02456182, 
    0.005135377, 0.01047908, 0.007186354, 0.03268987, 0.009154079, 0, 0, 0, 
    0, 0, 0, 0, -0.0002746487, -0.0002482854, 0, 0, 0, 0,
  0.01494445, 0.01241186, -1.000736e-05, 0, 1.399831e-05, 0, 0, 0, 
    -2.921213e-05, 0.01301552, 0.0006958214, 0, 0.02361177, 0.006930692, 
    0.007587413, -2.714939e-05, 0.0008376453, -4.914604e-06, -6.217674e-05, 
    -1.158191e-05, 0, 0, -3.917224e-06, 0.00839805, 0.008913366, 
    -2.986219e-05, 0.01370488, 0.002157208, 0.0003593566,
  2.62152e-05, 0, 0, 0.0003018248, 0, 0, 0, 0, -1.920877e-05, 0.03790845, 
    0.001824756, 0.01755791, 0.009505156, 0.0293139, -0.0002755883, 
    0.00399769, 0.0007434904, 0.000206558, -8.768735e-09, 7.100723e-05, 
    0.001065403, -0.0003420719, 0, -2.692673e-05, -4.202435e-05, 
    -8.968327e-05, 0, 0, -3.096219e-05,
  0, 0, 0, -2.147116e-06, 0, 0, 0, 0, 0, 0, 0.03135015, -5.324459e-05, 0, 0, 
    0, 0, 0, 6.7843e-05, -5.949689e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0.0006199971, 0.002398144, 0, 0, 0, -3.376394e-05, 0.01302032, 
    -0.0001835722, -5.113342e-05, 3.011298e-05, 0.0008623269, 0, 
    -2.566192e-05, 0, 0, 0, 0, 0, -0.0002606297, 0, -3.844117e-06, 0, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, -0.00011828, 0, 0, 0, 0, 0, 0.002042262, 0, 0.0004686103, 0, 
    0, 0, 0, 0, 0, 0, 0, -0.0001059384, 0, 0.0002789865, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0.0008605591, -8.354057e-06, 0, 0, -2.510617e-05, 4.000365e-06, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.0002505805, -1.393747e-06, 0, 0, 0, 0, 0.001500508, 0, 
    0, 0, 0, 0, 0, -1.732602e-06,
  0, -6.734195e-05, 0, 0.004326927, 0.00667494, 8.947947e-05, 0.0009574854, 
    0.003926392, 0, 0, 0, -1.091734e-05, 0, 0, -6.366228e-06, -2.080268e-05, 
    0.008620853, -3.215476e-05, 0.001445947, 7.295661e-05, 0.009777581, 
    0.005021774, 0.003852193, 0, 0.0005887425, 0.006550919, 0.004018346, 
    0.005331515, -4.480953e-05,
  0, 0, -6.944365e-05, 0.0005719227, 0.02864298, -0.0001366623, 0.01323318, 
    0, 0, 0, 0, 0, 0, 0, 0.001843787, 0.004516501, 0.001170703, 0, 
    0.000728571, 0.005430711, -5.163345e-05, -3.830855e-05, 0, 0, 
    1.807521e-05, 0.007179743, 0.002185031, 0.000308413, 0,
  0, 0, 0, 9.233873e-05, 0.004243927, 0.0006395575, -1.565072e-06, 
    -0.0003719507, -6.080178e-05, 0, 0, 0, -1.671494e-07, 3.946783e-06, 
    0.05067533, 0.002054731, 0.0001235543, 0, 0.004053671, 0, 0, 0, 0, 
    -3.7396e-10, -2.180472e-06, 0, 0, 0, 0,
  0, 0.003831314, -1.061314e-05, 0.003945898, -0.000168067, 0.01713665, 
    0.0174428, 0.007592541, 0.01780051, 0.0001128149, 0.04940473, 0.01384028, 
    0.01648192, 0.01203166, 0.05565523, 0.02702473, 0, 0, 0, 0, 0, 0, 0, 
    0.0005151124, 0.006913236, 0, -2.211696e-05, -4.914607e-06, 0,
  0.02697505, 0.01535512, 0.001777697, -4.124393e-07, 0.0009082974, 0, 0, 
    -3.188412e-05, 0.001496655, 0.02138242, 0.001270665, -1.426278e-06, 
    0.02673441, 0.01997919, 0.00910636, 1.985483e-05, 0.001391195, 
    0.000127146, 0.00192641, -7.159985e-05, 0, 1.873161e-05, -1.125263e-05, 
    0.01472712, 0.02030189, -0.00017237, 0.02518942, 0.009128652, 0.006088982,
  0.0004561086, 0, -5.242366e-06, 0.000582375, -1.810127e-05, 0, 0, 
    -4.486755e-06, -0.0002152129, 0.05477249, 0.00751919, 0.03457623, 
    0.02261993, 0.0540144, 0.0007623098, 0.008986806, 0.002878927, 
    0.001833734, -9.493358e-06, 0.001410768, 0.003692032, 0.0002920251, 
    1.924084e-05, 0.0003143541, 0.001420625, 0.0001753711, 0, 0, 0.0001317295,
  0, 0, 0, -4.748408e-06, 0, 0, 0, -8.917381e-06, -5.091181e-07, 0, 
    0.0368747, -0.0001514727, 0, 0, 0, 0, 0, 0.001549296, -4.872394e-05, 0, 
    0, 0, 0, 0, 0, -8.232159e-07, 0, 0, 0,
  0, 0, 0.0003717093, 0.001078414, 0.004227791, 0, 0, 0, -0.0001560431, 
    0.01974802, 0.004934358, 0.0001095321, 0.006185037, 0.002210234, 0, 
    -5.132384e-05, 0, -1.834372e-05, 0, 1.654297e-07, 0, 0.0006411933, 
    -9.390556e-06, 0.001743144, 0, 0, 0.005645258, 0, 0,
  0, 0, 0, -1.589139e-07, -1.288553e-05, -0.0002867905, 0, 0, 0, 0, 0, 
    0.005908914, 0.005218184, 0.001294466, 4.601962e-05, 0, 0, 0, 0, 0, 0, 
    -5.596443e-06, 0.001166897, 0, 0.0002539688, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -8.455451e-08, 0, -2.212089e-05, -1.061425e-05, 0.001087812, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0.001832415, -7.163129e-05, 0, -1.029801e-05, 0.001370152, 0.001121301, 
    0.002078601, 0, 0, 0, 0, 0, 0, 0, 0, 0.004312964, -7.645478e-05, 
    -6.541557e-06, 0, -2.205611e-06, -3.947485e-05, 0.003181144, 0, 0, 0, 
    -1.227662e-05, 0, -6.062209e-06, 0.002401964,
  0, 0.0005517245, 0, 0.009228114, 0.01690767, 0.003296239, 0.007375409, 
    0.01477937, 0, 0, 0, 0.0001238216, 0, 0, 0.002647444, -3.497853e-05, 
    0.02046312, 0.001767507, 0.005178944, 0.00161539, 0.02129912, 0.01446556, 
    0.0137994, 0.0002566043, 0.002897354, 0.009976864, 0.005129819, 
    0.01411301, -4.812844e-05,
  0, 0, -0.0001089056, 0.002170148, 0.03413879, -0.0001831596, 0.02183766, 0, 
    -1.791112e-06, 1.113641e-12, 3.699457e-07, 0, -7.836836e-10, 
    0.0003556473, 0.006706373, 0.02238922, 0.01441167, 0.0001443252, 
    0.01474492, 0.0237844, 0.001587276, -0.0001227072, 0, 1.972666e-09, 
    0.0003310708, 0.01994836, 0.007981393, 0.002815368, 0,
  0, 0, 0, 0.0007339661, 0.006910917, 0.001953179, -8.640204e-05, 
    0.0002631967, -0.0001772201, 1.709458e-09, 0, 0, -7.955138e-05, 
    0.005438363, 0.07153481, 0.007273617, 0.004157882, 0.001817481, 
    0.008594804, -7.377294e-06, -2.589516e-07, 0, -3.857784e-06, 3.5391e-07, 
    -5.595936e-06, 0, -1.021874e-07, 0, 0,
  -2.365269e-06, 0.008181665, 0.001086311, 0.01155117, 0.001920363, 
    0.0617155, 0.05849062, 0.01985634, 0.03572615, 0.008319759, 0.0878821, 
    0.04094813, 0.02809045, 0.02796626, 0.09674023, 0.0678897, 0.000283957, 
    -4.265833e-09, 1.565543e-07, 0, -7.822975e-08, 0, 0, 0.02110818, 
    0.01046217, -2.351547e-06, -5.305473e-05, -7.204604e-05, 0,
  0.05316807, 0.02430665, 0.02248266, 0.0004908755, 0.00706775, 
    -5.797777e-06, 0, -5.252028e-05, 0.009249443, 0.04854469, 0.007096507, 
    -6.208576e-05, 0.05020528, 0.02968183, 0.02399783, 0.0007614003, 
    0.01057759, -0.0001920134, 0.003274313, -6.505081e-05, -5.134847e-05, 
    0.000273074, -5.320879e-06, 0.06389647, 0.04276419, 0.001072992, 
    0.03749079, 0.01837029, 0.04424541,
  0.001216216, -4.440796e-05, 0.0005424439, 0.0005059032, 0.0008592319, 0, 
    0.003544352, 0.0003892779, 0.0008216852, 0.0755078, 0.01308253, 
    0.05178412, 0.03690717, 0.09381501, 0.003034194, 0.02818525, 0.0116188, 
    0.00929178, 0.0006345097, 0.001545449, 0.00988194, 0.001860778, 
    0.001346628, 0.003055366, 0.005006394, 0.00819176, 0, -3.234512e-06, 
    0.009205833,
  0, 2.499222e-09, 0, -7.280634e-06, 0, -7.300382e-07, 0, -1.80957e-05, 
    0.0005526905, 3.173953e-06, 0.03718868, -0.0002393756, 0.0006954528, 
    3.970617e-10, 0, 0, 0, 0.01508037, 0.004020706, 0.0001867255, 
    -5.70028e-08, 0.0002829022, 3.649755e-08, 0.0004174918, 0, -0.0001049341, 
    -1.424629e-06, 0, 0,
  0, 0, 0.002809711, 0.001672066, 0.009842223, 0.000607847, 0, 0, 
    -0.000247355, 0.03243436, 0.01052169, 0.01297801, 0.01340229, 
    0.008759907, -0.0002259337, -0.0001021323, 0, 0.001689503, 0, 0.00049987, 
    0, 0.0009297416, -0.0001505778, 0.006525411, 0.001291612, 0.0001881294, 
    0.01156979, 0, 0,
  0, 0, 0, 0.001657908, 0.0008164713, -0.000355754, -4.749696e-06, 
    -6.112869e-06, 0, 0, 0, 0.00998715, 0.01137755, 0.002591424, 0.001188069, 
    0, -7.692752e-06, 0, 0, 0, 0, 0.0003874642, 0.004697956, 0.001392732, 
    0.0002777064, 8.530817e-05, 0, 0, 0,
  4.829667e-05, 0.0005673529, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2.054878e-07, 
    0, 0, 0, 0, 0, 0, 0, -6.565943e-07, -0.0001368888, 0.0001936881, 
    0.0001313262, 0.005879998, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -7.405687e-06, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0.000504401, -4.494144e-06, 0, 0, 0, 0, 0, 2.946901e-05, 0, 0, 0, 
    2.450956e-05, 0, 0, 0.001068521, 0, 0, 0, 0, 0, 0, 0, 0.0005241013, 
    -1.056037e-05, 0, 0, 0.0002218823, 0, 0,
  0.00896461, 0.0005544128, -1.353416e-05, -3.102846e-05, 0.006116876, 
    0.005395088, 0.009029546, 1.31635e-05, -2.900153e-05, 0, -1.4982e-06, 
    0.0007569898, 0, 0, -2.890509e-05, 0.008137245, 0.002408421, 0.002125217, 
    0.001312866, 0.001623137, 0.004475052, 0.01129177, -2.439055e-05, 
    -1.413126e-05, 0, 0.002049374, 0.0002716628, 0.001216451, 0.006577052,
  -6.785305e-05, 0.01113104, -4.061624e-05, 0.01937399, 0.02880709, 
    0.01240411, 0.01686432, 0.02495234, 0.0005474638, 4.796321e-05, 0, 
    0.01080353, 0, 0.0005099109, 0.01140061, 0.004065244, 0.03238818, 
    0.01139837, 0.006859142, 0.0152697, 0.02865592, 0.01837116, 0.03529184, 
    0.004315457, 0.004646607, 0.02324433, 0.007351408, 0.0283805, 0.00511194,
  0, -2.01124e-10, -0.0001472486, 0.006256898, 0.04757745, 0.005128006, 
    0.04575488, -7.356735e-05, 0.007637811, 0.003167843, 1.673546e-05, 
    -3.202983e-13, 7.520646e-05, 0.001129694, 0.01685162, 0.06070823, 
    0.05016324, 0.002061745, 0.03402235, 0.05100402, 0.01554456, 0.000864534, 
    -2.561754e-05, 0.002445187, 0.001839101, 0.03044284, 0.03918719, 
    0.008963953, 0,
  2.40416e-07, 2.573639e-07, -1.292302e-07, 0.03803949, 0.04012176, 
    0.01156686, 0.01013515, 0.005493165, 0.0004622239, 0.0004274354, 
    1.05845e-05, -7.537937e-06, -0.0003296828, 0.01152376, 0.1107256, 
    0.04002096, 0.06229652, 0.008569621, 0.0150968, 0.001504758, 
    3.093983e-05, -2.636496e-05, 0.0003125276, 0.0003982202, 0.005007178, 
    -5.147751e-08, 0.001911174, 0.0001036121, -1.334326e-08,
  0.001011789, 0.06824489, 0.008642633, 0.02851228, 0.02600357, 0.1612099, 
    0.1521917, 0.1155074, 0.1599273, 0.0861189, 0.139749, 0.2158626, 
    0.1091645, 0.1381934, 0.2057198, 0.2250432, 0.01351618, -2.497086e-05, 
    2.723731e-05, 0.0001991338, 7.936072e-06, 1.022395e-05, -3.505074e-05, 
    0.1373772, 0.05157817, -5.220815e-06, -0.0003458699, -0.000348963, 
    -3.572994e-05,
  0.2991182, 0.06301809, 0.1004698, 0.002200934, 0.05144094, 0.002346498, 
    2.865627e-06, 0.01852399, 0.04760653, 0.1381435, 0.1277449, 0.0308187, 
    0.2465031, 0.1119991, 0.1422703, 0.02797311, 0.07877807, 0.02346565, 
    0.0130195, 0.008276524, 0.004629199, 0.0008634896, 0.00145493, 0.2311821, 
    0.1608185, 0.01232483, 0.07501426, 0.05687558, 0.192779,
  0.0202057, 0.0004718538, 0.003538148, 0.001225299, 0.006341041, 
    7.318793e-05, 0.05001408, 0.001999622, 0.03949272, 0.09553009, 
    0.03012675, 0.11697, 0.1371301, 0.1671207, 0.03284737, 0.0641353, 
    0.03635518, 0.02311275, 0.004423831, 0.005396176, 0.02683633, 
    0.008782548, 0.007978025, 0.05789044, 0.02682489, 0.02332865, 0.00031873, 
    0.003591566, 0.05667882,
  -1.46569e-05, -6.398008e-05, -1.67794e-06, 0.004538621, -5.315573e-05, 
    0.001681611, 0.0002033853, -5.332021e-05, 0.003620659, 0.001531904, 
    0.03923855, 0.006178081, 0.01987912, 0.0004213536, -0.0001363811, 
    -0.0001551816, 1.033054e-05, 0.0342324, 0.02324943, 0.004328499, 
    0.004469668, 0.01336334, -2.06204e-05, 0.001534397, -9.567992e-06, 
    0.0003276509, -0.0002382681, 4.340587e-05, -4.623928e-06,
  -8.169286e-07, -4.779033e-05, 0.01273106, 0.004139863, 0.01696984, 
    0.003351108, -1.138512e-05, 0, 0.002964255, 0.04471789, 0.03583845, 
    0.02490882, 0.02386953, 0.02399231, 0.00244035, -0.0001293331, 
    -8.696942e-10, 0.00958133, 0, 0.002386072, 0.0001692979, 0.001295618, 
    8.778933e-05, 0.01139742, 0.006280018, 0.003695384, 0.01836212, 
    -4.075874e-05, -2.704354e-08,
  -3.242837e-05, 0, -1.376238e-05, 0.005270919, 0.006286095, 0.001786092, 
    -3.303966e-05, 0.0003332589, -2.855598e-06, 5.809221e-07, -1.167363e-05, 
    0.01361365, 0.01586903, 0.005624825, 0.01209395, -8.67401e-05, 
    -8.694665e-05, 0.0009218593, 4.738098e-06, -1.466124e-05, -1.065656e-05, 
    0.001157201, 0.01324783, 0.01018207, 0.002446618, 0.001896897, 
    5.186121e-05, 0, -1.324424e-06,
  0.008774659, 0.005015138, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2.3219e-05, 
    -6.316977e-05, 0.005044964, -6.890241e-11, 0, 0.0008804626, 0, 
    -3.69438e-06, -7.618759e-05, -1.873847e-08, -1.60032e-06, 0.003589638, 
    0.007910272, 0.007884699, 0.007934527, 0, 0, -8.355e-05,
  0.0006245762, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.0001813744, 0, 0.002624543, -6.042284e-05, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1.85715e-05, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, -3.627869e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0.001719716, 0.0004236297, -2.492111e-06, 0.00012753, 9.387113e-05, 
    -7.978234e-06, 0, 0.002098314, 0.001577525, 0, 0, 0.0001065564, 
    9.313166e-05, 0, 0.004719855, 0.002575801, -0.0001044207, -1.250728e-07, 
    0.0003552886, -2.242361e-05, 0, -1.148877e-05, 0.004331343, 0.0011048, 0, 
    0, 0.003032741, 0, -0.0001042359,
  0.02074496, 0.003254474, -0.0001193348, -5.296335e-05, 0.01987031, 
    0.02081593, 0.01574687, 0.005553368, 0.0038468, -1.964511e-05, 
    0.0009764109, 0.006335957, -1.988093e-06, 0.00449082, -9.422489e-05, 
    0.0110431, 0.01340961, 0.01278684, 0.003812225, 0.005265498, 0.01293311, 
    0.01937898, 0.0001254363, 0.007165156, -5.704856e-06, 0.007648535, 
    0.005149343, 0.003826285, 0.01987452,
  0.003050089, 0.01967924, 0.00199496, 0.03206787, 0.04378416, 0.04053603, 
    0.03141245, 0.04610103, 0.007163129, 0.01200897, 0.0009198699, 
    0.01783441, 0.001790427, 0.003109039, 0.03131367, 0.01152456, 0.05288342, 
    0.03895262, 0.02169613, 0.04964054, 0.04607668, 0.02687129, 0.05165787, 
    0.01531568, 0.0111693, 0.03785107, 0.01565362, 0.04758227, 0.01797865,
  2.976202e-05, 7.936978e-06, 0.0006498915, 0.009656497, 0.06352312, 
    0.02370105, 0.08158856, 0.02294386, 0.08296838, 0.02614061, 0.004086713, 
    0.009010417, 0.001061497, 0.004307762, 0.02403689, 0.0918386, 0.1294439, 
    0.05962888, 0.08035504, 0.09654655, 0.03656025, 0.0006003267, 
    0.002022231, 0.01697566, 0.01239539, 0.04892825, 0.06789168, 0.04114982, 
    0.005982073,
  4.206369e-07, 1.174385e-05, 0.006655701, 0.05377364, 0.08160265, 
    0.07141373, 0.05174294, 0.04164391, 0.0626605, 0.0687028, 0.01194302, 
    0.005993511, 0.002750216, 0.02070685, 0.1585015, 0.1651559, 0.1807143, 
    0.1171861, 0.09509544, 0.045087, 0.006090802, 0.02142427, 0.02727868, 
    0.03852866, 0.09200606, 0.008169126, 0.01392152, 0.01814851, 0.01053379,
  0.0001004195, 0.09263495, 0.1165295, 0.09726865, 0.03652372, 0.1969442, 
    0.1695325, 0.1206386, 0.1649957, 0.09615687, 0.1675934, 0.2277037, 
    0.08753914, 0.1021641, 0.1805339, 0.2285437, 0.09067725, 0.007412391, 
    0.004993804, 0.01998378, 0.0008603896, 9.650569e-06, 0.0098277, 
    0.3638569, 0.09108534, 0.006369027, 0.01536951, 0.003975058, 0.001588949,
  0.2835001, 0.2399744, 0.3685946, 0.03353384, 0.1282386, 0.01296944, 
    0.0005250932, 0.08135837, 0.1874584, 0.3460194, 0.09823646, 0.06111802, 
    0.2259191, 0.101498, 0.1146467, 0.0321523, 0.06393399, 0.01650501, 
    0.02361373, 0.01139232, 0.01287191, 0.006618246, 0.05028001, 0.3568667, 
    0.2549966, 0.04576068, 0.1055153, 0.1092929, 0.2159514,
  0.1094941, 0.01529379, 0.03399253, 0.002374887, 0.07817114, 0.004690565, 
    0.05809782, 0.008993426, 0.05079728, 0.1055871, 0.03370516, 0.1092411, 
    0.108123, 0.1571791, 0.06479858, 0.2363725, 0.1169955, 0.04514096, 
    0.0520312, 0.0611755, 0.07455485, 0.08486226, 0.05592026, 0.1606525, 
    0.1042077, 0.05233735, 0.006324608, 0.01024373, 0.295434,
  0.07418928, 0.04827154, 0.0004475804, 0.03251142, 0.0460759, 0.06977884, 
    0.02894149, 0.003396588, 0.01579294, 0.03319268, 0.07594857, 0.01132256, 
    0.06340131, 0.01355314, 0.0245376, 0.01262822, 0.00662748, 0.07301914, 
    0.1362691, 0.119628, 0.1199579, 0.05871488, 0.004890037, 0.04232278, 
    0.01997633, 0.1089971, 0.07110238, 0.05289512, 0.01102786,
  -0.000157258, 4.885659e-05, 0.01849276, 0.009739655, 0.03857717, 
    0.007068204, 0.0001126045, -2.483272e-05, 0.01570908, 0.08493996, 
    0.1256352, 0.07041358, 0.08212195, 0.0593584, 0.02519302, 0.001848849, 
    0.0002998454, 0.01848198, -0.0001632932, 0.005340901, 0.004949583, 
    0.002517242, 0.01026317, 0.01720828, 0.01817173, 0.01987331, 0.04476723, 
    0.02798715, 9.680786e-07,
  -8.762319e-05, 0.001046337, 0.0004826572, 0.010606, 0.01516362, 
    0.004034884, 0.0003322771, 0.0006869686, -1.552114e-05, 1.218025e-05, 
    -6.478207e-05, 0.01796983, 0.03254544, 0.01853133, 0.032253, 0.002850401, 
    0.001722498, 0.004843021, 0.002717461, -0.0001922476, -2.880131e-05, 
    0.00257198, 0.03218203, 0.03263935, 0.01681249, 0.008056053, 
    0.0004904818, -9.280921e-06, -3.392663e-06,
  0.01371108, 0.005915142, 0, 0, 0, 0, 0, 0, 0, 0, 0, -5.481541e-05, 
    -9.523079e-05, 0.007426496, 0.0002027959, -2.8602e-06, 0.004693905, 
    7.061888e-06, -2.595939e-05, -0.0001181257, 0.0009143057, -2.732617e-06, 
    0.009159112, 0.02576689, 0.02363854, 0.0123737, 2.066482e-09, 0, 
    0.006381097,
  0.002025428, 0, -5.121936e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.0003920632, 0.004381639, 0, 0.004666669, -0.0001183006, 0, 0, 0,
  0, -7.633042e-07, 0.0001394916, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.001381619, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, -5.243908e-05, 2.804558e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, -2.768275e-05, 0, 0, 0, 0, 0, 0, 0,
  0.007324206, 0.007459636, 0.0006285456, 0.002272924, 0.00334147, 
    -0.0001045634, 0, 0.002134401, 0.005684812, -0.0001126364, 0, 
    0.002336171, 0.002295388, 0, 0.005961976, 0.006965575, 0.001242308, 
    0.0006885449, 0.00325072, 0.002701975, 0.004496641, 0.0067015, 
    0.006936726, 0.004353053, 0, -7.583236e-05, 0.004766051, -9.927411e-05, 
    0.002355921,
  0.03178818, 0.01713583, 0.01188799, 0.001205356, 0.03581921, 0.03782704, 
    0.02510489, 0.01058664, 0.0194196, 0.003536004, 0.009851453, 0.01148489, 
    0.004394504, 0.01851405, 0.0176809, 0.02449756, 0.03359567, 0.05098374, 
    0.02057594, 0.04353046, 0.06272226, 0.0762938, 0.01294294, 0.01197126, 
    0.0003191511, 0.01745965, 0.01529336, 0.0110917, 0.04432958,
  0.03259528, 0.03654108, 0.01008701, 0.05286333, 0.08590945, 0.07825587, 
    0.05713717, 0.104939, 0.05744297, 0.05264597, 0.05012758, 0.08940992, 
    0.01938083, 0.01674147, 0.06090065, 0.03424526, 0.06909211, 0.08301276, 
    0.04264544, 0.1363433, 0.1265634, 0.06983947, 0.07567073, 0.02334861, 
    0.0353713, 0.05042663, 0.04014454, 0.1235651, 0.09093092,
  0.02776895, 0.009985065, 0.002208407, 0.06752288, 0.1191022, 0.04483494, 
    0.1389637, 0.0657906, 0.1498646, 0.1484307, 0.09493315, 0.04200402, 
    0.01566136, 0.020165, 0.03277637, 0.13749, 0.1332328, 0.09380779, 
    0.1470376, 0.1991854, 0.1301146, 0.04958544, 0.05334891, 0.06981612, 
    0.02772585, 0.09273873, 0.1756832, 0.1120795, 0.09591331,
  1.818586e-07, 0.0002374647, 0.002743512, 0.04767008, 0.07239056, 
    0.05001732, 0.04453577, 0.03273097, 0.09626973, 0.06479824, 0.01151206, 
    0.001153417, 0.01139489, 0.03454142, 0.1581745, 0.1380608, 0.1428861, 
    0.1004277, 0.07763826, 0.02502834, 0.004385532, 0.008875084, 0.00428826, 
    0.02936966, 0.06386311, 0.0259461, 0.0136666, 0.01416632, 0.003850047,
  8.326273e-06, 0.04812429, 0.09479146, 0.07794187, 0.02170414, 0.1433683, 
    0.1476416, 0.08325918, 0.119287, 0.06103558, 0.1577551, 0.1776386, 
    0.06946214, 0.0844936, 0.1650239, 0.1847006, 0.05139557, 0.002758204, 
    0.001688397, 0.01063828, 0.001086132, 3.022404e-06, 0.0003986188, 
    0.3167776, 0.05525741, 0.0001475525, 0.002931016, 0.000101925, 
    5.544402e-05,
  0.2291987, 0.2067606, 0.2778881, 0.02175191, 0.08901443, 0.007579349, 
    0.0002430683, 0.07069012, 0.140869, 0.2963663, 0.05528639, 0.03888178, 
    0.1819309, 0.08455697, 0.08530507, 0.01412918, 0.04008984, 0.01020329, 
    0.01456815, 0.01100171, 0.005958407, 0.001995313, 0.01544608, 0.3100827, 
    0.2191202, 0.03145559, 0.0949211, 0.08142093, 0.1513982,
  0.1214169, 0.009876684, 0.02470936, 0.03860088, 0.08623426, 0.001186468, 
    0.0418521, 0.005561118, 0.04027615, 0.09649146, 0.02443165, 0.08657344, 
    0.08765719, 0.1450048, 0.04297187, 0.1932079, 0.129951, 0.03607433, 
    0.03309292, 0.04625092, 0.0566787, 0.06309813, 0.02169003, 0.08101914, 
    0.08449619, 0.04301755, 0.003847915, 0.002208665, 0.2382303,
  0.091039, 0.1222361, 0.0143304, 0.05206025, 0.1348371, 0.08579034, 
    0.04260812, 0.01343909, 0.01070962, 0.02041536, 0.06657209, 0.009419953, 
    0.04573962, 0.003533858, 0.04043715, 0.02104981, 0.01388947, 0.09154126, 
    0.1642118, 0.117834, 0.08196545, 0.06926294, 0.01213229, 0.04984584, 
    0.01478478, 0.1261875, 0.0986641, 0.04913408, 0.05744314,
  0.07226073, 0.01294035, 0.04868202, 0.01810253, 0.05619031, 0.04067004, 
    0.04629013, -3.299189e-05, 0.03737769, 0.1114135, 0.156347, 0.1087271, 
    0.1260511, 0.1438028, 0.09665528, 0.04641368, 0.0231822, 0.02880031, 
    0.007422396, 0.02115549, 0.02497735, 0.07940903, 0.105981, 0.05899728, 
    0.05333924, 0.07676504, 0.08556158, 0.01421109, 0.03832415,
  0.0006397339, 0.005973626, 0.004613355, 0.01852861, 0.03421607, 0.05227431, 
    0.004291846, 0.001763214, 0.01748783, -7.146173e-05, 0.01186593, 
    0.03073069, 0.07106463, 0.07519946, 0.09195442, 0.1295688, 0.06263789, 
    0.0403701, 0.00655693, 0.000147996, -8.775486e-05, 0.009359371, 
    0.05376424, 0.05633878, 0.03546571, 0.02543612, 0.004128518, 
    0.0005564768, 0.0006131512,
  0.01848978, 0.006655731, -2.362099e-05, -0.0001125253, -1.43095e-05, 
    -3.569922e-05, 0, 0, 0, -1.909267e-05, -2.45833e-06, 0.001684093, 
    -0.0001860632, 0.01535152, 0.006478408, 0.001144127, 0.02763442, 
    0.01618596, 0.006948598, 0.0001245764, 0.003405484, 0.0001265169, 
    0.01340427, 0.04109509, 0.03606394, 0.03124357, -3.360639e-07, 0, 
    0.009395168,
  0.002150491, -0.000104382, -0.000163306, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 6.508102e-10, -3.245129e-05, -6.492697e-09, 0, -6.478943e-05, 
    0.005057988, 0.005462627, 0, 0.008179553, 3.674993e-05, 0, 0, 5.198526e-05,
  -8.73032e-05, -1.266373e-06, 0.000698957, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.003325772, -2.713197e-06, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  -4.179824e-06, 0.0001055372, -0.0001393975, 0.0004914865, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.001422856, 0, 0, 0, 0, 0, -3.752529e-05, 0, 0.0003266075, 
    -8.017907e-06, -1.378101e-05, -1.134971e-05, 0, 0, 0, 0,
  0.01264136, 0.01342613, 0.00803567, 0.004450716, 0.00884947, 0.005291946, 
    -4.547349e-06, 0.005950163, 0.01659412, 0.009592486, 0.001104554, 
    0.006273317, 0.01308254, 0.0007009372, 0.01119135, 0.01339345, 
    0.007180624, 0.01565879, 0.02553865, 0.02047142, 0.02532958, 0.02588641, 
    0.02545813, 0.01201613, 6.753958e-08, -7.763236e-05, 0.01096849, 
    0.002900204, 0.006061798,
  0.1034232, 0.0818456, 0.05768172, 0.05233718, 0.06308832, 0.08916205, 
    0.08901396, 0.07276807, 0.08995485, 0.06294569, 0.07021541, 0.04942197, 
    0.0561998, 0.08242198, 0.03658298, 0.05223727, 0.07912408, 0.1196178, 
    0.1316554, 0.1014873, 0.1531517, 0.2053016, 0.1418574, 0.0369986, 
    0.02593426, 0.06527942, 0.0534435, 0.03554199, 0.09672712,
  0.07928399, 0.08908115, 0.07528343, 0.1234696, 0.1401296, 0.1348007, 
    0.09394938, 0.1594958, 0.1167401, 0.1067202, 0.1582784, 0.1805315, 
    0.09680185, 0.0655249, 0.06688875, 0.08904403, 0.1580038, 0.1214524, 
    0.04730415, 0.1507222, 0.1423872, 0.1059801, 0.1192221, 0.07946684, 
    0.1674763, 0.1845712, 0.1025774, 0.2110706, 0.1874073,
  0.0175945, 0.01137903, 0.05634645, 0.03646101, 0.1101203, 0.06445696, 
    0.1345451, 0.07801422, 0.1616903, 0.1364408, 0.09497838, 0.04794733, 
    0.01681324, 0.02458534, 0.03853716, 0.1368201, 0.1081738, 0.07007724, 
    0.1272054, 0.1838284, 0.1136597, 0.04184606, 0.06085145, 0.05952464, 
    0.02422778, 0.0784706, 0.1654746, 0.09509567, 0.04337986,
  7.740432e-08, 0.0006680656, 0.0002661039, 0.05768767, 0.06720496, 
    0.04485235, 0.03123281, 0.02660167, 0.1245918, 0.04619635, 0.003264255, 
    0.0002055132, 0.0155438, 0.04346234, 0.1594661, 0.1226408, 0.1031702, 
    0.08761597, 0.05781164, 0.005028426, 3.283922e-05, 0.001209178, 
    -0.0001137937, 0.03283126, 0.05118684, 0.01949469, 0.008075486, 
    0.003965197, 0.0018448,
  2.136411e-06, 0.02820924, 0.07281467, 0.06455278, 0.01664428, 0.1138441, 
    0.1323146, 0.07163201, 0.1105008, 0.06042059, 0.1499487, 0.1341579, 
    0.05889723, 0.07262771, 0.164998, 0.1518529, 0.04492796, 0.004764285, 
    0.0003716572, 0.002937891, 0.007014609, 3.634765e-06, -8.873332e-05, 
    0.2786169, 0.04775139, 0.0002911832, -0.0003424091, 0.0001145639, 
    1.373183e-05,
  0.1907382, 0.1827853, 0.2120823, 0.01070352, 0.05714756, 0.009723875, 
    0.001359176, 0.05342241, 0.09995244, 0.2566678, 0.04701228, 0.03478696, 
    0.1550711, 0.08821654, 0.09382863, 0.01234098, 0.02115484, 0.01330701, 
    0.008559303, 0.01385162, 0.005036418, 0.002937893, 0.01222279, 0.2881849, 
    0.2041831, 0.02759022, 0.08017216, 0.06659023, 0.1067065,
  0.1140384, 0.005618643, 0.0192394, 0.0291394, 0.08048809, 0.001372965, 
    0.03653305, 0.004350438, 0.03058977, 0.09497509, 0.02408654, 0.07416447, 
    0.07737126, 0.1416496, 0.02492908, 0.1585294, 0.1231597, 0.04111248, 
    0.01857542, 0.03762944, 0.05040697, 0.0390108, 0.01125778, 0.05873874, 
    0.06385487, 0.03091456, 0.002063558, 0.001509365, 0.2039657,
  0.1146323, 0.1118117, 0.009617831, 0.0474317, 0.09954332, 0.07329303, 
    0.04768112, 0.009462855, 0.0120299, 0.02170336, 0.04298545, 0.008405658, 
    0.03561126, 0.005737253, 0.02886397, 0.005519716, 0.006882086, 
    0.08354117, 0.1003578, 0.09838706, 0.05698664, 0.0545052, 0.01747037, 
    0.04381368, 0.01173702, 0.09869649, 0.09080581, 0.04012273, 0.04588583,
  0.09687225, 0.06350286, 0.09770133, 0.07184373, 0.09435741, 0.07457323, 
    0.1023166, -0.0001106369, 0.06261776, 0.1304416, 0.1623939, 0.1142693, 
    0.1127508, 0.1408482, 0.1140778, 0.06912623, 0.06401389, 0.08024669, 
    0.03762919, 0.04571725, 0.07280361, 0.1253423, 0.1473465, 0.08148932, 
    0.04578273, 0.1086497, 0.1392968, 0.04413593, 0.08663696,
  0.01059688, 0.02948009, 0.05075033, 0.04185419, 0.09665449, 0.1375837, 
    0.008615499, 0.02477767, 0.04379665, 0.02470593, 0.04192962, 0.08413464, 
    0.1348719, 0.16409, 0.191749, 0.2176912, 0.1474917, 0.1031218, 
    0.03668735, 0.004746942, -4.750659e-05, 0.02338131, 0.1515613, 0.1560136, 
    0.1326758, 0.07907415, 0.1193648, 0.02798367, 0.03051395,
  0.03739175, 0.007570957, 0.006000089, -0.0002645401, 0.0070344, 
    0.001933902, -9.312526e-06, 0.0001193977, -4.823237e-07, -4.659391e-05, 
    2.953331e-05, 0.00257377, 0.009987588, 0.04762954, 0.06864351, 
    0.05220385, 0.09560518, 0.1226867, 0.08131982, 0.0008915557, 0.006910228, 
    0.01618376, 0.03682517, 0.07129085, 0.1306316, 0.1437792, 0.04720052, 
    0.001702658, 0.01994107,
  0.004831055, -0.0003490575, -0.0003216791, 0, 0.0009109629, 0, 0, 0, 0, 0, 
    0, 0, -8.878082e-06, -4.857796e-06, 0, 0, -7.940189e-07, 0.0007804846, 
    -5.049013e-05, 1.851586e-05, -0.0001285519, 0.007782228, 0.008086897, 
    0.00100896, 0.02451731, 0.009921918, 0.02240288, 8.819883e-05, 0.00463767,
  0.005635737, 0.0002515732, 0.0007848718, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, -5.083932e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0.005693488, -5.994624e-06, 0, 
    -8.129213e-06, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  -5.614308e-05, 0.006156448, 0.009396111, 0.003445134, -2.3101e-05, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.006232811, -0.0001112923, 0, 0, 0.001412444, 
    -0.0003044706, 0.01603663, 0.0002651878, 0.0006519195, 0.00170426, 
    0.0002106455, 0.002932733, 0, -3.246643e-07, 0, 4.915551e-05,
  0.05107898, 0.0805913, 0.06955564, 0.07755754, 0.05845676, 0.04486137, 
    0.02887248, 0.01110356, 0.03483314, 0.03628667, 0.04383483, 0.04500772, 
    0.06568928, 0.06837551, 0.09380043, 0.06369609, 0.0697612, 0.1090578, 
    0.1317776, 0.1071424, 0.09786823, 0.08196795, 0.1105544, 0.08453508, 
    0.03301128, 0.02068649, 0.02818632, 0.01566316, 0.03926874,
  0.1825992, 0.1434948, 0.1274021, 0.1404547, 0.1317614, 0.1691176, 
    0.1466234, 0.1789081, 0.1573003, 0.1302896, 0.1881115, 0.1561175, 
    0.1315717, 0.1178993, 0.08958257, 0.1308155, 0.1174154, 0.1782621, 
    0.1765341, 0.1300202, 0.2383736, 0.2251352, 0.1696547, 0.07736357, 
    0.08249146, 0.1455284, 0.1211811, 0.1131643, 0.1672001,
  0.07152206, 0.07994343, 0.1087531, 0.1206421, 0.1181775, 0.111724, 
    0.09259785, 0.1509728, 0.1188615, 0.1265394, 0.1451979, 0.1799606, 
    0.09806695, 0.05844259, 0.09321229, 0.1019181, 0.1648666, 0.1388018, 
    0.06297687, 0.1522333, 0.1152325, 0.09535769, 0.1270166, 0.07459208, 
    0.1617376, 0.1974261, 0.1247838, 0.2000803, 0.1695684,
  0.009228948, 0.01801256, 0.05243616, 0.01864506, 0.1087649, 0.07659471, 
    0.1134153, 0.07671526, 0.1495029, 0.1156126, 0.08410323, 0.03046268, 
    0.02277069, 0.01870508, 0.01912061, 0.1292712, 0.1075157, 0.07775501, 
    0.09586559, 0.1679489, 0.09377791, 0.0300356, 0.05454675, 0.04015873, 
    0.01927253, 0.06254682, 0.1381194, 0.07591609, 0.02118914,
  -2.012422e-09, 0.007838399, 0.0002496534, 0.04528962, 0.04706265, 
    0.04416229, 0.01991144, 0.02551198, 0.1150266, 0.02407506, 0.001201547, 
    5.125473e-05, 0.02463539, 0.04337257, 0.1688933, 0.1127102, 0.07712907, 
    0.07810969, 0.05044796, 0.0009168271, 3.102866e-06, 0.0001590327, 
    -0.0003388828, 0.02218307, 0.03339832, 0.01303796, 0.002760737, 
    9.826351e-05, 0.001042012,
  1.02295e-06, 0.03248569, 0.06435893, 0.05274682, 0.01102693, 0.08486374, 
    0.1086235, 0.05540821, 0.09773594, 0.04513916, 0.1493169, 0.1137335, 
    0.05491808, 0.05930272, 0.1513236, 0.1233441, 0.04037784, 0.005421798, 
    8.830904e-06, 0.0008868661, 4.959897e-05, 1.751668e-06, -3.126047e-06, 
    0.2039793, 0.04125998, 0.0002878684, -0.0002017892, 4.88703e-05, 
    2.961262e-06,
  0.1475705, 0.1663916, 0.1246291, 0.007640994, 0.04026484, 0.007018188, 
    0.004300165, 0.03037005, 0.06488521, 0.19303, 0.02916438, 0.02890128, 
    0.1195862, 0.07943866, 0.08378646, 0.01364984, 0.01022721, 0.0148864, 
    0.008405614, 0.006220451, 0.003285763, 0.002101029, 0.01736826, 
    0.2472125, 0.1814609, 0.03222292, 0.07810801, 0.04648542, 0.07679415,
  0.07153292, 0.004295032, 0.01663069, 0.01438243, 0.06297593, 0.001581691, 
    0.0241525, 0.004053062, 0.01978139, 0.09295499, 0.02175415, 0.06518136, 
    0.07860939, 0.1411578, 0.02097683, 0.1318227, 0.0969316, 0.04108574, 
    0.006649933, 0.02962631, 0.03603623, 0.02367055, 0.005856849, 0.06309594, 
    0.06282068, 0.02876059, 4.102407e-05, 0.000804477, 0.1624837,
  0.1279031, 0.09104253, 0.01665436, 0.05117794, 0.06561968, 0.05377612, 
    0.03116083, 0.002637417, 0.009292478, 0.02918431, 0.03000355, 0.00856759, 
    0.03241334, 0.01127357, 0.01268294, 0.002507623, 0.007167518, 0.05850583, 
    0.06369492, 0.08424416, 0.05203071, 0.04176009, 0.01400721, 0.039747, 
    0.002190246, 0.06346195, 0.07814774, 0.0548789, 0.04039903,
  0.09139159, 0.08869048, 0.1083266, 0.1356554, 0.1212844, 0.08445226, 
    0.08054414, 0.0007701885, 0.100796, 0.1230956, 0.1481641, 0.1403025, 
    0.1068293, 0.1258314, 0.1076824, 0.05181519, 0.05517889, 0.06369194, 
    0.04090594, 0.04857563, 0.07313234, 0.1004267, 0.1284594, 0.07468013, 
    0.03602479, 0.1260439, 0.1366131, 0.03992221, 0.0910389,
  0.0743368, 0.09326429, 0.1208522, 0.09152249, 0.1746226, 0.1608463, 
    0.02374225, 0.106364, 0.0941004, 0.06310103, 0.05698168, 0.103538, 
    0.1616872, 0.1801126, 0.2055607, 0.2372179, 0.1495102, 0.1387988, 
    0.06601261, 0.0437049, 0.009166561, 0.03252453, 0.133284, 0.1458366, 
    0.1521864, 0.1104522, 0.1484774, 0.05898366, 0.06852347,
  0.144207, 0.01985681, 0.07992438, 0.02117134, 0.2011176, 0.02031871, 
    9.525865e-05, -1.854093e-06, -9.773878e-06, 0.0001293067, 0.00761758, 
    0.009755235, 0.05632309, 0.08438339, 0.1038973, 0.06286988, 0.1182247, 
    0.2501203, 0.2123432, 0.02985667, 0.06742132, 0.1047799, 0.09990517, 
    0.1227192, 0.172943, 0.1900679, 0.08356243, 0.02701928, 0.06116819,
  0.01677794, 0.001910079, 0.04405684, 0.03776489, 0.00949946, 2.255913e-05, 
    0, -9.01308e-06, 0, 0, 0, 0, -0.0001093944, 0.001226331, 0.00277872, 
    0.007174597, 0.003615522, 0.02501533, 5.804877e-05, 0.004926946, 
    0.006277621, 0.02426677, 0.0263242, 0.02314757, 0.1134567, 0.07234654, 
    0.04160067, 0.005426034, 0.01648089,
  0.008030042, 0.0009461922, 0.001814733, -4.713836e-08, 0, -3.243926e-06, 0, 
    0, 0, 0, 0, 0, 0, 0.006910919, 0.002711352, 0.001021756, 9.936821e-06, 
    4.746675e-05, -1.664288e-08, 3.565986e-05, 0, 0, -1.902443e-08, 
    -0.003069693, 0.06108709, -0.0001452704, -1.650453e-08, 0.001072535, 
    0.0001531207,
  -2.407608e-05, 0, 0, 0.000561723, 0.003190051, 0, 0, 0, 0, -1.454637e-07, 
    9.782382e-09, 2.321069e-09, 0, 0, 0, 0, -3.297771e-06, 0.0005868859, 
    -2.412304e-05, 0, -3.177709e-05, 0.000964721, -6.12572e-05, 
    -0.0003152189, -0.0002545643, 0, 0, -8.798275e-05, 3.10766e-07,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0.001120835, 0.01415301, 0.0138426, 0.01172546, -0.0004055325, 0, 
    1.260819e-06, 0.0002196484, 0, -1.483687e-05, 0, -7.775296e-06, 
    0.0003325238, 0.01122479, 0.00517018, 0.01362498, 0.01928833, 0.01807209, 
    0.03080921, 0.05957486, 0.03612249, 0.07755239, 0.05463078, 0.01320715, 
    0.0196242, 0.003033089, 0.0006127497, 0.009103234, 0.006029642,
  0.08256079, 0.123414, 0.1248598, 0.1243284, 0.1323984, 0.1151649, 
    0.09692306, 0.0869955, 0.1008624, 0.08350546, 0.07231648, 0.1519632, 
    0.186127, 0.1711124, 0.1882253, 0.1669765, 0.1561189, 0.1852494, 
    0.221739, 0.1243081, 0.138258, 0.1465825, 0.1745204, 0.1963698, 
    0.08103527, 0.07810465, 0.09443704, 0.06443729, 0.07071201,
  0.2055492, 0.1613826, 0.1278244, 0.1531865, 0.1278996, 0.1822909, 0.152984, 
    0.1747849, 0.1869864, 0.1896468, 0.2159566, 0.1808927, 0.1246149, 
    0.126192, 0.1049553, 0.1186202, 0.1230994, 0.1766682, 0.1769563, 
    0.1233658, 0.2389286, 0.210398, 0.1646586, 0.1002005, 0.1173686, 
    0.1631032, 0.1427398, 0.1142739, 0.1794809,
  0.06104015, 0.06547532, 0.08911201, 0.09102186, 0.09603614, 0.104801, 
    0.09511077, 0.1293967, 0.1030521, 0.1104845, 0.1141501, 0.1545479, 
    0.07975736, 0.04866463, 0.09396012, 0.09638152, 0.1484003, 0.1164024, 
    0.07613874, 0.1499062, 0.1055709, 0.0818067, 0.1484041, 0.06972704, 
    0.1230583, 0.1584749, 0.08729391, 0.1753552, 0.1657219,
  0.001128101, 0.009357265, 0.03176513, 0.01173923, 0.1027968, 0.1115176, 
    0.1091546, 0.09197693, 0.1240119, 0.06869219, 0.06590997, 0.01968537, 
    0.01050208, 0.01719944, 0.004310766, 0.1200666, 0.1209295, 0.05508426, 
    0.09747321, 0.1557494, 0.09570093, 0.02856154, 0.02813868, 0.01241043, 
    0.01221467, 0.05471168, 0.1114813, 0.07391512, 0.00848535,
  2.00226e-07, 0.00136094, 0.0003945403, 0.024122, 0.03960688, 0.04444914, 
    0.01487375, 0.02556885, 0.08424527, 0.00589129, 0.0005908022, 
    4.00676e-05, 0.03221907, 0.04184021, 0.1563261, 0.09752315, 0.0476489, 
    0.05356731, 0.04408881, 0.0009239116, 1.312609e-06, 0.001841814, 
    -2.64421e-05, 0.02224887, 0.02221613, 0.002006973, 0.001628547, 
    1.114712e-05, 1.720209e-05,
  3.599753e-07, 0.05083441, 0.05500944, 0.04431483, 0.008816586, 0.05936936, 
    0.08225826, 0.04453624, 0.08777599, 0.03554113, 0.1568708, 0.1097529, 
    0.04874486, 0.04333825, 0.1336424, 0.09771965, 0.0263649, 0.004833188, 
    3.592171e-05, 0.000155491, -9.208824e-06, 4.342144e-07, 9.208037e-05, 
    0.1274693, 0.03843605, 0.0003762303, 5.488558e-06, 8.5771e-06, 
    1.354766e-06,
  0.1021786, 0.1337023, 0.08061551, 0.008212561, 0.03158435, 0.005108132, 
    0.008101196, 0.01380922, 0.04140306, 0.1449332, 0.02263587, 0.01724024, 
    0.08651756, 0.06278536, 0.07331812, 0.00998046, 0.007172502, 0.02036014, 
    0.009878651, 0.001501613, 0.00176023, 0.002198457, 0.02357062, 0.2181719, 
    0.1740524, 0.05829396, 0.08920727, 0.03682103, 0.05446503,
  0.04730333, 0.002409216, 0.01323316, 0.01250906, 0.05155092, 0.001642531, 
    0.01302545, 0.002411408, 0.01173506, 0.0863986, 0.01951164, 0.05854158, 
    0.06973716, 0.1239807, 0.02981501, 0.1055527, 0.08727443, 0.04440101, 
    0.003348738, 0.01762679, 0.02302392, 0.01149782, 0.004263484, 0.05379948, 
    0.06319924, 0.03415536, -1.209658e-05, 0.006149249, 0.1246106,
  0.1543853, 0.06336799, 0.01531853, 0.05358284, 0.04542554, 0.04063035, 
    0.01107686, 0.001102805, 0.005347623, 0.02592348, 0.02847841, 
    0.006539878, 0.02055936, 0.005710225, 0.004052818, 0.002379678, 
    0.008768751, 0.03773636, 0.06856314, 0.07533504, 0.03361133, 0.02847069, 
    0.008357523, 0.03767849, 0.001821172, 0.04585389, 0.06874869, 0.04787751, 
    0.04367317,
  0.0647961, 0.08889006, 0.09708988, 0.1227844, 0.1360984, 0.08170533, 
    0.06532343, 0.00228575, 0.1382, 0.1229889, 0.1427035, 0.1822373, 
    0.1283206, 0.1059877, 0.09220605, 0.04587105, 0.04292039, 0.04570346, 
    0.04128942, 0.03356326, 0.07547237, 0.08603441, 0.1043763, 0.07759699, 
    0.03392378, 0.1129252, 0.1483952, 0.03470397, 0.06493039,
  0.1006422, 0.1162251, 0.1263998, 0.1265592, 0.1713461, 0.1354164, 
    0.05032754, 0.1370988, 0.1303584, 0.09657411, 0.05222629, 0.1269477, 
    0.1522171, 0.1611138, 0.201891, 0.2546, 0.1561416, 0.1063241, 0.06450582, 
    0.09467965, 0.05571976, 0.03607986, 0.1159141, 0.1463125, 0.1465014, 
    0.09978963, 0.1552243, 0.0481572, 0.06425802,
  0.2373, 0.07572108, 0.1777593, 0.1053115, 0.2387879, 0.1109204, 0.0259704, 
    0.003116411, 0.0008328678, 0.008135786, 0.02392633, 0.01682485, 
    0.1151309, 0.09633289, 0.1296811, 0.06758436, 0.1218046, 0.2950459, 
    0.219738, 0.1682656, 0.1081331, 0.1496549, 0.149565, 0.12716, 0.2329997, 
    0.1946236, 0.09633191, 0.04068384, 0.1307462,
  0.1717832, 0.06017806, 0.1047237, 0.08352526, 0.1233549, 0.03101553, 
    0.02026385, 0.0002338341, 0.0005822468, 0, 0, 0, 0.0002460495, 
    0.05074258, 0.03294237, 0.0349919, 0.04197147, 0.06193686, 0.03181138, 
    0.05726078, 0.07584892, 0.09928209, 0.1304644, 0.04392903, 0.2225539, 
    0.08790111, 0.05516829, 0.02739932, 0.1232383,
  0.1556771, 0.07297411, 0.04970646, 0.03644826, 0.01975947, 0.01486258, 
    0.008063923, 7.154106e-05, -0.0002095989, 0, 0, 6.784497e-05, 
    0.0007182342, 0.04471959, 0.07041357, 0.02950645, 0.002600071, 
    0.01043468, -0.000344087, 0.0007479971, 0, -9.524189e-06, -0.0001717074, 
    0.0233, 0.1394941, 0.002890829, -2.967339e-06, 0.0177294, 0.06240155,
  0.02838635, 0.03069795, 0.03656008, 0.02694442, 0.01567135, 0.01448704, 
    0.0117675, 0.01159486, 0.000156126, 0.01720537, 0.04533059, 0.01967843, 
    0.01487334, 0.002340906, 0.008979877, 0.01069044, 0.01626655, 0.01599725, 
    0.01437249, 0.01549055, 0.01594925, 0.01730853, 0.009140717, 0.006852266, 
    0.01129357, 0.0004633841, -0.002197736, 0.01142613, 0.0140345,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -4.88426e-06, 0, 0, 
    0, 0.0005415035, 0.01545553, 0.009226584, -0.0001881763, 0, 0, 0,
  0.09931701, 0.07465268, 0.04812003, 0.0279037, 0.001233795, -0.0001187167, 
    0.004368075, -3.160882e-05, -5.783755e-05, -0.0005115357, -3.55869e-06, 
    -0.000204233, 0.004307369, 0.06779032, 0.09088241, 0.127015, 0.09064893, 
    0.1127516, 0.1561528, 0.1286318, 0.1259168, 0.1758373, 0.1358983, 
    0.1254769, 0.1026207, 0.04337125, 0.04074739, 0.05093401, 0.06270502,
  0.1547572, 0.1256939, 0.1518, 0.1998855, 0.1949332, 0.1525642, 0.112411, 
    0.1814415, 0.1812413, 0.1443555, 0.1009417, 0.2060532, 0.2486013, 
    0.2244551, 0.2224649, 0.2016592, 0.1624594, 0.2030956, 0.2459007, 
    0.16325, 0.1628541, 0.1925629, 0.2556156, 0.224695, 0.1668576, 0.1452926, 
    0.155983, 0.1197711, 0.1262978,
  0.2232855, 0.2028952, 0.1417469, 0.1392335, 0.1290042, 0.1758274, 
    0.1424821, 0.1633961, 0.199466, 0.1930982, 0.2006598, 0.1792229, 
    0.1240501, 0.1336507, 0.09931345, 0.09912273, 0.1023968, 0.1823505, 
    0.1429847, 0.1294702, 0.2401219, 0.2068955, 0.1625415, 0.104319, 
    0.1265392, 0.1489373, 0.1292214, 0.1243983, 0.1863751,
  0.0502944, 0.06347876, 0.0460966, 0.07562222, 0.08386534, 0.1012676, 
    0.1102193, 0.1068303, 0.0951925, 0.08793429, 0.1104685, 0.161841, 
    0.06579404, 0.04697631, 0.09035657, 0.08994909, 0.1229314, 0.1007421, 
    0.0874222, 0.1380249, 0.1051217, 0.07701454, 0.163075, 0.07396836, 
    0.1071936, 0.1073813, 0.07898781, 0.160261, 0.1735215,
  2.097539e-05, 0.01306128, 0.01759072, 0.01117912, 0.09721406, 0.1180584, 
    0.08447253, 0.1006142, 0.07332712, 0.04762242, 0.0583467, 0.02307624, 
    0.003140352, 0.01417974, 0.002103258, 0.1100794, 0.1045331, 0.04760987, 
    0.08325824, 0.1385225, 0.09000086, 0.02028347, 0.02370379, 0.002624288, 
    0.01396225, 0.05111462, 0.09611063, 0.05450326, 0.003679215,
  7.92599e-07, 0.0003824135, 0.001203324, 0.01547542, 0.04089098, 0.04765286, 
    0.01132884, 0.01617998, 0.04776045, 0.002085541, 0.0005334026, 
    7.124509e-05, 0.06496824, 0.04473119, 0.1427587, 0.08669554, 0.02319716, 
    0.03805747, 0.04276881, 0.001230014, 2.011453e-05, 0.0007405372, 
    8.689596e-07, 0.004049693, 0.01347728, 0.0002985813, 0.0009252461, 
    3.256755e-06, 2.149168e-06,
  9.181565e-09, 0.05584344, 0.04145299, 0.0419629, 0.007525207, 0.05122887, 
    0.06882023, 0.04310513, 0.08550297, 0.02399149, 0.1488715, 0.09356535, 
    0.05283743, 0.03853117, 0.1264284, 0.08971722, 0.02115752, 0.004767832, 
    2.596106e-05, 6.418262e-05, 3.274574e-06, 1.623124e-07, 0.003564853, 
    0.08293546, 0.0374437, 0.0004232091, 0.0004002115, -4.064978e-06, 
    1.171917e-06,
  0.09394617, 0.1189968, 0.05461603, 0.008300295, 0.02948148, 0.00365962, 
    0.004141211, 0.007934275, 0.02522609, 0.118422, 0.01688088, 0.01241445, 
    0.06434221, 0.05252418, 0.0589065, 0.007859393, 0.006357267, 0.02172667, 
    0.0189393, 0.0004985183, 0.001750052, 0.001524731, 0.04525347, 0.2013416, 
    0.1833382, 0.085033, 0.09917971, 0.03545075, 0.04653433,
  0.03383209, 0.003134173, 0.008674284, 0.009756085, 0.03223217, 0.001143994, 
    0.007613987, 0.000960372, 0.007768382, 0.08060177, 0.01986622, 
    0.06279773, 0.0645621, 0.1242968, 0.02071833, 0.08000959, 0.07701884, 
    0.04484169, 0.009110729, 0.01768132, 0.01504119, 0.005450311, 
    0.003765565, 0.0483194, 0.05767903, 0.036978, -1.71121e-06, 0.002814531, 
    0.09874777,
  0.1624935, 0.03737767, 0.01072046, 0.04541799, 0.02873497, 0.0273346, 
    0.001071449, 0.0005402902, 0.002653714, 0.01871975, 0.02724234, 
    0.004788645, 0.01782403, 0.006388654, 0.001521646, 0.002530796, 
    0.005171007, 0.02894107, 0.06865117, 0.05854765, 0.02364271, 0.02717124, 
    0.006302871, 0.04425605, 0.001159273, 0.03814543, 0.03624166, 0.02445412, 
    0.05372313,
  0.0573167, 0.08237997, 0.09361902, 0.1154131, 0.127541, 0.07281696, 
    0.05193962, 0.007454594, 0.1767322, 0.1298372, 0.1349977, 0.1690543, 
    0.1211505, 0.0731141, 0.08434435, 0.04114466, 0.03775087, 0.04738786, 
    0.02914722, 0.02587559, 0.06518145, 0.08733296, 0.07481591, 0.06652797, 
    0.03284062, 0.1184097, 0.1442068, 0.02957312, 0.04316325,
  0.09657709, 0.1159496, 0.1047139, 0.1437495, 0.1551983, 0.105814, 
    0.1361903, 0.1325467, 0.1146183, 0.08613303, 0.0547957, 0.123034, 
    0.1538419, 0.154199, 0.1906684, 0.2508409, 0.1574111, 0.07071009, 
    0.05660041, 0.09891576, 0.09261558, 0.03404161, 0.1030322, 0.1479398, 
    0.1332471, 0.09085206, 0.1610782, 0.03722301, 0.09631648,
  0.2379351, 0.1236494, 0.1780449, 0.1007937, 0.2349599, 0.1338716, 
    0.0874896, 0.01554501, 0.002960555, 0.0410089, 0.0529437, 0.09290221, 
    0.1379172, 0.1227805, 0.1609677, 0.09666497, 0.1802722, 0.2944234, 
    0.2143598, 0.1665221, 0.1114543, 0.1517188, 0.154446, 0.1249932, 
    0.2196985, 0.196744, 0.1088727, 0.04246137, 0.2132183,
  0.1966289, 0.1481387, 0.1224376, 0.1292212, 0.1252006, 0.0591673, 
    0.0659767, 0.04244369, 0.01893053, 0.002220899, 0.009564155, 
    -0.0002314769, 0.05318067, 0.1152813, 0.1191092, 0.1098146, 0.06978555, 
    0.1182407, 0.1042028, 0.1090954, 0.1269187, 0.144004, 0.1477769, 
    0.09471562, 0.2291489, 0.1013399, 0.05172168, 0.05621361, 0.1478015,
  0.1986922, 0.1359626, 0.1672083, 0.07228442, 0.1160659, 0.1092856, 
    0.04021576, 0.07419989, 0.02349283, 0.01166951, 0.01977198, 0.006141289, 
    0.06588156, 0.1102879, 0.08695395, 0.02535068, 0.0236287, 0.03183879, 
    0.02361254, 0.0120832, 0.001720803, 0.02541645, 0.005500013, 0.06356924, 
    0.194341, 0.03113136, -0.0001590926, 0.08961586, 0.1679375,
  0.1245905, 0.1185549, 0.1111978, 0.1023994, 0.09354677, 0.07178391, 
    0.04743868, 0.02733061, 0.02548821, 0.06779277, 0.09283412, 0.07821863, 
    0.06711199, 0.03978134, 0.03474339, 0.02683723, 0.03166469, 0.04066891, 
    0.04123987, 0.02392986, 0.02505466, 0.03477492, 0.03221816, 0.0230463, 
    0.04842671, 0.009705484, -0.006411176, 0.03200668, 0.08698686,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3.607196e-05, -0.000344528, 
    -0.0007423398, 0.01715222, 0.0197858, 0.002765066, -1.002459e-05, 0, 0, 
    0.005153663, 0.09494326, 0.04803894, 0.004862437, -0.001498703, 
    -2.518405e-05, 0,
  0.2433451, 0.1333924, 0.1447838, 0.07925199, 0.006651169, -0.001997265, 
    0.02906408, 0.00156921, 0.0006242954, 0.0009423997, -0.0003097588, 
    -0.0004254105, 0.01984185, 0.1553582, 0.2070917, 0.2276878, 0.1853454, 
    0.1898, 0.2374756, 0.2131804, 0.2271426, 0.2968397, 0.3307949, 0.1865853, 
    0.1743948, 0.07335581, 0.1148791, 0.1334677, 0.1282818,
  0.2056706, 0.1872952, 0.2256068, 0.2522543, 0.2671466, 0.2144614, 
    0.1798531, 0.2226476, 0.2488376, 0.1864856, 0.1409998, 0.2809294, 
    0.2823904, 0.2487904, 0.2410091, 0.1905701, 0.1589237, 0.1930684, 
    0.2431097, 0.1920735, 0.1846104, 0.2164541, 0.2871086, 0.2473386, 
    0.2384008, 0.2000383, 0.2067244, 0.2074405, 0.2406614,
  0.2109828, 0.2121153, 0.1487069, 0.1378302, 0.1322429, 0.163027, 0.1377046, 
    0.1523164, 0.1978798, 0.2070845, 0.1883513, 0.1673038, 0.1100079, 
    0.1406869, 0.09380756, 0.0813485, 0.07450677, 0.1940084, 0.1549141, 
    0.127113, 0.2193072, 0.1950569, 0.1230418, 0.1016911, 0.1224812, 
    0.1833909, 0.1522897, 0.1291207, 0.1726484,
  0.05241495, 0.07107794, 0.04140608, 0.07606109, 0.08632483, 0.09192143, 
    0.1217034, 0.1048585, 0.07506881, 0.07606584, 0.09091575, 0.1462544, 
    0.06553832, 0.04154451, 0.0866383, 0.1029142, 0.1164267, 0.09093788, 
    0.07920098, 0.1134752, 0.09799345, 0.0731907, 0.1491525, 0.08681439, 
    0.08525138, 0.07655796, 0.06602415, 0.1616393, 0.190172,
  9.910755e-06, 0.01457418, 0.01128551, 0.009127543, 0.0910948, 0.1114639, 
    0.06672736, 0.07950883, 0.02137448, 0.04220554, 0.05895758, 0.02294933, 
    0.002389909, 0.01083195, 0.00227567, 0.1113664, 0.111227, 0.05253169, 
    0.08645351, 0.1244816, 0.08763129, 0.0181, 0.007446696, 0.0003702978, 
    0.01360884, 0.04501655, 0.07912462, 0.04805427, 0.004954003,
  1.032443e-07, 0.0002822, 0.0006641077, 0.01208647, 0.0346817, 0.04782112, 
    0.01233237, 0.01742623, 0.02437335, 0.0003935327, 0.0007724682, 
    -2.260502e-05, 0.08496624, 0.04154544, 0.1210547, 0.07864261, 0.01391599, 
    0.03086455, 0.04880174, 0.001206403, 3.693384e-05, 1.265963e-05, 
    4.229306e-07, 0.0009315126, 0.008002133, 0.0003711728, 0.001784286, 
    1.058485e-06, 5.898449e-07,
  6.333353e-06, 0.06437685, 0.02492362, 0.03477748, 0.006614455, 0.05019683, 
    0.0653854, 0.04186366, 0.08115372, 0.0173634, 0.1549115, 0.07930099, 
    0.0538746, 0.04321755, 0.1184322, 0.0774713, 0.01830548, 0.003266528, 
    -4.64971e-06, 5.067206e-05, -1.391648e-06, 1.821249e-07, 0.0004256558, 
    0.05888132, 0.0368316, 0.0005603314, 0.0001377638, 1.164178e-06, 
    8.536831e-06,
  0.09007268, 0.1096167, 0.04278997, 0.00944306, 0.02764906, 0.004480235, 
    0.004238282, 0.006657038, 0.01363445, 0.1129684, 0.01339479, 0.009101129, 
    0.05377734, 0.0407557, 0.05467496, 0.00746497, 0.006249189, 0.01268777, 
    0.02558072, 0.0006089823, 0.001497403, 0.001545322, 0.07770316, 
    0.2147304, 0.1997041, 0.1074355, 0.1161267, 0.0407104, 0.03246583,
  0.03320389, 0.007790772, 0.007304857, 0.009583236, 0.01847309, 0.001095343, 
    0.006206112, 0.0008767336, 0.005103284, 0.07697492, 0.01649488, 
    0.06417727, 0.06523857, 0.1306316, 0.02807344, 0.05433304, 0.07689273, 
    0.0454669, 0.004464378, 0.01654298, 0.01173197, 0.003794555, 0.003748337, 
    0.04531898, 0.05027347, 0.03916418, -9.706786e-07, 3.379976e-05, 
    0.07526013,
  0.1639272, 0.02039436, 0.009084065, 0.03743058, 0.01845956, 0.0123688, 
    0.0001522688, 0.0001893168, 0.001898916, 0.01495756, 0.02885555, 
    0.005757876, 0.009638028, 0.007327782, 0.0009731416, 0.002003223, 
    0.001390638, 0.02053967, 0.06050822, 0.05458099, 0.01359838, 0.02574489, 
    0.003362828, 0.04919849, 0.001611618, 0.03100502, 0.02517625, 
    0.006465256, 0.03516735,
  0.051374, 0.08395775, 0.08946168, 0.09743892, 0.1103444, 0.06166628, 
    0.04415999, 0.02701038, 0.1972493, 0.1306832, 0.1414565, 0.156398, 
    0.1125236, 0.103207, 0.0821896, 0.02791185, 0.02600459, 0.0572702, 
    0.02013275, 0.01490978, 0.04479432, 0.07721019, 0.06033285, 0.05286011, 
    0.0268342, 0.1263088, 0.1049032, 0.0209941, 0.0295689,
  0.08294316, 0.1234274, 0.09956253, 0.1284966, 0.1317245, 0.07760356, 
    0.1508321, 0.1201684, 0.1080929, 0.06828779, 0.0533192, 0.1153676, 
    0.1566226, 0.147099, 0.1803015, 0.237004, 0.1576722, 0.06436105, 
    0.05225996, 0.09258334, 0.109698, 0.03464149, 0.1031512, 0.1738886, 
    0.114641, 0.09243894, 0.1514918, 0.04671952, 0.09857289,
  0.2007842, 0.1260348, 0.1735419, 0.09945887, 0.2238188, 0.1235785, 
    0.123424, 0.04734625, 0.03348396, 0.1343687, 0.1277566, 0.1432831, 
    0.2007053, 0.1555285, 0.1762985, 0.1475866, 0.209141, 0.2659257, 
    0.2068752, 0.1645009, 0.1047451, 0.1704151, 0.1647565, 0.1231806, 
    0.2301906, 0.2026339, 0.1086642, 0.05677986, 0.1778138,
  0.2088162, 0.1582081, 0.1594778, 0.2782302, 0.1835668, 0.06300586, 
    0.08253805, 0.07653335, 0.09115144, 0.03783181, 0.02764133, 0.03031223, 
    0.1705856, 0.2119393, 0.1730209, 0.1819771, 0.1345627, 0.1779365, 
    0.1548104, 0.1246463, 0.1651653, 0.2121198, 0.1602694, 0.1025684, 
    0.2166932, 0.1019029, 0.04547817, 0.07927673, 0.1833745,
  0.2576067, 0.1429515, 0.1997999, 0.160046, 0.1445468, 0.1104637, 
    0.04807972, 0.07590544, 0.05766023, 0.1014986, 0.1009943, 0.1240991, 
    0.1905716, 0.1738232, 0.1017276, 0.04302813, 0.0741563, 0.08039703, 
    0.078711, 0.06673241, 0.06550489, 0.07941164, 0.1001258, 0.1277678, 
    0.239055, 0.06202245, 0.004283862, 0.1571974, 0.2242241,
  0.1934884, 0.1582353, 0.1474522, 0.1774444, 0.1278755, 0.1117956, 
    0.1062426, 0.1135014, 0.06889636, 0.09391455, 0.08278146, 0.08833813, 
    0.09704391, 0.09320403, 0.06382446, 0.05107627, 0.04788378, 0.06555798, 
    0.06440824, 0.05034455, 0.04584889, 0.05642791, 0.0428621, 0.02399247, 
    0.06671381, 0.04238396, 0.02676105, 0.07334618, 0.1550607,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -6.20707e-06, 0.0017273, 0.0004732446, 
    0.04042052, 0.110558, 0.08972975, 0.02892072, 0.001870448, -0.002085367, 
    -0.001804236, 0.03723474, 0.2088697, 0.2091251, 0.0624221, 0.04153741, 
    -0.002127246, 0,
  0.3248349, 0.2288678, 0.2321513, 0.1667556, 0.01866001, 0.006710894, 
    0.07206269, 0.01150471, 0.009171933, 0.006199659, -0.0003700452, 
    0.001440266, 0.0384748, 0.19423, 0.298577, 0.3229113, 0.3044484, 
    0.3090466, 0.3619151, 0.333151, 0.2877263, 0.388528, 0.4072181, 
    0.3113367, 0.2603992, 0.1210533, 0.1710392, 0.1812009, 0.371453,
  0.2559932, 0.2488075, 0.2648483, 0.2672496, 0.2836701, 0.2816763, 
    0.2203031, 0.3169889, 0.3233402, 0.2414045, 0.2030092, 0.3250911, 
    0.3075923, 0.2569427, 0.2500349, 0.2234633, 0.150898, 0.1865714, 
    0.2587133, 0.2279372, 0.2014912, 0.216708, 0.2663219, 0.2580243, 
    0.2290948, 0.2101137, 0.2571262, 0.2625442, 0.3036952,
  0.2105801, 0.2162999, 0.1526772, 0.147812, 0.1393964, 0.1567532, 0.154549, 
    0.1506771, 0.2113194, 0.2327906, 0.1780139, 0.1648868, 0.1255956, 
    0.1361036, 0.09949271, 0.07913709, 0.05465158, 0.1826855, 0.1369019, 
    0.1213349, 0.2171636, 0.2223722, 0.124069, 0.09641883, 0.117034, 
    0.1919448, 0.1501288, 0.1353344, 0.1803533,
  0.07747962, 0.06156416, 0.03654202, 0.07351884, 0.09823459, 0.07093942, 
    0.1222761, 0.09891169, 0.07565682, 0.07410213, 0.08434669, 0.1138105, 
    0.0587646, 0.03933604, 0.08122034, 0.1141903, 0.1028733, 0.07822879, 
    0.07748347, 0.1052154, 0.1056064, 0.07079233, 0.1531131, 0.08931106, 
    0.07300679, 0.06540515, 0.06187705, 0.1553093, 0.1736324,
  2.713073e-06, 0.01793527, 0.0132702, 0.01085925, 0.08813071, 0.09979081, 
    0.05317501, 0.0573319, 0.005474774, 0.0355936, 0.05756887, 0.02198482, 
    0.00317972, 0.01285499, 0.00223194, 0.1007724, 0.1206406, 0.07021242, 
    0.07353562, 0.1059985, 0.1024816, 0.01785104, 0.004963455, 0.0005910004, 
    0.02030174, 0.042246, 0.08272125, 0.05811636, 0.01334185,
  2.099968e-09, 0.0002675311, 0.0004093423, 0.01046385, 0.03132254, 
    0.04141373, 0.01148049, 0.02919195, 0.02248128, 0.001555596, 0.000728461, 
    0.0006404741, 0.06912615, 0.03337157, 0.1176602, 0.06965273, 0.01268843, 
    0.03196027, 0.04784237, 0.001696113, 2.392871e-05, 2.764167e-06, 
    3.816603e-07, 0.0004512493, 0.008783583, 0.0003440314, 0.009880045, 
    8.145134e-07, 4.506614e-07,
  1.796962e-06, 0.05578338, 0.01473996, 0.02606417, 0.006733052, 0.0481648, 
    0.06151155, 0.0416345, 0.07727909, 0.01893733, 0.1505061, 0.09693527, 
    0.06377615, 0.03980529, 0.1185774, 0.05733204, 0.0142805, 0.002921903, 
    9.510655e-06, 0.0003023302, -1.126287e-06, 6.685858e-08, 0.001226657, 
    0.04414374, 0.0362752, 0.001411384, 0.001728854, 9.924132e-06, 
    1.189474e-05,
  0.09049097, 0.1163222, 0.04298593, 0.008511314, 0.02069052, 0.00383141, 
    0.003434914, 0.006430732, 0.009820191, 0.09741154, 0.01296597, 
    0.006858687, 0.04571339, 0.03675263, 0.05009951, 0.00799437, 0.004743788, 
    0.007761652, 0.0264225, 9.323459e-05, 0.001946264, 0.001585969, 
    0.09993704, 0.2052787, 0.1756798, 0.09442568, 0.1081474, 0.05022345, 
    0.03524208,
  0.03393504, 0.008485347, 0.005641979, 0.01878088, 0.01065195, 0.001222384, 
    0.006031242, 0.001120604, 0.004256911, 0.0747285, 0.01499068, 0.06110797, 
    0.06932297, 0.1215184, 0.03856595, 0.03693255, 0.08547376, 0.04941719, 
    0.001627832, 0.01682491, 0.008822764, 0.003360535, 0.002979753, 
    0.03750087, 0.04069468, 0.02227514, 1.020475e-06, 0.005009152, 0.04567061,
  0.1591167, 0.01652958, 0.01779243, 0.02381477, 0.01883811, 0.006094123, 
    0.0004370472, 0.0001552715, 0.001769669, 0.01035603, 0.03032087, 
    0.00534798, 0.006889537, 0.005609327, 0.001040073, 0.002298481, 
    0.0009097287, 0.01686877, 0.05042005, 0.03211958, 0.004828056, 
    0.02909486, 0.0009979655, 0.04860872, -3.256382e-05, 0.03360119, 
    0.02016496, 0.0006691647, 0.05940953,
  0.04270547, 0.08869594, 0.08573578, 0.08615542, 0.1039642, 0.05543895, 
    0.04813123, 0.03846603, 0.1942407, 0.1292828, 0.1439342, 0.150042, 
    0.1117513, 0.126297, 0.06054037, 0.03332784, 0.02256685, 0.06015468, 
    0.01872811, 0.008063915, 0.03962794, 0.0665647, 0.04554531, 0.03970435, 
    0.02859479, 0.1162579, 0.07614972, 0.02088606, 0.01571924,
  0.07210501, 0.1106099, 0.09741142, 0.1225906, 0.1131147, 0.0672947, 
    0.1339454, 0.1237152, 0.1022207, 0.04564098, 0.05207987, 0.1123339, 
    0.1473102, 0.1429016, 0.1683151, 0.21775, 0.1475552, 0.06010506, 
    0.05428824, 0.08274115, 0.08017708, 0.0374775, 0.1137761, 0.1920084, 
    0.1029274, 0.09424697, 0.1188498, 0.04442765, 0.08571495,
  0.1991782, 0.1175003, 0.1689381, 0.1061028, 0.2122852, 0.1283369, 
    0.1204559, 0.1419554, 0.1100536, 0.2121445, 0.1566378, 0.1543848, 
    0.2260348, 0.1817675, 0.1848567, 0.1519699, 0.2237208, 0.2470421, 
    0.1664176, 0.1502572, 0.1184419, 0.1822298, 0.1737769, 0.1194202, 
    0.2407888, 0.2053145, 0.1059027, 0.051989, 0.159876,
  0.2273608, 0.1694848, 0.1613142, 0.308121, 0.2176667, 0.1018431, 0.1229697, 
    0.1039919, 0.2021906, 0.06850996, 0.02504465, 0.0871892, 0.2217121, 
    0.2042201, 0.2280409, 0.2457428, 0.2583311, 0.2520717, 0.1761197, 
    0.1463149, 0.1812308, 0.2937272, 0.1666168, 0.1043497, 0.2109619, 
    0.1091481, 0.05097868, 0.1103709, 0.20578,
  0.312449, 0.1443067, 0.2225763, 0.1576445, 0.1331836, 0.09780718, 
    0.04679732, 0.09860827, 0.08754411, 0.1335069, 0.1726887, 0.1712941, 
    0.2360721, 0.1951684, 0.1651947, 0.1103687, 0.09941682, 0.1197401, 
    0.179777, 0.1784957, 0.1495192, 0.1429849, 0.1665672, 0.1917357, 
    0.2492746, 0.09439145, 0.01563574, 0.2237955, 0.2835048,
  0.2080559, 0.1696065, 0.1623854, 0.2223993, 0.1517394, 0.1314788, 
    0.09768764, 0.114515, 0.08852038, 0.09327218, 0.1156434, 0.1501804, 
    0.1688457, 0.1850421, 0.1355486, 0.1048624, 0.1114141, 0.1122888, 
    0.07305346, 0.06269848, 0.07483646, 0.07977619, 0.05513972, 0.03147482, 
    0.1012049, 0.04675448, 0.04162536, 0.1252924, 0.1858697,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.411549e-05, 0.0311556, 0.0232667, 
    0.1068516, 0.1767631, 0.1971033, 0.08943354, 0.0338272, 0.02710926, 
    0.0135809, 0.1270018, 0.2339497, 0.2847499, 0.2425388, 0.254788, 
    0.008949728, 1.249239e-05,
  0.33623, 0.2601451, 0.3000686, 0.2720976, 0.05845487, 0.03926153, 
    0.1276925, 0.0202805, 0.01878878, 0.02267928, -0.000231666, 0.004121387, 
    0.09456847, 0.2264604, 0.3259406, 0.3996961, 0.3744535, 0.3420842, 
    0.4174215, 0.3666073, 0.3057509, 0.3824892, 0.463098, 0.3305807, 
    0.3118493, 0.182971, 0.2372753, 0.2612158, 0.3940327,
  0.2849452, 0.243222, 0.2776484, 0.2617484, 0.2624353, 0.3064843, 0.2288125, 
    0.3181808, 0.3974559, 0.2883908, 0.2371703, 0.3429981, 0.3111209, 
    0.2634742, 0.2491126, 0.2384137, 0.1844968, 0.1939791, 0.2661455, 
    0.2337108, 0.2040929, 0.2174466, 0.283634, 0.2459927, 0.2611086, 
    0.1984869, 0.2651604, 0.2639978, 0.3155021,
  0.2042443, 0.2215583, 0.1551669, 0.1666503, 0.1479544, 0.1687746, 
    0.1587362, 0.1635517, 0.215818, 0.2271305, 0.1900987, 0.1732754, 
    0.1115717, 0.1406106, 0.1116575, 0.0624596, 0.04213998, 0.1862148, 
    0.1533927, 0.1304716, 0.1930828, 0.1853627, 0.1248614, 0.09296889, 
    0.1151162, 0.1666724, 0.15997, 0.1470508, 0.1754248,
  0.08267146, 0.05821683, 0.02813526, 0.06777409, 0.08885522, 0.05635173, 
    0.1007308, 0.1074576, 0.06712601, 0.05420645, 0.06987935, 0.1024415, 
    0.05576199, 0.04515471, 0.06936506, 0.111514, 0.1066963, 0.07788157, 
    0.06934641, 0.09964386, 0.1141183, 0.06879152, 0.1314817, 0.08363798, 
    0.05438526, 0.05261273, 0.05970304, 0.1442339, 0.172948,
  9.565642e-05, 0.02261164, 0.01597629, 0.01058202, 0.09115391, 0.08257371, 
    0.04239421, 0.03973571, 0.002537102, 0.02960939, 0.0511819, 0.01421564, 
    0.008083987, 0.01322298, 0.002229913, 0.1041332, 0.1298098, 0.08003326, 
    0.07274491, 0.09944196, 0.09472835, 0.01539898, 0.005716885, 
    0.0004808204, 0.02180902, 0.03877028, 0.07790237, 0.0565942, 0.01077998,
  5.124263e-08, 0.0001972642, 0.0006131512, 0.01048745, 0.03008837, 
    0.02605795, 0.008524098, 0.03366829, 0.01086124, 0.005443344, 
    0.0006131849, 0.0001178626, 0.04753289, 0.02273671, 0.1087397, 
    0.07388513, 0.01477528, 0.0374909, 0.03836092, 0.001540597, 
    -9.363704e-07, 2.613336e-06, 5.723915e-08, 0.001283962, 0.01665998, 
    0.000245409, 0.01840294, 1.45626e-06, 3.609099e-07,
  -0.0001043801, 0.05565876, 0.01313047, 0.02176127, 0.008968506, 0.05330215, 
    0.07174905, 0.05105599, 0.08361934, 0.02663533, 0.1568431, 0.1149133, 
    0.07169318, 0.03893147, 0.1095741, 0.05340926, 0.01490678, 0.003212467, 
    5.938326e-05, 0.0007168748, -6.826637e-07, 2.420563e-08, 0.01130645, 
    0.05401293, 0.0373533, 0.001854587, 0.0004860443, 4.167058e-05, 
    1.450363e-06,
  0.09208201, 0.1261857, 0.06153209, 0.007348231, 0.01305215, 0.003678368, 
    0.003799884, 0.003547521, 0.01072187, 0.09212479, 0.01249342, 
    0.006287286, 0.04893152, 0.03708821, 0.04676073, 0.008306814, 
    0.005048953, 0.00673089, 0.02256746, 0.0005682789, 0.002502665, 
    0.003454736, 0.1078306, 0.1983131, 0.1644528, 0.08557563, 0.094835, 
    0.05052555, 0.05077291,
  0.02644398, 0.02437936, 0.00400931, 0.04185923, 0.007126774, 0.001706601, 
    0.006930747, 0.0005184053, 0.006881568, 0.07988819, 0.01328044, 
    0.06456151, 0.07542364, 0.1168584, 0.05764233, 0.04343806, 0.1083485, 
    0.05326274, 0.001323681, 0.02280079, 0.008689255, 0.004261455, 
    0.005584436, 0.02373492, 0.03707668, 0.01176028, 1.012434e-06, 
    0.003128335, 0.04144299,
  0.1177225, 0.01436437, 0.01933141, 0.0121951, 0.03156921, 0.003003962, 
    0.008202968, 0.0003001865, 0.001973021, 0.005063144, 0.03053518, 
    0.004446805, 0.008713856, 0.00278599, 0.001154687, 0.002898126, 
    0.00125558, 0.01907195, 0.02140972, 0.02444649, 2.200365e-05, 0.03342308, 
    0.0007566107, 0.04768233, 5.038396e-05, 0.04701871, 0.007218054, 
    0.0005504929, 0.07955595,
  0.03552832, 0.09455672, 0.06572893, 0.07998669, 0.1063156, 0.04983723, 
    0.07864913, 0.05910992, 0.1791905, 0.1562062, 0.1456472, 0.1545812, 
    0.1181556, 0.1119909, 0.05316987, 0.02083954, 0.01804169, 0.05914164, 
    0.01691682, 0.003997687, 0.03548714, 0.05573545, 0.02814681, 0.04766859, 
    0.0154409, 0.09976178, 0.06636366, 0.01906107, 0.006147902,
  0.06831622, 0.1164551, 0.1008197, 0.1351822, 0.1076136, 0.06473867, 
    0.137151, 0.1234193, 0.09447666, 0.04187519, 0.05142084, 0.1173046, 
    0.1407923, 0.1287374, 0.1434047, 0.211625, 0.1401743, 0.08616745, 
    0.04941195, 0.08209791, 0.07515339, 0.03413583, 0.1262165, 0.1651563, 
    0.1043006, 0.08891601, 0.1157345, 0.04561822, 0.08794299,
  0.2017903, 0.1088043, 0.1650702, 0.1121272, 0.1926086, 0.1357331, 
    0.1254666, 0.1676906, 0.1506176, 0.2188659, 0.1751424, 0.1902417, 
    0.2506493, 0.1986291, 0.1941418, 0.1481446, 0.2257275, 0.2197263, 
    0.1518478, 0.1476763, 0.1287997, 0.1791779, 0.1870071, 0.1261292, 
    0.2250537, 0.1821562, 0.1174799, 0.04754353, 0.1455632,
  0.2388977, 0.1808576, 0.1531048, 0.3081775, 0.2224173, 0.09702145, 
    0.1407461, 0.1502045, 0.2326007, 0.2086989, 0.06862788, 0.1531869, 
    0.3036038, 0.2176102, 0.1966423, 0.2515551, 0.2987384, 0.2855916, 
    0.2552195, 0.1870911, 0.2023553, 0.3197578, 0.2008752, 0.1016012, 
    0.2242558, 0.1013468, 0.06278446, 0.1303382, 0.23486,
  0.3224726, 0.1874938, 0.2148973, 0.1373868, 0.1266468, 0.07611504, 
    0.04485984, 0.09909533, 0.1072859, 0.118149, 0.1767513, 0.1871101, 
    0.2187169, 0.2103225, 0.1694832, 0.1160538, 0.1522955, 0.16454, 
    0.1982301, 0.2542645, 0.2302694, 0.1534953, 0.1602113, 0.1939951, 
    0.251201, 0.1194209, 0.03012294, 0.283535, 0.2816983,
  0.2135518, 0.1764499, 0.1729502, 0.2195469, 0.1615443, 0.1340134, 
    0.0866398, 0.11536, 0.09331579, 0.09490489, 0.1382019, 0.1804146, 
    0.2090987, 0.248712, 0.2241281, 0.1884765, 0.1455286, 0.1321954, 
    0.1388147, 0.08760034, 0.1118584, 0.1476962, 0.05390365, 0.027866, 
    0.1400723, 0.08280563, 0.06823508, 0.149889, 0.1861266,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  -9.199804e-05, 0, 0, 0, 0, -5.081648e-06, 0, 0, 0, 0, 0, 1.141168e-07, 
    -1.44412e-05, 0.07856443, 0.06061438, 0.147903, 0.2996903, 0.2459341, 
    0.1615899, 0.1174462, 0.0942426, 0.07908651, 0.2349443, 0.2397521, 
    0.2571678, 0.3062764, 0.2955657, 0.1495133, 0.004549465,
  0.319661, 0.274495, 0.3169506, 0.3071428, 0.1021514, 0.08156389, 0.1539581, 
    0.03100802, 0.04380734, 0.05630139, 0.004235995, 0.008105135, 0.1486942, 
    0.2221895, 0.330509, 0.4126244, 0.3913977, 0.3388112, 0.4544415, 
    0.4130686, 0.3113656, 0.3732005, 0.4392842, 0.2990823, 0.3309956, 
    0.2145334, 0.2239732, 0.2580552, 0.397448,
  0.286788, 0.2478988, 0.297697, 0.2726582, 0.2764938, 0.3413007, 0.2489793, 
    0.3119553, 0.410486, 0.3086882, 0.2188875, 0.333436, 0.2932069, 
    0.2817966, 0.2434224, 0.2265515, 0.206128, 0.2107377, 0.2881633, 
    0.2462145, 0.2025539, 0.1944126, 0.2775088, 0.2008317, 0.241884, 
    0.1869874, 0.2620444, 0.2773327, 0.3052775,
  0.2270094, 0.2123895, 0.1578225, 0.1334251, 0.1382587, 0.162738, 0.1593107, 
    0.1639265, 0.1971669, 0.2319976, 0.1999748, 0.1764497, 0.1157127, 
    0.143427, 0.1084005, 0.05971983, 0.0403306, 0.1741136, 0.1729388, 
    0.1345081, 0.1940624, 0.2012271, 0.1251034, 0.08884691, 0.1000603, 
    0.2440358, 0.140044, 0.1459751, 0.168586,
  0.07932018, 0.06844868, 0.03474239, 0.05669169, 0.07351888, 0.05155498, 
    0.100822, 0.09878664, 0.06783978, 0.05711932, 0.0600617, 0.1065592, 
    0.05208637, 0.03954578, 0.07039572, 0.1130992, 0.1004392, 0.07971754, 
    0.07096905, 0.09769992, 0.1165162, 0.06606787, 0.1141188, 0.07744304, 
    0.03894945, 0.04965007, 0.05456501, 0.141341, 0.1640935,
  0.003095504, 0.03030329, 0.02393135, 0.01541986, 0.08801346, 0.07723414, 
    0.04086613, 0.03080598, -0.0001950415, 0.02248982, 0.06382692, 
    0.02155877, 0.01222647, 0.01306288, 0.003525655, 0.09895623, 0.1204659, 
    0.09044085, 0.07366402, 0.08990789, 0.09650337, 0.01894674, 0.005771617, 
    0.001206578, 0.02074916, 0.03852651, 0.09075657, 0.06585289, 0.01065866,
  8.020839e-07, 0.0002383876, 0.001335615, 0.01329779, 0.03648841, 
    0.02071353, 0.01220962, 0.05865465, 0.009122248, 0.02594231, 
    0.0004788484, 0.0001275646, 0.04071704, 0.0212261, 0.1105455, 0.07950295, 
    0.0283929, 0.04873385, 0.03590352, 0.002877078, 1.909488e-05, 
    5.688627e-06, 1.686799e-07, 0.002231791, 0.03074291, 0.0009342115, 
    0.02168021, 2.819096e-06, 2.254084e-07,
  9.234011e-06, 0.06804724, 0.01247261, 0.02141335, 0.01106862, 0.08201325, 
    0.1011459, 0.06822657, 0.09843451, 0.0345123, 0.1593854, 0.157414, 
    0.09244848, 0.04432119, 0.1113403, 0.05920364, 0.01840332, 0.003818842, 
    9.254739e-05, 0.0008517414, 4.975976e-06, 3.377904e-07, 0.003942729, 
    0.08471875, 0.04554055, 0.004433593, 0.002822859, 5.113137e-05, 
    7.303574e-06,
  0.1153774, 0.1483608, 0.09478842, 0.007357087, 0.01965754, 0.003640004, 
    0.003557538, 0.003923076, 0.01472013, 0.1113632, 0.01881717, 0.007896317, 
    0.07844266, 0.04430901, 0.060787, 0.009113013, 0.00584826, 0.009957299, 
    0.02497641, 0.003573818, 0.01849874, 0.008892863, 0.08504767, 0.2291085, 
    0.1863701, 0.08772344, 0.1083014, 0.07127327, 0.06870642,
  0.02403276, 0.07302269, 0.01245757, 0.09887197, 0.007019041, 0.002262798, 
    0.008392671, 0.0004851945, 0.01403675, 0.08606593, 0.0188757, 0.08131474, 
    0.08262441, 0.1319479, 0.06615929, 0.05371283, 0.1201251, 0.04744919, 
    0.002854097, 0.02573741, 0.009865977, 0.004303815, 0.01076835, 
    0.02484966, 0.03463305, 0.006995551, 0.0003037553, 0.03199899, 0.05740745,
  0.0287635, 0.01146903, 0.02320614, 0.00810669, 0.07118996, 0.003355986, 
    0.01687859, 0.0005045667, 0.01066795, 0.003078252, 0.02911181, 
    0.004611961, 0.01024516, 0.001843741, 0.001529424, 0.002998848, 
    0.002708332, 0.02058953, 0.005516964, 0.02388446, 2.325334e-05, 
    0.03426307, 0.001627039, 0.04986647, 0.0008958547, 0.07425455, 
    0.006468187, 3.659146e-06, 0.1097516,
  0.02966788, 0.08534174, 0.04463, 0.05394556, 0.1118183, 0.04111965, 
    0.1131473, 0.06687752, 0.1782299, 0.1764807, 0.1510775, 0.138855, 
    0.1324697, 0.09936406, 0.07176494, 0.02435992, 0.01376969, 0.0690606, 
    0.01999274, 0.004915162, 0.03828658, 0.05040744, 0.02288053, 0.04107058, 
    0.02118289, 0.0824215, 0.07407881, 0.01876044, 0.003822781,
  0.07014067, 0.1047117, 0.1052486, 0.1343556, 0.1116627, 0.0670831, 
    0.1255258, 0.1181023, 0.07669038, 0.04773786, 0.04749721, 0.1187304, 
    0.1324178, 0.1244708, 0.1213079, 0.1878318, 0.1169325, 0.078914, 
    0.06316812, 0.078807, 0.08272026, 0.02774113, 0.1317233, 0.1647362, 
    0.100685, 0.09378245, 0.1029364, 0.03730515, 0.1045497,
  0.1839358, 0.1097875, 0.1674932, 0.122486, 0.1829164, 0.1452338, 0.1321725, 
    0.1729621, 0.1897604, 0.213257, 0.193973, 0.2070932, 0.2690876, 0.174367, 
    0.2007561, 0.1253625, 0.2103719, 0.187066, 0.1287338, 0.1562189, 
    0.1315842, 0.1601187, 0.1873973, 0.1368409, 0.2312663, 0.1999439, 
    0.09871241, 0.05599962, 0.1327113,
  0.2079463, 0.1748208, 0.1413548, 0.2978292, 0.2092835, 0.1051736, 0.114116, 
    0.1579733, 0.2304061, 0.2188303, 0.1656554, 0.1825847, 0.3592863, 
    0.2196367, 0.1777654, 0.2531821, 0.2878093, 0.2864792, 0.2702198, 
    0.1933109, 0.1934123, 0.3206232, 0.1787544, 0.1435183, 0.2466201, 
    0.09804331, 0.0848581, 0.1388623, 0.2213852,
  0.3066614, 0.1636849, 0.210782, 0.1255746, 0.1350726, 0.06728856, 
    0.03462934, 0.1037596, 0.1073704, 0.105618, 0.1691878, 0.1910298, 
    0.200869, 0.2161181, 0.1617028, 0.109074, 0.1906022, 0.1679907, 
    0.1923892, 0.2237162, 0.2224367, 0.1576482, 0.1630962, 0.1844805, 
    0.2367673, 0.1676554, 0.05539611, 0.3086548, 0.2518296,
  0.213711, 0.1891439, 0.1728123, 0.2073047, 0.1780375, 0.1272239, 
    0.08579301, 0.1261336, 0.09097639, 0.09365758, 0.1328766, 0.168132, 
    0.1990797, 0.2419093, 0.2264581, 0.2062414, 0.1627585, 0.1187268, 
    0.1389886, 0.1738467, 0.2376838, 0.1940487, 0.08378932, 0.03273685, 
    0.1885061, 0.1110158, 0.1103336, 0.1532678, 0.1786651,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0.001440697, 0, 0, 0, 0, -0.000156291, 3.984829e-05, 0, 0, 0, 0.0007115821, 
    0.004165045, 0.001936256, 0.1232784, 0.06293794, 0.1553627, 0.3012421, 
    0.2911307, 0.1989333, 0.2572852, 0.2263542, 0.2290438, 0.3628592, 
    0.2455058, 0.2593192, 0.2928458, 0.3129973, 0.2187396, 0.07492073,
  0.2933173, 0.2953966, 0.3455881, 0.3236325, 0.1705321, 0.1072776, 
    0.1995955, 0.09275684, 0.06861757, 0.1322025, 0.04611737, 0.02083618, 
    0.157333, 0.2265595, 0.3248171, 0.4184071, 0.3373279, 0.3524812, 
    0.490228, 0.4555937, 0.368899, 0.3780994, 0.4621594, 0.313392, 0.370192, 
    0.2286316, 0.2169114, 0.2841562, 0.3868741,
  0.3090249, 0.2140288, 0.2738636, 0.2732592, 0.2497733, 0.3167926, 0.258963, 
    0.3528992, 0.3906443, 0.3363798, 0.2677017, 0.3196674, 0.2893792, 
    0.2713848, 0.251258, 0.2563039, 0.2231635, 0.2188987, 0.261505, 
    0.2094282, 0.2072435, 0.193756, 0.2777447, 0.2262559, 0.2830575, 
    0.2540288, 0.2770455, 0.2920028, 0.3107138,
  0.1954177, 0.2078493, 0.1740606, 0.1340628, 0.1484915, 0.1612695, 
    0.1428517, 0.1450937, 0.2042736, 0.2456825, 0.2233206, 0.1833633, 
    0.1163119, 0.158052, 0.09686213, 0.0563835, 0.03440098, 0.1884417, 
    0.158316, 0.1321873, 0.1885262, 0.1658756, 0.1360587, 0.08303364, 
    0.1044619, 0.1891243, 0.143123, 0.1615571, 0.1699344,
  0.07620607, 0.08182399, 0.03033839, 0.05933557, 0.07079067, 0.06404616, 
    0.1054408, 0.0986952, 0.06907839, 0.05375085, 0.05563681, 0.1167461, 
    0.0631963, 0.03747539, 0.07118393, 0.1149895, 0.09645066, 0.0934919, 
    0.07239217, 0.1006896, 0.1174957, 0.06008508, 0.1078164, 0.07475496, 
    0.03338127, 0.0442243, 0.0485629, 0.1312503, 0.170875,
  0.004201786, 0.0390056, 0.03925181, 0.01375151, 0.1145264, 0.0776879, 
    0.04152487, 0.04059684, -0.0001836346, 0.01617819, 0.08731788, 
    0.03533576, 0.01733521, 0.01402218, 0.008056567, 0.1045371, 0.1201734, 
    0.09825342, 0.06831297, 0.09202106, 0.130027, 0.02253337, 0.009456141, 
    0.002797932, 0.02705714, 0.04070503, 0.09718537, 0.06916988, 0.01319798,
  1.649403e-06, 0.0006210912, 0.001650754, 0.02172372, 0.04376485, 
    0.02192126, 0.0342732, 0.05777385, 0.01801668, 0.03993622, 0.001024493, 
    0.0003630992, 0.04024783, 0.0117281, 0.1112893, 0.08794111, 0.04541011, 
    0.0812187, 0.03658182, 0.004118375, 0.0002108286, -4.345511e-06, 
    1.45572e-07, 0.001234866, 0.03134772, 0.001406257, 0.01955133, 
    9.021183e-06, 1.604697e-07,
  0.0001552612, 0.07926105, 0.02376926, 0.02395594, 0.01820963, 0.09265693, 
    0.1334803, 0.07131291, 0.1035172, 0.04984412, 0.1713166, 0.1875213, 
    0.08957826, 0.04096791, 0.1147435, 0.0634907, 0.01608191, 0.004508308, 
    0.0007312488, 0.0003550408, 6.331491e-06, 1.141915e-06, 0.005115624, 
    0.1188996, 0.06061657, 0.003718957, 0.005515205, 6.022213e-05, 
    0.0001082205,
  0.1216804, 0.1939775, 0.1129196, 0.01203135, 0.02157639, 0.00276076, 
    0.002416596, 0.004674905, 0.01910461, 0.1477265, 0.03184082, 0.008370066, 
    0.08934056, 0.05265221, 0.06729235, 0.00937422, 0.006066401, 0.01023362, 
    0.0212277, 0.01611697, 0.01491219, 0.01542823, 0.0914919, 0.2626059, 
    0.2238769, 0.09222437, 0.1326765, 0.08215926, 0.09101236,
  0.02938821, 0.05376877, 0.02831756, 0.1662494, 0.008347148, 0.002022434, 
    0.008815238, 0.0005692252, 0.01660267, 0.08407851, 0.02437201, 
    0.08326935, 0.08381671, 0.1407447, 0.07132106, 0.07076286, 0.1318475, 
    0.04314919, 0.007350778, 0.03712449, 0.009453443, 0.00428575, 0.01864279, 
    0.03062703, 0.0361025, 0.00391044, -1.238952e-05, 0.0203093, 0.08662309,
  0.009716133, 0.004567123, 0.01718455, 0.006600268, 0.09050353, 0.00321247, 
    0.02598157, 0.0008064656, 0.0402773, 0.004797111, 0.02881787, 
    0.004435581, 0.01099711, 0.00238121, 0.003052162, 0.002655437, 
    0.003020191, 0.01201639, 0.0009699124, 0.01173819, 6.195566e-06, 
    0.03160578, 0.003334726, 0.05677047, 0.004842179, 0.08806626, 0.01764436, 
    9.286699e-06, 0.07818433,
  0.01831353, 0.07032239, 0.03773867, 0.02978718, 0.1109155, 0.03570781, 
    0.08416556, 0.07012071, 0.1687533, 0.2078662, 0.1663881, 0.1385957, 
    0.1522014, 0.08772732, 0.09648754, 0.0218521, 0.01104559, 0.06707623, 
    0.02424962, 0.008692668, 0.04566897, 0.04097737, 0.021354, 0.03501263, 
    0.03679219, 0.07086597, 0.06511752, 0.02704632, 0.002492554,
  0.06968537, 0.0793899, 0.09740613, 0.1253981, 0.1179587, 0.07674594, 
    0.1229237, 0.1023261, 0.04415849, 0.05443307, 0.05145996, 0.1180297, 
    0.1305404, 0.1146392, 0.1119269, 0.1766964, 0.123824, 0.08597396, 
    0.08223728, 0.07826518, 0.06674081, 0.02418367, 0.1406703, 0.1561789, 
    0.1083541, 0.09646182, 0.1271148, 0.0348814, 0.09872731,
  0.190622, 0.1002877, 0.1593303, 0.1248052, 0.1907257, 0.1526304, 0.1350241, 
    0.175283, 0.1927711, 0.1937205, 0.2071784, 0.20211, 0.2840301, 0.1827583, 
    0.2054096, 0.1219347, 0.2076748, 0.1830424, 0.1407302, 0.1607126, 
    0.1207596, 0.1490245, 0.1697609, 0.1471921, 0.2307626, 0.1982026, 
    0.1005035, 0.0604042, 0.126258,
  0.1859605, 0.1568729, 0.1208304, 0.2565331, 0.1914253, 0.1151223, 
    0.1049027, 0.1624908, 0.2611787, 0.2198046, 0.1786099, 0.1740997, 
    0.3701259, 0.2289765, 0.1788552, 0.255991, 0.2904722, 0.2960441, 
    0.2614088, 0.1768294, 0.1744242, 0.316788, 0.1654169, 0.1541654, 
    0.2607938, 0.1129669, 0.08322612, 0.1743748, 0.2014511,
  0.2981442, 0.1552664, 0.2125046, 0.1413713, 0.1287921, 0.07740139, 
    0.02205799, 0.1013392, 0.1084319, 0.09492389, 0.1663701, 0.1825052, 
    0.1982557, 0.220272, 0.1474021, 0.102604, 0.1718474, 0.1729211, 
    0.1949791, 0.1978867, 0.2141232, 0.1391918, 0.1595734, 0.181611, 
    0.2385683, 0.1979047, 0.09876557, 0.334507, 0.2538909,
  0.2186487, 0.2010707, 0.1731165, 0.1929404, 0.175665, 0.1082872, 
    0.08523028, 0.1282481, 0.07914422, 0.09771183, 0.1289203, 0.1585749, 
    0.1971958, 0.2217041, 0.2119453, 0.2174465, 0.1655202, 0.1037786, 
    0.1369874, 0.2435515, 0.2554759, 0.2114482, 0.09821018, 0.07571092, 
    0.1958112, 0.1424542, 0.1793912, 0.1478771, 0.1723129,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0.0004796693, -0.0004109319, 
    -0.0003421945, -0.0002734571, -0.0002047197, -0.0001359823, 
    -6.724492e-05, -0.0001668321, -0.0002355695, -0.0003043069, 
    -0.0003730443, -0.0004417817, -0.0005105191, -0.0005792565, 0,
  0.091052, -0.003702047, 0, 0, 0, -6.380077e-05, -0.0003387099, 
    -0.0004212306, 1.475076e-05, -3.762858e-06, 8.742549e-05, 0.004192709, 
    0.01516068, 0.149519, 0.1479686, 0.2326324, 0.3435913, 0.3140776, 
    0.26061, 0.3321851, 0.4068741, 0.37934, 0.4008817, 0.2593724, 0.2810874, 
    0.3247309, 0.3218784, 0.2327225, 0.2391496,
  0.2863562, 0.2964241, 0.4033196, 0.3667484, 0.2411851, 0.1568422, 
    0.2277108, 0.2010981, 0.129247, 0.1952742, 0.1912207, 0.06729232, 0.1626, 
    0.2267439, 0.3067571, 0.4208558, 0.3780719, 0.3840889, 0.4691329, 
    0.4526656, 0.3586104, 0.3751433, 0.4325138, 0.3354571, 0.385247, 
    0.2456249, 0.2120049, 0.2751813, 0.3419236,
  0.351602, 0.2810505, 0.2932602, 0.3100518, 0.3160634, 0.375979, 0.2831545, 
    0.3790285, 0.3979025, 0.317245, 0.2339999, 0.3163906, 0.3076033, 
    0.2993588, 0.2386876, 0.2534797, 0.2369376, 0.225703, 0.270861, 
    0.2360044, 0.2347778, 0.2113257, 0.2870405, 0.1723067, 0.259407, 
    0.2342899, 0.3063633, 0.302963, 0.3712885,
  0.1893951, 0.1908168, 0.1779237, 0.1402915, 0.1561664, 0.1709016, 
    0.1480132, 0.1559603, 0.2212249, 0.2430685, 0.2397893, 0.1825432, 
    0.1302985, 0.1640303, 0.08445287, 0.0719365, 0.04073319, 0.1829056, 
    0.160281, 0.1385005, 0.1639656, 0.1807178, 0.147392, 0.08307943, 
    0.09445877, 0.1675215, 0.1380105, 0.1583043, 0.1540519,
  0.07498901, 0.08836406, 0.04285064, 0.06660487, 0.06888551, 0.07632113, 
    0.09516738, 0.1056726, 0.08061237, 0.04957159, 0.05599321, 0.1288983, 
    0.05262973, 0.03933959, 0.09141064, 0.117988, 0.1026172, 0.1091973, 
    0.09466583, 0.1012824, 0.1123581, 0.05567237, 0.1010598, 0.07568251, 
    0.0529807, 0.05151634, 0.05476744, 0.127613, 0.1744535,
  0.004254196, 0.04343797, 0.08402892, 0.01445982, 0.128796, 0.08785398, 
    0.04482177, 0.04968132, -0.000240803, 0.01300297, 0.07022913, 0.03165801, 
    0.04591986, 0.01709394, 0.01816893, 0.1152093, 0.1107064, 0.09606043, 
    0.07824874, 0.1025238, 0.157941, 0.03073557, 0.01360196, 0.002720114, 
    0.04063423, 0.04618789, 0.09069233, 0.07978828, 0.02266379,
  4.238167e-05, 0.003479521, 0.00313111, 0.0307704, 0.03818576, 0.02415121, 
    0.02891334, 0.07217406, 0.01477884, 0.02910807, 0.001345759, 0.005387236, 
    0.03589188, 0.02003711, 0.1261752, 0.07575849, 0.04531658, 0.08227684, 
    0.04144846, 0.003776069, 0.004699719, -1.163324e-05, 1.00877e-07, 
    0.0002738696, 0.02945183, 0.004671511, 0.02281988, -2.301593e-08, 
    1.869805e-07,
  0.002302527, 0.07364939, 0.03871677, 0.03163949, 0.01307974, 0.07616664, 
    0.1030622, 0.05977428, 0.08567459, 0.04975777, 0.1703244, 0.1646693, 
    0.0837567, 0.04014822, 0.1000522, 0.05830346, 0.01556884, 0.007213499, 
    0.001412571, 0.001161531, 5.647465e-06, 9.318461e-07, 0.005923149, 
    0.1175507, 0.07879899, 0.003840389, 0.005867049, 2.948615e-05, 
    0.0001010102,
  0.08242279, 0.1999876, 0.1070953, 0.01592102, 0.01508052, 0.003353611, 
    0.00288251, 0.00634788, 0.02124721, 0.1706799, 0.03377731, 0.007637559, 
    0.07749265, 0.03770201, 0.0521482, 0.009573279, 0.007626974, 0.00959597, 
    0.02166243, 0.006240543, 0.01426672, 0.01223833, 0.07831472, 0.2496974, 
    0.2438008, 0.07540455, 0.1379148, 0.07040327, 0.0626788,
  0.03748258, 0.02626206, 0.03433706, 0.1865142, 0.007287847, 0.002027208, 
    0.0106067, 0.0003003863, 0.01852385, 0.07187648, 0.01893921, 0.071775, 
    0.06594472, 0.1164947, 0.07351936, 0.07118347, 0.1122225, 0.05145406, 
    0.009156632, 0.04871691, 0.01167186, 0.006152213, 0.02485106, 0.03742227, 
    0.02815984, 0.006498925, -1.998782e-05, 0.007284819, 0.0990136,
  0.001728082, 0.001456321, 0.01319775, 0.008000985, 0.06641848, 
    0.0009496745, 0.004777416, 0.0007595979, 0.06443558, 0.003960503, 
    0.03025343, 0.004172391, 0.008666267, 0.005133376, 0.005637381, 
    0.004292435, 0.006229627, 0.0006075411, 0.0004640133, 0.001234254, 
    3.656608e-06, 0.02661905, 0.006775026, 0.05827314, 0.007189289, 
    0.09241911, 0.01483851, 1.510122e-05, 0.02278484,
  0.01013747, 0.04776758, 0.01975659, 0.0241486, 0.1151191, 0.03318167, 
    0.0326978, 0.06236341, 0.1564942, 0.2285722, 0.1900245, 0.147002, 
    0.1595182, 0.07975152, 0.104586, 0.01718759, 0.01580431, 0.07539223, 
    0.02978487, 0.01380622, 0.03935185, 0.0484186, 0.02394064, 0.04558711, 
    0.04888292, 0.07419328, 0.05490798, 0.03105224, 0.001736078,
  0.06571072, 0.05712481, 0.1079133, 0.12175, 0.1213722, 0.07354146, 
    0.1195809, 0.05913569, 0.0140624, 0.06825712, 0.05545842, 0.116722, 
    0.1236376, 0.1224366, 0.11794, 0.1774868, 0.1300685, 0.08453471, 
    0.07195549, 0.09013241, 0.06917202, 0.01668296, 0.1420275, 0.1605679, 
    0.116662, 0.08867618, 0.1103482, 0.03923179, 0.09827018,
  0.16691, 0.09042178, 0.188293, 0.1448422, 0.1856833, 0.1572174, 0.1509159, 
    0.1859748, 0.175921, 0.176335, 0.220985, 0.1906664, 0.2924325, 0.2035152, 
    0.2071602, 0.1308405, 0.2160704, 0.1721188, 0.1165363, 0.1749033, 
    0.1372621, 0.1621512, 0.1760579, 0.1659707, 0.220066, 0.1947649, 
    0.09884331, 0.07640129, 0.1185826,
  0.1939369, 0.1560166, 0.1234234, 0.2786029, 0.2016118, 0.1334626, 
    0.1149685, 0.1852974, 0.2830264, 0.2181114, 0.174403, 0.1651129, 
    0.369083, 0.2350877, 0.1813733, 0.2475658, 0.2914964, 0.3165894, 
    0.2603785, 0.1620581, 0.155853, 0.2876548, 0.1560784, 0.1557761, 
    0.2764232, 0.1062828, 0.1159468, 0.1740063, 0.2114735,
  0.2951039, 0.1530151, 0.2027164, 0.1532432, 0.1271364, 0.09013611, 
    0.01976618, 0.07743113, 0.1166321, 0.1048415, 0.1736681, 0.1803951, 
    0.1961107, 0.2056008, 0.1473709, 0.08341086, 0.1520101, 0.190339, 
    0.1843709, 0.1839843, 0.1924325, 0.1184644, 0.1869334, 0.1991236, 
    0.2059862, 0.2261856, 0.1350951, 0.3443438, 0.2517675,
  0.2238294, 0.2099248, 0.1946586, 0.1774443, 0.1575058, 0.09110097, 
    0.1006606, 0.1360859, 0.08217993, 0.09860101, 0.1322386, 0.1532084, 
    0.2099369, 0.2177105, 0.2206839, 0.2151279, 0.1708569, 0.0982945, 
    0.1611074, 0.3098105, 0.2612845, 0.2238172, 0.1173842, 0.07863697, 
    0.1870719, 0.1504751, 0.1949214, 0.1557091, 0.1834318,
  0.006848796, 0.006259379, 0.005669961, 0.005080544, 0.004491127, 
    0.003901709, 0.003312292, 0.008682395, 0.009661473, 0.01064055, 
    0.01161963, 0.01259871, 0.01357779, 0.01455687, 0.01856254, 0.0207809, 
    0.02299925, 0.02521761, 0.02743597, 0.02965432, 0.03187268, 0.0262738, 
    0.02366578, 0.02105776, 0.01844974, 0.01584172, 0.01323371, 0.01062569, 
    0.00732033,
  0.2699322, 0.02864366, -0.000281155, 0, -9.188779e-05, 0.005556292, 
    0.0006042884, 0.004044537, 0.006147102, -5.377518e-05, -0.001411897, 
    0.03541813, 0.05722738, 0.1719662, 0.1280348, 0.2612272, 0.3473936, 
    0.3290511, 0.2488641, 0.353452, 0.4539436, 0.468733, 0.3963569, 
    0.2430392, 0.2495214, 0.3342575, 0.3079009, 0.2591784, 0.3208508,
  0.333887, 0.354328, 0.4797998, 0.4044922, 0.2772494, 0.167419, 0.2383108, 
    0.2553239, 0.1892669, 0.2399204, 0.2183578, 0.1010364, 0.1517974, 
    0.2292067, 0.3255537, 0.4288259, 0.3438408, 0.3854291, 0.4743629, 
    0.4075792, 0.3745576, 0.4030818, 0.4621537, 0.3441494, 0.4230103, 
    0.2941749, 0.2441011, 0.3470403, 0.3505793,
  0.2886316, 0.23229, 0.2771162, 0.2865805, 0.3099514, 0.3872813, 0.2698128, 
    0.4064927, 0.4386332, 0.3730983, 0.2783757, 0.3109043, 0.3041774, 
    0.2817131, 0.2538853, 0.2448935, 0.2507131, 0.2337333, 0.2957231, 
    0.2326337, 0.2399483, 0.2162555, 0.2871836, 0.1894576, 0.2670576, 
    0.2517398, 0.3509896, 0.2872457, 0.3359383,
  0.2205237, 0.1851523, 0.1888319, 0.1449421, 0.1499316, 0.1760708, 
    0.1496267, 0.1617197, 0.2372629, 0.2404351, 0.2321826, 0.1910643, 
    0.1273709, 0.1637065, 0.09262437, 0.07296693, 0.06123772, 0.2105109, 
    0.1770982, 0.1330473, 0.1614297, 0.1687863, 0.1523699, 0.08487589, 
    0.09689534, 0.1763942, 0.1519402, 0.1845665, 0.1658302,
  0.07358932, 0.09682265, 0.05042983, 0.06813538, 0.07191543, 0.09746312, 
    0.08684836, 0.1082226, 0.08210243, 0.0468419, 0.06298875, 0.1152005, 
    0.05211677, 0.04964681, 0.09608316, 0.1423116, 0.1261465, 0.1423789, 
    0.1077743, 0.1045908, 0.1086327, 0.05952243, 0.09586032, 0.07663938, 
    0.05507654, 0.0543543, 0.06871549, 0.1256927, 0.1919344,
  0.001771269, 0.03293379, 0.09769413, 0.01684733, 0.141209, 0.06041063, 
    0.04600509, 0.03740141, 0.0003241312, 0.01071048, 0.04670751, 0.01675179, 
    0.06891725, 0.02483088, 0.0276895, 0.1160877, 0.07758763, 0.09538461, 
    0.07825685, 0.09705191, 0.1638428, 0.05271962, 0.01999371, 0.005896096, 
    0.04679929, 0.05822638, 0.08539087, 0.09075364, 0.0189161,
  -3.363038e-06, 0.007295681, 0.003862923, 0.01532649, 0.03051735, 
    0.02691968, 0.02864126, 0.08471714, 0.003256176, 0.009363793, 0.01223863, 
    0.0423478, 0.03733964, 0.02161051, 0.1077642, 0.06768952, 0.04145576, 
    0.07952157, 0.03654834, 0.007450514, 0.003529233, 9.988229e-05, 
    5.869496e-08, 0.0001067764, 0.0238819, 0.01647483, 0.03016657, 
    0.0009168221, 3.881679e-07,
  0.0005050123, 0.07141244, 0.046248, 0.04390327, 0.01308013, 0.06388751, 
    0.09053521, 0.05258395, 0.07549284, 0.05061274, 0.150679, 0.1441569, 
    0.1023437, 0.0387559, 0.08174596, 0.05208743, 0.01669526, 0.007097273, 
    0.001465216, 0.0007380823, 4.103705e-06, 6.852304e-07, 0.008453959, 
    0.08121203, 0.08156218, 0.005869597, 0.0107912, 2.907483e-05, 2.649882e-05,
  0.06658754, 0.1344447, 0.03090619, 0.01766064, 0.01016216, 0.003643396, 
    0.003609337, 0.005869055, 0.01794099, 0.1431676, 0.03407437, 0.006946793, 
    0.06982926, 0.03057669, 0.04058928, 0.01231665, 0.01183219, 0.01288739, 
    0.0240535, 0.006249624, 0.01987563, 0.007073674, 0.06190074, 0.1910607, 
    0.2261292, 0.0686316, 0.1309307, 0.06080459, 0.04690286,
  0.02281479, 0.01188384, 0.01931251, 0.2116409, 0.005254185, 0.0024729, 
    0.009441985, 0.0001748786, 0.01800131, 0.0576551, 0.01753986, 0.06820653, 
    0.06004816, 0.104302, 0.06970195, 0.06236906, 0.08590241, 0.04707415, 
    0.01468196, 0.0470078, 0.01309007, 0.01158448, 0.02446392, 0.03788231, 
    0.02623118, 0.004907225, 2.221788e-05, 0.001066548, 0.03988285,
  4.700403e-05, 0.0001443427, 0.002165213, 0.002754976, 0.0248397, 
    0.0002827136, 0.001409499, 0.0001160221, 0.03019968, 0.0004719867, 
    0.02880009, 0.004790311, 0.01172617, 0.01402916, 0.01035732, 0.008834954, 
    0.007281641, 0.002382766, -5.391008e-05, -0.0004019723, 2.299638e-06, 
    0.02420575, 0.01201631, 0.05396209, 0.009330322, 0.09637152, 0.01259968, 
    1.167649e-05, 0.000928456,
  0.002442014, 0.03296333, 0.02214084, 0.01879192, 0.114644, 0.03301596, 
    0.006274831, 0.04724517, 0.1557803, 0.2648171, 0.1851821, 0.1526454, 
    0.1706354, 0.06956162, 0.1024458, 0.0157503, 0.02111344, 0.07853867, 
    0.030713, 0.0199399, 0.01955956, 0.06416956, 0.02819126, 0.05823316, 
    0.05573778, 0.08989915, 0.04620505, 0.03295702, 0.0005155771,
  0.05952256, 0.04430592, 0.1298325, 0.1252614, 0.1221472, 0.0602625, 
    0.1179694, 0.03621851, 0.005506099, 0.05868334, 0.06256291, 0.1167605, 
    0.1269268, 0.1342815, 0.1123848, 0.1829568, 0.1360354, 0.1031421, 
    0.06372412, 0.09869387, 0.08401782, 0.01928329, 0.170348, 0.1688616, 
    0.1400428, 0.09476221, 0.1111601, 0.05669852, 0.1110171,
  0.1722657, 0.1039928, 0.1601119, 0.1890129, 0.1739263, 0.1494769, 
    0.1528085, 0.1966668, 0.1413027, 0.1593001, 0.2492229, 0.1842432, 
    0.2885387, 0.213537, 0.2115236, 0.152943, 0.2348569, 0.1744018, 
    0.1083141, 0.1847853, 0.1259707, 0.1468769, 0.1636467, 0.159863, 
    0.2270067, 0.1932632, 0.1020407, 0.1040534, 0.1189919,
  0.2015092, 0.1573363, 0.1396117, 0.2730599, 0.2067081, 0.1497218, 
    0.1397998, 0.2115685, 0.3179844, 0.2180586, 0.1608498, 0.163699, 
    0.3762666, 0.2189552, 0.1841253, 0.2623788, 0.3069331, 0.3221514, 
    0.2462952, 0.1633199, 0.1631671, 0.2717133, 0.1388264, 0.1449176, 
    0.2823781, 0.1109649, 0.125025, 0.160291, 0.1948782,
  0.2883601, 0.1299787, 0.186845, 0.1643364, 0.1612662, 0.09859104, 
    0.03198851, 0.07452247, 0.1206041, 0.08649497, 0.1696612, 0.1792536, 
    0.1870051, 0.2153485, 0.1538756, 0.09806109, 0.1365436, 0.2066697, 
    0.1730893, 0.1696846, 0.1852891, 0.1160387, 0.2056133, 0.1991471, 
    0.1922858, 0.232047, 0.1580108, 0.3649442, 0.2542513,
  0.2284709, 0.2417182, 0.2202862, 0.1926712, 0.1649659, 0.09572067, 
    0.1053974, 0.1368414, 0.08651114, 0.10598, 0.1429285, 0.1630085, 
    0.224192, 0.2165187, 0.2385261, 0.201287, 0.1713974, 0.09805408, 
    0.1805247, 0.3121052, 0.2616375, 0.2250848, 0.1386107, 0.07173748, 
    0.1896577, 0.1342854, 0.1761285, 0.1520587, 0.1865824,
  0.04017341, 0.03704654, 0.03391966, 0.03079279, 0.02766591, 0.02453904, 
    0.02141216, 0.03379101, 0.03665895, 0.03952688, 0.04239482, 0.04526275, 
    0.04813069, 0.05099862, 0.03930668, 0.0437601, 0.04821353, 0.05266696, 
    0.05712039, 0.06157381, 0.06602724, 0.06355434, 0.05935985, 0.05516537, 
    0.05097087, 0.04677639, 0.0425819, 0.03838741, 0.04267491,
  0.40229, 0.186595, -0.002108173, 0, 8.578198e-05, 0.01520209, 0.002618985, 
    0.007108769, 0.009761464, 7.190612e-05, 0.01484056, 0.05661578, 
    0.1252711, 0.2050893, 0.07171436, 0.1571394, 0.3076282, 0.2957495, 
    0.2734566, 0.3792392, 0.4989912, 0.5132489, 0.4020608, 0.2234834, 
    0.2015386, 0.318346, 0.3298547, 0.3026949, 0.3914731,
  0.3801156, 0.3832706, 0.4708665, 0.4331467, 0.3112447, 0.1605769, 
    0.2561464, 0.2593534, 0.244888, 0.2603164, 0.1962408, 0.1229936, 
    0.1830666, 0.2650557, 0.3310875, 0.4412895, 0.3509265, 0.3607351, 
    0.5034703, 0.4251978, 0.3264602, 0.3686408, 0.4416969, 0.332798, 
    0.4165117, 0.2890919, 0.1951584, 0.3193401, 0.34831,
  0.3742395, 0.3154884, 0.3059918, 0.3367526, 0.2603694, 0.3819907, 0.313166, 
    0.405661, 0.4200714, 0.3459066, 0.2823684, 0.3231673, 0.3389232, 
    0.3044186, 0.2685681, 0.2498865, 0.2555501, 0.2396811, 0.2334041, 
    0.2356808, 0.2328085, 0.2244974, 0.2581032, 0.2082535, 0.3073318, 
    0.2616298, 0.381899, 0.2893736, 0.3853806,
  0.2367996, 0.2258363, 0.2064557, 0.1609273, 0.1534316, 0.1858546, 
    0.1592255, 0.1815341, 0.2428853, 0.2550634, 0.2387426, 0.1880983, 
    0.1155426, 0.1646134, 0.09549282, 0.08570313, 0.07204653, 0.2181741, 
    0.1913924, 0.1562799, 0.1965409, 0.2007182, 0.1968141, 0.09969945, 
    0.1039305, 0.1664882, 0.1727394, 0.1914082, 0.1957417,
  0.08105159, 0.114555, 0.05255811, 0.07903843, 0.08467331, 0.1121596, 
    0.09778119, 0.1166321, 0.0924632, 0.06766544, 0.05747208, 0.08408576, 
    0.05262117, 0.06351519, 0.1400068, 0.1563644, 0.1568003, 0.157975, 
    0.110081, 0.1115857, 0.1028064, 0.08593361, 0.09749169, 0.08450428, 
    0.05534372, 0.06887161, 0.0955331, 0.1299874, 0.2055919,
  0.0001825236, 0.03396944, 0.09325624, 0.01503941, 0.1337364, 0.03163289, 
    0.0512024, 0.03338797, 0.001325717, 0.008650838, 0.03702617, 0.007052106, 
    0.1066394, 0.04116111, 0.03527915, 0.1294003, 0.05879712, 0.1026613, 
    0.08360698, 0.08538733, 0.1570238, 0.09012321, 0.02539843, 0.005970488, 
    0.05270306, 0.07955595, 0.08766069, 0.08396327, 0.03091234,
  1.880537e-07, 0.005029492, 0.009160286, 0.02112629, 0.03606011, 0.03054137, 
    0.03666599, 0.09569727, 0.003416603, 0.005845692, 0.005819473, 
    0.06056638, 0.04286491, 0.02635813, 0.09570064, 0.06199607, 0.04762206, 
    0.08663174, 0.04136256, 0.0151801, 0.008514645, 0.002067322, 
    6.870556e-08, 5.624709e-05, 0.02392626, 0.06137304, 0.0653344, 
    0.009519376, 4.430171e-07,
  4.975922e-05, 0.0678956, 0.03387973, 0.04879085, 0.01939236, 0.05575319, 
    0.08472081, 0.05087476, 0.07303457, 0.04847009, 0.1535217, 0.1358807, 
    0.1140506, 0.03541215, 0.07039502, 0.04931833, 0.02014822, 0.0102423, 
    0.003299769, 0.001327122, 2.961021e-05, 4.460138e-07, 0.00485521, 
    0.08175287, 0.0899625, 0.01359155, 0.02153051, 5.394104e-05, 6.147708e-06,
  0.05563794, 0.1097813, 0.01549679, 0.03097481, 0.00883599, 0.005533477, 
    0.004626086, 0.005622962, 0.02089092, 0.1350091, 0.03020582, 0.007437775, 
    0.05527635, 0.0263167, 0.03986495, 0.01711763, 0.01460214, 0.01481538, 
    0.03097191, 0.0107188, 0.02777423, 0.01300673, 0.05496924, 0.1724953, 
    0.2249227, 0.06155741, 0.1293929, 0.05733353, 0.03571999,
  0.009494859, 0.0065491, 0.01059995, 0.1911626, 0.00444523, 0.002574709, 
    0.006391737, 0.000224049, 0.01900012, 0.05318546, 0.02125101, 0.06340563, 
    0.06039905, 0.102915, 0.07175984, 0.04806467, 0.0818942, 0.05386807, 
    0.02952132, 0.04843278, 0.01943406, 0.01485085, 0.02578812, 0.0413321, 
    0.03040425, 0.00194862, 4.071121e-05, 0.0003126511, 0.01812634,
  1.027719e-05, 1.516752e-05, 4.687827e-05, 0.0006874294, 0.008724757, 
    0.0001532925, 0.0001182716, 5.640208e-05, 0.009763177, 0.001972817, 
    0.02728276, 0.009150297, 0.02412286, 0.01660383, 0.02543992, 0.01516639, 
    0.01151186, 0.001210999, -7.904676e-06, -0.0001737882, 2.330958e-06, 
    0.0251711, 0.01648597, 0.05511195, 0.01376911, 0.1049936, 0.02292935, 
    8.70516e-06, 2.237876e-05,
  0.008835557, 0.01664495, 0.01991971, 0.01973886, 0.1060749, 0.0184113, 
    -0.002528061, 0.03511867, 0.1356525, 0.3038665, 0.2074322, 0.1482819, 
    0.1553231, 0.06608795, 0.1188728, 0.01761803, 0.02763597, 0.07969055, 
    0.04660294, 0.02631605, 0.006696116, 0.0825728, 0.0340789, 0.07587721, 
    0.0562253, 0.1087203, 0.04410914, 0.02844889, -0.0002404379,
  0.04466205, 0.03600759, 0.1609107, 0.1441651, 0.1227605, 0.05126937, 
    0.1171993, 0.02593419, 0.003231444, 0.04549679, 0.06780215, 0.1156351, 
    0.1202688, 0.1263506, 0.1125713, 0.1901703, 0.1374861, 0.1222656, 
    0.06508432, 0.1113858, 0.08450633, 0.02961925, 0.1902789, 0.185951, 
    0.13495, 0.09595687, 0.1090459, 0.08148361, 0.1304713,
  0.18966, 0.1292283, 0.2079141, 0.2027099, 0.182813, 0.1632899, 0.1613814, 
    0.213902, 0.1096142, 0.1418857, 0.2259794, 0.1801609, 0.3125327, 
    0.2331418, 0.2637126, 0.1740357, 0.2507062, 0.1819739, 0.1276644, 
    0.1886051, 0.1200021, 0.1384186, 0.215404, 0.1984701, 0.2504035, 
    0.1939519, 0.1212648, 0.1539176, 0.1399916,
  0.2033812, 0.1715776, 0.1985865, 0.2815826, 0.238332, 0.1622528, 0.1976803, 
    0.2123895, 0.3494507, 0.2265581, 0.1677581, 0.1839627, 0.390124, 
    0.3006702, 0.2036275, 0.2784088, 0.3116853, 0.3323288, 0.2275228, 
    0.1798684, 0.1742652, 0.2661692, 0.1511422, 0.1634811, 0.2956404, 
    0.1173916, 0.1421439, 0.1938158, 0.1885872,
  0.2938768, 0.1388738, 0.1873788, 0.2228494, 0.262069, 0.08162958, 
    0.06535005, 0.1059122, 0.1422816, 0.08464099, 0.1815507, 0.2291574, 
    0.1996567, 0.214302, 0.1737962, 0.08468866, 0.1224004, 0.1868207, 
    0.1800038, 0.2173237, 0.1846525, 0.1139352, 0.2274408, 0.1878643, 
    0.179029, 0.2539622, 0.2021358, 0.3588114, 0.2784275,
  0.2472348, 0.2789651, 0.2371365, 0.2195513, 0.2081537, 0.1306442, 
    0.1513912, 0.1693962, 0.1198793, 0.1589612, 0.1775219, 0.1965377, 
    0.2443281, 0.2377677, 0.2149169, 0.185141, 0.1625215, 0.08157328, 
    0.1376015, 0.3058629, 0.2554346, 0.2385896, 0.1706084, 0.07568558, 
    0.193434, 0.1304751, 0.1630176, 0.1435859, 0.240595,
  0.1169933, 0.1078761, 0.09875884, 0.08964161, 0.08052438, 0.07140715, 
    0.06228992, 0.08570375, 0.08965667, 0.09360959, 0.09756251, 0.1015154, 
    0.1054684, 0.1094213, 0.09465557, 0.1035216, 0.1123877, 0.1212537, 
    0.1301198, 0.1389859, 0.1478519, 0.1482278, 0.1445261, 0.1408243, 
    0.1371226, 0.1334208, 0.1297191, 0.1260173, 0.1242871,
  0.5538808, 0.3293002, 0.04856, -0.0005271481, 0.005646944, 0.01970991, 
    0.005593826, 0.01192736, 0.009984158, 0.001646099, 0.03114156, 
    0.09389131, 0.1607619, 0.2176062, 0.09034681, 0.1547715, 0.2632856, 
    0.2687154, 0.2783857, 0.3876369, 0.5271809, 0.5494518, 0.3918305, 
    0.2307128, 0.1445971, 0.3042737, 0.3249002, 0.3446721, 0.3919607,
  0.325624, 0.3772706, 0.3996572, 0.4112785, 0.3279595, 0.1542867, 0.2794936, 
    0.2864128, 0.2725925, 0.2637297, 0.1759839, 0.1210417, 0.1889392, 
    0.3019607, 0.3528544, 0.3660712, 0.3095816, 0.3191683, 0.4220919, 
    0.3830742, 0.3058196, 0.3986778, 0.390577, 0.353658, 0.32796, 0.2553097, 
    0.1577866, 0.3061038, 0.3859589,
  0.3944489, 0.3062814, 0.3038987, 0.3155543, 0.3224296, 0.3999326, 
    0.3272637, 0.4063388, 0.4051819, 0.3534524, 0.2730792, 0.3101884, 
    0.3462252, 0.3090309, 0.2701214, 0.248683, 0.2857173, 0.2583807, 
    0.2286507, 0.2180814, 0.2542473, 0.2378417, 0.261091, 0.2118567, 
    0.2895693, 0.2490264, 0.3514675, 0.3051063, 0.3626663,
  0.2508758, 0.2476875, 0.2318596, 0.157536, 0.1557704, 0.1827657, 0.187512, 
    0.1984042, 0.2557181, 0.2619049, 0.2511693, 0.216897, 0.1337107, 
    0.1905366, 0.09154235, 0.1045973, 0.1250889, 0.2378625, 0.2131342, 
    0.1871074, 0.2322784, 0.2033271, 0.2238905, 0.1011611, 0.1232702, 
    0.1917972, 0.165859, 0.2323814, 0.2198855,
  0.09522162, 0.1269959, 0.06088392, 0.09007616, 0.08360704, 0.1176461, 
    0.1130633, 0.1409233, 0.09037562, 0.08540111, 0.08168835, 0.06673446, 
    0.05012621, 0.07316907, 0.1555103, 0.1838861, 0.1733606, 0.1799879, 
    0.117586, 0.1352123, 0.1000902, 0.09305149, 0.1114109, 0.0909329, 
    0.05380133, 0.0912944, 0.1184923, 0.1359165, 0.20456,
  0.005047156, 0.03493559, 0.07349013, 0.0233691, 0.1173218, 0.02203818, 
    0.05397956, 0.03321935, 0.003848059, 0.01283931, 0.0295152, 0.0002148113, 
    0.06915597, 0.04030154, 0.04337961, 0.147765, 0.05995653, 0.1162638, 
    0.09519453, 0.09247088, 0.1544519, 0.09632803, 0.03699782, 0.006929717, 
    0.05427207, 0.09339621, 0.103532, 0.08924468, 0.03816434,
  4.895251e-05, 0.001938752, 0.02242179, 0.03705579, 0.03841763, 0.0386437, 
    0.04743096, 0.1104652, 0.004244187, 0.003920954, 0.003062487, 0.08091155, 
    0.05520542, 0.03027046, 0.09305289, 0.05916735, 0.05147087, 0.0993629, 
    0.03621571, 0.02420458, 0.02721729, 0.009649489, -9.496764e-08, 
    2.785916e-05, 0.0218526, 0.06469094, 0.07181536, 0.02827664, 3.524066e-05,
  5.671194e-06, 0.0546704, 0.03908024, 0.05598611, 0.02233738, 0.05289884, 
    0.08147381, 0.05447115, 0.07031112, 0.04588244, 0.1589118, 0.1222252, 
    0.1183062, 0.03764302, 0.0634001, 0.04624065, 0.02300238, 0.01721451, 
    0.006874707, 0.004726166, 0.0002759424, 2.598197e-06, 0.001433676, 
    0.08455426, 0.09574918, 0.0383951, 0.03930688, 0.0002493479, 1.98048e-06,
  0.04868275, 0.09051051, 0.01377212, 0.0388526, 0.009946599, 0.007580139, 
    0.008468488, 0.008745113, 0.02673926, 0.1331459, 0.02996029, 0.008943261, 
    0.04916038, 0.02392946, 0.03722934, 0.02155155, 0.02008934, 0.02098138, 
    0.035174, 0.02584841, 0.03419292, 0.02790953, 0.0480421, 0.1686717, 
    0.219275, 0.05473679, 0.1275753, 0.06165616, 0.04231774,
  0.004095177, 0.002011625, 0.00789417, 0.1139343, 0.005528782, 0.003004572, 
    0.006728937, 0.0003974886, 0.01988102, 0.05020872, 0.02997182, 
    0.06133121, 0.05560673, 0.09840132, 0.07317737, 0.04059037, 0.08569167, 
    0.06602927, 0.0457885, 0.0594344, 0.02346041, 0.01952846, 0.03666718, 
    0.05215289, 0.03899356, 0.002200444, 3.119908e-05, 7.150926e-06, 
    0.01073632,
  5.874059e-06, 8.02678e-06, 6.682028e-06, 0.000260986, 0.006987066, 
    0.0001868533, 1.33073e-05, 0.0001150603, 0.002606302, 0.00314805, 
    0.02793469, 0.02145581, 0.03067913, 0.03475169, 0.03820872, 0.02352695, 
    0.0214712, 0.003214387, 3.088563e-05, 0.001471989, 8.347553e-07, 
    0.03760311, 0.02307518, 0.04830214, 0.02064996, 0.1124105, 0.03097627, 
    4.737258e-06, 1.754255e-05,
  0.00686295, 0.003795156, 0.01896454, 0.01632906, 0.09463257, 0.006188106, 
    -0.004004423, 0.02372777, 0.1179982, 0.3392008, 0.2240836, 0.1553776, 
    0.1442105, 0.06584039, 0.1142708, 0.02251758, 0.0345214, 0.07330266, 
    0.07147625, 0.03312157, 0.002677958, 0.1038812, 0.03491022, 0.08965923, 
    0.06351651, 0.1201837, 0.05137037, 0.02044651, 3.20661e-05,
  0.03506112, 0.0366432, 0.1699494, 0.1523577, 0.08990484, 0.02359654, 
    0.1277834, 0.01766853, 0.0003427301, 0.04115698, 0.07330438, 0.1148989, 
    0.1212833, 0.1478334, 0.1111498, 0.1871628, 0.1445214, 0.1276205, 
    0.07743752, 0.1393354, 0.07878859, 0.01894862, 0.1829326, 0.2001648, 
    0.1564569, 0.1087874, 0.1158057, 0.1152857, 0.1656618,
  0.2282304, 0.156214, 0.2044485, 0.2091093, 0.1757292, 0.1451475, 0.1534559, 
    0.23027, 0.08440547, 0.111521, 0.2012903, 0.1750224, 0.3202668, 
    0.2482363, 0.2603073, 0.1673598, 0.2560064, 0.2031246, 0.1232479, 
    0.183288, 0.1069073, 0.138421, 0.1976521, 0.234135, 0.2807753, 0.1970322, 
    0.1430664, 0.192292, 0.1737969,
  0.235295, 0.1885064, 0.2073577, 0.2774172, 0.2473083, 0.2064943, 0.1968825, 
    0.1891222, 0.383291, 0.2256195, 0.1541019, 0.2107038, 0.3850185, 
    0.2577252, 0.2510175, 0.3093493, 0.3337261, 0.325849, 0.2374972, 
    0.1854535, 0.2015532, 0.245642, 0.1333314, 0.1518988, 0.2703907, 
    0.1369165, 0.1548669, 0.2072841, 0.1858916,
  0.3085258, 0.1602823, 0.1901717, 0.1589581, 0.2055193, 0.09210708, 
    0.07573362, 0.0861166, 0.1597585, 0.1104694, 0.1665467, 0.1562969, 
    0.163803, 0.1752986, 0.1717681, 0.07478321, 0.1415054, 0.1496632, 
    0.1802965, 0.1617557, 0.1864307, 0.1225932, 0.2321394, 0.1585544, 
    0.1722527, 0.2916111, 0.2089291, 0.356163, 0.3708278,
  0.2795347, 0.2722609, 0.2518266, 0.2648332, 0.2123935, 0.104269, 0.165501, 
    0.1563035, 0.1074042, 0.1437935, 0.1753053, 0.2122858, 0.2479158, 
    0.2578669, 0.2480279, 0.1813594, 0.1529448, 0.1158609, 0.1275219, 
    0.2789582, 0.2752964, 0.255544, 0.1755649, 0.08385728, 0.1827865, 
    0.1374448, 0.1492248, 0.1784102, 0.232174,
  0.2205237, 0.2104179, 0.2003121, 0.1902063, 0.1801005, 0.1699947, 
    0.1598889, 0.1828387, 0.18822, 0.1936013, 0.1989826, 0.2043639, 
    0.2097452, 0.2151265, 0.2040007, 0.2164378, 0.2288748, 0.2413119, 
    0.2537489, 0.266186, 0.278623, 0.2846336, 0.276921, 0.2692085, 0.2614959, 
    0.2537834, 0.2460709, 0.2383583, 0.2286083,
  0.6179182, 0.4483205, 0.1781649, 0.01605432, 0.008395975, 0.02374589, 
    0.008914863, 0.01439551, 0.01278175, 0.001936666, 0.06074015, 0.119456, 
    0.1795517, 0.2324824, 0.1273945, 0.1650071, 0.2689712, 0.2416615, 
    0.2524445, 0.3822384, 0.5688695, 0.5698454, 0.3899612, 0.2259736, 
    0.1880053, 0.2295097, 0.3203169, 0.411457, 0.4285446,
  0.3261971, 0.4056633, 0.4153458, 0.3941153, 0.3271745, 0.1432957, 
    0.3369895, 0.2957531, 0.3012005, 0.289309, 0.1861544, 0.1185931, 
    0.1865718, 0.3206176, 0.3680847, 0.3540044, 0.3245296, 0.3225639, 
    0.3906106, 0.3319013, 0.3126172, 0.4241525, 0.4116008, 0.3423983, 
    0.310576, 0.2497376, 0.1642465, 0.3050645, 0.3845214,
  0.3320287, 0.2721376, 0.2965947, 0.2812997, 0.2995644, 0.3813345, 0.300116, 
    0.3741493, 0.4131684, 0.3430623, 0.2743886, 0.3258307, 0.3407758, 
    0.3109372, 0.2799066, 0.2589041, 0.2861434, 0.2596664, 0.2639985, 
    0.2513619, 0.2657996, 0.2374027, 0.2784072, 0.228559, 0.3104407, 
    0.2292242, 0.3043327, 0.3184443, 0.370432,
  0.2431315, 0.2367587, 0.239966, 0.1775661, 0.1959622, 0.2052132, 0.204123, 
    0.215636, 0.2766466, 0.2717312, 0.2639014, 0.2307116, 0.1376021, 
    0.2095581, 0.1025741, 0.1301069, 0.144146, 0.2414335, 0.2429814, 
    0.2071947, 0.2609807, 0.2019577, 0.2153218, 0.1121393, 0.1411657, 
    0.1982747, 0.1879629, 0.2607354, 0.2115071,
  0.1030461, 0.1455828, 0.08629886, 0.09719928, 0.08025033, 0.1316321, 
    0.1156228, 0.1777833, 0.1006395, 0.09933562, 0.08173252, 0.07487237, 
    0.05400263, 0.07402629, 0.156586, 0.1673623, 0.1894723, 0.1991943, 
    0.1125343, 0.1511736, 0.1090849, 0.1251526, 0.1359976, 0.09319661, 
    0.04871425, 0.100913, 0.1466343, 0.1543586, 0.2018643,
  0.01202275, 0.0281001, 0.043961, 0.02205091, 0.1068137, 0.02883404, 
    0.06411041, 0.04635258, 0.01183607, 0.009124653, 0.02387282, 
    2.875052e-05, 0.02021831, 0.07829179, 0.0461491, 0.1362214, 0.0797867, 
    0.1438426, 0.1156239, 0.07824446, 0.1423796, 0.1145149, 0.04581206, 
    0.0066409, 0.05077297, 0.1001427, 0.1174232, 0.1076505, 0.03637585,
  1.806596e-05, -0.0001257182, 0.01815809, 0.04441912, 0.03956257, 
    0.04165645, 0.04924916, 0.1090019, 0.005146269, 0.003062118, 0.005444707, 
    0.01132952, 0.06943296, 0.04233535, 0.07872813, 0.05784787, 0.04467822, 
    0.08964166, 0.03708693, 0.02643601, 0.05651541, 0.03687186, 0.0002703784, 
    4.528037e-06, 0.0228857, 0.0653325, 0.06579383, 0.07423659, 0.004550135,
  1.640954e-06, 0.04406854, 0.04344735, 0.06020252, 0.02291347, 0.04805177, 
    0.07343486, 0.05280358, 0.06575835, 0.04158937, 0.1293376, 0.09628508, 
    0.1411815, 0.04136736, 0.0564359, 0.03868601, 0.02286254, 0.01857677, 
    0.01114051, 0.01032901, 0.001391945, 0.0002571037, 8.882909e-05, 
    0.08873167, 0.1011005, 0.02148391, 0.05211325, 0.003867983, 3.568862e-05,
  0.04426683, 0.07106043, 0.01601792, 0.04488419, 0.01122546, 0.009848578, 
    0.01178122, 0.01019851, 0.03666194, 0.1409028, 0.03012695, 0.01153638, 
    0.04574398, 0.02238867, 0.03467008, 0.02029204, 0.02369365, 0.02649496, 
    0.03386666, 0.02364059, 0.04418429, 0.03547418, 0.04396825, 0.1671282, 
    0.2069987, 0.04490691, 0.1130074, 0.07693467, 0.05301557,
  0.001818354, 0.0004844391, 0.001853884, 0.0531711, 0.007467266, 0.00414044, 
    0.009174674, 0.002367796, 0.02227854, 0.05554195, 0.03652692, 0.05553216, 
    0.0515243, 0.08782312, 0.06438114, 0.03398706, 0.08605174, 0.08362663, 
    0.06095003, 0.07012442, 0.02499185, 0.02220111, 0.05100958, 0.08162211, 
    0.04686762, 0.003254809, 1.324673e-05, 2.973149e-06, 0.006351274,
  4.683643e-06, 3.343793e-06, 1.683306e-06, 8.58505e-05, 0.00439661, 
    0.000236889, 1.497631e-05, 0.000194037, 0.002172649, 0.006295104, 
    0.03032045, 0.02718054, 0.02509759, 0.03068435, 0.04197128, 0.02415492, 
    0.03666172, 0.009340513, 0.001509548, -0.0002420873, 2.46531e-07, 
    0.05677133, 0.03157559, 0.0514043, 0.02411089, 0.09405176, 0.0484707, 
    8.913925e-07, 8.818392e-06,
  0.003169202, 0.0007495738, 0.01914413, 0.01119075, 0.07473987, 0.001394798, 
    -0.003454921, 0.01672824, 0.1078724, 0.355013, 0.1924829, 0.1680782, 
    0.1552378, 0.06216654, 0.1128503, 0.03314075, 0.0353302, 0.06587168, 
    0.08056356, 0.0458259, 0.0007285251, 0.1111069, 0.03994619, 0.07979273, 
    0.08878341, 0.1281116, 0.06999649, 0.04433936, 0.005138705,
  0.01894783, 0.03348457, 0.1492845, 0.1441925, 0.06578483, 0.01219914, 
    0.1400758, 0.01093766, -0.0001355017, 0.03264794, 0.07488344, 0.114846, 
    0.1253045, 0.147198, 0.1192014, 0.1842623, 0.1773033, 0.122773, 
    0.09889975, 0.1581323, 0.04448368, 0.02552898, 0.1931894, 0.1983754, 
    0.1581193, 0.129334, 0.1098547, 0.1306549, 0.1711037,
  0.2677126, 0.1631743, 0.2114607, 0.1987057, 0.1220685, 0.1239799, 
    0.1349162, 0.2349525, 0.06048119, 0.09505696, 0.1613732, 0.1792852, 
    0.3039023, 0.2908744, 0.2485185, 0.1884063, 0.2879164, 0.2224871, 
    0.1279321, 0.1922867, 0.1076039, 0.1208467, 0.1403117, 0.2520011, 
    0.2947323, 0.1957205, 0.1835369, 0.2068392, 0.1954861,
  0.2434296, 0.2130029, 0.2477174, 0.2411904, 0.2354937, 0.2092583, 
    0.1731906, 0.1220187, 0.3394985, 0.2323988, 0.09889686, 0.2264758, 
    0.3985921, 0.2391028, 0.2235067, 0.2742014, 0.3064459, 0.3279447, 
    0.2196099, 0.1663779, 0.2231779, 0.2228793, 0.1118697, 0.1659061, 
    0.2832392, 0.1818469, 0.1974004, 0.223329, 0.205538,
  0.3186479, 0.208417, 0.201332, 0.1403318, 0.1489479, 0.07164678, 
    0.02940569, 0.07977063, 0.1451738, 0.1084989, 0.1360497, 0.1724212, 
    0.1192684, 0.1552866, 0.1679778, 0.07377987, 0.1220879, 0.1526829, 
    0.1806903, 0.149325, 0.2077628, 0.112785, 0.2008084, 0.1322196, 
    0.1744273, 0.3143045, 0.2037565, 0.3281804, 0.3183136,
  0.2891538, 0.3247292, 0.2998435, 0.204067, 0.16213, 0.100245, 0.1359921, 
    0.1403162, 0.0878632, 0.09626106, 0.1187932, 0.2139428, 0.2245789, 
    0.2103616, 0.223995, 0.1952882, 0.1538531, 0.1070411, 0.211884, 
    0.3483037, 0.3056254, 0.274979, 0.1869123, 0.09299737, 0.1802599, 
    0.1322994, 0.1426421, 0.1965088, 0.1867135,
  0.2861318, 0.281342, 0.2765522, 0.2717624, 0.2669725, 0.2621827, 0.2573929, 
    0.3132749, 0.3223349, 0.331395, 0.3404551, 0.3495151, 0.3585752, 
    0.3676352, 0.3353816, 0.3435131, 0.3516446, 0.3597761, 0.3679076, 
    0.3760391, 0.3841707, 0.3896434, 0.3772417, 0.3648399, 0.3524382, 
    0.3400364, 0.3276347, 0.3152329, 0.2899636,
  0.6023822, 0.5506296, 0.3264333, 0.05232674, 0.02271631, 0.0443468, 
    0.0367104, 0.0191578, 0.01295203, 0.006810752, 0.1197627, 0.1233925, 
    0.2146273, 0.2193871, 0.1407278, 0.1548963, 0.2455087, 0.2023983, 
    0.2440083, 0.3466075, 0.5758526, 0.6032737, 0.410514, 0.2304513, 
    0.2425251, 0.1982517, 0.3145659, 0.4080475, 0.4654171,
  0.3256164, 0.3786667, 0.4250607, 0.3767467, 0.3106177, 0.1454703, 
    0.3693519, 0.2978273, 0.3112699, 0.2907693, 0.1909888, 0.1192969, 
    0.1751135, 0.349823, 0.382323, 0.3689353, 0.3312255, 0.3231371, 
    0.4266857, 0.3501873, 0.401642, 0.429273, 0.4655522, 0.3759191, 
    0.3330653, 0.3097045, 0.2043139, 0.3338259, 0.368193,
  0.3956598, 0.2947649, 0.3304054, 0.2915055, 0.2984191, 0.3912158, 
    0.3796447, 0.4057784, 0.4441905, 0.3641081, 0.2979666, 0.3513277, 
    0.3643533, 0.363317, 0.33429, 0.2954217, 0.2835942, 0.2747265, 0.3167152, 
    0.3267798, 0.3496299, 0.3235134, 0.3067652, 0.2885202, 0.3410954, 
    0.2618589, 0.4038239, 0.3792021, 0.4494617,
  0.2596773, 0.2689041, 0.2789986, 0.2362198, 0.2340943, 0.2476644, 
    0.2218271, 0.2625897, 0.2986335, 0.3146545, 0.3046729, 0.2638791, 
    0.1799895, 0.2563156, 0.1667047, 0.2319982, 0.1851414, 0.3043445, 
    0.2632238, 0.2473008, 0.2859605, 0.218536, 0.2626084, 0.1212295, 
    0.1767831, 0.2399738, 0.233136, 0.3280728, 0.2363286,
  0.1316399, 0.1768172, 0.1050424, 0.10727, 0.108764, 0.155438, 0.1222766, 
    0.200774, 0.1435465, 0.1549993, 0.1292465, 0.09816828, 0.07518136, 
    0.1363291, 0.1719689, 0.1665559, 0.2208352, 0.2340226, 0.1208938, 
    0.1577437, 0.1522697, 0.1585632, 0.1634699, 0.09868576, 0.06868897, 
    0.1133108, 0.1483458, 0.1792142, 0.220179,
  0.0274095, 0.02956616, 0.03730597, 0.04771729, 0.09539469, 0.05689178, 
    0.07481786, 0.07007772, 0.02948144, 0.006104686, 0.01984102, 1.31353e-05, 
    0.004475096, 0.1059467, 0.06544962, 0.1281181, 0.07452622, 0.1427992, 
    0.1223411, 0.07082187, 0.1201715, 0.1572471, 0.06591761, 0.005708626, 
    0.04702817, 0.1052392, 0.1249964, 0.09849102, 0.05582771,
  0.02240219, 1.101653e-05, 0.02213539, 0.04778847, 0.03530876, 0.05258882, 
    0.0424959, 0.1145884, 0.009271106, 0.002239428, 0.004172268, 0.001099295, 
    0.0560353, 0.04964074, 0.07163348, 0.0738333, 0.05254099, 0.07679185, 
    0.03497601, 0.02212692, 0.0517641, 0.05259807, 0.01090641, -3.937114e-06, 
    0.02670744, 0.08140133, 0.05860199, 0.07142942, 0.04757775,
  7.276027e-05, 0.02860043, 0.04551689, 0.06904163, 0.02287015, 0.04051073, 
    0.06372783, 0.04675349, 0.05118518, 0.03465188, 0.09994786, 0.08020262, 
    0.1314965, 0.04067105, 0.04621881, 0.03227174, 0.02198447, 0.01804712, 
    0.01523895, 0.01746452, 0.003408711, 0.002852149, 4.82973e-05, 0.0829917, 
    0.1003132, 0.0192528, 0.04996912, 0.01485454, 0.002431433,
  0.04627781, 0.05662144, 0.01789363, 0.03750851, 0.01311598, 0.01153219, 
    0.01470294, 0.01245444, 0.05090914, 0.1587526, 0.03365479, 0.01461087, 
    0.04216107, 0.0187564, 0.02865021, 0.02024122, 0.01848565, 0.02396498, 
    0.03200191, 0.02599561, 0.04857555, 0.03860066, 0.03405302, 0.1524546, 
    0.192945, 0.03620934, 0.09626244, 0.06770736, 0.05331756,
  0.0008621891, 0.0001613326, 0.0001891263, 0.02825549, 0.01186753, 
    0.01152474, 0.01438741, 0.006220996, 0.02433585, 0.0540624, 0.04292258, 
    0.04806287, 0.04458834, 0.07647757, 0.05866389, 0.03730278, 0.08895936, 
    0.1026887, 0.07967018, 0.07328366, 0.02681688, 0.02106902, 0.06553687, 
    0.09320785, 0.04784404, 0.005456672, 0.0003515623, 1.378019e-06, 
    0.003928877,
  3.548062e-06, 1.54616e-06, 6.675071e-07, 0.0001399413, 0.002637646, 
    0.0004086919, 9.841429e-06, 0.0001507279, 0.0008106263, 0.01919336, 
    0.03227734, 0.03024443, 0.02296167, 0.02734961, 0.03339513, 0.02825183, 
    0.0428601, 0.04755442, 0.01730287, -0.0001045916, 1.643351e-07, 
    0.07765998, 0.05171765, 0.05677572, 0.03486162, 0.06928091, 0.04883054, 
    1.214368e-05, 5.880343e-06,
  0.0007289879, 0.0004981167, 0.02312365, 0.00855435, 0.05839467, 
    0.000692016, -0.002843133, 0.01590074, 0.09878944, 0.3452969, 0.173175, 
    0.2197959, 0.1977548, 0.1092185, 0.1195634, 0.03746084, 0.05980506, 
    0.1190487, 0.09758618, 0.05249106, 0.0001141468, 0.1099146, 0.04685944, 
    0.07459902, 0.09154515, 0.1278175, 0.08931082, 0.09276366, 0.01329383,
  0.01018338, 0.03515282, 0.1214086, 0.1499557, 0.0507869, 0.005970448, 
    0.143938, 0.006998509, -0.0001559339, 0.01875421, 0.07078885, 0.1097009, 
    0.1417797, 0.1747109, 0.1568561, 0.2203351, 0.2310838, 0.1514608, 
    0.1500984, 0.1438097, 0.03134886, 0.01769054, 0.2137426, 0.2543134, 
    0.1825605, 0.1518862, 0.1303717, 0.150339, 0.1629989,
  0.2586038, 0.1603524, 0.2058087, 0.1714305, 0.07974294, 0.09764871, 
    0.1147093, 0.2372653, 0.04134663, 0.06550083, 0.1271171, 0.1853414, 
    0.3413436, 0.3228854, 0.2994676, 0.2366126, 0.2556998, 0.2654688, 
    0.1443645, 0.2398011, 0.08226546, 0.114263, 0.1334427, 0.2604341, 
    0.304739, 0.2155029, 0.2502016, 0.2511297, 0.2316802,
  0.2423833, 0.2556085, 0.2692041, 0.2750505, 0.1950413, 0.1545924, 
    0.1055522, 0.1047286, 0.332312, 0.2478679, 0.07396203, 0.1892008, 
    0.411417, 0.3189432, 0.2319053, 0.2467584, 0.2998013, 0.3249345, 
    0.2221185, 0.1364759, 0.2182512, 0.2180183, 0.09688096, 0.1919359, 
    0.3206656, 0.2377881, 0.1721386, 0.268192, 0.2255224,
  0.3073373, 0.1783373, 0.243706, 0.1703891, 0.2080271, 0.06194662, 
    0.02050116, 0.122155, 0.1429824, 0.112945, 0.1297457, 0.1546242, 
    0.1201115, 0.1112544, 0.1651545, 0.07666325, 0.08292851, 0.1662494, 
    0.1748559, 0.1522072, 0.2343954, 0.09687489, 0.1776554, 0.1419538, 
    0.1738232, 0.3298562, 0.1739364, 0.3119135, 0.2971464,
  0.2572759, 0.2626201, 0.2941162, 0.2060798, 0.1228997, 0.09706719, 
    0.1280691, 0.1260803, 0.05259524, 0.09040591, 0.1238986, 0.204204, 
    0.2262095, 0.1960329, 0.2037655, 0.1966062, 0.1541224, 0.1390079, 
    0.1937142, 0.2857245, 0.2772999, 0.285132, 0.2309102, 0.1285075, 
    0.172788, 0.1285111, 0.1596997, 0.1785653, 0.2232821,
  0.3371134, 0.3364006, 0.3356878, 0.334975, 0.3342622, 0.3335494, 0.3328366, 
    0.3375599, 0.3492414, 0.3609229, 0.3726044, 0.3842859, 0.3959673, 
    0.4076488, 0.4114118, 0.4163554, 0.421299, 0.4262426, 0.4311861, 
    0.4361297, 0.4410733, 0.4533367, 0.4374245, 0.4215122, 0.4055999, 
    0.3896876, 0.3737753, 0.357863, 0.3376836,
  0.5823221, 0.5602188, 0.434901, 0.09154928, 0.05511614, 0.08526134, 
    0.07810929, 0.03629498, 0.007700712, 0.01325878, 0.1429703, 0.1614545, 
    0.2379062, 0.1700835, 0.1695635, 0.119827, 0.2286618, 0.2213123, 
    0.2530093, 0.3337774, 0.5891625, 0.6193313, 0.4055758, 0.2472238, 
    0.2685213, 0.2025325, 0.3468735, 0.3241856, 0.5024651,
  0.4259211, 0.4045502, 0.396821, 0.3540475, 0.2952707, 0.1455652, 0.3695027, 
    0.3576289, 0.3101053, 0.2991098, 0.1946914, 0.1150275, 0.1692117, 
    0.3572885, 0.4191093, 0.3939825, 0.3660303, 0.381403, 0.5260168, 
    0.455859, 0.4530977, 0.4711032, 0.4958373, 0.4038863, 0.3582901, 
    0.3180166, 0.2099918, 0.3864194, 0.3884945,
  0.3927085, 0.3086151, 0.3526536, 0.3424405, 0.301518, 0.3939391, 0.3577256, 
    0.4285025, 0.5059641, 0.3775549, 0.3479042, 0.3393328, 0.4208928, 
    0.3842896, 0.3389614, 0.3344246, 0.3173298, 0.2848792, 0.3818525, 
    0.3816165, 0.3742451, 0.3991759, 0.371541, 0.3478671, 0.4151998, 
    0.3287398, 0.4297612, 0.4495263, 0.4338447,
  0.3051157, 0.3317886, 0.2976239, 0.2425038, 0.2555167, 0.2563585, 
    0.2667214, 0.2759517, 0.3066324, 0.3358943, 0.3103803, 0.3204418, 
    0.2520922, 0.2851869, 0.2600906, 0.2490363, 0.1988827, 0.3071178, 
    0.2747024, 0.3159668, 0.3526414, 0.2882194, 0.3673958, 0.1377643, 
    0.1931823, 0.2942497, 0.2309499, 0.3870969, 0.3121203,
  0.1666393, 0.1731569, 0.1421856, 0.1593322, 0.1427069, 0.1684356, 
    0.1694965, 0.2702274, 0.1903004, 0.2386835, 0.1550454, 0.1505146, 
    0.05915124, 0.1639599, 0.2125572, 0.1894991, 0.2354032, 0.2858142, 
    0.1687174, 0.2359675, 0.1844666, 0.1406042, 0.168312, 0.1150083, 
    0.08270941, 0.1257618, 0.1340764, 0.180024, 0.2320104,
  0.06982013, 0.06066338, 0.03572807, 0.1147783, 0.08167886, 0.06375922, 
    0.13153, 0.09481687, 0.07786537, 0.02248793, 0.02132342, 2.245789e-06, 
    -0.0002962416, 0.09889618, 0.07072633, 0.1434194, 0.09786293, 0.1561867, 
    0.1343216, 0.07577839, 0.1296409, 0.1446608, 0.1175468, 0.005381629, 
    0.0488992, 0.1236998, 0.1224159, 0.1118023, 0.07199299,
  0.07747311, 1.106547e-05, 0.005000594, 0.05955567, 0.0372266, 0.0562629, 
    0.04497733, 0.1026253, 0.02389356, 0.001702454, 0.001435655, 
    0.0002444777, 0.06176344, 0.0613634, 0.09138346, 0.07284728, 0.06785718, 
    0.07159635, 0.03745064, 0.02641402, 0.04542907, 0.0968295, 0.0709582, 
    0.0001159747, 0.03779997, 0.1337963, 0.06087656, 0.04944893, 0.1114624,
  0.002769695, 0.01756424, 0.0539034, 0.07508152, 0.0241417, 0.03859161, 
    0.05399344, 0.03818993, 0.0433187, 0.02872252, 0.07828134, 0.07140712, 
    0.1176751, 0.03819538, 0.04371085, 0.03038132, 0.02380135, 0.02191759, 
    0.02106616, 0.03130154, 0.01498791, 0.02337606, 0.0004683153, 0.07234076, 
    0.1057391, 0.01304572, 0.05471135, 0.04022359, 0.03138422,
  0.04693865, 0.04242255, 0.01824043, 0.03230681, 0.01997421, 0.01639515, 
    0.01766415, 0.0184443, 0.05640225, 0.1770838, 0.04035877, 0.01928081, 
    0.04160754, 0.01835384, 0.02590488, 0.02148241, 0.01633442, 0.02351084, 
    0.03100059, 0.02590905, 0.04473565, 0.03153779, 0.0313822, 0.1391323, 
    0.1812333, 0.03512451, 0.08210796, 0.06239581, 0.05583489,
  0.0004298471, 6.021297e-05, 2.583219e-05, 0.01647118, 0.02096127, 
    0.04244429, 0.02541366, 0.011269, 0.02554672, 0.06431346, 0.04587549, 
    0.04662029, 0.03674738, 0.06693451, 0.05652555, 0.03898777, 0.09060508, 
    0.147274, 0.1224053, 0.07122885, 0.02972728, 0.02485707, 0.07503837, 
    0.09892184, 0.0543269, 0.01786591, 0.003477228, 7.012499e-07, 0.002963444,
  2.415111e-06, 8.087521e-07, 2.494034e-07, 0.0001194232, 0.001150271, 
    0.0005607267, 2.0121e-06, 7.138386e-05, 0.0001361562, 0.03737808, 
    0.05061403, 0.03485888, 0.0252904, 0.03019984, 0.03721177, 0.04450487, 
    0.0728452, 0.08998297, 0.05565432, 0.008323723, 2.762257e-07, 0.08285156, 
    0.1010794, 0.07292128, 0.05270885, 0.0741223, 0.08325858, 0.01327667, 
    3.58275e-06,
  9.333836e-05, 0.008268972, 0.02372118, 0.00744601, 0.04452277, 
    0.0001910735, -0.002535789, 0.01061161, 0.09713434, 0.3351379, 0.1856755, 
    0.2602742, 0.2073939, 0.1540148, 0.1395005, 0.1079543, 0.1606256, 
    0.1649213, 0.1481571, 0.06936679, 1.785649e-05, 0.1131865, 0.04758753, 
    0.1112574, 0.09259719, 0.1761045, 0.0909755, 0.09558625, 0.01511851,
  0.007118557, 0.02258075, 0.09390283, 0.1480685, 0.03428879, 0.00246735, 
    0.1508687, 0.004398873, -0.0001324315, 0.01087699, 0.06526014, 0.1195035, 
    0.1692796, 0.2192347, 0.2149122, 0.2649019, 0.2664774, 0.2511532, 
    0.2094159, 0.1540276, 0.02249411, 0.02020191, 0.2325601, 0.237959, 
    0.2338313, 0.1494496, 0.1789449, 0.1298311, 0.1711611,
  0.2248134, 0.2469894, 0.1796388, 0.1494469, 0.06949974, 0.08836477, 
    0.09411695, 0.235519, 0.03275252, 0.04269779, 0.107682, 0.2008186, 
    0.3805222, 0.3369663, 0.3864441, 0.2245406, 0.269236, 0.2822143, 
    0.1785468, 0.2403913, 0.0721809, 0.1237912, 0.1442577, 0.2731167, 
    0.3312726, 0.2651151, 0.3707098, 0.3048729, 0.2677487,
  0.2593898, 0.2955227, 0.2625618, 0.2387281, 0.2509707, 0.1690442, 
    0.0492883, 0.08766255, 0.2453675, 0.1614926, 0.06166648, 0.1613665, 
    0.3968471, 0.3454547, 0.3202086, 0.2444195, 0.3145058, 0.333683, 
    0.2235975, 0.08587121, 0.1717458, 0.1946229, 0.1379553, 0.1951484, 
    0.3754242, 0.2708048, 0.2201812, 0.2635484, 0.253443,
  0.3128164, 0.1758321, 0.200014, 0.198339, 0.2256141, 0.04386944, 
    0.02128415, 0.117493, 0.1796043, 0.1287933, 0.1192266, 0.1723527, 
    0.1129783, 0.1101296, 0.1708131, 0.07366621, 0.08865739, 0.1702435, 
    0.1958769, 0.1723511, 0.2244028, 0.08310352, 0.2010981, 0.1521638, 
    0.1678053, 0.3412074, 0.1544182, 0.3088399, 0.359232,
  0.3300809, 0.349151, 0.2990876, 0.2450792, 0.1788821, 0.1145417, 0.1263641, 
    0.1019452, 0.05162209, 0.1291299, 0.1606461, 0.233765, 0.2313426, 
    0.2164184, 0.2020198, 0.2212877, 0.2204186, 0.1500511, 0.2225678, 
    0.3036979, 0.2927701, 0.2852561, 0.2238157, 0.1645195, 0.1532342, 
    0.1315727, 0.1389146, 0.1809932, 0.288963,
  0.3471834, 0.348908, 0.3506327, 0.3523573, 0.3540819, 0.3558066, 0.3575312, 
    0.378454, 0.3931156, 0.4077773, 0.422439, 0.4371007, 0.4517624, 
    0.4664241, 0.474622, 0.4748942, 0.4751664, 0.4754387, 0.4757109, 
    0.4759831, 0.4762553, 0.4683029, 0.4516444, 0.4349859, 0.4183273, 
    0.4016688, 0.3850103, 0.3683517, 0.3458037,
  0.5693925, 0.5608546, 0.4706399, 0.1669296, 0.09277254, 0.1198408, 
    0.1312543, 0.08887268, 0.01142782, 0.02870624, 0.1706661, 0.2208254, 
    0.2955889, 0.09088869, 0.2025909, 0.1107021, 0.2246828, 0.28951, 
    0.2338106, 0.3709175, 0.621072, 0.6517121, 0.3900177, 0.2615368, 
    0.2681248, 0.324702, 0.3246202, 0.301428, 0.4890436,
  0.4648865, 0.4269652, 0.404251, 0.2941037, 0.2756695, 0.1526049, 0.301145, 
    0.3793885, 0.3150566, 0.3044678, 0.1935268, 0.1106295, 0.1620469, 
    0.3487433, 0.4370874, 0.4155684, 0.3991629, 0.4511695, 0.6069814, 
    0.5227067, 0.5416932, 0.5494766, 0.495382, 0.426005, 0.3967694, 0.251329, 
    0.2789904, 0.3864241, 0.4644841,
  0.4124039, 0.3200386, 0.3719275, 0.3812131, 0.3357616, 0.4153531, 
    0.3794311, 0.4010366, 0.4724759, 0.3671384, 0.3101779, 0.3603545, 
    0.4371967, 0.401212, 0.3167206, 0.3368163, 0.322723, 0.350666, 0.3806558, 
    0.3601436, 0.339816, 0.3677263, 0.4126244, 0.3197759, 0.4965564, 
    0.4270324, 0.4498451, 0.4186094, 0.3862968,
  0.3473135, 0.358568, 0.3356568, 0.2553719, 0.2964864, 0.2862859, 0.3207812, 
    0.2752461, 0.3255048, 0.3398152, 0.3000726, 0.3181809, 0.238461, 
    0.2623547, 0.2163959, 0.2605205, 0.2517634, 0.2981952, 0.2857231, 
    0.3681575, 0.3724052, 0.3879451, 0.3356517, 0.1686216, 0.1651242, 
    0.2567869, 0.2880627, 0.4098249, 0.326611,
  0.1965362, 0.2297022, 0.1512962, 0.2601781, 0.2345537, 0.2681704, 
    0.2789858, 0.2968476, 0.2218699, 0.2740804, 0.14339, 0.1152364, 
    0.06782427, 0.2105843, 0.2542672, 0.2426391, 0.225915, 0.2983758, 
    0.2305855, 0.2729146, 0.2534757, 0.1842265, 0.1936191, 0.1607435, 
    0.05988229, 0.1364746, 0.1117801, 0.1712048, 0.2523026,
  0.1553848, 0.04682474, 0.0263728, 0.160553, 0.1084122, 0.1206284, 
    0.1948804, 0.1229831, 0.1758357, 0.04132599, 0.02432233, -5.059228e-06, 
    -0.002227372, 0.07956808, 0.04131804, 0.1150454, 0.1232733, 0.155446, 
    0.1548022, 0.07908718, 0.1589148, 0.1257509, 0.1035995, 0.006909608, 
    0.08966, 0.1426289, 0.1244653, 0.112813, 0.1170229,
  0.1440536, -8.360719e-05, 0.003173824, 0.05634202, 0.05713417, 0.06225748, 
    0.0610708, 0.1183335, 0.04586462, 0.01403101, 0.000461248, 0.0001298769, 
    0.07720915, 0.06683889, 0.0905128, 0.07943309, 0.06123172, 0.06746715, 
    0.06950264, 0.0351811, 0.05591349, 0.1348042, 0.2886128, 0.0003094901, 
    0.04589744, 0.104495, 0.06645831, 0.05465473, 0.172405,
  0.02302519, 0.01668715, 0.01785836, 0.1034549, 0.02851354, 0.04512978, 
    0.0543909, 0.04391248, 0.04112966, 0.02929912, 0.06937367, 0.07394297, 
    0.1043658, 0.03756402, 0.04604899, 0.03445396, 0.03756703, 0.03641804, 
    0.03621233, 0.05128085, 0.0584112, 0.124658, 0.01824487, 0.0645612, 
    0.09503578, 0.004046554, 0.07678851, 0.08200491, 0.1121994,
  0.05387935, 0.02823154, 0.01416296, 0.02604027, 0.02722269, 0.02744014, 
    0.03177835, 0.02555021, 0.06830798, 0.185405, 0.04526849, 0.02630481, 
    0.04322128, 0.02129041, 0.02875654, 0.02706685, 0.01723133, 0.02429308, 
    0.0359646, 0.0278965, 0.0371455, 0.0304429, 0.0221159, 0.1287275, 
    0.158853, 0.03762344, 0.07683863, 0.05591867, 0.05953567,
  0.0002508613, 2.425917e-05, 3.913134e-06, 0.007563326, 0.01985396, 
    0.1122584, 0.03925215, 0.03498772, 0.03334109, 0.09096635, 0.06721982, 
    0.05016796, 0.03870286, 0.0669304, 0.05187515, 0.04535712, 0.1028092, 
    0.1916901, 0.1386727, 0.0757967, 0.03925573, 0.06064088, 0.07361613, 
    0.09910785, 0.06402614, 0.08596347, 0.0279789, 1.051653e-05, 0.001817493,
  1.409986e-06, 4.706775e-07, 1.271398e-07, 0.0001742778, 0.0004423805, 
    0.001163079, 3.876456e-07, 3.147665e-05, 6.289992e-05, 0.05747607, 
    0.08208057, 0.04506343, 0.04466133, 0.04667002, 0.05496229, 0.05733902, 
    0.05771401, 0.0940792, 0.1541321, 0.03970457, 7.500944e-07, 0.1003696, 
    0.05251365, 0.07400924, 0.1135042, 0.09908979, 0.07075166, 0.03716126, 
    2.360474e-06,
  -6.524708e-06, 0.02553051, 0.02227176, 0.005997111, 0.03700772, 
    3.045412e-05, -0.00215706, 0.004172032, 0.08075204, 0.3419419, 0.2055964, 
    0.2699791, 0.2508491, 0.1921537, 0.2270945, 0.2374343, 0.2303292, 
    0.1803621, 0.2278834, 0.1540074, 8.876234e-06, 0.1151868, 0.0402389, 
    0.0944005, 0.09799415, 0.140507, 0.1074347, 0.08056632, 0.0163564,
  0.008490562, 0.01110318, 0.08138211, 0.134296, 0.03024145, 0.0004975611, 
    0.1538508, 0.002821974, -9.984944e-05, 0.01021867, 0.0622534, 0.1127737, 
    0.1528518, 0.191087, 0.200685, 0.2568619, 0.2484259, 0.3031121, 0.247723, 
    0.1565759, 0.01892154, 0.02591904, 0.242333, 0.2197669, 0.244384, 
    0.1612859, 0.2092858, 0.2152723, 0.1692015,
  0.1955034, 0.2137724, 0.1619932, 0.1762884, 0.04316091, 0.0891733, 
    0.09118964, 0.233325, 0.02455543, 0.03104235, 0.1036277, 0.1907409, 
    0.3971259, 0.332463, 0.3119179, 0.1859011, 0.2795279, 0.2921072, 
    0.2724599, 0.2393975, 0.06788387, 0.1238404, 0.1784324, 0.2865675, 
    0.3525181, 0.4212941, 0.3525454, 0.208755, 0.2613523,
  0.2440819, 0.2756445, 0.2435272, 0.2210732, 0.2010783, 0.1351198, 
    0.06366967, 0.1048733, 0.1348161, 0.0752859, 0.04194191, 0.1320915, 
    0.3327439, 0.33569, 0.4037957, 0.2681006, 0.3379218, 0.3493082, 
    0.2514795, 0.0517379, 0.1738527, 0.1808291, 0.1736154, 0.2312818, 
    0.4996634, 0.1839704, 0.2406567, 0.3142215, 0.2645036,
  0.3130127, 0.2244792, 0.2161088, 0.2507469, 0.1812102, 0.0422856, 
    0.03735284, 0.08852302, 0.2319658, 0.1582626, 0.122972, 0.2376002, 
    0.1180075, 0.1161808, 0.1841183, 0.06782755, 0.08283464, 0.1616958, 
    0.1944563, 0.178169, 0.187369, 0.07667103, 0.2151267, 0.1458591, 
    0.1336384, 0.3574693, 0.1417942, 0.2693658, 0.4158732,
  0.3221321, 0.4440823, 0.2942811, 0.2534737, 0.2105801, 0.1323939, 
    0.1520561, 0.09078053, 0.05702674, 0.1697875, 0.1993188, 0.2734157, 
    0.2878298, 0.269962, 0.2393553, 0.2739284, 0.2521797, 0.2128823, 
    0.3299905, 0.3631679, 0.278115, 0.2801409, 0.2042626, 0.1906956, 
    0.1519344, 0.1269599, 0.1125579, 0.2071961, 0.3529726,
  0.3724307, 0.3750005, 0.3775703, 0.38014, 0.3827098, 0.3852796, 0.3878493, 
    0.41316, 0.4284772, 0.4437945, 0.4591117, 0.474429, 0.4897462, 0.5050635, 
    0.5318683, 0.5308102, 0.5297521, 0.528694, 0.5276359, 0.5265778, 
    0.5255197, 0.4870991, 0.4702702, 0.4534413, 0.4366124, 0.4197835, 
    0.4029545, 0.3861256, 0.3703749,
  0.5662165, 0.5662276, 0.4790339, 0.2348443, 0.1309006, 0.1517714, 
    0.1488106, 0.1062872, 0.016646, 0.04534533, 0.2027789, 0.2667472, 
    0.3075009, 0.04166638, 0.2001164, 0.1314519, 0.1948223, 0.3172575, 
    0.2423796, 0.3593377, 0.6427475, 0.6990807, 0.4008445, 0.267877, 
    0.2693143, 0.3717885, 0.3404381, 0.2827556, 0.5024597,
  0.3789795, 0.3520156, 0.3960967, 0.2577792, 0.2836628, 0.1440327, 
    0.1988752, 0.4059387, 0.3038955, 0.3038404, 0.1842571, 0.1133279, 
    0.1630651, 0.3095369, 0.3902486, 0.456431, 0.4432085, 0.5035564, 
    0.5934067, 0.5888906, 0.6084205, 0.5615901, 0.5012516, 0.4745071, 
    0.4080073, 0.2348986, 0.3240828, 0.4188572, 0.4502113,
  0.4516222, 0.3646456, 0.3496361, 0.381172, 0.3281594, 0.4435076, 0.4078042, 
    0.371379, 0.4224533, 0.3398765, 0.2930687, 0.403233, 0.4401041, 
    0.3821638, 0.351216, 0.3636177, 0.3829612, 0.3811933, 0.3698268, 
    0.3295476, 0.3677711, 0.3623381, 0.3938096, 0.3026938, 0.4773696, 
    0.4152974, 0.4416863, 0.3980022, 0.39878,
  0.3731249, 0.3703199, 0.4028799, 0.295427, 0.2968039, 0.3658464, 0.3399584, 
    0.3155086, 0.3421406, 0.3667673, 0.3095283, 0.2866869, 0.2122512, 
    0.2185677, 0.253744, 0.2194277, 0.2816324, 0.3375404, 0.3204565, 
    0.3955171, 0.378221, 0.3320785, 0.2814819, 0.1760431, 0.1202006, 
    0.2377058, 0.2774002, 0.3841198, 0.3742442,
  0.2846537, 0.3381273, 0.1394604, 0.2564531, 0.2990438, 0.2343508, 
    0.2353977, 0.2134777, 0.2227357, 0.2207777, 0.1366472, 0.08609958, 
    0.03395367, 0.1294264, 0.2846819, 0.2214048, 0.2126661, 0.3034123, 
    0.2267212, 0.2590183, 0.1843321, 0.1891554, 0.2131441, 0.1837399, 
    0.04867579, 0.1145605, 0.118727, 0.1620324, 0.2683931,
  0.1973382, 0.1375811, 0.02311085, 0.1143223, 0.1396098, 0.09010912, 
    0.1794518, 0.1765974, 0.2412692, 0.03046621, 0.06666898, -2.334163e-05, 
    -0.00426064, 0.0585146, 0.06932436, 0.1448495, 0.08509777, 0.1126347, 
    0.1286083, 0.08501814, 0.1327197, 0.09919503, 0.1246032, 0.01291861, 
    0.105402, 0.1424512, 0.1190824, 0.1097554, 0.1370049,
  0.3176119, -0.0004214969, 0.001073611, 0.07245685, 0.09947364, 0.07708581, 
    0.09542635, 0.1130227, 0.05822473, 0.002654211, 0.0001496215, 
    5.614283e-05, 0.02403321, 0.04618429, 0.08436199, 0.1117956, 0.08675674, 
    0.08654228, 0.06661215, 0.07858538, 0.09533652, 0.07836875, 0.3534154, 
    0.0001970885, 0.05162141, 0.1038978, 0.1326136, 0.05154856, 0.1015349,
  0.317014, 0.01770307, 0.006997305, 0.07060116, 0.07234577, 0.05197684, 
    0.06292611, 0.05708584, 0.04741336, 0.0403276, 0.0624442, 0.0733036, 
    0.1169303, 0.09997032, 0.05815095, 0.05637307, 0.04860985, 0.08733612, 
    0.1252048, 0.1516135, 0.1659391, 0.1529021, 0.2729204, 0.04318876, 
    0.05277951, 0.0007203787, 0.08957091, 0.08552132, 0.156872,
  0.05717785, 0.02187245, 0.006976508, 0.04088987, 0.06453183, 0.2144472, 
    0.1896081, 0.1987283, 0.05078093, 0.1192978, 0.09457516, 0.1322133, 
    0.05305059, 0.02920059, 0.04595156, 0.07534239, 0.04504935, 0.0323827, 
    0.08710404, 0.04081861, 0.03600166, 0.04472423, 0.01789804, 0.1090504, 
    0.1128642, 0.05062666, 0.08586852, 0.05533711, 0.06444091,
  0.0001989073, 4.559624e-06, 1.3544e-06, 0.002476928, 0.0323393, 0.1919734, 
    0.09256149, 0.2170237, 0.06180506, 0.1862409, 0.09032524, 0.0792657, 
    0.05262929, 0.06787197, 0.04622287, 0.05301592, 0.1022794, 0.176009, 
    0.1586202, 0.1198539, 0.07434692, 0.1023933, 0.1213066, 0.09863786, 
    0.09366447, 0.2613336, 0.3334871, 0.000778252, 0.0005077688,
  8.30524e-07, 3.173168e-07, 7.075873e-08, 0.0003386264, 0.0001905765, 
    0.007948067, 3.908817e-07, -0.0003539108, 2.709474e-05, 0.1060658, 
    0.1021719, 0.07140506, 0.06033681, 0.04317632, 0.03433959, 0.04900278, 
    0.09006803, 0.07905206, 0.2133425, 0.2348242, -1.884968e-06, 0.09700029, 
    0.04166171, 0.05235035, 0.05593168, 0.1006753, 0.1837709, 0.170997, 
    1.275864e-06,
  -1.310298e-05, 0.02742616, 0.0172706, 0.005061412, 0.03190465, 
    -3.341888e-05, -0.001787204, 7.386979e-05, 0.082189, 0.3430145, 
    0.2192133, 0.2654265, 0.300424, 0.2560713, 0.3043999, 0.2183522, 
    0.2998734, 0.1754231, 0.2747001, 0.1331453, 4.723353e-06, 0.1242116, 
    0.03332502, 0.09190248, 0.07307492, 0.1023214, 0.1076414, 0.06218389, 
    0.01953906,
  0.009691822, 0.010608, 0.06929008, 0.1321066, 0.03202294, 0.0003121316, 
    0.1516126, 0.002535321, -7.261486e-05, 0.007453125, 0.06157098, 
    0.1119673, 0.1315151, 0.1582149, 0.1836011, 0.2747558, 0.2964782, 
    0.2548565, 0.2531397, 0.1469678, 0.01401902, 0.02196285, 0.2009498, 
    0.2332365, 0.294888, 0.2246143, 0.1964485, 0.3039392, 0.1643789,
  0.2123765, 0.1837107, 0.09794684, 0.1625761, 0.03723489, 0.07981001, 
    0.1062762, 0.2103818, 0.01706729, 0.03051259, 0.08578009, 0.1861015, 
    0.4014577, 0.3624331, 0.2694627, 0.159142, 0.2685356, 0.2980791, 
    0.2787296, 0.2329977, 0.06668641, 0.1246832, 0.1704901, 0.2994835, 
    0.324778, 0.3494404, 0.3108742, 0.1299582, 0.2440324,
  0.216642, 0.2167842, 0.2438636, 0.1999422, 0.2078322, 0.1152754, 0.0880315, 
    0.1034324, 0.09411968, 0.03423332, 0.02181515, 0.07310728, 0.2822155, 
    0.2698647, 0.5852088, 0.3545682, 0.3577961, 0.3395077, 0.3114327, 
    0.04267612, 0.1803796, 0.1791877, 0.1452834, 0.2127776, 0.577027, 
    0.1514524, 0.1741335, 0.2770357, 0.2162563,
  0.3642725, 0.182029, 0.2116583, 0.2515882, 0.1640778, 0.04459452, 
    0.04208131, 0.1489265, 0.225313, 0.2131527, 0.1471232, 0.2578838, 
    0.1814655, 0.1444393, 0.17403, 0.0806298, 0.07308971, 0.1629711, 
    0.152511, 0.1827571, 0.1819112, 0.09548671, 0.2162226, 0.1456743, 
    0.1076438, 0.3559638, 0.141572, 0.2132404, 0.4098287,
  0.3117957, 0.4044545, 0.2728188, 0.2236578, 0.1934696, 0.141996, 0.169734, 
    0.06888378, 0.07237775, 0.1891696, 0.2185399, 0.2924055, 0.3039023, 
    0.3196349, 0.3447287, 0.3355916, 0.2909009, 0.2630728, 0.3107047, 
    0.3399584, 0.2935647, 0.2753002, 0.2278095, 0.220869, 0.1550205, 
    0.1369125, 0.1054275, 0.2068316, 0.3267946,
  0.400697, 0.4055333, 0.4103696, 0.4152059, 0.4200422, 0.4248785, 0.4297149, 
    0.4753662, 0.4882526, 0.5011389, 0.5140252, 0.5269115, 0.5397978, 
    0.5526841, 0.5704615, 0.5648255, 0.5591894, 0.5535535, 0.5479175, 
    0.5422814, 0.5366455, 0.4737275, 0.4616409, 0.4495542, 0.4374676, 
    0.425381, 0.4132943, 0.4012077, 0.3968279,
  0.5854999, 0.590511, 0.5116244, 0.2670159, 0.1652751, 0.1600591, 0.1585655, 
    0.1197709, 0.02356232, 0.05592716, 0.2384969, 0.3189031, 0.3778411, 
    0.01979633, 0.1472318, 0.1831571, 0.2102417, 0.2928362, 0.2228798, 
    0.3592697, 0.6999745, 0.7352333, 0.3870534, 0.2675512, 0.237005, 
    0.3859385, 0.360519, 0.294137, 0.5537022,
  0.3059804, 0.2592359, 0.3643665, 0.2135236, 0.2737982, 0.1400495, 
    0.1399567, 0.3935828, 0.289658, 0.2999572, 0.1678215, 0.1088462, 
    0.1519121, 0.2457511, 0.3619898, 0.5542757, 0.3925484, 0.4628535, 
    0.5334187, 0.5967301, 0.5637803, 0.5300074, 0.5296947, 0.4602857, 
    0.4168006, 0.2456345, 0.2950379, 0.3737166, 0.4537948,
  0.4675535, 0.337883, 0.3327096, 0.3920953, 0.3365681, 0.4145658, 0.4002344, 
    0.3455261, 0.3679758, 0.3012212, 0.2851698, 0.372674, 0.4480841, 
    0.3655551, 0.3591886, 0.392873, 0.3949856, 0.4019602, 0.3832594, 
    0.3590398, 0.3582488, 0.3746502, 0.3658597, 0.272159, 0.4375901, 
    0.3552805, 0.4560367, 0.3713041, 0.3962772,
  0.3607172, 0.3892066, 0.3956989, 0.3309072, 0.3279077, 0.4120106, 
    0.3296544, 0.3042712, 0.3266368, 0.3339997, 0.2892686, 0.2488516, 
    0.1471737, 0.2373609, 0.2413854, 0.1745829, 0.249154, 0.3275919, 
    0.3591386, 0.3883862, 0.3019151, 0.2515139, 0.2637918, 0.170924, 
    0.09893485, 0.2287444, 0.2551698, 0.3412284, 0.4115556,
  0.217857, 0.2520027, 0.08997001, 0.1908588, 0.2246656, 0.1725495, 
    0.2126976, 0.1748813, 0.219587, 0.143868, 0.06943096, 0.05198759, 
    0.02275859, 0.07879571, 0.3118803, 0.1985815, 0.1849752, 0.2384146, 
    0.1838622, 0.2035818, 0.1189448, 0.1219116, 0.1472191, 0.1945773, 
    0.05451363, 0.1330153, 0.08276772, 0.1661268, 0.3076799,
  0.1427665, 0.124963, 0.01691188, 0.1363313, 0.08941333, 0.06462423, 
    0.1404291, 0.1287372, 0.1322345, 0.01543435, 0.05627895, -7.519507e-05, 
    -0.002593558, 0.01955467, 0.02038228, 0.1107685, 0.0970196, 0.133606, 
    0.08753663, 0.05146681, 0.06969143, 0.05044935, 0.07822301, 0.02113122, 
    0.0873004, 0.1175153, 0.06148765, 0.07216721, 0.08521277,
  0.1701481, -0.0003523872, 0.0003069143, 0.09793316, 0.07248507, 0.04783413, 
    0.04516511, 0.09373915, 0.05940311, 0.005137687, 5.327752e-05, 
    2.18418e-05, 0.007652255, 0.02244187, 0.06047299, 0.05765992, 0.07085539, 
    0.03519338, 0.02724013, 0.08840719, 0.01455642, 0.05936561, 0.1451677, 
    0.07931641, 0.04878731, 0.1093706, 0.035166, 0.01612755, 0.04079447,
  0.4314995, 0.06621658, 0.002199772, 0.06985973, 0.1679877, 0.04635907, 
    0.06711365, 0.07773837, 0.05388958, 0.02492272, 0.04949196, 0.03562891, 
    0.09824371, 0.06505494, 0.07050541, 0.02502935, 0.02357233, 0.05758641, 
    0.05031402, 0.03511658, 0.04204499, 0.05059019, 0.3819516, 0.03114313, 
    0.02715198, 0.0001274633, 0.01738469, 0.01852473, 0.08730973,
  0.08757304, 0.01818103, 0.001832175, 0.03953791, 0.02045881, 0.04112485, 
    0.05184079, 0.03760494, 0.07376977, 0.06426563, 0.031256, 0.05832285, 
    0.03317708, 0.03201634, 0.04837864, 0.09438933, 0.08053201, 0.07834103, 
    0.05222226, 0.07413512, 0.04541832, 0.2213066, 0.03340686, 0.0802607, 
    0.07756377, 0.03261549, 0.09881094, 0.07376293, 0.101316,
  0.0001567966, -7.640172e-07, 9.350643e-07, -0.001268749, 0.02979789, 
    0.07308087, 0.0819289, 0.1061134, 0.02119794, 0.08848146, 0.03324798, 
    0.05584235, 0.04780196, 0.05029591, 0.02231862, 0.0236879, 0.0631587, 
    0.1100975, 0.1292721, 0.1168853, 0.03764762, 0.01406642, 0.2408205, 
    0.09944032, 0.05035609, 0.07236289, 0.3210713, 0.08253906, 0.0001385507,
  5.534122e-07, 2.488196e-07, 4.958748e-08, 0.0008211631, 0.0001168658, 
    0.01539435, -9.735459e-07, 0.01551934, 4.5193e-05, 0.1876625, 0.1945386, 
    0.05760373, 0.03038929, 0.02015226, 0.01205637, 0.01088176, 0.02768216, 
    0.04860171, 0.2302599, 0.2227067, -7.367014e-05, 0.08936537, 0.01599666, 
    0.02429328, 0.01190851, 0.05389709, 0.134256, 0.1043563, 7.430194e-07,
  4.052784e-06, 0.01965279, 0.01957708, 0.004112773, 0.02850824, 
    -3.075067e-05, -0.001482574, -0.0002949706, 0.0846331, 0.3252893, 
    0.2304896, 0.2618116, 0.3229286, 0.3038781, 0.1768573, 0.1570403, 
    0.2749575, 0.1000776, 0.2326223, 0.1452288, 2.66179e-06, 0.1429707, 
    0.02203362, 0.07687893, 0.09027898, 0.08504483, 0.0750275, 0.04156176, 
    0.02190439,
  0.007730834, 0.006407435, 0.06251296, 0.1434935, 0.03701556, 6.531338e-05, 
    0.1426307, 0.002722902, -6.077571e-05, 0.004307389, 0.0579159, 
    0.09903172, 0.123942, 0.1499536, 0.1390672, 0.233862, 0.316817, 
    0.2028498, 0.3406034, 0.1372167, 0.01085394, 0.013575, 0.1857987, 
    0.2823642, 0.3094236, 0.1726882, 0.160521, 0.2070392, 0.1548368,
  0.1746296, 0.1613345, 0.07167234, 0.1330726, 0.02842936, 0.0603516, 
    0.08678138, 0.1899546, 0.01504566, 0.03267377, 0.071427, 0.1842504, 
    0.3339144, 0.352386, 0.2225513, 0.1341293, 0.2943532, 0.2813012, 
    0.290199, 0.220949, 0.06675772, 0.09455853, 0.1379816, 0.2841851, 
    0.3127123, 0.2884257, 0.2730693, 0.0875689, 0.2031229,
  0.1516172, 0.2018142, 0.2427112, 0.191995, 0.198905, 0.116993, 0.1122914, 
    0.104035, 0.07027755, 0.02030948, 0.009669647, 0.03152475, 0.2146081, 
    0.1710567, 0.5324667, 0.4719647, 0.3618481, 0.3233139, 0.2589491, 
    0.05130353, 0.1839993, 0.2090151, 0.122473, 0.1856467, 0.5045471, 
    0.140588, 0.1299166, 0.1770928, 0.1330546,
  0.3156311, 0.1566968, 0.2657332, 0.2590777, 0.1499677, 0.03177695, 
    0.06056502, 0.1338013, 0.2056106, 0.2067479, 0.1482979, 0.2417878, 
    0.2244398, 0.1354438, 0.1773484, 0.1075054, 0.08739701, 0.1357647, 
    0.1945055, 0.1714389, 0.1927269, 0.1175422, 0.2093608, 0.142561, 
    0.09477037, 0.3627465, 0.1577344, 0.1609404, 0.3750496,
  0.3282431, 0.3480545, 0.2572994, 0.2137221, 0.2832974, 0.1882038, 
    0.1715876, 0.09300348, 0.1158173, 0.2100458, 0.3008223, 0.3299985, 
    0.3119141, 0.3647925, 0.4406454, 0.430931, 0.3433463, 0.2605776, 
    0.3007306, 0.375489, 0.3671924, 0.2723759, 0.2570975, 0.2835666, 
    0.1429419, 0.167835, 0.1223161, 0.1812262, 0.2901868,
  0.3868661, 0.3872755, 0.3876849, 0.3880943, 0.3885037, 0.3889131, 
    0.3893225, 0.4190341, 0.4321283, 0.4452226, 0.4583168, 0.471411, 
    0.4845053, 0.4975995, 0.5198265, 0.514377, 0.5089276, 0.5034781, 
    0.4980287, 0.4925792, 0.4871297, 0.4624291, 0.4543749, 0.4463207, 
    0.4382665, 0.4302123, 0.4221582, 0.414104, 0.3865386,
  0.5967954, 0.6180573, 0.5310461, 0.2824039, 0.1697249, 0.1667415, 
    0.1608173, 0.1238863, 0.01014222, 0.01467532, 0.2137813, 0.3536927, 
    0.4575853, 0.006450993, 0.127845, 0.2430119, 0.2720586, 0.287132, 
    0.2144484, 0.3691599, 0.7285258, 0.7646494, 0.3496532, 0.2467545, 
    0.2116727, 0.3863384, 0.3848662, 0.2787372, 0.6278208,
  0.2289199, 0.176787, 0.3305393, 0.1566954, 0.251713, 0.1417732, 0.09419365, 
    0.3652483, 0.2776855, 0.2711659, 0.1397203, 0.1173565, 0.1435534, 
    0.1967875, 0.3505678, 0.5160266, 0.3881235, 0.3902878, 0.4498214, 
    0.5061392, 0.4686661, 0.5279044, 0.511032, 0.4361054, 0.4064237, 
    0.2980188, 0.260257, 0.3089873, 0.3893101,
  0.4074221, 0.3090163, 0.3163529, 0.3648553, 0.3442417, 0.3553786, 
    0.3671269, 0.3139696, 0.3211505, 0.2588829, 0.2425383, 0.2983813, 
    0.4458742, 0.3528943, 0.3417213, 0.4025105, 0.3583047, 0.4052334, 
    0.4205056, 0.3573782, 0.311864, 0.3430329, 0.3202172, 0.2413907, 
    0.3732771, 0.3383733, 0.4373731, 0.3453569, 0.3670828,
  0.3702493, 0.4341972, 0.4038587, 0.3422149, 0.3668472, 0.4148256, 
    0.3115617, 0.247331, 0.280596, 0.2805841, 0.2547733, 0.2224709, 
    0.1436843, 0.2518852, 0.205504, 0.1641335, 0.2242413, 0.3684448, 
    0.3449963, 0.3554994, 0.262863, 0.215493, 0.2472245, 0.1502587, 
    0.07623211, 0.2169502, 0.2400758, 0.3317387, 0.3703287,
  0.1822146, 0.1399787, 0.08479806, 0.1393601, 0.1723253, 0.1326545, 
    0.1554665, 0.1671955, 0.1636291, 0.08977579, 0.04097634, 0.03171604, 
    0.006900489, 0.04349794, 0.3012375, 0.1951784, 0.1704552, 0.2066281, 
    0.1276903, 0.168195, 0.1034916, 0.06462875, 0.08896616, 0.1975673, 
    0.04304462, 0.1034649, 0.05116035, 0.1616241, 0.2742196,
  0.06414787, 0.07547474, 0.01093837, 0.04528914, 0.06167715, 0.03118066, 
    0.1170709, 0.07317582, 0.04330744, 0.005416066, 0.02965837, 
    -4.055192e-05, -2.198729e-05, 0.005714761, 0.01002105, 0.09761872, 
    0.04708151, 0.09264783, 0.06429154, 0.02056901, 0.05516566, 0.03455295, 
    0.02785426, 0.07016915, 0.07398061, 0.06616231, 0.03998451, 0.04365405, 
    0.02112217,
  0.1611694, -0.000177389, -3.299703e-06, 0.01760111, 0.01136887, 0.01516325, 
    0.01795247, 0.0545079, 0.01918618, 0.0003206765, 1.363951e-05, 
    6.028959e-06, 0.002780989, 0.008685705, 0.02633682, 0.02961403, 
    0.01790732, 0.01239316, 0.004247406, 0.01205016, 0.002532594, 0.01445989, 
    0.04697301, 0.1604489, 0.04717894, 0.09381983, 0.01432083, 0.001664261, 
    0.006989348,
  0.1717023, 0.06287311, 0.0003296088, 0.07950007, 0.02199456, 0.01290323, 
    0.0200483, 0.01773127, 0.02098137, 0.005697724, 0.04353537, 0.01380284, 
    0.05337871, 0.01729088, 0.02684998, 0.01192585, 0.003496038, 0.006450906, 
    0.01005772, 0.007290734, 0.0114353, 0.01201253, 0.119004, 0.01051418, 
    0.02024526, 5.386734e-05, -0.002729719, 0.004102722, 0.02840969,
  0.03696312, 0.01241999, 0.000687615, 0.03980977, 0.002763855, 0.00827192, 
    0.00958446, 0.007726877, 0.05567588, 0.03671801, 0.008569302, 
    0.008496485, 0.01808728, 0.007844293, 0.01171349, 0.01424715, 0.06881495, 
    0.06026355, 0.01657922, 0.04026143, 0.04628354, 0.1061231, 0.3326052, 
    0.06753087, 0.06166659, 0.01323187, 0.07279742, 0.03360272, 0.03447343,
  8.80271e-05, -1.208738e-06, 2.071996e-07, -0.002155392, 0.02578187, 
    0.01872027, 0.03331771, 0.02115575, 0.003781002, 0.02362042, 0.009429418, 
    0.009524378, 0.01930042, 0.02823911, 0.006715273, 0.006294591, 
    0.03626708, 0.0391387, 0.07032731, 0.03833904, 0.006591364, 0.002360299, 
    0.2746719, 0.09938236, 0.01462729, 0.01873719, 0.09273128, 0.1914459, 
    0.0001624051,
  4.311964e-07, 2.191132e-07, 3.784782e-08, 0.001561047, 0.0001117786, 
    0.01106387, -4.211149e-06, 0.005087048, 3.233287e-05, 0.2135565, 
    0.1217864, 0.01970358, 0.008671671, 0.004266018, 0.001062171, 
    0.001695534, 0.009532349, 0.02404126, 0.1212122, 0.0874887, 
    -1.906854e-05, 0.07577346, 0.005316191, 0.01155689, 0.005172541, 
    0.03699859, 0.03341366, 0.08233958, 4.800048e-07,
  -2.901185e-07, 0.01469016, 0.0229373, 0.004168265, 0.02448569, 
    -1.447304e-05, -0.001349217, -0.0006798996, 0.07853522, 0.3075356, 
    0.2431261, 0.2602131, 0.287953, 0.2829112, 0.1282658, 0.1519827, 
    0.1579218, 0.04391523, 0.1224147, 0.1200243, 1.74153e-06, 0.1396936, 
    0.01431565, 0.0496491, 0.04758791, 0.05483904, 0.03443964, 0.05409665, 
    0.02572285,
  0.004446277, 0.003267981, 0.04641763, 0.1781527, 0.03476167, -0.0001373461, 
    0.1353117, 0.004225449, -5.62688e-05, 0.002774441, 0.05386966, 
    0.08648805, 0.1502648, 0.1650245, 0.1226975, 0.2041814, 0.3001245, 
    0.1875741, 0.2754476, 0.135907, 0.009022516, 0.008189421, 0.1604919, 
    0.2893119, 0.2478094, 0.1135976, 0.09969614, 0.1045627, 0.1424921,
  0.1411476, 0.1330907, 0.07191851, 0.1072254, 0.02207168, 0.0501966, 
    0.06768364, 0.1615039, 0.01236608, 0.03557051, 0.06212122, 0.1755666, 
    0.2790059, 0.3165676, 0.1879417, 0.1088525, 0.2652026, 0.2679489, 
    0.2856475, 0.2208456, 0.06181019, 0.08007208, 0.1247541, 0.2422514, 
    0.2947213, 0.2933627, 0.2583452, 0.05705004, 0.1581446,
  0.1089734, 0.2041003, 0.2230698, 0.1734757, 0.2075204, 0.1079039, 
    0.1219481, 0.07988242, 0.05335139, 0.01465073, 0.004915211, 0.01105537, 
    0.1652008, 0.104496, 0.4046595, 0.5031984, 0.3394097, 0.2987782, 
    0.1779717, 0.06569092, 0.1705849, 0.1929061, 0.09522448, 0.1898334, 
    0.4179116, 0.1215488, 0.09907697, 0.1165448, 0.08667009,
  0.2968509, 0.1235933, 0.2405951, 0.2280152, 0.1649937, 0.05913199, 
    0.08199187, 0.1161805, 0.1944635, 0.2398939, 0.1348296, 0.238066, 
    0.2493907, 0.1462275, 0.1915444, 0.1112064, 0.1680625, 0.1505328, 
    0.1711535, 0.1975786, 0.2686697, 0.1644871, 0.2092104, 0.1758138, 
    0.08862657, 0.3777854, 0.1650854, 0.1056501, 0.340614,
  0.390929, 0.3513135, 0.2517692, 0.3204469, 0.3598093, 0.2483601, 0.2030892, 
    0.1329232, 0.1428963, 0.2946134, 0.3383702, 0.3794249, 0.3561896, 
    0.4375744, 0.4748904, 0.5497696, 0.4489938, 0.3223063, 0.3340993, 
    0.4335345, 0.3960966, 0.2535414, 0.2730901, 0.3520049, 0.1365873, 
    0.1872544, 0.1183801, 0.1586302, 0.3404497,
  0.1366692, 0.1245681, 0.1124669, 0.1003658, 0.08826464, 0.07616349, 
    0.06406234, 0.07104716, 0.09480055, 0.1185539, 0.1423073, 0.1660607, 
    0.1898141, 0.2135675, 0.3255659, 0.3311469, 0.3367279, 0.3423089, 
    0.3478899, 0.3534709, 0.3590519, 0.3851615, 0.3679282, 0.350695, 
    0.3334618, 0.3162285, 0.2989953, 0.281762, 0.1463502,
  0.5546175, 0.570996, 0.4306986, 0.2299035, 0.1370795, 0.1426233, 0.1472208, 
    0.1187859, 0.02657329, 0.004948268, 0.07612416, 0.2867902, 0.4811784, 
    0.001547172, 0.1508587, 0.2951824, 0.3788588, 0.2929019, 0.1968152, 
    0.3992746, 0.7624702, 0.7756107, 0.2855538, 0.2051668, 0.2029014, 
    0.3850449, 0.4064744, 0.2393332, 0.5903586,
  0.1736684, 0.1190422, 0.3000989, 0.1001301, 0.2178648, 0.1403626, 
    0.05702235, 0.3223978, 0.2617425, 0.2380124, 0.1117204, 0.1142212, 
    0.1317277, 0.1629499, 0.3315916, 0.4603607, 0.3230395, 0.3216162, 
    0.385313, 0.4392726, 0.3875728, 0.5006415, 0.4555319, 0.4051873, 
    0.3997321, 0.3154796, 0.3084629, 0.2840196, 0.3187017,
  0.3187394, 0.2584738, 0.27225, 0.3221678, 0.298521, 0.2883441, 0.3110335, 
    0.2640362, 0.2662438, 0.2187718, 0.1914789, 0.2521136, 0.4381309, 
    0.3343888, 0.2997338, 0.3602115, 0.3156775, 0.4020303, 0.3984152, 
    0.3088577, 0.2743774, 0.2983578, 0.2628768, 0.2050739, 0.3358454, 
    0.3291436, 0.3873765, 0.324987, 0.3409856,
  0.3615403, 0.4401399, 0.403384, 0.3301967, 0.3707223, 0.3785949, 0.282047, 
    0.1960268, 0.2314362, 0.2325921, 0.2040654, 0.1888408, 0.1138698, 
    0.2134725, 0.1697264, 0.141245, 0.2085743, 0.3727507, 0.3145449, 
    0.309444, 0.2399811, 0.1874102, 0.2209503, 0.1241656, 0.04817369, 
    0.1772576, 0.2421707, 0.3192454, 0.3420644,
  0.1616755, 0.09200358, 0.04724497, 0.1028908, 0.1203526, 0.1023015, 
    0.1162665, 0.1609949, 0.09617139, 0.05370147, 0.02128406, 0.02476311, 
    0.002556219, 0.02851595, 0.2609049, 0.1490767, 0.1736949, 0.1673684, 
    0.08567503, 0.1416806, 0.08946995, 0.04048672, 0.044565, 0.2098301, 
    0.03168551, 0.05996075, 0.02689922, 0.126167, 0.2261585,
  0.02782258, 0.04722205, 0.006533794, 0.0170273, 0.02978262, 0.01148873, 
    0.07143939, 0.02931383, 0.01670202, 0.002326103, 0.01532704, 
    -7.708542e-06, 0.0002330241, 0.001722664, 0.04644332, 0.04247399, 
    0.03502364, 0.04682528, 0.02535732, 0.006290744, 0.03020918, 0.02356208, 
    0.008857417, 0.05605876, 0.06266613, 0.03457566, 0.02658189, 0.01539463, 
    0.006702613,
  0.0929727, 4.178124e-05, -7.893025e-05, 0.006447508, 0.0005831187, 
    0.004820013, 0.00590006, 0.02700291, 0.004986127, 7.683779e-05, 
    4.044172e-06, 2.332472e-06, 0.0007480511, 0.001913077, 0.01194676, 
    0.01051291, 0.003276068, 0.004637456, 0.001072779, 0.004176397, 
    0.0009267705, 0.005745237, 0.01675349, 0.08829287, 0.03611661, 
    0.07647216, 0.004835494, 0.0002748912, 0.00232629,
  0.06892417, 0.03181875, 0.0001805126, 0.06450556, 0.005684912, 0.003513375, 
    0.005009008, 0.003797613, 0.007802206, -0.0007000663, 0.03938427, 
    0.005726291, 0.03141037, 0.004434557, 0.01138429, 0.007320492, 
    0.0003455428, 0.001574878, 0.004226288, 0.003121529, 0.004727256, 
    0.004151024, 0.04583094, 0.00680574, 0.01681736, 1.841887e-05, 
    -0.001785345, 0.001781942, 0.01082254,
  0.0107135, 0.02165769, 0.0004881376, 0.03428443, 0.0003058213, 0.003351281, 
    0.003382953, 0.002874516, 0.03031109, 0.02324463, 0.001266035, 
    0.003005345, 0.01369004, 0.0005376636, 0.001574275, 0.002765934, 
    0.009554631, 0.007825489, 0.002152703, 0.004684268, 0.0372281, 
    0.03105492, 0.2688411, 0.06782065, 0.04982321, 0.004633308, 0.02962156, 
    0.00899973, 0.003391171,
  6.581387e-05, -8.29311e-07, -1.564567e-07, -0.002255855, 0.0317818, 
    0.008155624, 0.009336517, 0.008861598, 0.0004360342, 0.01015082, 
    0.001830304, 0.001923556, 0.005098309, 0.01194763, 0.001743244, 
    0.0007147479, 0.01774875, 0.009515527, 0.02525085, 0.01046116, 
    0.001144769, 0.0006439073, 0.2220033, 0.08949316, 0.007841802, 
    0.00714292, 0.03513329, 0.08282938, 0.0001578891,
  3.758058e-07, 2.045504e-07, 3.741652e-08, 0.0008429088, 6.457178e-06, 
    0.002051317, -5.233876e-06, 0.0008881375, 2.785671e-05, 0.056448, 
    0.04016024, 0.006912253, 0.001625409, 0.000722479, 0.0002032628, 
    0.0002999008, 0.002643618, 0.004514895, 0.04416204, 0.04065963, 
    -3.568405e-06, 0.06499763, 0.0006296417, 0.009248625, 0.002057803, 
    0.02687505, 0.01411516, 0.02938636, 3.714864e-07,
  -5.830524e-06, 0.01070776, 0.01794296, 0.003987657, 0.02041784, 
    -6.988791e-06, -0.001309892, -0.0007647733, 0.06846549, 0.2628532, 
    0.2280936, 0.2352994, 0.2837472, 0.2114835, 0.08999248, 0.1108032, 
    0.09541459, 0.02074547, 0.06653688, 0.1252601, 1.652867e-06, 0.1309891, 
    0.006216933, 0.0385366, 0.02722696, 0.03314878, 0.01610431, 0.03521695, 
    0.03080881,
  0.003408117, 0.0009397332, 0.02883758, 0.1950036, 0.03383499, 
    -3.405505e-05, 0.1226254, 0.003118368, -4.625424e-05, 0.001961034, 
    0.04912305, 0.08478627, 0.1332669, 0.1746187, 0.1086961, 0.1831158, 
    0.290722, 0.1837411, 0.1783098, 0.1242649, 0.01052864, 0.006645109, 
    0.1269703, 0.2754238, 0.1818212, 0.07752416, 0.04895192, 0.06344434, 
    0.1148322,
  0.1128383, 0.1027319, 0.05521533, 0.08561042, 0.01833444, 0.04905526, 
    0.04722604, 0.1312663, 0.008794961, 0.02901126, 0.06014284, 0.157452, 
    0.2312121, 0.282887, 0.1539989, 0.07985944, 0.2451829, 0.2585782, 
    0.2482347, 0.2220438, 0.05163812, 0.0587549, 0.1165782, 0.2193419, 
    0.2841023, 0.2792572, 0.2007236, 0.03543537, 0.1185939,
  0.07604586, 0.1933302, 0.1963844, 0.1653537, 0.1886404, 0.1100279, 
    0.1006567, 0.06201896, 0.04263961, 0.01009034, 0.002102018, 0.00679906, 
    0.1415061, 0.06543532, 0.319658, 0.4605533, 0.2992047, 0.2694578, 
    0.1176867, 0.07000721, 0.1441316, 0.1824011, 0.07333808, 0.1891124, 
    0.3691871, 0.09061141, 0.07877937, 0.08645277, 0.05408802,
  0.2558227, 0.0888505, 0.2034932, 0.1894281, 0.1617574, 0.0999658, 
    0.08658471, 0.1164644, 0.1673188, 0.2397809, 0.1342701, 0.2169466, 
    0.2616602, 0.1976021, 0.2004718, 0.1266771, 0.2288313, 0.1415879, 
    0.1657391, 0.1726895, 0.3146902, 0.1930442, 0.2035577, 0.2310966, 
    0.1081874, 0.36223, 0.1619093, 0.0637842, 0.3413982,
  0.4435524, 0.3746348, 0.2836453, 0.3822385, 0.3655778, 0.2827495, 
    0.2273083, 0.1851686, 0.1707819, 0.3372749, 0.3708405, 0.4109408, 
    0.4410091, 0.485525, 0.4860115, 0.5932931, 0.5399023, 0.4155662, 
    0.3920709, 0.4891808, 0.447565, 0.2191344, 0.2540176, 0.3916091, 
    0.118161, 0.18297, 0.09678552, 0.1769518, 0.3981528,
  0.04669929, 0.04464187, 0.04258446, 0.04052704, 0.03846962, 0.03641221, 
    0.03435479, 0.04106007, 0.05144155, 0.06182302, 0.07220449, 0.08258597, 
    0.09296744, 0.1033489, 0.1027928, 0.1099694, 0.117146, 0.1243226, 
    0.1314991, 0.1386757, 0.1458523, 0.1209006, 0.1054, 0.08989932, 
    0.07439868, 0.05889804, 0.0433974, 0.02789677, 0.04834522,
  0.4912306, 0.4536555, 0.3137576, 0.1079977, 0.06432465, 0.09768672, 
    0.0645965, 0.08465902, 0.03463352, 0.01421878, 0.02539864, 0.2696905, 
    0.4634269, -0.002102675, 0.2415441, 0.4138453, 0.4000892, 0.304639, 
    0.1822037, 0.3831368, 0.7556778, 0.7791058, 0.2186845, 0.1862756, 
    0.288103, 0.4330613, 0.3862226, 0.2123121, 0.5097831,
  0.1393964, 0.07909986, 0.2491326, 0.06358835, 0.1860197, 0.1416361, 
    0.03949773, 0.2615415, 0.2485128, 0.2057794, 0.09998048, 0.1096793, 
    0.1166846, 0.1325134, 0.2875498, 0.4005707, 0.2565379, 0.2586477, 
    0.3181577, 0.3695373, 0.3136559, 0.4414572, 0.421733, 0.3699906, 
    0.3520645, 0.304841, 0.3748538, 0.2230119, 0.2302601,
  0.2526255, 0.1983533, 0.2080036, 0.2527999, 0.2092029, 0.2153101, 
    0.2330913, 0.2052524, 0.2241244, 0.1725029, 0.1607425, 0.2100371, 
    0.3840042, 0.2899555, 0.2320008, 0.3022275, 0.2712725, 0.353304, 
    0.3373331, 0.2507719, 0.2283474, 0.2441535, 0.2075971, 0.1541435, 
    0.2958907, 0.2853069, 0.3025494, 0.2586468, 0.2797675,
  0.3038476, 0.3859706, 0.3512415, 0.2837285, 0.3132989, 0.296975, 0.2306774, 
    0.1456898, 0.1824852, 0.1711685, 0.1537958, 0.1457986, 0.08580692, 
    0.1569756, 0.1465901, 0.1198498, 0.1856494, 0.3068666, 0.2606566, 
    0.2585641, 0.1859525, 0.1494647, 0.1839235, 0.1038141, 0.03504819, 
    0.1352423, 0.2079567, 0.2921377, 0.2969101,
  0.1254338, 0.05693943, 0.02422313, 0.07330021, 0.0795316, 0.06781065, 
    0.08892027, 0.1355789, 0.06462168, 0.02921676, 0.009932306, 0.01978206, 
    0.001445099, 0.01964592, 0.2293761, 0.1075432, 0.1200788, 0.1363018, 
    0.05339723, 0.1183469, 0.06855981, 0.02420762, 0.02268804, 0.200309, 
    0.02082861, 0.0367004, 0.01273175, 0.0902034, 0.1848605,
  0.01217568, 0.02504938, 0.005025957, 0.006888161, 0.01588545, 0.0051502, 
    0.03851344, 0.01923859, 0.007724905, 0.001349975, 0.01215447, 
    -2.269172e-06, -0.0001499291, 0.0006475517, 0.02873293, 0.02091343, 
    0.02603429, 0.02771256, 0.007999038, 0.001534194, 0.01231139, 0.01264019, 
    0.00433774, 0.03738214, 0.05059116, 0.01445091, 0.01457093, 0.005520091, 
    0.003341875,
  0.04623142, 0.000101426, 5.200832e-05, 0.003048812, -0.0008725672, 
    0.001330347, 0.001335384, 0.01261555, 0.002160114, 3.452924e-05, 
    1.532366e-06, 2.148647e-06, 0.0001692899, 0.0002634184, 0.004926814, 
    0.003134692, 0.0005140304, 0.001922008, 0.0002633197, 0.002303093, 
    0.0004940914, 0.003299037, 0.008706909, 0.04512462, 0.02611252, 
    0.05872563, 0.001895333, 0.000116202, 0.001200401,
  0.03457422, 0.02046271, 5.158478e-05, 0.03833337, 0.00250085, 0.00175404, 
    0.000816801, 0.001209936, 0.002979553, -0.001048357, 0.02868796, 
    0.00205673, 0.01536499, 0.001928112, 0.005105497, 0.003463037, 
    0.0001360924, 0.000730999, 0.002390261, 0.001817794, 0.002612831, 
    0.002067082, 0.02411729, 0.004015022, 0.01597191, 6.708951e-06, 
    -0.0007341806, 0.000985119, 0.005658293,
  0.005657854, 0.03885091, 0.0003030811, 0.02294236, 0.0001256934, 
    0.001848497, 0.001897414, 0.001598482, 0.02185018, 0.02049695, 
    0.0005441346, 0.001630604, 0.008130427, 0.0001030353, 0.0004304802, 
    0.001110558, 0.003282576, 0.002134333, 0.0004277694, 0.0008988015, 
    0.005939312, 0.009113747, 0.1323436, 0.07744411, 0.04698871, 0.001598705, 
    0.0179939, 0.004249461, 0.0004231552,
  4.270136e-05, -5.211791e-07, -3.405769e-08, -0.002174405, 0.02750665, 
    0.004700947, 0.003348909, 0.005120366, 0.0001219629, 0.004838212, 
    0.0005875069, 0.0009525694, 0.001047123, 0.003642514, 0.0004882584, 
    9.840104e-05, 0.006483674, 0.0029005, 0.005739999, 0.003953763, 
    0.0004741463, 0.0003879759, 0.1584857, 0.07732122, 0.003795565, 
    0.003842625, 0.01836928, 0.04064098, 4.481175e-05,
  3.428096e-07, 1.948308e-07, 3.688557e-08, 5.886533e-05, 0.0001008314, 
    0.0007478498, -3.661644e-05, 0.0002885475, 1.82648e-05, 0.01682802, 
    0.01644126, 0.001529567, 0.000343801, 0.0002297383, 0.0001078099, 
    0.0001503164, 0.001036576, 0.00211312, 0.02331459, 0.02361911, 
    -1.457585e-06, 0.05362201, 0.0001747284, 0.006034104, 0.0009065344, 
    0.0148284, 0.008279296, 0.01629535, 3.377955e-07,
  -4.334032e-06, 0.007355702, 0.009806258, 0.002552367, 0.01850079, 
    -2.580601e-06, -0.001303466, -0.0007305923, 0.05774375, 0.1976555, 
    0.2069221, 0.1928456, 0.2164699, 0.1486953, 0.06712515, 0.04313133, 
    0.07334169, 0.010413, 0.03945074, 0.1045455, 1.478641e-06, 0.1217574, 
    0.002004172, 0.02764023, 0.01817399, 0.01876166, 0.009903775, 0.01720348, 
    0.02082394,
  0.002608731, 9.332199e-05, 0.01628972, 0.1908945, 0.06849387, 
    -3.860011e-05, 0.107039, 0.003032042, -3.598214e-05, 0.001242119, 
    0.04413839, 0.08158624, 0.1161523, 0.1378353, 0.08496312, 0.1517305, 
    0.2443135, 0.1670894, 0.1111516, 0.1050932, 0.007280317, 0.004874869, 
    0.0963175, 0.2541898, 0.123511, 0.05137047, 0.02661161, 0.03612797, 
    0.08475085,
  0.09395405, 0.07921567, 0.03644624, 0.06247954, 0.01752135, 0.0371365, 
    0.03326576, 0.1057739, 0.003393189, 0.02318723, 0.05671892, 0.1377982, 
    0.1872097, 0.2342027, 0.1213018, 0.06497594, 0.2171726, 0.206693, 
    0.2028613, 0.2145398, 0.04359614, 0.03751092, 0.09647661, 0.2024736, 
    0.2665686, 0.2993231, 0.1384473, 0.01820058, 0.07167652,
  0.0622895, 0.170955, 0.1652343, 0.1518163, 0.1706905, 0.1003162, 
    0.08109493, 0.05090775, 0.02919854, 0.007758127, 0.001792842, 
    0.007033916, 0.1376458, 0.04114921, 0.2524833, 0.4172658, 0.2650206, 
    0.232703, 0.07202008, 0.06253156, 0.127966, 0.1744424, 0.08110694, 
    0.1809216, 0.3213566, 0.07140458, 0.05144648, 0.06233873, 0.03076472,
  0.199945, 0.06582359, 0.1754264, 0.1422201, 0.1600922, 0.1052838, 
    0.09028181, 0.1065489, 0.1316581, 0.1840271, 0.1214114, 0.1895271, 
    0.271938, 0.2307149, 0.1943363, 0.1953976, 0.2175426, 0.1601988, 
    0.1747518, 0.1696155, 0.3649729, 0.2056698, 0.1933049, 0.2584982, 
    0.1274298, 0.3349516, 0.1670916, 0.03354951, 0.325166,
  0.5024199, 0.3926893, 0.3359887, 0.3919246, 0.3464511, 0.3091357, 
    0.2973044, 0.2405604, 0.208392, 0.3609673, 0.368824, 0.4247763, 0.511663, 
    0.5444506, 0.5889716, 0.6636182, 0.6018517, 0.4871856, 0.37857, 
    0.4776992, 0.4943277, 0.2083266, 0.2295734, 0.431006, 0.117876, 
    0.1485007, 0.07187954, 0.1622259, 0.3683443,
  0.04971619, 0.04916412, 0.04861207, 0.04806, 0.04750795, 0.04695588, 
    0.04640383, 0.04022042, 0.04619131, 0.0521622, 0.05813309, 0.06410398, 
    0.07007487, 0.07604576, 0.09058465, 0.09546646, 0.1003483, 0.1052301, 
    0.1101119, 0.1149937, 0.1198756, 0.08464182, 0.07434118, 0.06404053, 
    0.05373988, 0.04343923, 0.03313858, 0.02283793, 0.05015783,
  0.4878913, 0.3927369, 0.216169, 0.02814543, 0.01713998, 0.04129656, 
    0.02323254, 0.02381752, 0.03803113, 0.01198893, 0.008742523, 0.2059198, 
    0.3339315, -0.003765488, 0.3427715, 0.412407, 0.3990667, 0.2991568, 
    0.1527921, 0.3835275, 0.7413929, 0.7824572, 0.1775316, 0.1663821, 
    0.4015885, 0.4839799, 0.3971413, 0.2033151, 0.4412237,
  0.1085602, 0.05826522, 0.1965514, 0.03511035, 0.1385245, 0.133267, 
    0.03048375, 0.2205079, 0.2294991, 0.1677837, 0.08454663, 0.1008927, 
    0.08695863, 0.1165828, 0.2501473, 0.3474893, 0.2061364, 0.2127306, 
    0.2495111, 0.2994276, 0.2459822, 0.3601897, 0.3499897, 0.3369482, 
    0.3306885, 0.2802011, 0.3353658, 0.158035, 0.1802032,
  0.1918594, 0.1475721, 0.1559683, 0.185347, 0.146326, 0.1573622, 0.1602837, 
    0.1432668, 0.169313, 0.128204, 0.1287332, 0.1666881, 0.2974455, 
    0.2151944, 0.1646831, 0.2456561, 0.2224315, 0.2798587, 0.262889, 
    0.2000233, 0.168348, 0.181355, 0.1448867, 0.1095117, 0.2459718, 
    0.2403479, 0.2260595, 0.1906173, 0.2140943,
  0.2352052, 0.3139885, 0.2733156, 0.2260187, 0.2353886, 0.2264607, 
    0.1822736, 0.1140072, 0.1397436, 0.1140468, 0.1055797, 0.09543508, 
    0.05973415, 0.1038891, 0.1096655, 0.09544518, 0.139343, 0.2201654, 
    0.1837585, 0.1975295, 0.1413605, 0.1121668, 0.1288099, 0.08433529, 
    0.02104454, 0.09025602, 0.1557249, 0.2403598, 0.2419218,
  0.08948363, 0.03176253, 0.01343388, 0.04699716, 0.04989695, 0.03776328, 
    0.06654116, 0.1053703, 0.03737638, 0.01307435, 0.004095179, 0.01181273, 
    0.001043835, 0.01133774, 0.1910196, 0.07420176, 0.05803272, 0.0990868, 
    0.03279302, 0.08769377, 0.0454896, 0.0130655, 0.01226179, 0.1795036, 
    0.01365885, 0.02052973, 0.005534501, 0.05730499, 0.1277065,
  0.007756336, 0.01504498, 0.005137758, 0.004225933, 0.009339567, 0.00212856, 
    0.01627694, 0.009283164, 0.004827093, 0.0009481166, 0.01312476, 
    -1.027422e-06, 0.0001318521, 0.0003499367, 0.01340705, 0.009441144, 
    0.01609082, 0.01605646, 0.003005924, 0.0008857744, 0.005331506, 
    0.006259212, 0.002765592, 0.0255395, 0.03505456, 0.006502266, 
    0.007655505, 0.002154941, 0.002218239,
  0.02779736, -9.763212e-05, -5.664914e-05, 0.001827912, -0.0007814015, 
    0.0004972756, 0.0005448901, 0.005139705, 0.001338422, 2.021083e-05, 
    2.992847e-07, 1.50834e-06, 9.61778e-05, 0.0001328468, 0.00210096, 
    0.001151858, 0.0002224658, 0.0007993444, 0.0001413757, 0.001514132, 
    0.0003161868, 0.002248729, 0.005670882, 0.0293858, 0.01857907, 0.0435206, 
    0.001046153, 7.055712e-05, 0.0007542616,
  0.02131565, 0.01037478, 1.653731e-05, 0.03060602, 0.001493413, 
    0.0008460351, 0.0002244744, 0.0005843724, 0.001303748, -0.0006159008, 
    0.01721172, 0.0006428341, 0.006304568, 0.0008970161, 0.001922616, 
    0.001260024, 8.345771e-05, 0.0004379931, 0.001585479, 0.001229095, 
    0.001696572, 0.00126976, 0.01550728, 0.003948333, 0.01402909, 
    1.938455e-06, -0.0002080985, 0.0006370024, 0.003630159,
  0.002804705, 0.03709131, 0.0001525621, 0.01419304, 7.128515e-05, 
    0.001198193, 0.001260392, 0.001048037, 0.01528614, 0.02140327, 
    0.0003432813, 0.001043368, 0.003662464, 5.712729e-05, 0.0002544796, 
    0.0006336007, 0.001865024, 0.001046587, 0.000227148, 0.0004708833, 
    0.002029585, 0.005101695, 0.06973653, 0.07821234, 0.04736141, 
    0.0004548845, 0.009007943, 0.002202519, 0.0001862113,
  2.9285e-05, -2.021287e-07, 2.343172e-08, -0.000953224, 0.01697395, 
    0.003180095, 0.000898009, 0.003479062, 9.455247e-05, 0.00218168, 
    0.000437191, 0.0004702172, 0.0003894544, 0.001140336, 0.0001744915, 
    3.498597e-05, 0.002042384, 0.00131418, 0.002238594, 0.002041454, 
    0.0003269887, 0.0003075321, 0.1211509, 0.06554385, 0.001692217, 
    0.002498856, 0.01177982, 0.0245856, -1.560639e-05,
  3.245385e-07, 1.89968e-07, 3.515853e-08, 2.122683e-05, 2.890907e-06, 
    0.0004049449, -2.313362e-05, 0.0001281712, 1.060905e-05, 0.008272082, 
    0.007602103, 0.0005318208, 0.0001916144, 0.0001497335, 7.077853e-05, 
    9.28058e-05, 0.0006802416, 0.001299544, 0.01516938, 0.01612348, 
    -8.373365e-07, 0.04496678, 0.0001151419, 0.00246993, 0.0006004354, 
    0.007474673, 0.00573607, 0.01086302, 3.222754e-07,
  -1.558204e-06, 0.005044578, 0.005375572, 0.001841592, 0.01509955, 
    -9.244254e-07, -0.00123711, -0.0008037159, 0.05229297, 0.1250653, 
    0.172909, 0.1288427, 0.1288226, 0.09336036, 0.04429061, 0.02369734, 
    0.05383423, 0.005784828, 0.02493565, 0.08073492, 1.311936e-06, 0.1018424, 
    0.001312663, 0.01718142, 0.01107179, 0.01157743, 0.00492664, 0.009955936, 
    0.01499368,
  0.00224824, 2.998999e-05, 0.008980094, 0.1742226, 0.06722017, 
    -2.968998e-05, 0.09385318, 0.002897103, -2.764257e-05, 0.0008749511, 
    0.0406164, 0.07432184, 0.09418421, 0.1046222, 0.05406227, 0.111004, 
    0.1963512, 0.1329164, 0.0683516, 0.08537554, 0.006917385, 0.003397249, 
    0.07167426, 0.2330318, 0.08130938, 0.03271849, 0.01494934, 0.02086575, 
    0.06288514,
  0.06968576, 0.0586543, 0.02628991, 0.04259299, 0.01773965, 0.0287595, 
    0.02450615, 0.08754051, 0.002480187, 0.01775198, 0.04515968, 0.1113995, 
    0.138754, 0.1829493, 0.09385496, 0.049853, 0.16794, 0.1400176, 0.1382334, 
    0.2018763, 0.0341641, 0.02369117, 0.07993595, 0.1815703, 0.2384506, 
    0.2863602, 0.1017866, 0.009260396, 0.03813672,
  0.03980131, 0.1492545, 0.1414312, 0.1324173, 0.1471984, 0.08627123, 
    0.0676498, 0.03480349, 0.01682267, 0.00503649, 0.001427446, 0.01152367, 
    0.1303411, 0.03248832, 0.2055504, 0.3621122, 0.2346966, 0.1987179, 
    0.05408423, 0.05035159, 0.1065261, 0.1578798, 0.09091601, 0.1796324, 
    0.2731537, 0.05211116, 0.02851768, 0.04257276, 0.01861971,
  0.1565951, 0.04481646, 0.1531345, 0.1072504, 0.1558663, 0.1292764, 
    0.1554692, 0.1212955, 0.1210748, 0.1881226, 0.1231163, 0.1524064, 
    0.2316539, 0.1938767, 0.15498, 0.1966124, 0.2068571, 0.1645096, 0.218498, 
    0.1976957, 0.3391359, 0.238473, 0.1748982, 0.2974452, 0.145646, 
    0.2821214, 0.1599049, 0.01483007, 0.2699271,
  0.5049919, 0.3172886, 0.3092412, 0.3372289, 0.3259493, 0.3132712, 0.299918, 
    0.2311957, 0.2533845, 0.3471058, 0.3311507, 0.3719122, 0.4790092, 
    0.5438417, 0.5395377, 0.5789079, 0.4692301, 0.4352635, 0.3752363, 
    0.4383796, 0.4366187, 0.1790143, 0.2315667, 0.442724, 0.1033584, 
    0.1299354, 0.05697004, 0.1519416, 0.3290025,
  0.04410319, 0.04345647, 0.04280975, 0.04216303, 0.04151631, 0.04086959, 
    0.04022286, 0.03754795, 0.04262602, 0.04770409, 0.05278216, 0.05786023, 
    0.0629383, 0.06801636, 0.08061361, 0.08337748, 0.08614135, 0.08890522, 
    0.09166908, 0.09443295, 0.09719682, 0.08114171, 0.0739465, 0.06675129, 
    0.05955607, 0.05236086, 0.04516564, 0.03797043, 0.04462057,
  0.4162822, 0.281952, 0.09486887, 0.003934475, 0.008187909, 0.01647861, 
    0.01613661, 0.003103761, 0.002065618, 0.01029987, 0.00929933, 0.1433271, 
    0.2807586, -0.003192288, 0.4157841, 0.3947799, 0.3884391, 0.2945652, 
    0.1148707, 0.4244578, 0.7239621, 0.7710384, 0.1754263, 0.1620592, 
    0.3867792, 0.5038946, 0.4019568, 0.1805334, 0.4255804,
  0.09733959, 0.04712917, 0.1562055, 0.02264513, 0.1081978, 0.1100992, 
    0.024899, 0.1962952, 0.2261189, 0.1232366, 0.07890379, 0.08968244, 
    0.06693931, 0.1000506, 0.2296348, 0.305291, 0.1747802, 0.1864109, 
    0.2011954, 0.2433047, 0.1994237, 0.2954361, 0.3010508, 0.297881, 
    0.2923414, 0.2624362, 0.2999553, 0.1159572, 0.153493,
  0.1527623, 0.1177439, 0.1240408, 0.1474661, 0.1101485, 0.1237229, 
    0.1260394, 0.1086647, 0.1324783, 0.1028988, 0.1072199, 0.1403913, 
    0.2412501, 0.1693965, 0.1204197, 0.1989143, 0.1918315, 0.2257621, 
    0.2116954, 0.1689722, 0.1289759, 0.1361557, 0.1092022, 0.08112194, 
    0.2102774, 0.1988453, 0.1792532, 0.1504927, 0.169353,
  0.1915206, 0.2605893, 0.2171506, 0.1769364, 0.1782861, 0.1830737, 
    0.1492748, 0.09325937, 0.1103242, 0.08112352, 0.07466674, 0.06383798, 
    0.04287963, 0.07094596, 0.08223066, 0.07076915, 0.1039551, 0.1504068, 
    0.1277575, 0.1523884, 0.1032824, 0.08219658, 0.08849638, 0.0757443, 
    0.01054954, 0.06045827, 0.118815, 0.186215, 0.2040687,
  0.06640002, 0.01948038, 0.009223147, 0.02851379, 0.03015621, 0.02180817, 
    0.04996385, 0.07072953, 0.02191491, 0.00747754, 0.002573366, 0.008096527, 
    0.0008423801, 0.006026867, 0.1655879, 0.04703633, 0.03413476, 0.06947443, 
    0.02017872, 0.0598045, 0.02591275, 0.007548041, 0.007642276, 0.1607568, 
    0.009430845, 0.01103458, 0.002947427, 0.03437377, 0.09026436,
  0.005815357, 0.0106931, 0.004999818, 0.00310912, 0.004762749, 0.001256078, 
    0.007904101, 0.005104685, 0.003635787, 0.0007426564, 0.007837522, 
    -6.744634e-07, 0.0003047964, 0.000268347, 0.006524154, 0.005751045, 
    0.009220564, 0.008976769, 0.001880245, 0.000699772, 0.002643758, 
    0.003209351, 0.002060134, 0.01948058, 0.02638203, 0.003647916, 
    0.003868004, 0.001159746, 0.001676327,
  0.02003696, -0.0001996465, -0.0001063627, 0.001301013, -0.0004446701, 
    0.0002454253, 0.0003178351, 0.002413875, 0.0009629593, 1.394806e-05, 
    6.374413e-08, -1.494962e-06, 6.996935e-05, 0.000114624, 0.001187355, 
    0.000599865, 0.0001807355, 0.0004072682, 0.0001140563, 0.001116219, 
    0.0002286984, 0.001708305, 0.004226343, 0.02194701, 0.01500368, 
    0.03334195, 0.000744577, 5.043562e-05, 0.0005477165,
  0.01523919, 0.005821596, 0.0005946003, 0.03266374, 0.001041887, 
    0.000515399, 0.0001624535, 0.0002880051, 0.0006052442, -0.0005026071, 
    0.01155582, 0.0002696124, 0.002871637, 0.0004868432, 0.0008338455, 
    0.0005149401, 6.129082e-05, 0.0003078728, 0.001183995, 0.0009309906, 
    0.001248534, 0.0009010425, 0.01137036, 0.00492859, 0.01662207, 
    6.567293e-08, -2.602635e-05, 0.0004664383, 0.002660524,
  0.001378375, 0.02772894, -5.693694e-05, 0.009724294, 4.852692e-05, 
    0.000873754, 0.0009395134, 0.0007343218, 0.01078833, 0.02241893, 
    0.0002555977, 0.0007641857, 0.001576569, 3.704835e-05, 0.0001714341, 
    0.0004308156, 0.001277627, 0.0006599284, 0.0001507533, 0.0003136952, 
    0.001259685, 0.003607174, 0.0453308, 0.06004861, 0.03811159, 
    0.0001976942, 0.004366263, 0.00113302, 0.0001259356,
  2.263628e-05, -1.235084e-07, 3.308953e-08, -0.0001133217, 0.01093102, 
    0.002416684, -0.0005527924, 0.002629624, 8.220183e-05, 0.001213635, 
    0.0003881913, 0.0003184145, 0.0002008542, 0.000441014, 9.655308e-05, 
    2.209474e-05, 0.0007793674, 0.0008665615, 0.001358774, 0.001277595, 
    0.0002403786, 0.0002452628, 0.08592592, 0.05052159, 0.0006801714, 
    0.00183317, 0.008623874, 0.01756812, 0.0009859182,
  3.15916e-07, 1.827167e-07, 3.286185e-08, 1.630617e-05, 3.453957e-06, 
    0.0002682235, -1.344048e-05, 7.335584e-05, 5.337992e-06, 0.005108817, 
    0.004298318, 0.0003452421, 0.0001360624, 0.000113464, 5.319068e-05, 
    6.725469e-05, 0.0005145576, 0.0009528908, 0.01125661, 0.01236126, 
    -5.802736e-07, 0.03893166, 9.18048e-05, 0.0004402446, 0.0004641264, 
    0.003446964, 0.004421237, 0.008152222, 3.119866e-07,
  -1.424884e-07, 0.003254038, 0.003789922, 0.001216959, 0.01289914, 
    -3.728852e-07, -0.001217326, -0.001189125, 0.05353396, 0.07770526, 
    0.1280701, 0.07946851, 0.08010594, 0.0602176, 0.02912818, 0.01435259, 
    0.03650562, 0.004019868, 0.01597621, 0.05337017, 1.199725e-06, 
    0.08537455, 0.003684948, 0.007460559, 0.005249737, 0.006175629, 
    0.003054053, 0.005555319, 0.01041934,
  0.001630255, -4.208718e-05, 0.005298852, 0.167497, 0.05879648, 
    -2.496682e-05, 0.08412757, 0.002757424, -2.377751e-05, 0.0007085086, 
    0.04222902, 0.06178613, 0.07760579, 0.08641309, 0.03797869, 0.08083598, 
    0.1468697, 0.09403344, 0.04685861, 0.07113077, 0.006813584, 0.002645919, 
    0.05353952, 0.2145841, 0.05488286, 0.01951672, 0.009678438, 0.0137906, 
    0.04544024,
  0.05054822, 0.04349288, 0.02105985, 0.02815726, 0.01499602, 0.02281302, 
    0.02030685, 0.07816918, 0.00249866, 0.01506815, 0.03957067, 0.09070406, 
    0.1070934, 0.1468066, 0.07525162, 0.03977479, 0.1318114, 0.103153, 
    0.09055673, 0.1915687, 0.02793867, 0.01783922, 0.07831197, 0.1650272, 
    0.2066081, 0.2653264, 0.07444666, 0.005824801, 0.02193411,
  0.02174984, 0.1376304, 0.1286786, 0.1411206, 0.1287469, 0.07921115, 
    0.05926293, 0.02927733, 0.01339476, 0.004527696, 0.001316886, 0.0497536, 
    0.1359579, 0.03005739, 0.1743915, 0.3078662, 0.2172251, 0.1737277, 
    0.05019642, 0.04156168, 0.08965448, 0.1440732, 0.08417539, 0.2024123, 
    0.2316965, 0.04013091, 0.01903361, 0.03043215, 0.01306839,
  0.1225814, 0.03364301, 0.1427332, 0.0847814, 0.1736813, 0.128787, 
    0.2459982, 0.1689232, 0.1571129, 0.208695, 0.1439224, 0.1325044, 
    0.2442854, 0.1572366, 0.1091433, 0.1505504, 0.2038067, 0.1415138, 
    0.2224116, 0.1649784, 0.3072793, 0.2379681, 0.2341427, 0.3125414, 
    0.1852233, 0.253383, 0.1734404, 0.009821991, 0.2261498,
  0.465789, 0.2861094, 0.2799534, 0.2939342, 0.2912748, 0.260639, 0.2430173, 
    0.1713635, 0.2207707, 0.2259009, 0.2297377, 0.2821181, 0.3408364, 
    0.3800872, 0.3897265, 0.3811986, 0.3000226, 0.2890104, 0.2551006, 
    0.3339245, 0.3199081, 0.1443312, 0.2157252, 0.4752583, 0.1006243, 
    0.09447647, 0.05420959, 0.1391256, 0.2702056,
  0.0358117, 0.03473014, 0.03364859, 0.03256703, 0.03148547, 0.03040392, 
    0.02932236, 0.01993156, 0.02369464, 0.02745772, 0.0312208, 0.03498388, 
    0.03874695, 0.04251003, 0.0493119, 0.05231174, 0.05531157, 0.0583114, 
    0.06131123, 0.06431106, 0.06731089, 0.07037184, 0.06469048, 0.05900913, 
    0.05332777, 0.04764642, 0.04196506, 0.03628371, 0.03667695,
  0.3148237, 0.2041708, 0.02222653, 0.004553586, 0.00273609, 0.008481689, 
    0.01450041, 0.002558272, 0.00149582, 0.004938014, 0.007365971, 0.126764, 
    0.265945, -0.002362208, 0.407178, 0.3577735, 0.383374, 0.3242823, 
    0.1155092, 0.434729, 0.7123053, 0.7564479, 0.1888811, 0.1664669, 
    0.3132206, 0.4989768, 0.4142755, 0.1950515, 0.3942465,
  0.09352481, 0.04193753, 0.1378149, 0.01871812, 0.07899155, 0.09489914, 
    0.02215217, 0.1882085, 0.2149388, 0.1119769, 0.07067185, 0.08357164, 
    0.05799197, 0.09259711, 0.2250809, 0.2811872, 0.1630645, 0.1735318, 
    0.1735635, 0.2138793, 0.1734621, 0.2591896, 0.2711095, 0.2704697, 
    0.265344, 0.2439045, 0.2856686, 0.1005609, 0.13992,
  0.1307168, 0.1023448, 0.1054112, 0.1274978, 0.09310675, 0.1070369, 
    0.1105288, 0.09056245, 0.113596, 0.08981843, 0.09263074, 0.1214881, 
    0.2084045, 0.1427554, 0.09986626, 0.1655391, 0.1654737, 0.1952759, 
    0.1799624, 0.1432357, 0.1071468, 0.1142761, 0.0922729, 0.06766424, 
    0.1737635, 0.1722843, 0.1541924, 0.1286307, 0.1476099,
  0.1630696, 0.2154195, 0.1812598, 0.1429082, 0.1477967, 0.1560524, 0.127537, 
    0.08048102, 0.09122885, 0.0676443, 0.05892375, 0.04922612, 0.03264503, 
    0.05480658, 0.06536236, 0.0563746, 0.08388732, 0.1132497, 0.09568715, 
    0.1201443, 0.07592437, 0.06295442, 0.06813861, 0.0964866, 0.005728802, 
    0.04696752, 0.09459036, 0.1526026, 0.1682279,
  0.04849358, 0.01463144, 0.007264787, 0.01882955, 0.02064257, 0.01445281, 
    0.03696315, 0.04771626, 0.0156992, 0.005382494, 0.002077549, 0.006657519, 
    0.0007525893, 0.004204372, 0.1681164, 0.02900664, 0.0244809, 0.05068983, 
    0.01328093, 0.04341808, 0.01647023, 0.005261591, 0.005795624, 0.161409, 
    0.006182709, 0.007608676, 0.001980375, 0.02360383, 0.06553547,
  0.004806913, 0.008592973, 0.009152737, 0.002585606, 0.003356971, 
    0.0009616851, 0.005124541, 0.003397863, 0.003053841, 0.0006384396, 
    0.004666715, -5.598396e-07, 0.003087356, 0.0002289204, 0.003755295, 
    0.004378279, 0.005660778, 0.005207144, 0.001487867, 0.0005918441, 
    0.001503256, 0.002086511, 0.001710778, 0.01587605, 0.02757002, 
    0.002620767, 0.002508421, 0.0008475062, 0.001401875,
  0.01596098, -0.0001062943, -0.0001031727, 0.001046793, -0.0006011935, 
    0.0001768896, 0.0002377574, 0.001670398, 0.0007687857, 1.114328e-05, 
    4.444299e-08, -5.060617e-05, 5.88287e-05, 0.000104136, 0.0008579049, 
    0.0004388983, 0.0001569744, 0.0002791226, 9.811996e-05, 0.000908562, 
    0.0001847219, 0.001422939, 0.003519384, 0.01809545, 0.03235358, 
    0.03370818, 0.0006044025, 4.097693e-05, 0.0004540374,
  0.01234933, 0.005127815, 0.003979652, 0.05937536, 0.0008225494, 
    0.0003885725, 0.0001420971, 0.0001967227, 0.0003841026, -0.0006120965, 
    0.009120646, 0.0001810923, 0.002182102, 0.0003503853, 0.0005283198, 
    0.0003210425, 5.076387e-05, 0.0002474043, 0.0009845662, 0.0007797171, 
    0.001032205, 0.0007302819, 0.009345134, 0.04012878, 0.05304395, 
    -4.275378e-05, 3.468041e-06, 0.0003869936, 0.002193614,
  0.0009180531, 0.02915362, 0.0005434752, 0.0100588, 3.867308e-05, 
    0.0007065633, 0.0007718512, 0.0005958523, 0.0133671, 0.06183758, 
    0.000211811, 0.0006299185, 0.000876496, 2.581078e-05, 9.661429e-05, 
    0.0003368796, 0.000978736, 0.0005158516, 0.0001228059, 0.0002341448, 
    0.0009560026, 0.002912304, 0.03358206, 0.06264969, 0.08849155, 
    0.0001420183, 0.002534901, 0.0007613914, 0.0001008896,
  0.0009749989, -2.276755e-06, 3.334445e-08, 0.002484643, 0.007519472, 
    0.002019273, -0.000884608, 0.002191358, 4.953386e-05, 0.0008615828, 
    0.000231873, 0.0002522838, 0.0001402363, 0.0002816887, 7.08003e-05, 
    1.767539e-05, 0.0004707282, 0.0006819291, 0.001040556, 0.0009641818, 
    0.0002033057, 0.0002114711, 0.1119355, 0.04705631, 0.0003872461, 
    0.001523463, 0.007088599, 0.01414851, 0.02094192,
  3.137193e-07, 1.813795e-07, 3.16226e-08, 1.353349e-05, -4.193639e-06, 
    0.0002028374, -8.471507e-06, 7.11262e-05, 2.321113e-06, 0.002839877, 
    0.003098437, 0.0002422143, 0.000112137, 8.370007e-05, 4.483883e-05, 
    5.60944e-05, 0.0004322431, 0.0007989751, 0.0093433, 0.01044378, 
    -4.709621e-07, 0.0369921, 7.933464e-05, -0.000231561, 0.0003951984, 
    0.002220623, 0.00373361, 0.00679942, 3.077596e-07,
  3.71146e-07, 0.002531228, 0.003604122, 0.0007703257, 0.01370411, 
    -1.332913e-07, -0.001297371, -0.001857722, 0.06567147, 0.06076205, 
    0.08988766, 0.05063333, 0.05727334, 0.04460006, 0.02063374, 0.01008111, 
    0.02669672, 0.003341356, 0.01195375, 0.03820882, 1.050483e-06, 
    0.09495625, 0.02848683, 0.003804237, 0.002947821, 0.00399195, 
    0.002123602, 0.002981933, 0.007578087,
  0.001576903, -0.0002489737, 0.003951957, 0.1637266, 0.05246269, 
    -1.979357e-05, 0.0751366, 0.002612564, -2.126429e-05, 0.0006796942, 
    0.0484203, 0.04664958, 0.06818753, 0.06569985, 0.03001179, 0.06550276, 
    0.1072792, 0.07188419, 0.03676539, 0.06697174, 0.007180512, 0.003506238, 
    0.04364186, 0.1901212, 0.04257551, 0.01258656, 0.007469077, 0.01093588, 
    0.03696728,
  0.0406485, 0.03770508, 0.01863948, 0.02112408, 0.01269706, 0.02028896, 
    0.01844035, 0.08362276, 0.0006500058, 0.01753078, 0.04554808, 0.09607149, 
    0.08589967, 0.1275374, 0.06518488, 0.03431809, 0.1140572, 0.08389733, 
    0.06701092, 0.1998139, 0.02793287, 0.02208081, 0.0857211, 0.1793547, 
    0.1902011, 0.2225751, 0.05338471, 0.004528142, 0.01603359,
  0.01639861, 0.1430628, 0.1315002, 0.1657685, 0.1467278, 0.08540869, 
    0.05930274, 0.03339732, 0.01815834, 0.008462771, 0.004030494, 0.1982172, 
    0.1720932, 0.0332906, 0.1559424, 0.2819626, 0.2459298, 0.1594069, 
    0.06951115, 0.04357939, 0.0887249, 0.1677491, 0.07232601, 0.2678009, 
    0.2058222, 0.03668398, 0.01488962, 0.0245828, 0.01084729,
  0.1038649, 0.02933553, 0.1647128, 0.06300677, 0.2152103, 0.1248952, 
    0.3416477, 0.2506973, 0.271262, 0.2760519, 0.2042397, 0.1626445, 
    0.3078758, 0.141524, 0.09849557, 0.1069328, 0.271039, 0.1467502, 
    0.2440698, 0.1624887, 0.3068599, 0.2225711, 0.3003099, 0.3402369, 
    0.1911805, 0.235783, 0.2142444, 0.0116649, 0.1939587,
  0.4240766, 0.2610314, 0.251304, 0.2627169, 0.2644277, 0.2209376, 0.2024382, 
    0.1370138, 0.1547272, 0.1725472, 0.1700522, 0.1929437, 0.2429715, 
    0.2732264, 0.2554131, 0.2770264, 0.2234904, 0.2311385, 0.1895527, 
    0.2334417, 0.2306476, 0.1342824, 0.2290425, 0.5121822, 0.08933163, 
    0.07361466, 0.05937312, 0.1438744, 0.2444025,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, -5.862915e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0002929461, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, -3.784163e-05, 0.0005665174, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, -2.304413e-05, 0, 0, -2.634399e-10, 0, 0, 0, 1.243703e-05, 0, 
    -1.418364e-10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, -4.931804e-06, 0.001811716, 0, -9.593207e-06, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.0002594731, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, -3.345096e-05, -0.0001306504, 0, -8.163258e-05, 
    0.0008497718, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, -9.010768e-05, 0, 0, 0.001228287, 0, 0, 0, 2.465658e-05, 
    0.0001875303, 1.321171e-05, 0, 0, -1.78845e-06, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, -3.12206e-06, 0, 0,
  0, 0, 0, 0, 0, 0, 0, -7.685249e-06, 0, -3.344151e-05, 0.0047882, 
    -2.588332e-05, -4.226278e-05, -1.960104e-05, 0, 0, 0, 0, 0, 0, 0, 
    0.001120088, 0.001352596, 0.0001064647, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4.087927e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -3.35912e-05, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0.00259812, 0.001023044, 0, -0.0001593335, 0.003002255, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0002178069, 0, 0, 0, 0, 0,
  0, 0, -1.201261e-05, 0, 0, 0.006174447, 0.002444618, 0, 0, 3.644114e-05, 
    0.001187145, 1.981766e-05, 0, 0, 4.781515e-05, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0001802935, 0, 0, -1.460812e-05, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0.0003406273, 0, -4.084218e-05, 0.009712369, 
    -6.919707e-05, -0.0002103639, -0.0001423693, 0, 0, 0, -2.759505e-05, 
    -2.491064e-05, -2.378213e-05, 0, 0.005706223, 0.002253368, 0.0001242088, 
    0, 0, 0, 0, -6.038068e-05,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0004066568, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, -4.631582e-05, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -5.440896e-06, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, -1.566946e-05, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0005069728, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0001385835, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, -4.022025e-06, 0, 0, 0, 0,
  0, 0, 0, 0, 0, -9.665681e-05, -9.575534e-06, -1.119205e-05, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, -3.307419e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, -1.537066e-05, -2.179487e-05, 0, 0, 0, 0.005845943, 0.002396834, 
    -7.495759e-06, -0.0002229146, 0.006010562, -8.677594e-06, 0, 0.000346578, 
    0, 0, -1.537748e-05, 0, 0, 0, 0, 0, 0, 0.001215004, 0, 0, 0, 0, 0,
  0, 0, 0.0001701052, 0, 0, 0.007871994, 0.004599601, 0, 2.121699e-06, 
    3.929982e-05, 0.003058517, 1.087029e-06, 0, 1.520171e-07, 0.001981335, 0, 
    0, 0, 0, 0, 0, 0, -1.310224e-08, 0.001008965, 0, 0, -5.047528e-05, 0, 0,
  0, 0, 0, -2.943848e-05, 0, 0, 0, 0.0006678515, -5.001743e-06, 0.0008134257, 
    0.01447005, -0.0001268638, 0.0001530322, 0.0003325126, -3.268726e-05, 
    -4.343673e-05, 0, -7.601836e-05, 0.0001015274, -0.0001597764, 0, 
    0.01174629, 0.003614269, 0.0001207041, 0, 0, 0, 0, -8.810026e-05,
  0, 0, 0, 0, 0, 0, 0, 0, 0, -6.440476e-06, 0.001493452, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, -0.0001610717, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0003424904, 0, 0, -5.662232e-06, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.002903268, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.385512e-05, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.0007241916, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.003509236, -3.672637e-05, 
    -4.658738e-05, 0, -1.192847e-06, 0, 0.0003364817, 0, 0, 0, -1.608502e-05, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, -0.0002465495, -9.733187e-05, -0.0001033444, 0, 0, 
    -9.382099e-05, 0, 0, 0, 0, 0, 0, -1.815862e-05, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0,
  0, -0.0001652362, 9.907984e-05, 0, 0, 0, 0.0100862, 0.01155272, 
    0.001723381, -0.0006638626, 0.008270103, -1.074234e-05, 0, 0.000406659, 
    -9.066099e-06, 0, -2.400762e-05, 0, 0, 0, 0, 0, 0, 0.002558374, 0, 0, 0, 
    0, 0,
  0, 3.74494e-05, 0.003112496, -1.877735e-05, 0, 0.01546314, 0.006354061, 0, 
    4.243374e-06, 6.015197e-05, 0.01019555, -0.000111024, 4.059317e-08, 
    2.700478e-06, 0.007039957, -2.215279e-05, 7.253941e-06, 0, 0, 0, 0, 0, 
    -4.585784e-08, 0.003819995, -3.617985e-05, 0, -0.0001533359, 0, 0,
  0, 0, 0, -3.284459e-05, 0, 0, 0.0003672462, 0.0007018446, 0.0005481232, 
    0.001065909, 0.02085712, 0.0009315335, 0.001983627, 0.000719043, 
    -0.0002056204, -0.0001544955, 0, 0.0009583046, 0.0003709505, 
    -0.0002048662, 0, 0.02392318, 0.006777318, 0.002949942, 0, 0, 0, 
    -4.904561e-06, -0.0001687493,
  0, 0, 0, 0, 0, 0, 0, 0, 0.0001958675, -6.440476e-06, 0.002411575, 0, 
    -2.001803e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0.0003168734, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001176484, 0.0001708068, -2.186126e-05, 
    1.879476e-05, 0, 0, -4.787686e-06, 0, 0, 0, 0, 0, 0, 0, 0.004211401, 0, 
    0.0005229578, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.567172e-05, 0.0003596045, 0.00164228, 
    0, 0, 0, 0, 0, 0, 0, 0.0001645724, 0.001057597, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.339278e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, -1.101431e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, -9.921234e-06, 0, 0, 0,
  0, 0, 0, -6.251582e-07, -1.362803e-05, 0.0002884573, -5.381211e-05, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.0006893559, 0, 0, -2.446401e-05, 0, 0, 0.0005851033, 
    0, 0, 0.00245679, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01128679, 0.002616933, 
    0.0004622402, -8.685356e-06, 0.0002665243, 0, 0.003476991, 0, 0, 0, 
    -1.611419e-05, -2.962841e-05, 0, 0, 0,
  0, 0, 0, 0, 0, 0.00165847, 0.001110366, -0.0003211516, 0, 0, 0.001054551, 
    0, 0, 0, 0, 0, -1.102166e-07, 0.0001161932, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -7.380314e-06,
  0, 0.0009249018, 0.001297515, 0, 0.0009257115, 6.926163e-05, 0.01614421, 
    0.03589895, 0.006531905, 0.0007990189, 0.01334523, 1.4251e-05, 
    -5.33444e-07, 0.0004580262, -2.987724e-05, 0, -5.238988e-05, 0, 0, 0, 0, 
    0, 0, 0.007454987, 0, 0, 0, 0, 0,
  0, 0.0001251125, 0.004577245, -7.785301e-05, -1.501635e-05, 0.04066259, 
    0.01014209, -7.062166e-06, 0.0004801356, 0.001378809, 0.01902615, 
    0.0003760762, -7.243145e-05, 3.75357e-05, 0.01654018, -2.390079e-05, 
    0.003485887, 0, -3.954756e-05, 0, 0, 0, -1.267386e-05, 0.006226389, 
    -5.368778e-05, 0, 0.0003795268, -1.507909e-06, 0,
  0.0004350794, 0, -1.241527e-06, -5.607641e-05, 0, 0, 0.002117877, 
    0.002662601, 0.001812617, 0.006882224, 0.03426128, 0.002575519, 
    0.0100263, 0.004629453, -0.0004251411, -0.0003441787, 0, 0.004107315, 
    0.006328436, 0.001621255, 0, 0.04971137, 0.0119833, 0.004557831, 
    3.018252e-06, -1.553535e-06, 0.0001660688, 1.55011e-05, 0.0002282638,
  0, 0, 0, 0, 0, 0, 0, 0, 0.001330314, -1.860153e-05, 0.008690393, 
    1.704055e-05, -1.118054e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0.0005046058, 0, 
    0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, -4.574964e-05, 0.003537969, 0.004140997, 
    0.00454505, 0.001931414, 0, 0, 0.0007373022, 0, 0, 0, 0, 0, 0, 0, 
    0.006951177, 0.001320998, 0.006190583, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.471029e-05, 0.0003006409, 0.002790685, 
    0.007033158, 0, 0, 0, 0, 0, 0, 0, 0.001355204, 0.005123973, 0, 
    -2.075387e-05, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2.635942e-05, 0.0009844544, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, -8.20127e-08, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, -3.662649e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -4.783789e-06, 0, 0, 0.0009904167, 0, 0, -6.735289e-05, 0, 0, 0,
  -5.064603e-05, 0, 0, 0.0002577172, 0.0007300055, 0.0005589064, 
    -8.81209e-05, 0, 0, 0, 0, 0, 0, 0, 0.000205341, 0.002284991, 0.00378403, 
    7.940417e-07, 0.0008357569, 3.541997e-05, -1.774305e-05, 0.003856421, 0, 
    0, 0.01263622, 0, 0, -1.688417e-05, 0.0003576383,
  0, 0, 0, 0.0001444533, 0, 6.32779e-05, 0, 0, 0, 0, 0, -7.075525e-09, 0, 
    0.005897518, 0.01944209, 0.01159974, 0.002412771, -6.96682e-05, 
    0.006371764, -4.639259e-05, 0.006952037, 0, 0, 0, -6.552818e-05, 
    0.0001497667, 0, 0, 0,
  0, 0, 0, 0, 0, 0.005576264, 0.006504793, -0.0007149756, -6.59647e-06, 0, 
    0.004097805, -3.445201e-08, 0, 0, -4.13562e-06, 0, 0.0004332694, 
    0.0002811952, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -7.845095e-06,
  0, 0.001895819, 0.005559853, 0, 0.002567226, 0.0001102925, 0.02544365, 
    0.06496668, 0.01132144, 0.005918616, 0.03177197, 0.0005764982, 
    -3.2155e-05, 0.005320259, -2.085547e-05, -3.5157e-05, 0.0008841115, 0, 0, 
    0, 0, 0, 0, 0.01424053, -4.662883e-05, 0, 0, -2.171637e-07, 0,
  -2.891155e-05, 0.001368433, 0.005510592, 0.001072462, -0.0001161865, 
    0.06359173, 0.01901267, 7.976382e-06, 0.001328623, 0.006375131, 
    0.03972727, 0.004808974, 0.000217273, 0.0004705106, 0.05475156, 
    -3.022642e-05, 0.007744813, -2.310059e-05, -0.0002099552, 0, 0, 0, 
    -5.797948e-05, 0.01808102, -0.0002708295, -4.763986e-05, 0.005054244, 
    0.0002305103, 2.769154e-06,
  0.0004596402, 0, -2.554853e-06, -0.0001215077, 0, 0, 0.004951072, 
    0.01083566, 0.006038941, 0.02421632, 0.0600617, 0.007646583, 0.02121232, 
    0.01367705, 0.001461937, 0.0002376802, -2.984643e-05, 0.009877913, 
    0.01164875, 0.003430788, 0.0002615819, 0.09259284, 0.03834537, 
    0.007300494, 0.000683391, -9.466788e-05, 0.001006213, 0.0007447624, 
    0.00044475,
  0, 0, 0, 0, 0, 0, 0, 0, 0.007307757, -0.0003082273, 0.01163587, 
    3.684374e-05, 0.006788079, -1.016989e-05, 0, 0, 0.0001133102, 
    0.0001533366, -7.772632e-06, 0, 0, 0, 0.0008542681, 0.0002005999, 0, 0, 
    0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0.002309522, 0.01277158, 0.01047569, 0.02259862, 
    0.008476041, 1.326161e-05, 0, 0.004485541, 0, 0, 0, 0, 0, 0, 
    0.0001439159, 0.01592539, 0.00247619, 0.009074608, 0, 0, 0,
  0, 0, 0, 0, -1.088805e-05, -6.041705e-05, 0.0002006764, 0, 0, 0, 
    0.0001042745, 0.005268177, 0.006832384, 0.01363483, 0, 0, 0, 
    -1.344822e-05, 0, 0, 0, 0.007681682, 0.008218293, -1.700048e-05, 
    0.0006211286, -5.544935e-05, 0, 0, 0,
  0, 0, 0, -5.505131e-05, 0, 0, 0, -3.754201e-06, 0, 0, 7.762132e-05, 
    0.002733604, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2.726743e-05, -5.083499e-05, 0, 
    0, -2.950701e-05, 0, 0, 0,
  0, 5.151124e-09, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 9.170188e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, -3.529941e-05, 0, 0, 0, 0, 0,
  0, -9.777605e-07, 8.293439e-05, 0, 0.002177911, 0, 0, 2.557785e-05, 0, 
    6.017731e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0.0001904321, 0.002242288, 0, 0, 
    0.002104744, 0, 0, -0.0001656613, 0.00140487, -6.722642e-05, -1.669429e-06,
  0.0007417147, 0, 0, 0.004110754, 0.00429506, 0.003765675, 0.002428867, 
    0.0007478084, 1.038238e-05, 0, 0, 0, 0, -1.252213e-05, 0.001802535, 
    0.006302501, 0.00853134, 0.001459826, 0.006724603, 0.003346919, 
    -3.609219e-05, 0.004793148, 0.001105407, -2.238042e-05, 0.01668829, 
    -6.98878e-06, 0, 0.0003559575, 0.002309723,
  0, 0, 0, 0.002099703, -1.853736e-05, 0.006442441, -0.0002884112, 0, 0, 0, 
    -7.805981e-10, -8.764412e-06, 0, 0.01371216, 0.02687222, 0.0242181, 
    0.01095184, 0.008664561, 0.02663708, -0.000299017, 0.009944524, 
    -1.159692e-05, 0, 0, -0.0001576487, 0.005340329, -2.688671e-06, 
    1.384259e-08, 0,
  0, 0, 0, 0, -2.840143e-08, 0.01156617, 0.02690781, -0.0001999425, 
    -3.893857e-05, 0, 0.007179351, -1.498054e-05, -1.172788e-12, 
    -1.592357e-06, 0.001836676, 0.003008259, 0.01107655, 0.009195822, 
    -1.789341e-05, 0, -3.9265e-06, 0, 0, 0, 0, 0, 4.729587e-05, 0, 
    -2.054713e-05,
  0, 0.005268826, 0.007547252, 0, 0.0035218, 0.0005551169, 0.04957143, 
    0.09542916, 0.0248682, 0.0232144, 0.05698805, 0.009489506, -9.932532e-05, 
    0.03551877, -0.0003384371, -0.0001000491, 0.001468482, -9.721548e-08, 
    -4.604391e-07, 0, 0, 0, 6.389348e-11, 0.02545519, 0.003374618, 
    -7.390846e-07, -1.261822e-06, -8.796406e-06, 0,
  0.0004062479, 0.00870438, 0.01948652, 0.007492996, 0.0006614621, 0.1201964, 
    0.03323554, 0.0002697373, 0.01536333, 0.02960075, 0.07584044, 0.02144107, 
    0.004699821, 0.007910656, 0.08874416, 0.006546862, 0.012871, 
    -0.0001340112, 0.001335555, -1.37725e-06, 7.676937e-08, -7.665823e-06, 
    0.0001143466, 0.06632328, 0.003948861, 0.003098888, 0.01952208, 
    0.004981361, 0.0007329608,
  0.001013647, -1.322256e-05, 9.068876e-05, 5.309498e-05, 0, -6.643082e-05, 
    0.0201562, 0.04018895, 0.026688, 0.07294058, 0.1149696, 0.05773948, 
    0.07324956, 0.04570264, 0.006089238, 0.01151244, 0.000387923, 0.02040778, 
    0.02239793, 0.00959056, 0.002040091, 0.1541622, 0.1045005, 0.02194649, 
    0.002555058, 0.0004704041, 0.0009355969, 0.002058106, 0.008986602,
  0, -7.553719e-07, 0, 0, 0, 0, 0, -3.056404e-05, 0.03815972, 0.0007212884, 
    0.01636808, 0.001265837, 0.01714652, -1.327707e-05, 0, 0.0008799126, 
    -6.23096e-06, 0.005234413, 9.130283e-05, 0.001022169, 1.802527e-07, 
    5.537376e-06, 0.004919256, 9.543254e-06, -2.348409e-05, 3.02426e-05, 
    1.045527e-07, 0, 0.0003918986,
  0, 0, 0, 0, 0, 0, 0, 0, 0.009538716, 0.03182886, 0.02077777, 0.04606021, 
    0.03243247, 0.001086442, -1.693079e-05, 0.008702743, -0.0001764545, 0, 0, 
    0, 0, -9.679139e-06, 0.0003629995, 0.03163905, 0.008778356, 0.009872857, 
    0.001101562, 0, 0,
  0, -2.257874e-07, 0, -5.854813e-06, 0.00259048, -0.00024536, 0.002532993, 
    0.0005206101, -9.235205e-06, 1.909136e-05, 0.003454527, 0.01508529, 
    0.03111237, 0.02292418, -3.510964e-07, 0, 0, 0.002394984, 0, 
    1.713412e-05, 0, 0.01071408, 0.0147504, 0.005393553, 0.01066041, 
    0.003887971, 2.764042e-05, 0.0008952454, 0,
  0, 0, -4.095387e-06, 0.0008002558, -1.346514e-05, 0, 0, -7.538998e-05, 0, 
    0, 0.0006585554, 0.00485676, -9.78363e-06, 0.002996452, -1.403458e-05, 0, 
    0, 0, 0, 0, 0, 0.001167654, 0.003102381, -2.659962e-05, 0, -6.209084e-05, 
    0, 0, 0,
  -0.0001252119, 6.037227e-05, 0, 0, 0.002572713, -2.11781e-05, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -4.865262e-06, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001702906, 
    0, -7.442204e-06, 0, 0, 0, 0, 0,
  0, -7.653002e-06, 0, 0, 0, 0.00144244, 0, 1.904605e-05, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001231724, 0, 0, 0, 0, 0,
  -1.515146e-05, 0.00113053, 0.003524444, -4.401652e-05, 0.01211032, 
    0.000391934, 0, 0.0006467344, 0, 0.0005679075, 0, 0, 0, 0.0001711499, 0, 
    0, 0, 0, 0.001964814, 0.001935271, 0.0009263224, 0, 0.004350326, 0, 0, 
    -0.000233189, 0.006330578, -0.0002194585, -3.80353e-05,
  0.008328277, 0.0003656567, 0, 0.01125887, 0.01578225, 0.01103107, 
    0.009339228, 0.003215046, 0.004572154, 0.0005540341, 0, 0, 0, 
    -0.0001187065, 0.004366941, 0.03023546, 0.01498618, 0.01669981, 
    0.02377151, 0.03735405, 0.00665298, 0.01779506, 0.00654741, 0.001880768, 
    0.0204665, 0.002552775, 0.001635862, 0.005987838, 0.007006163,
  -1.660038e-06, -4.873076e-06, 0, 0.005939899, 0.00144118, 0.01511252, 
    0.0008065415, -9.881547e-05, -2.014942e-05, -1.233324e-06, 0.001552879, 
    -7.487806e-05, 0, 0.02293904, 0.040551, 0.06396103, 0.0407216, 
    0.05106714, 0.05539024, 0.005148038, 0.0192264, 0.004882484, 
    0.0005372338, 0.0007839049, -0.0002968769, 0.01587306, 0.002990153, 
    0.002303106, -5.071073e-06,
  4.637002e-05, -4.024414e-06, 0, -1.325236e-10, -1.315325e-06, 0.01469789, 
    0.043393, 0.004006403, 0.00250873, 0.001900875, 0.009005317, 
    0.0001669448, 0.005649478, -2.587522e-05, 0.01563875, 0.01462123, 
    0.02322685, 0.03017273, 0.0005359931, 3.874083e-05, -3.883986e-05, 
    0.0007441542, -8.70591e-07, -4.812328e-10, 0.0004483798, -8.646137e-06, 
    0.001727282, -4.38263e-06, 0.0001871516,
  -2.099161e-05, 0.03355582, 0.01197966, -1.846334e-08, 0.01142746, 
    0.04209379, 0.08720304, 0.1243785, 0.1112172, 0.1021995, 0.1382023, 
    0.07789566, 0.02154969, 0.2567936, 0.04990688, 0.002479756, 0.0005159309, 
    0.001414313, 0.0009519018, 1.932141e-06, 4.475071e-07, -4.908948e-07, 
    -2.089436e-06, 0.04067603, 0.026212, 0.000276425, 3.489787e-07, 
    -3.172234e-05, -3.387268e-07,
  0.01512593, 0.02798138, 0.06748915, 0.0160901, 0.002047432, 0.2348344, 
    0.1399306, 0.1281917, 0.2102143, 0.1763125, 0.2206499, 0.1174994, 
    0.1109174, 0.07608574, 0.1805817, 0.1117064, 0.04619141, 0.007358029, 
    0.009554569, -1.755416e-06, -9.345158e-05, 0.001019769, 0.03000518, 
    0.2230108, 0.08755523, 0.05272824, 0.07545695, 0.02302667, 0.01107958,
  0.001855679, 0.001530222, 0.0004433119, 0.0003165433, -1.008729e-08, 
    -0.0005279905, 0.1436229, 0.2910633, 0.3056229, 0.3480675, 0.2831704, 
    0.2822846, 0.2812345, 0.191914, 0.1406721, 0.1856984, 0.02717153, 
    0.04737099, 0.03134253, 0.02380645, 0.01918409, 0.2439964, 0.2612742, 
    0.1758693, 0.01538006, 0.04359293, 0.001640827, 0.05727101, 0.050891,
  -0.0001037794, -1.646485e-06, 0, 0.001276904, -3.758818e-10, 0, 
    2.67893e-07, 0.007937889, 0.17472, 0.07832681, 0.0584763, 0.05045547, 
    0.1517411, 0.002980448, 0.0003992476, 0.005395411, 0.004078906, 
    0.01657628, 0.0134736, 0.003572223, 0.001188151, 0.00137916, 0.01196095, 
    0.06016149, 0.0009420217, 0.004683679, 0.006295239, 5.195862e-06, 
    -1.868459e-07,
  -4.22075e-09, 9.081232e-05, 9.873457e-05, -8.662109e-06, -5.275068e-05, 0, 
    4.381079e-09, -2.828453e-06, 0.02542524, 0.0807237, 0.07557114, 
    0.1002649, 0.1005566, 0.01325152, 2.698729e-05, 0.01314302, 0.005110434, 
    0, 4.307826e-07, 0, 0, 0.0005868559, 0.001907922, 0.05703535, 0.015693, 
    0.01053473, 0.007733322, -5.042178e-09, -1.767792e-10,
  0.0004062462, 0.003472796, -3.148492e-05, -6.719915e-05, 0.005382418, 
    -0.000350959, 0.005934563, 0.001546668, 2.734833e-06, 0.001595535, 
    0.006266327, 0.03409436, 0.06886081, 0.0476298, 0.00131338, 
    -7.307166e-06, -9.034378e-06, 0.008929888, 0, 0.001402012, 0.00019307, 
    0.0168551, 0.02838109, 0.01862726, 0.03211269, 0.01495748, 0.003451021, 
    0.002793343, 0,
  0.005724191, 0.0001535694, -0.0001230524, 0.001876312, 0.0007289973, 0, 
    -1.48404e-05, -8.988594e-05, 0, -1.198372e-05, 0.002216231, 0.007141638, 
    0.000422423, 0.005045776, 0.00508495, -1.622681e-06, 0, 0.000475103, 0, 
    0, 0, 0.002455225, 0.008933623, 0.0008377621, 0.003310794, 0.001699015, 
    0.0003993315, 0.0009621746, -0.000114425,
  -0.000322727, 0.0001197239, 3.835246e-05, 4.330706e-05, 0.005046974, 
    -1.269634e-05, 0.0002506438, -2.636905e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, -6.286911e-05, -2.642808e-05, 0, 0.003249164, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -4.266799e-06, 0.0003381183, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.005372598, 
    -1.123774e-05, 0.0001406357, 0.0001885667, 0, 0, 0, 0,
  0, -5.422806e-05, 0, -4.078933e-06, 0.0004397138, 0.002176317, 
    -9.324165e-05, 5.184579e-05, -1.57334e-05, 0, 0, -3.867824e-06, 0, 0, 0, 
    0, 0, 0, 0.0003502125, 1.730187e-05, 6.176804e-05, 0.0001971464, 
    0.001025854, 0.003777177, -0.0001612937, 0, 0, 0, -2.870656e-05,
  0.005036482, 0.003520237, 0.006704342, 0.007275262, 0.02842148, 
    0.004935055, 0.003588452, 0.001978798, -7.642344e-05, 0.001657482, 0, 0, 
    -4.42346e-06, 0.001660108, 0.0001894588, 2.695571e-05, 0, 0, 0.006002911, 
    0.009332569, 0.009622493, 9.46119e-05, 0.01452512, 0.002142314, 
    0.008133162, 0.002161891, 0.01060534, 0.002984717, 0.001244663,
  0.01685797, 0.003439947, 0.0001783669, 0.02463178, 0.02978777, 0.0220024, 
    0.01839826, 0.008436496, 0.01061287, 0.002128327, 0.00406519, 
    -4.230655e-05, -4.446242e-05, 0.004161267, 0.0163596, 0.05607182, 
    0.02764909, 0.0464235, 0.05253087, 0.07079221, 0.03105265, 0.04880281, 
    0.01004707, 0.009684541, 0.02138, 0.007205478, 0.003344657, 0.01877097, 
    0.01192582,
  0.0002947304, 0.0007541084, -1.821544e-05, 0.02120433, 0.007649674, 
    0.02263194, 0.009802788, 0.008448089, 0.0001894571, 0.003611324, 
    0.0007848293, 0.006806677, -1.768418e-05, 0.03049494, 0.06535082, 
    0.1637657, 0.1075614, 0.111916, 0.1133721, 0.05099582, 0.04550966, 
    0.01873916, 0.006152386, 0.01115393, -0.0003244338, 0.04817788, 
    0.02114598, 0.007803136, 0.004502325,
  0.005978545, 0.0004261315, 0.0002470645, 3.874643e-05, 0.0001582635, 
    0.01884808, 0.07094761, 0.02317629, 0.01170744, 0.007491047, 0.01462883, 
    9.948661e-05, 0.003056103, -0.0004191316, 0.07055067, 0.05442513, 
    0.07504996, 0.1332159, 0.1143343, 0.01010795, 0.003711342, 0.0004068103, 
    4.451318e-05, 0.001101676, 0.02216579, 0.004821898, 0.03436283, 
    0.001203601, 0.001264107,
  0.001670062, 0.05961173, 0.0354302, -2.386269e-05, 0.01752122, 0.05673871, 
    0.1204566, 0.1187691, 0.07284863, 0.0690845, 0.1346862, 0.04443162, 
    0.01443787, 0.1972342, 0.02751061, 0.001840567, 0.004050582, 0.01683206, 
    0.005681338, -2.926224e-06, 3.549676e-06, 1.707615e-05, 0.003108153, 
    0.2229501, 0.1290121, 0.1037674, 1.367413e-06, 0.001779308, 3.097209e-05,
  0.08782703, 0.2348882, 0.3529918, 0.05894224, 0.04105605, 0.2576094, 
    0.1189254, 0.1031036, 0.2935234, 0.3396846, 0.1948207, 0.08385109, 
    0.05078773, 0.06021303, 0.15396, 0.06988356, 0.05585622, 0.01741458, 
    0.006316857, 0.0004494618, 0.003827938, 0.001644309, 0.06855847, 
    0.329289, 0.103296, 0.08022969, 0.09997637, 0.03131941, 0.05223449,
  0.100212, 0.01170584, 0.03039135, 0.002096027, 0.0005527938, 0.0002140635, 
    0.1135762, 0.2124972, 0.2444637, 0.2670752, 0.2330692, 0.2032654, 
    0.224484, 0.1636286, 0.1552019, 0.2556444, 0.1204558, 0.1220572, 
    0.1217329, 0.07123619, 0.04290317, 0.3201602, 0.3887197, 0.2964791, 
    0.03690819, 0.08260427, 0.04398208, 0.03918495, 0.1542652,
  0.0570775, 0.007563244, -2.419202e-05, 0.04111405, -1.471293e-05, 0, 
    0.001972464, 0.004169314, 0.2047695, 0.05693552, 0.06404395, 0.02810082, 
    0.1588665, 0.07433596, 0.03403588, 0.05755792, 0.06353751, 0.08975919, 
    0.1529125, 0.05170007, 0.02720446, 0.005432466, 0.04972952, 0.2248662, 
    0.1151696, 0.1231765, 0.02527304, 0.02648086, 0.05041426,
  0.005354072, 0.001230411, 0.001331014, 3.093131e-05, 0.01099554, 
    0.0001484676, -5.354008e-05, -1.186071e-05, 0.05462466, 0.1850829, 
    0.1705022, 0.2648582, 0.2228563, 0.05959917, 0.01201792, 0.0251948, 
    0.01530075, 0.0009968609, 0.00650033, -7.668144e-06, 0.002645855, 
    0.004025479, 0.01636644, 0.1051466, 0.0784696, 0.02118889, 0.03395356, 
    0.00788508, -0.0001328673,
  0.002773602, 0.008346907, 0.006747989, 0.003927128, 0.01295753, 
    0.004582084, 0.01299755, 0.004820222, 0.0007241578, 0.006318243, 
    0.02902663, 0.08045276, 0.1633927, 0.1594057, 0.07599678, 0.03597426, 
    0.01595808, 0.02240834, -8.200235e-10, 0.001933286, 0.0004728912, 
    0.02438522, 0.04153534, 0.04359672, 0.05995622, 0.03749594, 0.007527156, 
    0.006487711, 0.0005742246,
  0.0170819, 0.001337506, -0.0002915024, 0.003158247, 0.002277717, 
    0.0002603912, 0.001418458, -3.856114e-05, 0, -2.615202e-05, 0.007668264, 
    0.01661492, 0.01197045, 0.03449613, 0.02846173, 0.002654555, 
    7.643014e-05, 0.01591584, -5.712173e-07, 0, 0, 0.006852045, 0.01850037, 
    0.003800742, 0.01104639, 0.007693076, 0.0007767986, 0.000618409, 
    0.005005195,
  0.0002040199, 0.0005601913, 7.385921e-05, 0.001594348, 0.009812087, 
    0.001896914, 0.001996813, -4.590267e-05, 0, 0, 0, -5.946794e-06, 
    0.0005090627, -2.413723e-06, -9.174016e-05, 0, 0, 0, 0, 0, 0.0007586008, 
    0.003571191, -3.153275e-06, 0.007207082, -1.623037e-05, 0, 0, 0, 
    -1.734461e-05,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0008056875, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.278691e-05, -1.027327e-05, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -4.266799e-06, 0.0003381183, -4.515333e-05, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.995017e-05, 
    6.467438e-06, 0.006849812, 0.009179909, 9.563259e-05, 0.001234218, 0, 0, 
    0, 0,
  0.001415224, 0.002694794, 0.001273124, 0.002279749, 0.001394774, 
    0.003210924, 2.146262e-05, 0.0007978583, 0.000259897, 0, 0.002136029, 
    0.0001083061, -7.817121e-05, 0, 0, -8.280325e-06, 0, 0, 0.001945013, 
    0.002068336, 0.006941023, 0.01218701, 0.005404088, 0.01501934, 
    0.006206817, 0.0007619853, 0, -6.551502e-08, -0.0001243493,
  0.02251133, 0.007370968, 0.01209711, 0.01709686, 0.04342137, 0.01766129, 
    0.01081469, 0.008262988, 0.006724662, 0.0070824, 0.003746006, 
    0.001570802, 0.003581606, 0.001593954, 0.002409408, 0.0004744793, 
    0.0009972784, 0.001657024, 0.009955501, 0.02802689, 0.02210588, 
    0.007490376, 0.03823483, 0.01860253, 0.01556986, 0.00836479, 0.02102604, 
    0.01291382, 0.01487105,
  0.03069286, 0.008670128, 0.009121034, 0.04194935, 0.05070809, 0.04890116, 
    0.03910338, 0.02810808, 0.02975039, 0.02029286, 0.0224734, 0.001820666, 
    0.002103192, 0.01691875, 0.05729996, 0.08405937, 0.04501367, 0.07857824, 
    0.09379466, 0.1377157, 0.09800512, 0.09786572, 0.03841545, 0.04110738, 
    0.02781272, 0.03452183, 0.03940465, 0.0620133, 0.03178459,
  0.02926483, 0.007533288, 0.0132109, 0.02496013, 0.03973574, 0.03915133, 
    0.03653245, 0.01280127, 0.01833016, 0.01896528, 0.02645309, 0.004922674, 
    -9.199283e-05, 0.03868975, 0.09582154, 0.2275359, 0.2095479, 0.16165, 
    0.2276151, 0.1827516, 0.1332323, 0.0586966, 0.04106519, 0.04328337, 
    0.0173514, 0.09613148, 0.05490724, 0.03307616, 0.02750601,
  0.0004926652, 0.007275471, 0.0008930076, 9.914991e-05, 0.0005405043, 
    0.01917553, 0.06547214, 0.02797745, 0.01332061, 0.01288989, 0.01637941, 
    1.732299e-06, 0.002016904, -0.0003908886, 0.08706728, 0.05730493, 
    0.07660104, 0.1434925, 0.05803249, 0.0006782589, 0.003167724, 
    8.999484e-05, 1.683938e-05, 6.011505e-05, 0.01269629, 0.0004119416, 
    0.01681936, 0.0009142332, 8.486034e-05,
  0.001131987, 0.05275257, 0.02640653, -3.660402e-05, 0.01310271, 0.03424377, 
    0.1000205, 0.1035166, 0.04948534, 0.04197135, 0.1170029, 0.02659103, 
    0.01023412, 0.1491354, 0.01711477, 0.002260871, 0.002347027, 0.01165977, 
    0.001242962, -1.78412e-06, 3.58132e-06, -1.497635e-07, 4.924011e-05, 
    0.1671248, 0.06597605, 0.06070164, 1.293691e-05, 0.0001000254, 1.49762e-05,
  0.07071988, 0.1974495, 0.2753873, 0.03973255, 0.02244343, 0.2003275, 
    0.09323899, 0.05086171, 0.2246793, 0.2494512, 0.1904038, 0.07416552, 
    0.0301043, 0.04552382, 0.1355894, 0.04857273, 0.04824369, 0.043555, 
    0.01836776, -8.382445e-05, 0.001545002, 5.061442e-05, 0.04451359, 
    0.2900735, 0.07311139, 0.04782503, 0.07313523, 0.02491174, 0.03493378,
  0.06419782, 0.00468121, 0.03436163, 0.02809922, 0.0001252936, 0.0002161373, 
    0.08438295, 0.1634827, 0.2157192, 0.2145306, 0.21141, 0.1505475, 
    0.1862434, 0.1410999, 0.09282129, 0.212422, 0.08043853, 0.09130326, 
    0.06090281, 0.05161076, 0.02914774, 0.2739551, 0.3284007, 0.2392233, 
    0.02571181, 0.05743829, 0.02510715, 0.03388501, 0.1138694,
  0.07400519, 0.006284474, 0.007065024, 0.03119617, 3.014965e-06, 
    -2.010392e-12, 0.01606343, 0.003305338, 0.1425613, 0.04383556, 0.0605919, 
    0.01655078, 0.1194474, 0.0465719, 0.01776982, 0.06988988, 0.07008298, 
    0.1062377, 0.1616847, 0.0251778, 0.01482965, 0.0105185, 0.05455345, 
    0.1993953, 0.1148754, 0.1312629, 0.02422725, 0.02187608, 0.03843193,
  0.04592355, 0.0928745, 0.04032381, 0.006858258, 0.08163142, 0.001253396, 
    0.008904921, -4.812552e-05, 0.097793, 0.1658237, 0.1603031, 0.2667505, 
    0.2284479, 0.0723419, 0.01231145, 0.1354437, 0.1066358, 0.08687515, 
    0.061474, 0.03470741, 0.01947198, 0.1251758, 0.04255306, 0.1289858, 
    0.1227921, 0.1331337, 0.1073076, 0.06283621, 0.04567726,
  0.0202287, 0.01573404, 0.01884501, 0.01340718, 0.02571305, 0.03247057, 
    0.01904725, 0.01106056, 0.0167328, 0.02863476, 0.06631668, 0.1299562, 
    0.2579281, 0.2576447, 0.166104, 0.1319166, 0.09137076, 0.1038252, 
    0.01631195, 0.009767759, 0.00153921, 0.03882058, 0.05671917, 0.09450044, 
    0.1307264, 0.07211743, 0.04846255, 0.03854413, 0.01981126,
  0.03185657, 0.005901882, 0.002784734, 0.01017507, 0.006546154, 0.009525521, 
    0.001570049, 0.001310565, -2.219555e-05, 0.0005724306, 0.02086127, 
    0.0279679, 0.06542019, 0.1068369, 0.1554236, 0.08877143, 0.02991483, 
    0.02805487, 0.01283413, -9.564083e-10, -2.683138e-06, 0.01656157, 
    0.0341157, 0.01124056, 0.02994003, 0.0289182, 0.02367149, 0.01325582, 
    0.01908801,
  0.0007874686, 0.004390724, 0.003936302, 0.00995683, 0.01587321, 
    0.008565912, 0.003265766, 0.001258391, 0, 0, 0, 2.488874e-05, 
    0.0006489341, 0.003233914, 0.007669693, 0.005406141, 0, 0.0003662588, 
    0.0009447563, -5.787135e-07, 0.001979206, 0.008162764, -0.0001408769, 
    0.01434734, 0.0008395493, 0.002560692, -4.533651e-09, 0, -0.0002235675,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5.699263e-05, -3.27545e-08, 0, 0, 
    -0.0001838835, 0.01019685, -1.836415e-06, 0, 0, -9.842427e-06, 
    3.047609e-05, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5.771628e-06, 0.0005582077, 
    0.002640487, 0.0009503114, 0.0001958353, 6.277384e-10, 1.482712e-09, 
    -4.370886e-07, -4.861209e-06, 0.0007456874, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0003089918, -5.669753e-05, 0.0004143931, -0.000232164, -3.07457e-05, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0.0001447018, 4.00252e-05, 0, 0, 
    0, 0.001193468, 0.000105122, 0.009317549, 0.013438, 0.00296782, 
    0.01103222, -7.515344e-05, 0, 0, 0,
  0.005853044, 0.005177211, 0.004053759, 0.009587852, 0.003557339, 
    0.006204456, 0.001261203, 0.001523937, 0.001316785, 0.003177798, 
    0.003793202, 0.00460206, 0.003318206, 0.0002224329, 0, 0.002172522, 
    0.001028574, 0, 0.009191571, 0.01032307, 0.01159055, 0.02084471, 
    0.024376, 0.03485622, 0.01961147, 0.004789511, 6.273625e-05, 
    -9.665253e-05, 0.0008024095,
  0.03685673, 0.01364301, 0.02365916, 0.03145637, 0.08778607, 0.06586646, 
    0.04343928, 0.03658065, 0.01659195, 0.0390098, 0.03174437, 0.02987403, 
    0.01103609, 0.002954973, 0.007143713, 0.02205717, 0.01316268, 0.02391479, 
    0.02882047, 0.05270171, 0.08195124, 0.06645287, 0.1127042, 0.05912204, 
    0.04725377, 0.03789164, 0.0501242, 0.03821737, 0.04354021,
  0.1252427, 0.09821371, 0.08511131, 0.1218542, 0.1325898, 0.1114689, 
    0.07457002, 0.07734947, 0.08148227, 0.07477597, 0.07766807, 0.04335796, 
    0.01789401, 0.02824141, 0.08616283, 0.134634, 0.0835933, 0.09651829, 
    0.1450195, 0.2171836, 0.1863171, 0.2535866, 0.1561218, 0.1032354, 
    0.1092563, 0.07680084, 0.1050908, 0.1211648, 0.0899654,
  0.05130042, 0.04020513, 0.01097819, 0.03322006, 0.08676869, 0.05314776, 
    0.06120545, 0.04058581, 0.03218101, 0.04182738, 0.0502606, 0.006914484, 
    0.0004001778, 0.0482642, 0.1267258, 0.2097, 0.2244741, 0.1501693, 
    0.2149051, 0.1537743, 0.1439798, 0.04035268, 0.02579594, 0.05032685, 
    0.02943714, 0.0968565, 0.07468197, 0.04527435, 0.05086341,
  6.167221e-06, 0.003592922, 0.0006350496, 0.001177549, 0.0009147294, 
    0.03839155, 0.06167163, 0.02114846, 0.01837114, 0.003845606, 0.02026546, 
    0.0001048517, 0.002590641, 0.002018676, 0.08373133, 0.04104349, 
    0.07105394, 0.1108945, 0.02267535, 2.649829e-05, 0.000363039, 
    -6.428864e-05, 2.615548e-07, 5.110264e-05, 0.005950949, 0.0005486747, 
    0.02024667, 0.0001604537, 3.299759e-06,
  0.0007197834, 0.06137316, 0.02481261, -7.759274e-06, 0.01563159, 
    0.02657511, 0.0835155, 0.101105, 0.04368586, 0.0336419, 0.1128301, 
    0.02093633, 0.008614266, 0.1242242, 0.01726459, 0.002009877, 0.003085448, 
    0.005895026, 7.036057e-05, 5.177823e-08, 1.516731e-06, 8.731166e-08, 
    1.178417e-05, 0.1102557, 0.02989988, 0.04179001, 0.0001249797, 
    -1.497768e-05, 8.300506e-06,
  0.05037476, 0.1766713, 0.2221206, 0.03685022, 0.02207444, 0.1761228, 
    0.08960681, 0.03100927, 0.1832067, 0.1986041, 0.1793606, 0.05753186, 
    0.03230669, 0.04752349, 0.1217291, 0.03621808, 0.03434762, 0.03828859, 
    0.02036598, -2.742859e-06, 0.0003332529, 1.575789e-05, 0.01682541, 
    0.2494188, 0.05584244, 0.03941847, 0.06317864, 0.02248872, 0.02360217,
  0.04257992, 0.00598912, 0.0476423, 0.02194362, 0.0006993827, 0.001041065, 
    0.07508728, 0.1334445, 0.1904107, 0.1762483, 0.1947161, 0.1109655, 
    0.1581438, 0.1200618, 0.06666305, 0.155827, 0.05256283, 0.08570776, 
    0.03185739, 0.03940317, 0.03213917, 0.2558286, 0.2539352, 0.2141497, 
    0.02433529, 0.05101954, 0.0114002, 0.02663141, 0.104977,
  0.07630706, 0.002809535, 0.00579681, 0.02164965, -1.509438e-06, 0, 
    0.01349607, 0.0004037052, 0.1188161, 0.03225556, 0.0436989, 0.0125089, 
    0.09861688, 0.02910793, 0.007049564, 0.03993525, 0.06369385, 0.08015841, 
    0.1319934, 0.01644457, 0.007500105, 0.007779307, 0.05709467, 0.1844539, 
    0.1149533, 0.1241694, 0.0213208, 0.02402464, 0.0127779,
  0.04137542, 0.1263498, 0.08103779, 0.04378766, 0.07525041, 0.0008083926, 
    0.01294572, 0.000344497, 0.160872, 0.1554305, 0.158758, 0.2384684, 
    0.2113818, 0.06760112, 0.01668002, 0.1189137, 0.1008968, 0.07070866, 
    0.06109161, 0.02644854, 0.1119595, 0.08204649, 0.0372673, 0.1304814, 
    0.1147923, 0.1152435, 0.09646851, 0.04651846, 0.04348616,
  0.1128821, 0.08579589, 0.07211921, 0.04499795, 0.08647716, 0.1178999, 
    0.02884382, 0.1212519, 0.08281426, 0.08526286, 0.1164528, 0.1538666, 
    0.2464881, 0.2510757, 0.1551392, 0.1640512, 0.157028, 0.2386869, 
    0.07573095, 0.0844342, 0.02111545, 0.1511329, 0.1142395, 0.187236, 
    0.1945909, 0.1249586, 0.09646517, 0.08591752, 0.0807386,
  0.08988914, 0.04318735, 0.01680407, 0.05978023, 0.06828622, 0.06209361, 
    0.02595128, 0.004994217, 0.0005187631, 0.008114262, 0.06224443, 
    0.1121303, 0.1109773, 0.1620527, 0.214669, 0.1641345, 0.06519385, 
    0.1113935, 0.1246685, 0.002413076, 0.01248099, 0.06585661, 0.07484204, 
    0.05257244, 0.1433284, 0.114084, 0.03164085, 0.02298368, 0.03252456,
  0.01815893, 0.004930125, 0.01010105, 0.02715664, 0.02684251, 0.03473804, 
    0.02770005, 0.01390536, -0.0002361943, 4.902017e-06, -2.66752e-05, 
    -0.0001765595, 0.004715648, 0.06467974, 0.07249943, 0.03847613, 
    -0.0004668521, 0.004918625, 0.001202467, 0.01103855, 0.007531898, 
    0.02247724, -0.0005469777, 0.03529585, 0.0404886, 0.01605888, 
    0.009467708, -5.048086e-05, 0.002928971,
  0, 0, 0, -3.439675e-06, 7.276883e-05, 4.615076e-05, 0, 0, 0, 0, 0, 0, 0, 
    0.005616536, 0.01765408, 0.01969902, 0.001619223, 0.007484592, 
    0.000764091, 0.01314784, -0.0001781768, -1.132411e-05, -8.630296e-06, 
    -2.840792e-05, 0.01396716, -9.203372e-06, 0, 2.767656e-10, -8.273613e-07,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.205662e-09, 7.757767e-06, 0.0003711626, 
    0.004311141, 0.02746938, 0.03043137, 0.01702536, 0.01684117, 0.01634952, 
    0.01107792, 0.0008953002, 0.00252878, 0.0003388115, -1.6426e-06, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.001869012, 0.004772467, 0.005803086, 0.0008850791, 0.000248435, 
    -7.996271e-05, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -4.189674e-05, -6.162477e-05, 
    0.001481465, 0.0003121323, 2.001786e-05, 0.0006609734, 0, 0.006090379, 
    0.01711934, 0.03633708, 0.05443341, 0.03852038, 0.02249469, 
    -0.0002281836, 0.001116347, -1.305144e-06, -1.266816e-06,
  0.01187747, 0.00812629, 0.01037668, 0.01605638, 0.01570806, 0.0127861, 
    0.01978233, 0.005713055, 0.01032299, 0.008133409, 0.009393812, 0.0133481, 
    0.02789558, 0.0009272852, 0.0001912184, 0.01831469, 0.02176932, 
    0.0001556893, 0.02469794, 0.0247591, 0.0161367, 0.04810289, 0.0502022, 
    0.0654704, 0.05459039, 0.02784479, 0.01599514, 0.006561932, 0.003234003,
  0.09454703, 0.07213517, 0.07974594, 0.1288233, 0.2302095, 0.164302, 
    0.1083804, 0.1074246, 0.1114733, 0.1102203, 0.1191672, 0.08949759, 
    0.05739373, 0.07405762, 0.1152513, 0.1094344, 0.1238777, 0.1029089, 
    0.09786421, 0.07790451, 0.1116877, 0.1246248, 0.1684426, 0.1172172, 
    0.1017945, 0.1509811, 0.1263264, 0.08472149, 0.1183982,
  0.1437045, 0.1246276, 0.1261347, 0.1768986, 0.1512588, 0.1220427, 
    0.07993986, 0.0902295, 0.1010519, 0.1041238, 0.1209452, 0.09311596, 
    0.06785582, 0.1142363, 0.1300623, 0.1797245, 0.1366433, 0.1103795, 
    0.1572186, 0.2406536, 0.1940464, 0.2590286, 0.1810993, 0.1748984, 
    0.1601521, 0.08301236, 0.129894, 0.1454726, 0.104878,
  0.03937437, 0.0145326, 0.01429251, 0.02800828, 0.07537034, 0.03716465, 
    0.06996407, 0.01784311, 0.02286352, 0.03367914, 0.05083151, 0.007888641, 
    0.0002533854, 0.05284659, 0.1341451, 0.2027273, 0.1860375, 0.1407313, 
    0.2013558, 0.1275891, 0.1245863, 0.03301789, 0.0181511, 0.03534262, 
    0.01833232, 0.1055221, 0.06848677, 0.0439491, 0.06878414,
  2.364206e-07, 0.000108183, 0.0001565218, 0.002681005, 0.0003495306, 
    0.0429622, 0.05417836, 0.01095641, 0.03277263, 0.004535479, 0.0323278, 
    0.00651444, 0.01570853, 0.02118186, 0.07767552, 0.0524802, 0.06847571, 
    0.08987769, 0.01522478, 1.310342e-05, 0.0001673857, 3.464692e-05, 
    -4.212117e-10, 0.0002819863, 0.00586259, 0.003199674, 0.02569232, 
    -6.378774e-05, 3.925992e-07,
  0.0002001707, 0.04893588, 0.02328044, 7.556118e-05, 0.02164226, 0.02303424, 
    0.07238454, 0.1001874, 0.0351731, 0.02503934, 0.1106929, 0.01742223, 
    0.01536092, 0.08292919, 0.01510222, 0.001751862, 0.002787714, 
    0.004315212, 1.800608e-05, 1.217376e-08, 1.187187e-06, -1.799811e-09, 
    -1.486979e-06, 0.08233611, 0.01269607, 0.01644356, 0.006348037, 
    1.740762e-05, 1.172813e-05,
  0.03725207, 0.1416534, 0.164917, 0.04845982, 0.01725186, 0.150039, 
    0.08110026, 0.02345256, 0.1205962, 0.1586691, 0.1691097, 0.04553578, 
    0.0332686, 0.04003091, 0.1081715, 0.03572011, 0.0309123, 0.03672977, 
    0.0189725, -2.774327e-05, 0.0001829461, 5.442641e-06, 0.003887124, 
    0.2142657, 0.04646179, 0.02882338, 0.04642018, 0.02211435, 0.01392562,
  0.04238673, 0.01033949, 0.03850053, 0.02032101, 0.0006958945, 0.001787778, 
    0.05724395, 0.1055768, 0.1668915, 0.1395718, 0.1892053, 0.08169104, 
    0.1483608, 0.09843317, 0.04731062, 0.1149156, 0.03892971, 0.07913418, 
    0.03570731, 0.03209517, 0.02594439, 0.2374693, 0.1850219, 0.1599538, 
    0.02650661, 0.0341318, 0.004923054, 0.01895702, 0.09324335,
  0.06523159, -0.0002473606, 0.001752441, 0.008951702, -2.848303e-06, 0, 
    0.01868564, 6.376731e-05, 0.100684, 0.02967789, 0.04880287, 0.00815666, 
    0.08288708, 0.01406835, 0.005451153, 0.03260089, 0.04283429, 0.06922692, 
    0.08458462, 0.005540533, 0.01477546, 0.008341097, 0.06045629, 0.1672899, 
    0.08102589, 0.1310934, 0.007152382, 0.028005, 0.005104747,
  0.04110883, 0.1061915, 0.07751643, 0.05137656, 0.05104537, 0.0003384585, 
    0.01270347, 0.00348521, 0.3021244, 0.1563121, 0.1647672, 0.2172945, 
    0.2083577, 0.05857165, 0.01522798, 0.088262, 0.08274329, 0.05620274, 
    0.05146923, 0.02224817, 0.09020861, 0.04680067, 0.02879423, 0.1280284, 
    0.1188264, 0.09721728, 0.08005365, 0.03428341, 0.02822696,
  0.1836772, 0.1059386, 0.08449969, 0.1032415, 0.07533076, 0.09195418, 
    0.04481957, 0.1501857, 0.0972587, 0.1416291, 0.104503, 0.1377145, 
    0.2073383, 0.2433204, 0.1549068, 0.1371971, 0.1581021, 0.2256471, 
    0.06685999, 0.09150009, 0.0944142, 0.1308051, 0.1159385, 0.1648914, 
    0.1994857, 0.162921, 0.1390919, 0.1306328, 0.119068,
  0.2118751, 0.0856773, 0.08439997, 0.09323494, 0.1135813, 0.1218213, 
    0.1015024, 0.0109536, 0.0150401, 0.05141466, 0.1096147, 0.1716792, 
    0.1474731, 0.1755003, 0.2072911, 0.2033722, 0.1145416, 0.1826164, 
    0.1788434, 0.04122009, 0.06598595, 0.111418, 0.1406463, 0.1081865, 
    0.1943874, 0.1362361, 0.07515837, 0.07460659, 0.1743068,
  0.03010242, 0.01532058, 0.02875744, 0.1029835, 0.1191166, 0.117234, 
    0.1032583, 0.1197583, 0.02793858, 0.003364761, 0.01362184, 0.02970291, 
    0.05275637, 0.2243925, 0.1305559, 0.08281086, 0.04490036, 0.04236171, 
    0.05362646, 0.04505927, 0.04739638, 0.07402528, 0.0634472, 0.07786927, 
    0.1000794, 0.1668675, 0.073843, 0.1087625, 0.08173792,
  0.03281168, 0.01639993, 0.0008774965, -0.0003374614, 0.01217033, 
    0.02771398, 0.04595648, 0.02132086, 0.01870543, 0.004202676, 0, 
    -3.998719e-10, 0.006316519, 0.01980687, 0.05880697, 0.06063254, 
    0.03355667, 0.03276532, 0.02925799, 0.06527701, 0.04633907, 0.03913224, 
    0.09155726, 0.05430514, 0.04599548, 2.606029e-05, -7.549871e-07, 
    0.03395024, 0.05712158,
  0, 7.406152e-05, 0.007276201, 0.009307562, 0.00714966, 5.307213e-05, 0, 
    -5.99493e-07, -4.421016e-05, 0.0008804296, 0.003563961, 0.00787927, 
    0.02260259, 0.02131884, 0.03119933, 0.03682186, 0.04193975, 0.01912495, 
    0.01994979, 0.02193593, 0.03070218, 0.02065302, 0.009020586, 0.000773965, 
    0.0004220028, -3.31741e-06, -4.765282e-07, -0.000163532, 3.565798e-05,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.476329e-05, 
    -2.716438e-05, 0.0091146, 0.0337289, 0.03339534, 0.03717099, 0.03926067, 
    -0.001791802, 0,
  0, 0, -1.561284e-05, -7.608485e-09, 0, 0, 0, 0, 0, 0, 0, -2.841594e-05, 
    8.935779e-05, 0.01063454, 0.02105582, 0.02037378, 0.01713352, 
    0.004686422, -1.029943e-05, 0.01105473, 0.02677125, 0.08115754, 
    0.08413538, 0.07192949, 0.05065918, 0.02179987, 0.009859974, 0.00928051, 
    0.0007812851,
  0.02957813, 0.02314796, 0.02312816, 0.03311711, 0.05870632, 0.03744538, 
    0.03897372, 0.03301378, 0.04347319, 0.03249791, 0.0559147, 0.07564201, 
    0.1269595, 0.1641503, 0.1081736, 0.1130037, 0.1164406, 0.04483631, 
    0.07270778, 0.06242573, 0.06722459, 0.1218713, 0.1205238, 0.1343676, 
    0.1067519, 0.07203393, 0.06042718, 0.07049274, 0.01975504,
  0.1320757, 0.1281118, 0.1520619, 0.2387755, 0.2616594, 0.2175901, 
    0.1660708, 0.1615972, 0.1523939, 0.1896041, 0.1991788, 0.1757062, 
    0.210505, 0.1327097, 0.1595709, 0.1582958, 0.1371424, 0.1431057, 
    0.1467029, 0.1048953, 0.1388936, 0.1454414, 0.2249632, 0.1634726, 
    0.1755587, 0.1828321, 0.175551, 0.1580158, 0.1700549,
  0.1313975, 0.1181869, 0.1193218, 0.1659189, 0.144235, 0.09698061, 
    0.07266088, 0.07204285, 0.1025884, 0.1117221, 0.1372054, 0.1210633, 
    0.08787385, 0.1007555, 0.1553664, 0.1879175, 0.132878, 0.1036539, 
    0.1853779, 0.2352612, 0.1941351, 0.2310443, 0.1776711, 0.1930152, 
    0.1794545, 0.09872068, 0.1280049, 0.1655646, 0.1040511,
  0.02034425, 0.003421297, 0.01250514, 0.02681572, 0.0695687, 0.03316952, 
    0.0681209, 0.02166583, 0.02991224, 0.02995116, 0.03008401, 0.001486682, 
    0.0001148876, 0.0589577, 0.1368516, 0.1867894, 0.1485234, 0.1432448, 
    0.1819029, 0.1098304, 0.1222856, 0.04845559, 0.006328794, 0.01813516, 
    0.01695568, 0.0895859, 0.0510646, 0.03793, 0.0477425,
  5.91714e-08, 8.557876e-06, 2.882526e-05, 0.004159197, 0.0001218659, 
    0.02796028, 0.05137458, 0.008747534, 0.01768376, 0.007834786, 0.04878459, 
    0.006284838, 0.001544176, 0.05067841, 0.07157364, 0.03864719, 0.06426167, 
    0.08737847, 0.01142239, 8.026397e-06, 0.0006715519, 2.745348e-05, 
    -4.788694e-09, 0.006279884, 0.0086266, 0.004834646, 0.03069792, 
    8.019846e-05, 9.628644e-08,
  3.6388e-05, 0.04342723, 0.01567395, 0.0001029272, 0.02352803, 0.02613754, 
    0.05828315, 0.09868614, 0.03057583, 0.02404818, 0.1258238, 0.01514872, 
    0.02095661, 0.05312982, 0.01309332, 0.002542031, 0.002740641, 
    0.002384756, 8.021657e-06, 6.166833e-07, 5.731007e-07, -2.983115e-09, 
    -1.157568e-06, 0.06114656, 0.004816032, 0.003411047, 0.01638143, 
    1.999502e-06, 1.033586e-05,
  0.02845703, 0.1489069, 0.1402895, 0.04891137, 0.01325362, 0.1265156, 
    0.0756752, 0.01876798, 0.0687335, 0.1299178, 0.1528686, 0.03612182, 
    0.02359567, 0.02615388, 0.0871581, 0.03044509, 0.02906607, 0.02493781, 
    0.00402606, -0.0001461807, 0.000146199, 1.37549e-06, 0.003830002, 
    0.1725157, 0.04931175, 0.02283852, 0.03838466, 0.01553986, 0.00892994,
  0.02875199, 0.01001385, 0.0206553, 0.02428734, 0.0009752823, 0.00137381, 
    0.03938318, 0.07718246, 0.1371523, 0.110325, 0.1851489, 0.06086628, 
    0.1282823, 0.07100774, 0.03011489, 0.07023016, 0.02276813, 0.06135123, 
    0.04854064, 0.0259611, 0.01471056, 0.2004438, 0.1361108, 0.1058655, 
    0.01274811, 0.02294123, 0.002172717, 0.01242, 0.08384389,
  0.04823508, -4.12955e-05, 8.714915e-05, 0.0009035158, -2.541248e-06, 0, 
    0.008230852, 0.0001782645, 0.08325798, 0.03200299, 0.05564378, 
    0.004971691, 0.05843593, 0.01068528, 0.004658243, 0.02730158, 0.03847094, 
    0.05187876, 0.03077752, 0.0005731269, 0.004475162, 0.007819954, 
    0.04707908, 0.1510401, 0.1064049, 0.1338421, 0.002725513, 0.01831635, 
    0.001152078,
  0.03087603, 0.07022006, 0.06179192, 0.03511488, 0.03011065, 0.0001055845, 
    0.01856507, 0.02573462, 0.3193566, 0.1627987, 0.165326, 0.2135309, 
    0.2084119, 0.04727521, 0.01776024, 0.07725938, 0.06889916, 0.0474674, 
    0.04068281, 0.02137879, 0.07308543, 0.02782631, 0.0197973, 0.1097046, 
    0.1144651, 0.07814761, 0.06004917, 0.02413299, 0.0170769,
  0.1855334, 0.1143648, 0.07774497, 0.1442967, 0.06157436, 0.07197071, 
    0.07861944, 0.1208215, 0.08409506, 0.1399046, 0.09048335, 0.1350334, 
    0.182358, 0.2423722, 0.1588503, 0.1271541, 0.1386061, 0.2137407, 
    0.04821624, 0.07571129, 0.09560252, 0.1181187, 0.1171265, 0.1473462, 
    0.1697137, 0.1437858, 0.1323947, 0.123082, 0.1087651,
  0.2395278, 0.1814972, 0.1260973, 0.1610936, 0.1251681, 0.1137735, 
    0.1131526, 0.04086701, 0.07625856, 0.1251025, 0.1473028, 0.215351, 
    0.1534629, 0.1797833, 0.2096641, 0.2265974, 0.1444973, 0.1876956, 
    0.1655455, 0.1295393, 0.1137327, 0.1306089, 0.2015506, 0.2017165, 
    0.1974746, 0.1316755, 0.1314919, 0.1543762, 0.2395075,
  0.06474217, 0.03387995, 0.04168298, 0.1578581, 0.2193433, 0.1597963, 
    0.1391303, 0.1569859, 0.1110171, 0.05191486, 0.09949507, 0.07437181, 
    0.1066167, 0.2626588, 0.1704566, 0.09166681, 0.1365982, 0.09253892, 
    0.07979873, 0.06911034, 0.08797096, 0.1233816, 0.1023597, 0.09946625, 
    0.1963615, 0.2340512, 0.1178183, 0.2650259, 0.1381785,
  0.08572858, 0.02070025, 0.0052752, 0.03383619, 0.04648617, 0.05630599, 
    0.1059066, 0.03189989, 0.01885249, 0.01591816, -1.145651e-05, 
    0.008331036, 0.03263065, 0.08871432, 0.10039, 0.07759563, 0.05182469, 
    0.06621016, 0.06873779, 0.1085545, 0.06781881, 0.05788482, 0.1300347, 
    0.1150287, 0.08252559, 0.003034226, -0.0001808801, 0.1599012, 0.1410694,
  0.00459586, 0.01208798, 0.01458671, 0.01090542, 0.02204622, 0.008559927, 
    0.01590589, 0.02606014, 0.02451649, 0.04355091, 0.03809865, 0.03188182, 
    0.02529166, 0.0228245, 0.02807791, 0.05164849, 0.06321775, 0.04963205, 
    0.05620573, 0.05995413, 0.05508516, 0.06111985, 0.03151641, 0.01780115, 
    0.01656298, 0.002974176, -0.00161633, 0.007508947, 0.01602805,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2.655457e-08, 0, 0, 0, 
    -7.38515e-05, -0.0003758019, -0.0002960888, 0.03050112, 0.08784648, 
    0.0926808, 0.05043873, 0.06609558, 0.03227606, 0.0002313635,
  0.001514661, 0.02146904, 0.0112709, 0.0006906966, -8.544294e-05, 0, 
    -2.338684e-06, 0, 0, -9.449675e-05, -1.120506e-05, -0.0003808655, 
    0.01714145, 0.1018233, 0.1050902, 0.06826509, 0.0625957, 0.04454807, 
    0.01615457, 0.03128723, 0.06285772, 0.1444839, 0.1373184, 0.1198068, 
    0.102987, 0.07419819, 0.06953707, 0.0557301, 0.02124373,
  0.08353992, 0.08098396, 0.08638802, 0.09160686, 0.1095775, 0.09427362, 
    0.07488181, 0.08626448, 0.09866283, 0.09628346, 0.147113, 0.1832454, 
    0.2681716, 0.2852505, 0.1839295, 0.243306, 0.2498759, 0.145698, 
    0.2342958, 0.1487505, 0.1306176, 0.1527068, 0.1830116, 0.1897949, 
    0.1754346, 0.1576559, 0.1368387, 0.1781712, 0.08066481,
  0.1694452, 0.1418911, 0.1751865, 0.2497823, 0.2579689, 0.199193, 0.1708544, 
    0.1701877, 0.1872537, 0.2159675, 0.2507124, 0.2354314, 0.1892949, 
    0.1088449, 0.1322619, 0.1524018, 0.1370106, 0.1588598, 0.1882354, 
    0.1245944, 0.1647689, 0.1826338, 0.2705885, 0.1939157, 0.1645335, 
    0.2083793, 0.1779565, 0.1604435, 0.1826046,
  0.1500911, 0.1273597, 0.1077011, 0.1484914, 0.1302832, 0.09177241, 
    0.06168259, 0.06010837, 0.09600204, 0.1070166, 0.1271042, 0.1163702, 
    0.09397212, 0.07237488, 0.1588151, 0.173446, 0.1424254, 0.08643428, 
    0.1669995, 0.2203951, 0.1683247, 0.218792, 0.1687252, 0.1920297, 
    0.1749285, 0.0984387, 0.1295972, 0.1495697, 0.09530318,
  0.006335171, 0.0009381395, 0.00690563, 0.02448881, 0.065018, 0.02678419, 
    0.07520121, 0.03160148, 0.02205458, 0.02091074, 0.01118471, 1.867666e-05, 
    0.001637362, 0.0521511, 0.1310486, 0.1759813, 0.1562233, 0.1487806, 
    0.1606735, 0.1048801, 0.1307941, 0.04126855, 0.001808157, 0.009742295, 
    0.01486035, 0.08049872, 0.04432417, 0.04138264, 0.03625752,
  2.698337e-08, 1.97208e-05, -7.562337e-06, 0.01089068, 0.0002838131, 
    0.0323945, 0.05640027, 0.007797432, 0.02306882, 0.006503233, 0.04595116, 
    0.01663188, 0.0002523605, 0.05344049, 0.06133645, 0.02980402, 0.05565074, 
    0.07643031, 0.007164956, 1.731207e-06, 0.0006372841, 1.772552e-05, 
    -3.78349e-09, 0.01978048, 0.01194084, 0.003581937, 0.02973729, 
    0.005175121, 1.747876e-08,
  -2.733972e-05, 0.03457861, 0.007700147, 0.0007508069, 0.03138652, 
    0.02323282, 0.04949347, 0.09728885, 0.02956969, 0.01635893, 0.119311, 
    0.0149767, 0.02849534, 0.02895223, 0.01174087, 0.0038345, 0.002516785, 
    0.001828648, 8.37581e-06, 1.372516e-06, 1.247447e-07, -2.478184e-10, 
    9.734559e-07, 0.05826806, 0.002924357, 0.002189212, 0.02540125, 
    -1.436521e-05, 6.150319e-07,
  0.02292289, 0.1301472, 0.1324922, 0.05673815, 0.01154332, 0.1179082, 
    0.08056181, 0.0158635, 0.05243287, 0.1171329, 0.1431746, 0.03081634, 
    0.01649638, 0.01908754, 0.07367889, 0.02637434, 0.02666004, 0.01695303, 
    -8.406497e-05, 0.0002903677, 0.0009893476, 1.4312e-07, 0.01587801, 
    0.1424904, 0.05298555, 0.01979986, 0.04442472, 0.01545482, 0.006390877,
  0.02890963, 0.007148436, 0.01672324, 0.02680802, 0.0007126377, 0.001934928, 
    0.03039306, 0.07808878, 0.1148512, 0.0967859, 0.1884076, 0.04731308, 
    0.1115771, 0.04989308, 0.02180529, 0.07060279, 0.01817137, 0.03040922, 
    0.04951769, 0.02402481, 0.008586399, 0.1718806, 0.09483199, 0.07360962, 
    0.008969892, 0.01344152, 0.006945667, 0.007680015, 0.07576995,
  0.04135722, -5.672996e-05, 6.305726e-06, 0.0001885391, -2.339742e-06, 
    -1.109461e-10, 0.00509367, 0.0002945468, 0.06453271, 0.03172158, 
    0.04137264, 0.003957956, 0.04808479, 0.01017714, 0.00329229, 0.02351732, 
    0.02546199, 0.04980679, 0.003094031, -4.996193e-06, 0.001986133, 
    0.006935457, 0.03559161, 0.1358246, 0.08238762, 0.06877854, 0.001490959, 
    0.0136479, 0.0003389565,
  0.01979648, 0.0580231, 0.05547825, 0.03170197, 0.02042532, 5.523727e-05, 
    0.02573544, 0.08303969, 0.3289415, 0.1574467, 0.1420446, 0.2078224, 
    0.1781568, 0.0393731, 0.01053776, 0.07378059, 0.06359942, 0.04856143, 
    0.02504105, 0.01224615, 0.05425817, 0.01735551, 0.0149262, 0.09417825, 
    0.08763877, 0.06183591, 0.04194298, 0.0131509, 0.009176234,
  0.1808862, 0.1104725, 0.05891339, 0.1370559, 0.06332164, 0.06823056, 
    0.123795, 0.09785096, 0.07362435, 0.1239927, 0.07996573, 0.1356111, 
    0.176208, 0.2414619, 0.1278153, 0.0976813, 0.1147496, 0.2186623, 
    0.04579053, 0.07467153, 0.0807115, 0.1127618, 0.1023787, 0.1266456, 
    0.1711521, 0.1348321, 0.1404076, 0.1097121, 0.1062182,
  0.2165508, 0.1828125, 0.1353866, 0.1406155, 0.1201756, 0.1162587, 
    0.0935427, 0.0571547, 0.1200163, 0.1474275, 0.2080262, 0.2344774, 
    0.1597674, 0.1684203, 0.2007069, 0.2245199, 0.1737879, 0.1975154, 
    0.1714936, 0.1359333, 0.1130156, 0.1210428, 0.185079, 0.2017419, 
    0.1902765, 0.1172934, 0.1279561, 0.1596106, 0.2312334,
  0.08581547, 0.08437101, 0.04584508, 0.1682381, 0.2208929, 0.2341422, 
    0.2153422, 0.2333916, 0.1419337, 0.1301261, 0.1510071, 0.09910913, 
    0.1469979, 0.3478086, 0.1568771, 0.09084703, 0.1732941, 0.1310116, 
    0.1244852, 0.1115255, 0.1410989, 0.2371607, 0.1425859, 0.09301641, 
    0.2170525, 0.239158, 0.1144547, 0.2677763, 0.1253718,
  0.1931261, 0.08546367, 0.02679104, 0.0662198, 0.094539, 0.09090029, 
    0.1279623, 0.05265261, 0.0420025, 0.05748068, 0.007786679, 0.08648852, 
    0.1215482, 0.1822498, 0.1024518, 0.1224851, 0.06262936, 0.09825404, 
    0.1299065, 0.08111063, 0.09653163, 0.06869034, 0.1732983, 0.123838, 
    0.1401815, 0.01441483, 8.878294e-06, 0.2337413, 0.2394523,
  0.05756544, 0.04143408, 0.04619626, 0.04602926, 0.1018548, 0.08205245, 
    0.06320742, 0.08851352, 0.08277626, 0.07916921, 0.07815447, 0.1369116, 
    0.1510104, 0.1820058, 0.162139, 0.1205098, 0.1151358, 0.09330016, 
    0.08563258, 0.08118147, 0.09505773, 0.1200559, 0.07426284, 0.04407058, 
    0.04358989, 0.02006502, 0.01565997, 0.02648291, 0.08493736,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  -0.0001745938, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.480566e-05, 
    8.709339e-05, -2.591956e-05, 0.0005456773, -6.792094e-05, -1.187588e-06, 
    -0.0005230905, 0.000937301, 0.002320423, 0.06132552, 0.1414251, 
    0.1673532, 0.1169502, 0.123111, 0.06615938, 0.001600671,
  0.02584411, 0.08001429, 0.05818302, 0.01468487, -0.0004825717, 
    -3.627155e-05, 0.01175418, 0, 0, -0.0003342082, -6.512018e-05, 
    0.001464939, 0.05399364, 0.1446712, 0.1872036, 0.1380393, 0.1266859, 
    0.08522649, 0.06566883, 0.05694528, 0.09469433, 0.1573804, 0.1938748, 
    0.2138817, 0.2052893, 0.1547167, 0.2360428, 0.1611918, 0.07343733,
  0.2177095, 0.1403262, 0.1249367, 0.1056089, 0.1443778, 0.1409672, 
    0.1288386, 0.1250184, 0.1450678, 0.1453568, 0.2126946, 0.2765053, 
    0.2917032, 0.3142907, 0.1856289, 0.2470951, 0.2611683, 0.1545703, 
    0.2658874, 0.2343015, 0.1903857, 0.2321509, 0.2213313, 0.2514974, 
    0.232421, 0.208626, 0.1671308, 0.2879563, 0.1823995,
  0.1705932, 0.1563895, 0.1951973, 0.2340592, 0.2454941, 0.1974137, 
    0.1584278, 0.1683751, 0.2043532, 0.2234043, 0.272252, 0.2572038, 
    0.1846628, 0.1090323, 0.1321606, 0.1561299, 0.1344779, 0.151615, 
    0.1939233, 0.148238, 0.1716403, 0.2047025, 0.2915055, 0.1836528, 
    0.1632281, 0.1983367, 0.1839997, 0.1637188, 0.187628,
  0.1795945, 0.1235381, 0.1096811, 0.1391659, 0.1126278, 0.08758723, 
    0.05813116, 0.0809122, 0.1039396, 0.08249788, 0.1117117, 0.1083799, 
    0.09135338, 0.06378304, 0.1361296, 0.1738273, 0.1466008, 0.08268024, 
    0.1509773, 0.2106349, 0.1488159, 0.2519288, 0.1416677, 0.1896727, 
    0.1810256, 0.08503129, 0.1290291, 0.1386828, 0.09333206,
  0.0003538854, 0.004022099, 0.00387437, 0.02610129, 0.05349766, 0.0170665, 
    0.07521802, 0.01652748, 0.03498841, 0.02735851, 0.008899691, 
    2.629376e-05, 0.00269591, 0.05480995, 0.1292361, 0.1754031, 0.1283021, 
    0.1437613, 0.1526716, 0.0883322, 0.1274747, 0.05649321, 0.007627395, 
    0.00493594, 0.01621196, 0.07180057, 0.04387768, 0.04325864, 0.03606845,
  9.845015e-09, 1.255438e-05, 0.0004065823, 0.01431521, 0.00274598, 
    0.03865303, 0.07514425, 0.005706235, 0.0189052, 0.009113857, 0.05727835, 
    0.02080001, 0.002695466, 0.06807564, 0.03650381, 0.02492201, 0.05955118, 
    0.06336213, 0.01024078, 5.622854e-06, 0.0006392903, 1.504541e-05, 
    -9.724465e-10, 0.02448428, 0.0127922, 0.001043776, 0.02705014, 
    0.005407254, 2.928447e-08,
  -6.185621e-05, 0.03287128, 0.003042422, 0.00430073, 0.02011249, 0.02401951, 
    0.044225, 0.09791417, 0.02943707, 0.0176596, 0.1187113, 0.02330983, 
    0.03290588, 0.0196088, 0.01105377, 0.005991744, 0.002533149, 0.001243314, 
    4.088434e-06, -4.940879e-08, 3.4739e-09, 0, 8.696481e-06, 0.04230839, 
    0.00256222, 0.001817297, 0.02726393, 3.450998e-06, 4.474793e-06,
  0.02282089, 0.1451682, 0.119176, 0.08112489, 0.01444045, 0.107685, 
    0.08643595, 0.01310679, 0.04188485, 0.1155447, 0.132349, 0.03218085, 
    0.01372851, 0.01554768, 0.06823866, 0.02755578, 0.02536372, 0.0171025, 
    0.01533449, -0.0003943311, 3.117665e-05, -3.309751e-08, 0.04260582, 
    0.1160301, 0.05777595, 0.0254376, 0.05936258, 0.01422219, 0.003848208,
  0.02178745, 0.0099455, 0.02581285, 0.03480887, 0.001570141, 0.004047011, 
    0.02439488, 0.06385904, 0.1023717, 0.09173324, 0.1870438, 0.04664904, 
    0.09409925, 0.04225366, 0.01587532, 0.09226543, 0.009967878, 0.01024267, 
    0.04764357, 0.02254686, 0.006296764, 0.1534301, 0.07952465, 0.06036135, 
    0.007649528, 0.01232689, 0.01166278, 0.00821962, 0.06828701,
  0.04777512, -8.251819e-05, 1.524107e-06, 0.0001171863, -9.414862e-07, 
    -3.38248e-10, 0.00443266, 0.0003953324, 0.07915934, 0.04265474, 
    0.03405111, 0.005120426, 0.03981017, 0.006774239, 0.003201009, 
    0.02516243, 0.03326119, 0.0538375, 0.00368788, -7.833579e-06, 
    0.0001330034, 0.005647107, 0.03108696, 0.1478785, 0.07515873, 0.04600505, 
    0.001624641, 0.02286637, 0.000107798,
  0.007630907, 0.05194176, 0.041993, 0.03415716, 0.0142728, -1.946487e-05, 
    0.03144891, 0.1399878, 0.3329817, 0.1548857, 0.1285119, 0.1958575, 
    0.1917708, 0.0306602, 0.004190712, 0.07056785, 0.05333816, 0.02677592, 
    0.01947295, 0.008007518, 0.02405089, 0.01197527, 0.01406423, 0.08701555, 
    0.07029074, 0.06413565, 0.03402093, 0.004187863, 0.00292419,
  0.1690063, 0.1215697, 0.0560826, 0.1249231, 0.05535027, 0.06185476, 
    0.1055248, 0.08889998, 0.06299438, 0.123341, 0.08725933, 0.1455933, 
    0.1754511, 0.2427001, 0.1133281, 0.08957766, 0.106679, 0.2024676, 
    0.05392444, 0.06332698, 0.07495928, 0.1158871, 0.08841018, 0.1135458, 
    0.1728109, 0.1162531, 0.129549, 0.1089908, 0.1206082,
  0.1879793, 0.1665776, 0.1218133, 0.1282264, 0.1155903, 0.09978877, 
    0.08021457, 0.07351843, 0.1334454, 0.1583978, 0.2183617, 0.2360006, 
    0.1555918, 0.153091, 0.2138635, 0.2005027, 0.1988718, 0.1842709, 
    0.1849137, 0.1452016, 0.1060101, 0.1295827, 0.1636282, 0.1965642, 
    0.2025424, 0.1232205, 0.1110596, 0.1342902, 0.2243602,
  0.09749251, 0.08884757, 0.06175184, 0.1590351, 0.2034375, 0.2343773, 
    0.1999499, 0.2194408, 0.2245328, 0.1809702, 0.1788949, 0.1039604, 
    0.1707182, 0.3515816, 0.1437967, 0.08663509, 0.2322148, 0.1853783, 
    0.1898405, 0.1451727, 0.2125117, 0.2373314, 0.1455479, 0.08369052, 
    0.2233702, 0.2284521, 0.1125709, 0.2524539, 0.1156534,
  0.178382, 0.1031771, 0.05464859, 0.07016979, 0.1028624, 0.1165752, 
    0.178226, 0.07590762, 0.07590034, 0.1469017, 0.08048593, 0.2003568, 
    0.1836442, 0.2017943, 0.09425092, 0.128083, 0.06849835, 0.1326882, 
    0.170146, 0.1020139, 0.1087749, 0.1051289, 0.192171, 0.1376043, 
    0.1386222, 0.08827244, 0.01617198, 0.2390693, 0.2267743,
  0.09641629, 0.09325118, 0.1198104, 0.1156732, 0.1580784, 0.1385573, 
    0.1204865, 0.1301313, 0.1264302, 0.1098467, 0.1208156, 0.1625672, 
    0.148191, 0.1673802, 0.1585661, 0.118362, 0.1185504, 0.09285255, 
    0.08473424, 0.1164069, 0.148091, 0.161457, 0.1279321, 0.05748278, 
    0.07070844, 0.03334059, 0.04134524, 0.08471525, 0.1380686,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  -0.002553057, -6.159259e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01379766, 
    0.01332147, 0.007513035, 0.008052507, 0.005879184, 0.001184591, 
    -0.001162861, 0.007866969, 0.0131064, 0.1220101, 0.3142819, 0.3012336, 
    0.2056593, 0.2036822, 0.07791577, 0.02392038,
  0.0591832, 0.1571008, 0.1227613, 0.06161075, -0.002042261, -0.001718344, 
    0.04515802, -1.993993e-06, -1.546441e-05, -0.001784125, 0.001770093, 
    0.005690958, 0.1116986, 0.1882676, 0.1988441, 0.171439, 0.1719459, 
    0.1552169, 0.1522184, 0.1835685, 0.2284312, 0.2093816, 0.2710133, 
    0.3497223, 0.3329568, 0.2755805, 0.3292598, 0.2752154, 0.2028872,
  0.2717995, 0.1885773, 0.1760275, 0.1642227, 0.2366697, 0.1705575, 
    0.1807822, 0.1902143, 0.2269957, 0.2436837, 0.2714758, 0.2994177, 
    0.3036246, 0.3125444, 0.1769361, 0.2339832, 0.24623, 0.1647912, 
    0.2888137, 0.2817949, 0.2552742, 0.290262, 0.2430073, 0.270225, 
    0.2581099, 0.2063193, 0.2151002, 0.343139, 0.2307356,
  0.1605538, 0.155186, 0.2179739, 0.2276415, 0.2288096, 0.1917019, 0.1572286, 
    0.1619217, 0.2281209, 0.2339156, 0.2953652, 0.2573563, 0.1830714, 
    0.08545044, 0.1086454, 0.1461527, 0.1296562, 0.1288992, 0.1797706, 
    0.1419893, 0.1629027, 0.2122948, 0.2692743, 0.1821875, 0.1539255, 
    0.1975965, 0.1733239, 0.1539641, 0.1885615,
  0.1689408, 0.100011, 0.09743305, 0.1142906, 0.1021634, 0.07877652, 
    0.06551193, 0.07855595, 0.08142653, 0.09364047, 0.1245686, 0.105848, 
    0.08501961, 0.06009496, 0.1307915, 0.1656741, 0.1455984, 0.09132832, 
    0.1342833, 0.1828418, 0.1261631, 0.2201053, 0.1311084, 0.1844537, 
    0.1455481, 0.07384674, 0.1300952, 0.1423248, 0.09620532,
  -1.267635e-05, 0.0004077101, 0.001373751, 0.0283932, 0.0394141, 0.01565687, 
    0.06717736, 0.005933686, 0.03511, 0.0156332, 0.01674324, 0.0003546328, 
    0.00747034, 0.0563819, 0.1135189, 0.1625387, 0.1214784, 0.1348875, 
    0.1412446, 0.08730096, 0.1080236, 0.06273735, 0.003156635, 0.004599852, 
    0.01868015, 0.06096601, 0.04489832, 0.04678919, 0.03234274,
  -3.142293e-07, 5.636783e-06, 0.004752477, 0.01694583, 0.005245968, 
    0.04779658, 0.07144526, 0.004580584, 0.03119551, 0.000929553, 0.07268625, 
    0.02181952, 0.001693241, 0.112367, 0.0252304, 0.0176103, 0.04164872, 
    0.05698716, 0.008132862, 1.541494e-05, 0.0006273528, 1.942364e-06, 
    -1.275721e-08, 0.01325209, 0.01548702, 0.0003367726, 0.02595833, 
    0.0002288082, 5.231083e-10,
  1.280677e-05, 0.03090116, 0.0009502261, 0.009064503, 0.02636429, 
    0.02863272, 0.03560434, 0.09895128, 0.03007912, 0.01439366, 0.1008955, 
    0.03142059, 0.03621637, 0.01718969, 0.0118156, 0.006026801, 0.002685021, 
    0.0009481185, 1.377343e-06, -1.94856e-09, -1.604071e-09, 3.185151e-11, 
    0.001557164, 0.04056584, 0.002410382, 0.005120666, 0.006453047, 
    1.295776e-05, 1.413403e-05,
  0.02045744, 0.1237313, 0.1185304, 0.08568744, 0.02121783, 0.1202388, 
    0.08880361, 0.01274359, 0.0329326, 0.09891102, 0.1270542, 0.033238, 
    0.01081068, 0.01603783, 0.06344131, 0.03355367, 0.02783311, 0.02201474, 
    0.007936972, 0.01042554, -0.000188205, -6.641063e-06, 0.04009199, 
    0.1164757, 0.0500962, 0.03378189, 0.04847058, 0.02379029, 0.004641478,
  0.01743816, 0.01701874, 0.041579, 0.0352836, 0.002853516, 0.004276535, 
    0.01679158, 0.067099, 0.09594718, 0.08976486, 0.1957784, 0.04613084, 
    0.08153033, 0.03501056, 0.0127669, 0.09476307, 0.01755311, 0.0129603, 
    0.02957225, 0.02276518, 0.00546873, 0.1438631, 0.07961039, 0.05333247, 
    0.006260792, 0.01687287, 0.01078603, 0.006637877, 0.07219433,
  0.01980904, -2.383678e-05, 1.134991e-06, 0.001252015, -1.800731e-08, 
    2.934336e-08, 0.003604572, 0.0005134442, 0.07408408, 0.05774368, 
    0.03468847, 0.007389383, 0.04114016, 0.003801659, 0.003148246, 
    0.03179875, 0.03216444, 0.05288223, -7.21137e-05, -1.089314e-05, 
    2.359271e-06, 0.006606096, 0.03800266, 0.1443236, 0.04842964, 0.03533887, 
    0.003738042, 0.01264807, -2.554475e-05,
  0.006012697, 0.02822496, 0.03143587, 0.03130201, 0.01224744, 6.359935e-05, 
    0.01019932, 0.1423381, 0.339525, 0.1439619, 0.1228482, 0.169482, 
    0.183148, 0.02611593, 0.002722146, 0.07561633, 0.05279556, 0.01612705, 
    0.01543762, 0.001407274, 0.006873287, 0.01118673, 0.01528441, 0.0796994, 
    0.05061468, 0.06582137, 0.03401034, 0.000585378, 0.0005364516,
  0.1387989, 0.1127004, 0.0529287, 0.1173263, 0.03969628, 0.0504837, 
    0.1013526, 0.07813303, 0.05371097, 0.1195904, 0.08815987, 0.1402641, 
    0.1650763, 0.2306596, 0.1024652, 0.0858214, 0.09664758, 0.175135, 
    0.04423173, 0.04546205, 0.0938447, 0.1195858, 0.08090471, 0.1022757, 
    0.1731561, 0.1179051, 0.1242954, 0.09768428, 0.1272278,
  0.1653489, 0.1406079, 0.1143062, 0.1213019, 0.1044933, 0.08465019, 
    0.07524489, 0.08824236, 0.1644273, 0.1546399, 0.2357655, 0.2177987, 
    0.1522457, 0.1370208, 0.2098966, 0.1822479, 0.2094409, 0.1791297, 
    0.1814206, 0.1605693, 0.1005358, 0.1339145, 0.1571932, 0.2028014, 
    0.2034566, 0.1260756, 0.1046593, 0.1118528, 0.2113735,
  0.1003705, 0.08926912, 0.06321723, 0.1641975, 0.1919979, 0.2423755, 
    0.1968222, 0.202601, 0.2454858, 0.2248819, 0.1953531, 0.1906601, 
    0.1721054, 0.3557221, 0.1373247, 0.08325783, 0.2379812, 0.2224529, 
    0.2481669, 0.1894864, 0.2142942, 0.2571231, 0.147276, 0.09760044, 
    0.2112424, 0.1950209, 0.1113497, 0.2344491, 0.1122119,
  0.1718679, 0.09570069, 0.07464442, 0.0689541, 0.1253012, 0.147535, 
    0.2299347, 0.1154595, 0.07582248, 0.1650349, 0.08850197, 0.3375444, 
    0.2071363, 0.2129925, 0.09302068, 0.1322667, 0.05612782, 0.1602697, 
    0.1898662, 0.1346503, 0.1113872, 0.1027622, 0.1837157, 0.138382, 
    0.1368913, 0.1708579, 0.03908591, 0.2408094, 0.2102624,
  0.08702307, 0.09273993, 0.1171746, 0.1707052, 0.1542735, 0.1365209, 
    0.1249523, 0.1255821, 0.1045424, 0.1041915, 0.1263768, 0.1460501, 
    0.1340316, 0.1448459, 0.1641038, 0.1088793, 0.1395684, 0.1659226, 
    0.08656464, 0.1137615, 0.136176, 0.1589544, 0.1337856, 0.05364098, 
    0.09761626, 0.0649578, 0.07001515, 0.1113618, 0.1396516,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -4.244298e-05, -4.244298e-05, 
    -4.244298e-05, -4.244298e-05, -4.244298e-05, -4.244298e-05, 
    -4.244298e-05, -3.596705e-05, -3.596705e-05, -3.596705e-05, 
    -3.596705e-05, -3.596705e-05, -3.596705e-05, -3.596705e-05, 0,
  0.01601959, -0.0001822365, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.000573932, 
    0.04693751, 0.05578991, 0.03803725, 0.05925771, 0.03081229, 0.0206854, 
    0.01409091, 0.03886132, 0.03464662, 0.2032936, 0.4647357, 0.3935527, 
    0.3014689, 0.2319496, 0.138545, 0.06523827,
  0.07355985, 0.1398278, 0.2770374, 0.1614577, 0.0005079767, -0.003523632, 
    0.09828272, -0.001435216, -0.001123633, 0.004013701, 0.008906585, 
    0.01425085, 0.1722704, 0.1912383, 0.2321765, 0.2141694, 0.2100096, 
    0.2228878, 0.2526041, 0.3220122, 0.3015819, 0.2964172, 0.3219176, 
    0.4283502, 0.351095, 0.2882567, 0.3380595, 0.3105213, 0.2500676,
  0.271158, 0.2234279, 0.2008055, 0.229295, 0.2931858, 0.1675016, 0.1812994, 
    0.1821202, 0.2451137, 0.2392657, 0.2908349, 0.3040343, 0.3016111, 
    0.3198636, 0.1782674, 0.2189143, 0.2475118, 0.1640445, 0.2970108, 
    0.2926607, 0.2881238, 0.2932099, 0.2470305, 0.2667256, 0.24647, 
    0.1991248, 0.2198228, 0.3554122, 0.2236268,
  0.1684355, 0.1578887, 0.230888, 0.2242367, 0.2343984, 0.1954811, 0.1591912, 
    0.1727355, 0.2453206, 0.2382597, 0.2956559, 0.2576351, 0.1675063, 
    0.09098164, 0.09531343, 0.1135325, 0.1104776, 0.1131417, 0.1704526, 
    0.1238419, 0.1845155, 0.2069212, 0.261938, 0.1659997, 0.1459915, 
    0.1864938, 0.1665829, 0.145447, 0.1945958,
  0.1559058, 0.09333962, 0.1013575, 0.106733, 0.1025928, 0.06805849, 
    0.05970205, 0.06682876, 0.06577867, 0.08379438, 0.09607176, 0.09362912, 
    0.0636102, 0.06302364, 0.1112064, 0.1619007, 0.1442511, 0.08845226, 
    0.1072552, 0.1776379, 0.1105681, 0.2100911, 0.1175864, 0.1736979, 
    0.1298371, 0.07163762, 0.1276718, 0.1217072, 0.09009843,
  -3.122277e-05, 0.000384413, 0.001458714, 0.03078771, 0.03562448, 
    0.01570494, 0.05383578, 0.004006556, 0.03434945, 0.01096041, 0.005943099, 
    0.001131889, 0.01903202, 0.05722648, 0.1028698, 0.1484256, 0.1069769, 
    0.1329129, 0.1389365, 0.08608948, 0.0985636, 0.06118569, 0.0002073087, 
    0.005935626, 0.02250816, 0.05576154, 0.0488039, 0.04922071, 0.02287694,
  -3.269217e-06, -3.95699e-05, 0.007377144, 0.0102716, 0.01548658, 
    0.05328546, 0.04955455, 0.02540918, 0.01744909, 0.002450643, 0.1007739, 
    0.01064317, 9.563567e-05, 0.1599201, 0.02146078, 0.01452372, 0.02252582, 
    0.04881385, 0.005227721, 2.043011e-05, 0.0003726335, -3.489375e-06, 
    -5.246573e-07, 0.001602289, 0.0252487, 0.0002119307, 0.02609567, 
    5.337976e-06, 1.025152e-08,
  0.0001252151, 0.03100198, 0.0002931538, 0.01234328, 0.03985411, 0.04768251, 
    0.0323149, 0.1049136, 0.03310608, 0.02102811, 0.1073877, 0.04513896, 
    0.04457775, 0.01637981, 0.01282017, 0.004941044, 0.003483635, 
    0.001063259, 1.888436e-06, 2.561154e-08, 7.090004e-09, 1.258205e-08, 
    0.01527704, 0.0310376, 0.003138729, 0.002250231, -0.0005116416, 
    3.17639e-05, 4.681607e-05,
  0.03023536, 0.11938, 0.1307196, 0.08289351, 0.01429894, 0.1240526, 
    0.09287193, 0.01405916, 0.02557227, 0.08835447, 0.1212649, 0.03282267, 
    0.01026553, 0.01620709, 0.05993063, 0.02831194, 0.02490943, 0.03092514, 
    0.004814387, 0.01822287, -0.0001364921, 0.002302572, 0.04540384, 
    0.1389904, 0.07900914, 0.03424023, 0.03999501, 0.02400127, 0.004231146,
  0.01511115, 0.02924458, 0.03668869, 0.04641941, 0.002506836, 0.003135312, 
    0.01616135, 0.07696518, 0.09982147, 0.1147452, 0.2067783, 0.04709596, 
    0.0926673, 0.03965633, 0.01293374, 0.1024821, 0.02646354, 0.01430726, 
    0.02401739, 0.02148189, 0.006747394, 0.1318625, 0.08960053, 0.05883582, 
    0.006194846, 0.01836459, 0.01498232, 0.00578147, 0.07907443,
  0.01006771, 6.029787e-07, 3.524495e-07, 0.001789378, -2.410684e-08, 
    3.916168e-08, 0.00446833, 0.001573364, 0.0845664, 0.06805563, 0.04889747, 
    0.01393852, 0.04252401, 0.004165447, 0.002654635, 0.03669634, 0.02916525, 
    0.02421302, 0.0004121571, -1.661794e-05, 3.553857e-06, 0.006069948, 
    0.04340809, 0.1642132, 0.02589194, 0.02497892, 0.0001641955, 0.01679608, 
    -3.585068e-05,
  0.005832251, 0.009420888, 0.02828068, 0.0267909, 0.01776537, 0.0006283487, 
    -0.001762996, 0.1630271, 0.3435711, 0.148477, 0.1062061, 0.1413514, 
    0.1780332, 0.04076025, 0.003574112, 0.0642109, 0.03395607, 0.02118636, 
    0.00391152, -2.695467e-05, 0.009787577, 0.01018383, 0.01572786, 
    0.07912319, 0.04368491, 0.04387705, 0.02517422, 0.000764381, 2.811134e-07,
  0.1123152, 0.08583416, 0.04850344, 0.1129193, 0.02701644, 0.03757503, 
    0.09643301, 0.06441277, 0.04037014, 0.1215529, 0.0934452, 0.1164314, 
    0.1581696, 0.2204274, 0.1038786, 0.0801191, 0.07361849, 0.1611907, 
    0.04164401, 0.02959903, 0.1044118, 0.1020508, 0.0938698, 0.1010505, 
    0.1677247, 0.09538073, 0.1141177, 0.08877908, 0.1136927,
  0.1614281, 0.1236029, 0.1230133, 0.113711, 0.1066405, 0.07685432, 
    0.07503281, 0.1301318, 0.1776379, 0.1522808, 0.2378003, 0.198544, 
    0.1488709, 0.1254912, 0.1934652, 0.1741813, 0.1625588, 0.1772049, 
    0.1727686, 0.1607003, 0.1039099, 0.1284237, 0.1449514, 0.199271, 
    0.1948681, 0.1209137, 0.1039977, 0.1009847, 0.1778233,
  0.09048088, 0.1047613, 0.06889021, 0.1690298, 0.1798897, 0.2395357, 
    0.2024538, 0.1933584, 0.2382079, 0.2219581, 0.1978264, 0.2065435, 
    0.1626864, 0.3626189, 0.1497153, 0.08360343, 0.2341161, 0.2344151, 
    0.2799395, 0.1894464, 0.211902, 0.2815849, 0.157204, 0.1134023, 
    0.2014561, 0.1726843, 0.1037817, 0.2125924, 0.1013973,
  0.1686541, 0.08113898, 0.07713945, 0.07279033, 0.1289268, 0.1430481, 
    0.259553, 0.1445096, 0.1180357, 0.2254355, 0.1809783, 0.2961342, 
    0.1925989, 0.199089, 0.09822704, 0.1263133, 0.04319124, 0.1611095, 
    0.1920384, 0.1438424, 0.1184287, 0.1088095, 0.1652234, 0.1433427, 
    0.1325361, 0.2466142, 0.0834604, 0.2383004, 0.1816935,
  0.08202026, 0.09417141, 0.1185185, 0.1734591, 0.1455225, 0.1230201, 
    0.09810022, 0.07715023, 0.06835882, 0.08622117, 0.1361697, 0.1522596, 
    0.1355894, 0.1388501, 0.1609911, 0.1139491, 0.14899, 0.1579731, 
    0.08476886, 0.0842803, 0.1188384, 0.1539539, 0.1339594, 0.03834279, 
    0.09143137, 0.09383149, 0.1433782, 0.1066533, 0.1410936,
  8.814842e-05, 5.609445e-05, 2.404048e-05, -8.013493e-06, -4.006747e-05, 
    -7.212144e-05, -0.0001041754, -0.0005092011, -0.0003581718, 
    -0.0002071424, -5.6113e-05, 9.491637e-05, 0.0002459457, 0.0003969751, 
    -0.0004035154, -0.0004713947, -0.000539274, -0.0006071533, -0.0006750326, 
    -0.0007429118, -0.0008107912, -9.495707e-05, -0.0001460532, 
    -0.0001971493, -0.0002482454, -0.0002993415, -0.0003504376, 
    -0.0004015337, 0.0001137916,
  0.04672474, 0.0002231111, -0.0001033206, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.003535937, 0.1037379, 0.07858134, 0.09224063, 0.1827515, 0.09055749, 
    0.05368462, 0.04281919, 0.07536374, 0.08893699, 0.3031337, 0.4887273, 
    0.3788674, 0.2996314, 0.2213732, 0.1933131, 0.08047409,
  0.06800518, 0.07889978, 0.3037197, 0.2662957, 0.01321153, 0.01964866, 
    0.1322938, 0.004954875, 0.01424451, 0.02897521, 0.05636514, 0.04360618, 
    0.2081704, 0.2003055, 0.2433421, 0.2167252, 0.2137663, 0.2383571, 
    0.2717915, 0.332931, 0.3105803, 0.3160695, 0.3632104, 0.4301904, 
    0.3337905, 0.2859251, 0.3269928, 0.32965, 0.2469736,
  0.2831956, 0.2270004, 0.2080722, 0.2466971, 0.2788047, 0.1875215, 
    0.2122929, 0.2158305, 0.3016666, 0.268575, 0.2970393, 0.3080422, 
    0.3012839, 0.3055849, 0.1948313, 0.2088935, 0.2554062, 0.1817219, 
    0.3249871, 0.2850609, 0.2657157, 0.2606224, 0.2244216, 0.2715023, 
    0.2515072, 0.2065872, 0.2356338, 0.3480773, 0.2387452,
  0.1647903, 0.1610099, 0.2310974, 0.2270679, 0.2283129, 0.1913559, 
    0.1621381, 0.1937178, 0.2483787, 0.2509909, 0.2853206, 0.2432351, 
    0.1508694, 0.06392469, 0.08055842, 0.1127518, 0.1134611, 0.0971121, 
    0.1733345, 0.1416964, 0.2026074, 0.1989888, 0.2327503, 0.1524037, 
    0.1421147, 0.168995, 0.1803683, 0.1537142, 0.1863136,
  0.1393335, 0.07738797, 0.09893984, 0.1034186, 0.09924879, 0.06648058, 
    0.06053367, 0.0579748, 0.05592743, 0.06768047, 0.08883593, 0.08323717, 
    0.0596129, 0.05234121, 0.1043001, 0.1575886, 0.1152107, 0.09485049, 
    0.1099411, 0.1666327, 0.1014334, 0.2083152, 0.09279878, 0.1625806, 
    0.13641, 0.07966655, 0.1262253, 0.1185066, 0.1002229,
  -3.21525e-05, 0.00117354, 0.003404152, 0.03235066, 0.03002797, 0.02064799, 
    0.03155271, 0.005873309, 0.03202768, 0.01063318, 0.01530563, 0.004021269, 
    0.02672295, 0.06243619, 0.09964848, 0.1468655, 0.1008017, 0.1213596, 
    0.1362466, 0.0918747, 0.09844939, 0.06348916, 0.001300817, 0.006480769, 
    0.02721653, 0.0549013, 0.04882167, 0.04920035, 0.01931332,
  -2.446989e-07, -3.431803e-05, 0.01076819, 0.003738285, 0.0254226, 
    0.06631913, 0.02674774, 0.0253302, 0.004828865, 0.003219809, 0.1043539, 
    0.003783764, 4.956113e-05, 0.1739675, 0.02270165, 0.01250178, 0.01550569, 
    0.0436648, 0.005565577, 2.353067e-05, 0.0004058009, -6.321287e-07, 
    -7.443579e-08, 5.894376e-06, 0.03272794, 0.0004890292, 0.027762, 
    4.797736e-06, 2.483874e-07,
  0.0005244485, 0.03361551, 0.002231274, 0.01486432, 0.04345133, 0.05803461, 
    0.0362904, 0.1213702, 0.04367764, 0.03757515, 0.1236156, 0.05022652, 
    0.0589511, 0.02068608, 0.01256367, 0.00392956, 0.00613222, 0.00130034, 
    2.385965e-06, 5.116743e-07, 1.315122e-08, 1.630454e-07, 0.002384244, 
    0.03864006, 0.005597583, 0.002370934, -0.0004193808, 0.0003111163, 
    0.001659095,
  0.0440154, 0.1579455, 0.1668951, 0.05396704, 0.02263329, 0.1451099, 
    0.09641449, 0.01670504, 0.03884685, 0.09125648, 0.1445995, 0.03965839, 
    0.01543999, 0.01752027, 0.05760836, 0.02822959, 0.0228557, 0.02957728, 
    0.02462637, 0.0268393, 0.00697252, 0.01525169, 0.06775822, 0.1521151, 
    0.0953834, 0.0343543, 0.04608101, 0.02316695, 0.00438353,
  0.01184236, 0.03695054, 0.03258954, 0.1557551, 0.002687633, 0.002848848, 
    0.02004571, 0.1088924, 0.1209211, 0.1460781, 0.238612, 0.0577003, 
    0.123952, 0.05547344, 0.01907192, 0.1095766, 0.01950958, 0.01547647, 
    0.01821653, 0.02183747, 0.010357, 0.1523466, 0.1182893, 0.07738899, 
    0.008406861, 0.02710947, 0.01993941, 0.01566019, 0.07430987,
  0.01322695, 5.60629e-07, 9.42196e-08, -0.000250701, -3.50443e-06, 
    5.313538e-08, 0.004570476, 0.001312768, 0.09678537, 0.08533579, 
    0.06952106, 0.02135397, 0.05093348, 0.006297741, 0.004965233, 0.04826055, 
    0.02124869, 0.01697397, 0.002952323, -2.295946e-05, 4.997889e-06, 
    0.007651723, 0.05763847, 0.18861, 0.0108279, 0.01879011, -0.000308726, 
    0.01539601, 0.001910898,
  0.00288317, 0.001587648, 0.01370679, 0.009976274, 0.02427549, 
    -6.116246e-05, -0.002131278, 0.1857195, 0.3473388, 0.1564503, 0.1097123, 
    0.1186106, 0.1743306, 0.05072387, 0.00530794, 0.06021542, 0.03939019, 
    0.0255705, 4.514814e-05, 6.264487e-07, 0.02064946, 0.01001782, 
    0.01500858, 0.07806375, 0.04879158, 0.03564903, 0.02721541, 3.670649e-05, 
    -3.635335e-05,
  0.08766457, 0.06044321, 0.03897139, 0.1119648, 0.03005917, 0.03631762, 
    0.1023793, 0.05798975, 0.03497872, 0.119711, 0.1033527, 0.1050389, 
    0.1476088, 0.1983765, 0.09471348, 0.07322443, 0.09376325, 0.1435398, 
    0.03121283, 0.0186845, 0.113654, 0.09888069, 0.1003883, 0.09988005, 
    0.1614379, 0.1002068, 0.105601, 0.07769861, 0.1203364,
  0.1466318, 0.1115923, 0.1286031, 0.1000777, 0.1226318, 0.0780695, 
    0.06989543, 0.1567794, 0.1797005, 0.1479712, 0.2398039, 0.1873372, 
    0.1531095, 0.1207914, 0.1870618, 0.1504034, 0.1839457, 0.1780924, 
    0.1779469, 0.1330608, 0.1042162, 0.1359855, 0.1249005, 0.2123849, 
    0.1938356, 0.1177769, 0.09631009, 0.09726951, 0.1807816,
  0.06048711, 0.147129, 0.07190051, 0.1814662, 0.1875264, 0.2553535, 
    0.2135132, 0.1866727, 0.2423798, 0.214742, 0.2108767, 0.193755, 
    0.1693401, 0.3748859, 0.1504823, 0.0910923, 0.2105887, 0.2440182, 
    0.2576906, 0.1792124, 0.2174997, 0.3038512, 0.1526894, 0.1128564, 
    0.1867025, 0.1792534, 0.1057236, 0.1872365, 0.08583231,
  0.158875, 0.06437605, 0.08038951, 0.0781729, 0.1237273, 0.1411263, 
    0.2662141, 0.1480602, 0.1453455, 0.2318427, 0.1876507, 0.2395635, 
    0.1834662, 0.1821463, 0.09547859, 0.1217664, 0.04191003, 0.156761, 
    0.1995225, 0.1476598, 0.1375919, 0.1658637, 0.1459713, 0.1455465, 
    0.1325389, 0.2675971, 0.1404737, 0.2139059, 0.1527246,
  0.08344642, 0.09431665, 0.1155216, 0.1531743, 0.1409722, 0.1174622, 
    0.1065126, 0.09290607, 0.09578916, 0.1138333, 0.1396963, 0.1721496, 
    0.1605056, 0.156851, 0.1480175, 0.1016924, 0.1517762, 0.1503738, 
    0.07324341, 0.06897573, 0.1043561, 0.1423711, 0.1411625, 0.04235678, 
    0.0905301, 0.1051226, 0.136798, 0.1109391, 0.1415544,
  0.005642292, 0.003587275, 0.001532259, -0.0005227569, -0.002577773, 
    -0.004632789, -0.006687805, -0.0009969, -0.0002765243, 0.0004438515, 
    0.001164227, 0.001884603, 0.002604979, 0.003325355, 0.005319286, 
    0.006514162, 0.007709039, 0.008903915, 0.01009879, 0.01129367, 
    0.01248854, 0.004779135, 0.004918899, 0.005058663, 0.005198427, 
    0.00533819, 0.005477954, 0.005617718, 0.007286305,
  0.06294678, 0.02191081, 0.001731903, 0, 0, 0, 0, 0, 0, 0, -7.768503e-07, 
    0.0006785445, 0.0227967, 0.1594812, 0.0782114, 0.1052274, 0.162822, 
    0.1966653, 0.07937913, 0.06575346, 0.111928, 0.1583623, 0.4052019, 
    0.4988033, 0.394619, 0.2907325, 0.2245533, 0.2144149, 0.1079954,
  0.07024279, 0.06569334, 0.3148741, 0.2950011, 0.04408375, 0.0386277, 
    0.1948638, 0.02934717, 0.03669312, 0.1031501, 0.08270751, 0.1200392, 
    0.2170734, 0.1698509, 0.2621185, 0.2167499, 0.21373, 0.2539669, 
    0.2850874, 0.2964388, 0.3196517, 0.3188445, 0.3476117, 0.4375051, 
    0.3197599, 0.2679376, 0.3107935, 0.3078696, 0.239168,
  0.2912906, 0.2178491, 0.208261, 0.2754405, 0.2966354, 0.2056531, 0.199884, 
    0.2244113, 0.3156046, 0.2951139, 0.2801236, 0.3195074, 0.3249366, 
    0.2902366, 0.1842396, 0.181081, 0.2429532, 0.2081008, 0.3216821, 
    0.2663026, 0.266016, 0.2445865, 0.2069199, 0.2523715, 0.2363725, 
    0.1911702, 0.2390956, 0.307117, 0.2258146,
  0.1950861, 0.1432881, 0.213311, 0.2172148, 0.2235033, 0.1896632, 0.1578342, 
    0.1971931, 0.2583631, 0.2354546, 0.2787751, 0.2217004, 0.1356581, 
    0.09442394, 0.07862426, 0.08874497, 0.1097336, 0.1082633, 0.169176, 
    0.1676583, 0.2105448, 0.1889646, 0.2173606, 0.1426395, 0.1265869, 
    0.1763351, 0.1645747, 0.1367452, 0.2095155,
  0.1356552, 0.08593973, 0.1009609, 0.1071757, 0.104002, 0.06626429, 
    0.06045343, 0.0481592, 0.05847916, 0.08276659, 0.08288396, 0.07796555, 
    0.0570201, 0.05325345, 0.1057121, 0.1375688, 0.1186628, 0.1051839, 
    0.1071562, 0.154868, 0.104349, 0.201796, 0.08501735, 0.161962, 0.1174374, 
    0.09638704, 0.1263383, 0.1186145, 0.1090633,
  -8.958319e-05, 0.0014905, 0.006952763, 0.03756842, 0.03146835, 0.03670479, 
    0.02072301, 0.01006179, 0.03310023, 0.01581281, 0.0297606, 0.008883002, 
    0.02765064, 0.06230999, 0.09765123, 0.1469098, 0.1095618, 0.122674, 
    0.121643, 0.1096145, 0.1059002, 0.07191439, 0.005219297, 0.008449067, 
    0.02995941, 0.0545805, 0.05499103, 0.05209961, 0.0235654,
  -7.702663e-06, 5.632711e-05, 0.02008457, 0.002433478, 0.05155895, 
    0.1025162, 0.01761773, 0.01951246, 0.0002915568, 0.01331305, 0.08369164, 
    0.001978617, 0.0002473413, 0.1672381, 0.02323961, 0.01178814, 
    0.009792616, 0.04220214, 0.01353744, 0.0002172943, 0.0009312959, 
    -1.828155e-06, 3.015211e-08, 1.413357e-06, 0.06282227, 0.002254612, 
    0.02901912, 7.761701e-06, 3.644828e-07,
  0.001759809, 0.03760351, 0.001491506, 0.02836538, 0.05038125, 0.0693322, 
    0.0448485, 0.1317041, 0.05665389, 0.03860249, 0.1316792, 0.05353676, 
    0.04953583, 0.02594109, 0.01079218, 0.004701583, 0.006782765, 
    0.001563678, 0.0001548667, -3.624762e-06, 6.804601e-07, -2.837038e-06, 
    0.007014844, 0.06419061, 0.006093074, 0.004636246, 0.002108122, 
    0.0002075485, 0.001484129,
  0.06280221, 0.2130808, 0.2030601, 0.02583293, 0.02225181, 0.1527777, 
    0.09050559, 0.01861621, 0.04936101, 0.1243019, 0.1540713, 0.04657574, 
    0.02497006, 0.01669721, 0.06069873, 0.02716678, 0.02441483, 0.02991744, 
    0.03121334, 0.03090686, 0.002015557, 0.016258, 0.07112611, 0.2087179, 
    0.1219481, 0.03441131, 0.04619275, 0.02389889, 0.01885184,
  0.0147595, 0.03631323, 0.02814117, 0.2408519, 0.003452783, 0.002138167, 
    0.018701, 0.1450615, 0.1250301, 0.1534591, 0.2847469, 0.07118522, 
    0.1530694, 0.05725333, 0.02568015, 0.106553, 0.01946785, 0.01789463, 
    0.01537102, 0.0205652, 0.01459751, 0.1556981, 0.1443475, 0.08939988, 
    0.01198882, 0.03672161, 0.02202738, 0.01732333, 0.07754549,
  0.006203042, 3.745174e-07, 2.929511e-07, -0.0001210379, -1.035822e-05, 
    3.467792e-08, 0.003627651, 0.001436621, 0.1374962, 0.1006503, 0.09671489, 
    0.02774227, 0.05553321, 0.009068897, 0.00800873, 0.05256001, 0.02289267, 
    0.01323847, 0.00122395, 5.6205e-07, 2.451666e-06, 0.008567543, 
    0.06255868, 0.2598712, 0.005169259, 0.01144716, -0.0004017409, 
    0.001838224, 0.00118795,
  0.0001266372, 2.145023e-05, 0.002178192, 0.005351375, 0.03396238, 
    -0.0001099505, -0.001444074, 0.1796129, 0.3230428, 0.1578346, 0.1283583, 
    0.1166507, 0.1778192, 0.05087486, 0.007426282, 0.05410491, 0.04831162, 
    0.02951109, -5.590207e-06, 7.732636e-06, 0.006542501, 0.009567054, 
    0.009886077, 0.07770541, 0.05643224, 0.03241576, 0.03329945, 
    0.0001598805, -4.809811e-05,
  0.08494714, 0.0407005, 0.03942543, 0.10522, 0.03842929, 0.03392613, 
    0.1049346, 0.04425011, 0.01964698, 0.1134065, 0.1177398, 0.08907076, 
    0.1296063, 0.182062, 0.1017593, 0.09241783, 0.1128086, 0.1366588, 
    0.03881163, 0.01337747, 0.08784081, 0.0964389, 0.09611378, 0.1109291, 
    0.1687811, 0.09260523, 0.09684958, 0.07582431, 0.1317996,
  0.1649048, 0.1054223, 0.1348686, 0.09794374, 0.1304929, 0.08433008, 
    0.06943251, 0.1552467, 0.1692963, 0.1296905, 0.2214738, 0.1905603, 
    0.154385, 0.1400211, 0.1695724, 0.1498539, 0.2079636, 0.1958889, 
    0.193106, 0.1216037, 0.1050823, 0.1418028, 0.1153736, 0.2613308, 0.20598, 
    0.126237, 0.1157785, 0.1050599, 0.1851157,
  0.042911, 0.1597925, 0.08407983, 0.1890437, 0.2059676, 0.2700537, 
    0.2105718, 0.2167766, 0.2442397, 0.2228068, 0.2193751, 0.1901072, 
    0.1656626, 0.3506547, 0.1572764, 0.1239135, 0.205987, 0.260065, 
    0.2358204, 0.190233, 0.2272087, 0.2847901, 0.1857766, 0.123887, 
    0.1966705, 0.1668015, 0.08857619, 0.1779685, 0.07750469,
  0.1465164, 0.06423219, 0.09183294, 0.09223869, 0.1259729, 0.1516931, 
    0.2730944, 0.1367527, 0.1377824, 0.2121281, 0.1889892, 0.1992064, 
    0.1789272, 0.159035, 0.0934873, 0.1166089, 0.04642384, 0.1447247, 
    0.1834139, 0.1751876, 0.1351475, 0.1660129, 0.1579729, 0.1690014, 
    0.1429697, 0.2803377, 0.1659385, 0.2015364, 0.136755,
  0.08370005, 0.100197, 0.1057831, 0.1510691, 0.1439228, 0.1354977, 
    0.1169879, 0.09785411, 0.1053011, 0.1224713, 0.1414721, 0.1610538, 
    0.1814311, 0.1716226, 0.1392394, 0.111332, 0.1962661, 0.1775676, 
    0.06510075, 0.07298338, 0.09683584, 0.1461559, 0.1636506, 0.05708149, 
    0.1045776, 0.1004935, 0.1279466, 0.1203495, 0.1431007,
  0.06900441, 0.06432658, 0.05964874, 0.05497091, 0.05029308, 0.04561525, 
    0.04093742, 0.05002916, 0.05053296, 0.05103676, 0.05154056, 0.05204437, 
    0.05254817, 0.05305197, 0.04584217, 0.05011861, 0.05439505, 0.0586715, 
    0.06294794, 0.06722438, 0.07150082, 0.07976355, 0.07966114, 0.07955872, 
    0.07945631, 0.07935391, 0.0792515, 0.07914908, 0.07274668,
  0.08861378, 0.04432161, 0.004712058, -6.735918e-05, 0, 0, 0, 0, 0, 0, 
    0.008292622, 0.02326497, 0.02564719, 0.1755757, 0.03892656, 0.07879442, 
    0.1304956, 0.2032844, 0.1898441, 0.1066707, 0.2222444, 0.3096268, 
    0.4823674, 0.52098, 0.3957564, 0.2825142, 0.2335537, 0.2051996, 0.1731979,
  0.06683649, 0.07600702, 0.3096097, 0.3077621, 0.105863, 0.04580741, 
    0.2391419, 0.08345288, 0.0944775, 0.1867333, 0.1532381, 0.2199288, 
    0.2186052, 0.1811073, 0.2559302, 0.2144292, 0.2375335, 0.2803506, 
    0.2914705, 0.3184585, 0.3355806, 0.3217577, 0.3814472, 0.4475594, 
    0.3227267, 0.2563418, 0.2922719, 0.3211093, 0.2329101,
  0.2898984, 0.2449955, 0.2421068, 0.2783967, 0.3098271, 0.2083243, 0.242897, 
    0.2276499, 0.3559664, 0.2885895, 0.2938932, 0.2916513, 0.2946526, 
    0.2859188, 0.1939013, 0.1922167, 0.2191866, 0.2065995, 0.2982525, 
    0.2725289, 0.295166, 0.2383686, 0.1932885, 0.2238807, 0.203662, 
    0.2036098, 0.2271917, 0.308474, 0.2119261,
  0.2217005, 0.1687643, 0.2510109, 0.2210898, 0.2394276, 0.1893439, 
    0.1632929, 0.2007477, 0.2513631, 0.2327328, 0.2899855, 0.2355279, 
    0.1369968, 0.08515663, 0.07839698, 0.08621693, 0.1101619, 0.1191199, 
    0.1919188, 0.1684561, 0.1928347, 0.170655, 0.1901173, 0.1407438, 
    0.1230099, 0.1750017, 0.1661173, 0.1414554, 0.1840676,
  0.1349077, 0.09923232, 0.1075251, 0.1277968, 0.1011479, 0.06809159, 
    0.06816977, 0.0426834, 0.07672796, 0.0815651, 0.08577319, 0.08914912, 
    0.05569236, 0.0581621, 0.1063941, 0.1252004, 0.1215375, 0.1023237, 
    0.09495061, 0.1342512, 0.09707683, 0.1970495, 0.09707823, 0.1549733, 
    0.1282834, 0.1140782, 0.1252245, 0.126431, 0.1260041,
  0.001363794, 0.0015058, 0.009956568, 0.03586738, 0.03330978, 0.05289412, 
    0.01624944, 0.01343407, 0.03132695, 0.0226761, 0.02383047, 0.002930658, 
    0.04990742, 0.06338212, 0.1002953, 0.1518176, 0.103184, 0.1164418, 
    0.102356, 0.1449098, 0.1297424, 0.08199344, 0.01140043, 0.009047482, 
    0.0380722, 0.05538384, 0.05981698, 0.04868148, 0.02636296,
  1.457591e-07, 0.0001130421, 0.02206569, 0.005685469, 0.06324206, 0.1184178, 
    0.01726188, 0.01804229, 1.199865e-05, 0.02196359, 0.06839653, 
    0.0002278691, 0.0006590887, 0.1624597, 0.02686362, 0.008837393, 
    0.008478549, 0.04756935, 0.02249638, 0.001207229, 0.00233361, 
    -4.910392e-06, 3.305852e-08, 1.701292e-06, 0.08063508, 0.003527769, 
    0.03666384, 2.365079e-05, 3.840101e-07,
  0.002427679, 0.03078406, 0.002837989, 0.03648112, 0.05539062, 0.07044822, 
    0.04103438, 0.138323, 0.06173731, 0.03274263, 0.1183149, 0.04189348, 
    0.04019825, 0.02681411, 0.01093167, 0.008372525, 0.008239494, 
    0.002000497, 0.0006296368, 6.460596e-05, 0.0002129758, 3.561003e-05, 
    0.00466746, 0.06337316, 0.006580441, 0.007947351, 0.003277622, 
    6.649565e-05, 0.0001728343,
  0.04473663, 0.245434, 0.2222592, 0.03625462, 0.02026445, 0.1194532, 
    0.06716163, 0.0147391, 0.04911268, 0.1377567, 0.1078444, 0.03385074, 
    0.02249229, 0.01329387, 0.05555376, 0.02178574, 0.02095756, 0.02481832, 
    0.01898394, 0.02332743, 0.002319202, 0.004968188, 0.06131799, 0.2381705, 
    0.1273977, 0.03507839, 0.05125543, 0.02611915, 0.01447098,
  0.01202186, 0.02053004, 0.02655043, 0.2179164, 0.007234227, 0.002016317, 
    0.01423945, 0.08392739, 0.08748644, 0.1005427, 0.2508317, 0.05095907, 
    0.09991515, 0.05009589, 0.02189654, 0.07446612, 0.019455, 0.02914252, 
    0.01237672, 0.01731708, 0.0130561, 0.1243212, 0.1442384, 0.08953534, 
    0.01017847, 0.03448275, 0.01455495, 0.005480611, 0.07115727,
  0.004633479, 1.738185e-07, 3.853513e-07, 6.612565e-06, -1.954725e-05, 
    9.920829e-09, 0.00476206, 0.0005981694, 0.1591647, 0.09992313, 
    0.09630974, 0.02849766, 0.05055489, 0.009030188, 0.01220671, 0.05521432, 
    0.02700735, 0.0006383297, 0.0002627261, 1.120274e-06, 1.111721e-06, 
    0.008218465, 0.05664282, 0.2111143, 0.006149982, 0.00756058, 
    -0.0003084615, 3.681162e-05, 0.0004046269,
  5.410829e-05, 3.873193e-06, 0.0001721333, 0.007298272, 0.04488464, 
    -1.516863e-05, -0.000936061, 0.174225, 0.3232069, 0.1481594, 0.1203041, 
    0.1021226, 0.1771269, 0.05406084, 0.006749151, 0.04704292, 0.0558523, 
    0.02694855, -3.712437e-05, 3.242307e-06, 0.001918765, 0.01011506, 
    0.009126253, 0.08252664, 0.07253253, 0.03822875, 0.03915313, 0.006338228, 
    -0.000166978,
  0.08694343, 0.03528228, 0.03661151, 0.104491, 0.04804358, 0.02761088, 
    0.1034292, 0.03200851, 0.01059217, 0.09079622, 0.1253488, 0.07834593, 
    0.1231619, 0.1659379, 0.1003416, 0.1060429, 0.116666, 0.1353845, 
    0.03766214, 0.0185686, 0.0559299, 0.08864421, 0.1024898, 0.1190143, 
    0.1714935, 0.1045012, 0.1099067, 0.08244019, 0.1360314,
  0.1691251, 0.09830957, 0.150415, 0.1002658, 0.1277246, 0.07956451, 
    0.0792867, 0.1633196, 0.162382, 0.1188576, 0.2149568, 0.2067295, 
    0.1569972, 0.1325049, 0.1655478, 0.1583904, 0.2332662, 0.1825598, 
    0.1614135, 0.1159501, 0.1148558, 0.1457157, 0.1393687, 0.2823232, 
    0.2425769, 0.121483, 0.1333599, 0.09566953, 0.2024979,
  0.04260974, 0.1649168, 0.1265216, 0.1850084, 0.1942113, 0.2721373, 
    0.2105641, 0.2370302, 0.2309537, 0.2321977, 0.2479333, 0.188382, 
    0.1658833, 0.3902964, 0.1301526, 0.1384331, 0.2389001, 0.2776491, 
    0.2497365, 0.2005265, 0.2222731, 0.2734747, 0.1644174, 0.142729, 
    0.1968309, 0.1652734, 0.1050931, 0.1827708, 0.06504171,
  0.1455882, 0.07779133, 0.1113135, 0.1146275, 0.1285812, 0.1415684, 
    0.2651088, 0.1137137, 0.1411798, 0.2124226, 0.1851413, 0.1927333, 
    0.1615787, 0.1505928, 0.09258529, 0.1322039, 0.0754452, 0.1503858, 
    0.1887169, 0.1651185, 0.1735504, 0.1503289, 0.1513282, 0.1881955, 
    0.1704298, 0.2949882, 0.1572245, 0.1754496, 0.1431359,
  0.08865984, 0.0919676, 0.1081847, 0.1166605, 0.1369678, 0.1466814, 
    0.1421205, 0.1213094, 0.1455773, 0.1704198, 0.1915934, 0.1627684, 
    0.1931996, 0.1656748, 0.1350284, 0.08779524, 0.2042818, 0.1476518, 
    0.06488656, 0.06903649, 0.09307846, 0.1600907, 0.1799656, 0.07550391, 
    0.1063135, 0.09383323, 0.1229599, 0.1544161, 0.146601,
  0.1122268, 0.1080231, 0.1038194, 0.09961574, 0.09541204, 0.09120834, 
    0.08700465, 0.09266038, 0.09299001, 0.09331963, 0.09364926, 0.09397888, 
    0.09430851, 0.09463813, 0.08772534, 0.09126218, 0.09479902, 0.09833586, 
    0.1018727, 0.1054095, 0.1089464, 0.1192497, 0.119587, 0.1199242, 
    0.1202614, 0.1205987, 0.1209359, 0.1212731, 0.1155898,
  0.1294441, 0.07652675, 0.02995579, -9.06508e-05, 0, -2.377305e-05, 
    -9.1993e-05, 0, 0.0001488482, 0.01934848, 0.04651782, 0.02678821, 
    0.0446581, 0.1947602, 0.04119647, 0.06533609, 0.1224169, 0.1789974, 
    0.1898866, 0.184098, 0.2997724, 0.4445584, 0.5462326, 0.5247528, 
    0.4280493, 0.2883664, 0.2553138, 0.2106736, 0.2037999,
  0.1071867, 0.1020561, 0.2935805, 0.3080359, 0.1653518, 0.0556767, 
    0.2143407, 0.1634104, 0.1834546, 0.273221, 0.2347447, 0.2581334, 
    0.2314297, 0.1832382, 0.2907927, 0.2356734, 0.2617117, 0.2869401, 
    0.3421075, 0.3369735, 0.3462534, 0.3480457, 0.4161554, 0.5152439, 
    0.3242114, 0.2753285, 0.4427462, 0.3537995, 0.2556845,
  0.3010775, 0.3078235, 0.2900239, 0.3202747, 0.3060026, 0.210037, 0.2160009, 
    0.258003, 0.3917795, 0.2809311, 0.3047318, 0.2837913, 0.2757697, 
    0.2771753, 0.2030534, 0.2249784, 0.2406875, 0.2259253, 0.3166219, 
    0.2905487, 0.2883455, 0.2502265, 0.2266651, 0.245252, 0.2312481, 
    0.2494625, 0.2484721, 0.315437, 0.298954,
  0.2460727, 0.2244185, 0.2716286, 0.2382991, 0.252561, 0.1926847, 0.1664867, 
    0.2242671, 0.2667612, 0.2427088, 0.2824802, 0.2270733, 0.143964, 
    0.08779597, 0.09739425, 0.1042507, 0.1132574, 0.1246936, 0.19606, 
    0.1701099, 0.2091106, 0.1847833, 0.1713457, 0.1396672, 0.114838, 0.17408, 
    0.1676215, 0.147753, 0.2061552,
  0.1399966, 0.1093452, 0.1116171, 0.137278, 0.1057534, 0.07177882, 
    0.07189383, 0.0420831, 0.09878714, 0.08493884, 0.08742894, 0.08097573, 
    0.05785538, 0.06298873, 0.1133009, 0.1185031, 0.1213027, 0.115105, 
    0.1044947, 0.1252489, 0.09534809, 0.2028231, 0.1063987, 0.1540347, 
    0.1344732, 0.112564, 0.1226579, 0.1268385, 0.1258002,
  0.001487538, 0.003827501, 0.02240674, 0.02905501, 0.03579981, 0.08097769, 
    0.01676933, 0.01647385, 0.02688783, 0.02269039, 0.02178114, 0.002976041, 
    0.0671089, 0.071643, 0.104411, 0.1665497, 0.1212236, 0.1117953, 
    0.09938918, 0.1580735, 0.1499703, 0.09482187, 0.02226746, 0.008740212, 
    0.04537856, 0.06495275, 0.07380156, 0.05953026, 0.02863141,
  2.909406e-07, 1.161748e-05, 0.03866284, 0.01328636, 0.07099754, 0.1149193, 
    0.05404312, 0.01605011, 0.001450562, 0.01477219, 0.06207322, 
    3.824364e-05, 0.004366247, 0.1664085, 0.02478896, 0.02234301, 0.02110822, 
    0.05140818, 0.03076055, 0.009129026, 0.00358339, -4.136128e-05, 
    2.996705e-08, 1.247338e-06, 0.07000583, 0.005936157, 0.05191454, 
    3.342779e-05, 9.872724e-07,
  0.003542137, 0.03117827, 0.003165955, 0.06028118, 0.06044127, 0.06065106, 
    0.03591049, 0.1358234, 0.06182561, 0.03871311, 0.1026847, 0.03625881, 
    0.04421778, 0.02925921, 0.01267594, 0.009302901, 0.01051518, 0.003543566, 
    0.000300612, 4.08341e-05, 0.000372382, 0.0004106846, 0.0009508897, 
    0.0605033, 0.008256817, 0.005812912, 0.003566273, 8.590185e-05, 
    1.522731e-06,
  0.01934872, 0.1813831, 0.170035, 0.04637267, 0.01757647, 0.09626183, 
    0.06285661, 0.01215753, 0.03909943, 0.1197514, 0.08502916, 0.02737769, 
    0.02020888, 0.01278761, 0.04734369, 0.0222781, 0.01841857, 0.02174433, 
    0.0159361, 0.02001357, 0.008467634, 0.006890381, 0.05743718, 0.2261777, 
    0.1228666, 0.03886028, 0.05669398, 0.03161365, 0.01019841,
  0.005913181, 0.01120866, 0.01684573, 0.1766929, 0.005303528, 0.001846784, 
    0.01139009, 0.02088225, 0.06955177, 0.07118481, 0.2132651, 0.03862515, 
    0.07105549, 0.05006704, 0.02091399, 0.06311295, 0.01750851, 0.02409888, 
    0.01228368, 0.01612475, 0.009693968, 0.1068233, 0.1434376, 0.07288542, 
    0.01194999, 0.03527173, 0.01134704, 0.002925233, 0.03437148,
  1.654142e-05, 6.093993e-08, 1.751252e-07, 4.191528e-06, -1.195312e-06, 
    1.502037e-09, 0.002286445, 0.0002414653, 0.1383091, 0.1041997, 
    0.09825259, 0.02396189, 0.04411363, 0.01416391, 0.01860093, 0.05262828, 
    0.01256383, 2.906969e-05, 2.166876e-05, 1.688666e-06, -5.69936e-08, 
    0.01054938, 0.04324538, 0.1401941, 0.008376574, 0.006217144, 
    0.0001324183, 1.479877e-05, 0.0007963851,
  -8.746039e-05, 1.583791e-06, 1.778511e-05, 0.01271201, 0.04345697, 
    2.827193e-06, -0.0007101392, 0.1365734, 0.3288917, 0.1277677, 0.1019904, 
    0.08190519, 0.1834893, 0.0617891, 0.006684707, 0.05728099, 0.08956268, 
    0.03069944, -9.720932e-06, 1.864959e-06, 0.0002640783, 0.01178316, 
    0.008270071, 0.08850597, 0.08976025, 0.04106386, 0.04696738, 0.006801494, 
    0.0001314461,
  0.08868415, 0.0329558, 0.0382162, 0.1169153, 0.05436205, 0.02142189, 
    0.09553801, 0.02821046, 0.00553118, 0.08181521, 0.1270245, 0.07611556, 
    0.1212827, 0.1678366, 0.1028057, 0.1104233, 0.1180637, 0.1373608, 
    0.04115799, 0.01667746, 0.04530498, 0.08317089, 0.1303928, 0.1152652, 
    0.176858, 0.1094291, 0.1295017, 0.0945172, 0.1438861,
  0.156301, 0.09235034, 0.1435174, 0.1123925, 0.1469995, 0.0716584, 
    0.09505442, 0.1739466, 0.159381, 0.1115193, 0.2224418, 0.2248008, 
    0.1708424, 0.1306107, 0.1635179, 0.1972909, 0.1989231, 0.2029902, 
    0.1602168, 0.1174491, 0.1078499, 0.1170975, 0.179748, 0.2966599, 
    0.2264274, 0.129798, 0.1202631, 0.09780134, 0.1994487,
  0.05439727, 0.2079215, 0.1276325, 0.1968727, 0.2046006, 0.3121427, 
    0.2185885, 0.2586087, 0.2423429, 0.2580232, 0.3448513, 0.2125022, 
    0.1662115, 0.3737434, 0.2285427, 0.1836825, 0.2507699, 0.3027104, 
    0.2984881, 0.202347, 0.2068122, 0.2513969, 0.1636159, 0.1514472, 
    0.2222616, 0.1504841, 0.07601554, 0.1753934, 0.09935719,
  0.1339812, 0.105946, 0.1287686, 0.138098, 0.1072397, 0.1574015, 0.2440431, 
    0.1034883, 0.1393007, 0.2780142, 0.2121683, 0.1871097, 0.1553161, 
    0.1555236, 0.08873126, 0.1083464, 0.107356, 0.1542821, 0.1529601, 
    0.2024278, 0.2109395, 0.2141468, 0.1677825, 0.1906067, 0.136408, 
    0.3522131, 0.1672361, 0.1614039, 0.1152189,
  0.1043177, 0.1450219, 0.1304341, 0.09234878, 0.126363, 0.1658761, 0.166126, 
    0.1647223, 0.206196, 0.2072616, 0.2286244, 0.2492954, 0.2359376, 
    0.163955, 0.09888133, 0.06719977, 0.1552271, 0.1103544, 0.0652302, 
    0.05038045, 0.1043134, 0.1840213, 0.223983, 0.1117964, 0.1521262, 
    0.1095338, 0.1475226, 0.1884055, 0.1808005,
  0.155934, 0.1508025, 0.145671, 0.1405396, 0.1354081, 0.1302767, 0.1251452, 
    0.13361, 0.1339737, 0.1343375, 0.1347013, 0.135065, 0.1354288, 0.1357926, 
    0.1309391, 0.1379399, 0.1449407, 0.1519415, 0.1589424, 0.1659432, 
    0.172944, 0.1810158, 0.1787827, 0.1765496, 0.1743164, 0.1720833, 
    0.1698502, 0.167617, 0.1600391,
  0.1624188, 0.09191135, 0.08390933, 0.005914688, -0.0001307829, 
    0.0004473477, -0.001550001, -0.0009997531, 0.020148, 0.05443624, 
    0.05756528, 0.06580382, 0.1023645, 0.1753785, 0.03746751, 0.07375005, 
    0.1274218, 0.171899, 0.2011277, 0.225464, 0.3608024, 0.5434153, 
    0.5887195, 0.5472072, 0.3971507, 0.275968, 0.2468445, 0.2135454, 0.2362551,
  0.08073701, 0.1268638, 0.3037608, 0.3453552, 0.2068187, 0.08943986, 
    0.220962, 0.2172945, 0.2324921, 0.3277431, 0.3218749, 0.2628563, 
    0.2284046, 0.1605223, 0.3075806, 0.2563478, 0.2963084, 0.3359758, 
    0.3649351, 0.3133433, 0.311171, 0.3842302, 0.3999154, 0.5232787, 
    0.3212573, 0.2657836, 0.3632875, 0.3029864, 0.2296466,
  0.2868147, 0.300976, 0.3324503, 0.3281531, 0.2940852, 0.2422294, 0.2598703, 
    0.3140126, 0.4138225, 0.3459766, 0.3467525, 0.2950174, 0.3137816, 
    0.2997641, 0.21681, 0.2258168, 0.2364247, 0.2689509, 0.379485, 0.3162563, 
    0.3361121, 0.2935348, 0.2611822, 0.2922054, 0.2417957, 0.244713, 
    0.2874189, 0.3253652, 0.2580212,
  0.2555459, 0.2398041, 0.2808314, 0.2492443, 0.2609375, 0.2017406, 
    0.1665933, 0.2652172, 0.269745, 0.2648717, 0.3093311, 0.2392195, 
    0.1479858, 0.1043942, 0.1131183, 0.1306523, 0.1165342, 0.1506714, 
    0.2045829, 0.1890729, 0.2206525, 0.1976364, 0.1664703, 0.1310581, 
    0.1046784, 0.1756335, 0.1616963, 0.1418194, 0.2277254,
  0.1655779, 0.1196403, 0.1190185, 0.139144, 0.1274271, 0.08615295, 
    0.07645492, 0.07318029, 0.1302902, 0.1002397, 0.0970749, 0.08303212, 
    0.06827657, 0.09567958, 0.1245689, 0.115768, 0.1114443, 0.1295432, 
    0.1112232, 0.1299083, 0.1017903, 0.2347766, 0.127126, 0.1565407, 
    0.1527412, 0.1202847, 0.1308988, 0.1366842, 0.1295739,
  0.006612862, 0.005532304, 0.04195162, 0.02165898, 0.04136278, 0.09729028, 
    0.01948471, 0.02391874, 0.02322203, 0.02659776, 0.005145712, 0.01562232, 
    0.07502443, 0.07463615, 0.1076494, 0.1700916, 0.1620245, 0.1049285, 
    0.1160041, 0.15505, 0.1448079, 0.09968597, 0.02578111, 0.009607607, 
    0.05294738, 0.08453485, 0.08035849, 0.06900655, 0.03743459,
  1.090256e-06, 0.005256375, 0.0308247, 0.01643874, 0.09628592, 0.1175591, 
    0.06105418, 0.02260526, 0.002631801, 0.002744689, 0.02612088, 
    0.0008462106, 0.0118258, 0.1603329, 0.02562565, 0.03752328, 0.02374126, 
    0.05271066, 0.07284078, 0.04482833, 0.01696654, 5.651571e-05, 
    2.859722e-08, 9.074133e-07, 0.06755272, 0.006613082, 0.06188682, 
    0.001451235, 0.0001833979,
  0.007244446, 0.0455093, 0.002452548, 0.08650629, 0.05919732, 0.05129917, 
    0.0341872, 0.1301035, 0.08523557, 0.04336454, 0.1002697, 0.04286295, 
    0.05028185, 0.03439406, 0.01739044, 0.01388079, 0.02017614, 0.008719887, 
    0.0003490298, 0.0004675993, 0.0001335268, 2.683621e-06, 0.0001368959, 
    0.06495506, 0.01619132, 0.01891257, 0.007096344, 0.000121318, 3.55745e-07,
  0.00815065, 0.1611864, 0.1436563, 0.0478624, 0.01394101, 0.09250295, 
    0.05630923, 0.01196364, 0.02810253, 0.1161841, 0.07792396, 0.02368196, 
    0.01974883, 0.01708054, 0.05795447, 0.02664217, 0.02067308, 0.02148915, 
    0.01405238, 0.007351081, 0.004265318, 0.002377488, 0.0351929, 0.2355648, 
    0.1308399, 0.03473813, 0.06277218, 0.03073687, 0.01025711,
  0.003850423, 0.006348851, 0.005177464, 0.1273082, 0.01156219, 0.00218379, 
    0.008134564, 0.01021555, 0.05670831, 0.05723299, 0.1836988, 0.03415399, 
    0.05893459, 0.05307838, 0.02404217, 0.0568202, 0.02172513, 0.02466645, 
    0.02023348, 0.01449847, 0.008385273, 0.09416388, 0.1410354, 0.06865511, 
    0.01602696, 0.03741776, 0.01321989, 0.00122135, 0.02269026,
  5.471796e-06, 3.769605e-08, 7.581365e-08, 2.210954e-06, -1.48945e-07, 
    3.92004e-10, 0.001251136, 0.0001293717, 0.1259955, 0.1308081, 0.09935047, 
    0.0214216, 0.04171355, 0.02134265, 0.03201891, 0.04577865, 0.01154669, 
    0.0003650304, 1.475995e-05, 1.717235e-06, 1.297145e-06, 0.01595135, 
    0.03812032, 0.1069995, 0.01285209, 0.0119689, 0.0027683, 3.167421e-06, 
    -6.028384e-05,
  -2.241312e-05, 7.542254e-07, 7.131661e-06, 0.005447781, 0.03141584, 
    1.692738e-06, -0.000466825, 0.09493285, 0.3160285, 0.1219044, 0.08957271, 
    0.09211989, 0.1812682, 0.06986791, 0.007330093, 0.05384366, 0.1126169, 
    0.0435949, 2.588503e-07, 1.031946e-06, 0.0008218996, 0.02431643, 
    0.008951772, 0.07056636, 0.09426781, 0.03098036, 0.04366257, 0.006165569, 
    0.002347863,
  0.08431974, 0.03499551, 0.04452419, 0.1431689, 0.05756273, 0.007161276, 
    0.09358977, 0.02482591, 0.002325446, 0.07575581, 0.1357625, 0.08466648, 
    0.1198024, 0.1782546, 0.104652, 0.1038781, 0.1393992, 0.1338856, 
    0.05204292, 0.02764088, 0.0296568, 0.08091344, 0.1507964, 0.1263953, 
    0.1829132, 0.1161554, 0.1455371, 0.1155285, 0.1586603,
  0.1751305, 0.1018159, 0.1602105, 0.1116394, 0.1238475, 0.08922386, 
    0.1025083, 0.1856716, 0.1502792, 0.1078373, 0.2367948, 0.2708378, 
    0.1757425, 0.1436286, 0.1721957, 0.1832238, 0.2171907, 0.2214251, 
    0.1697746, 0.1215592, 0.07503244, 0.09934007, 0.179766, 0.301662, 
    0.2331559, 0.1573996, 0.115956, 0.09963622, 0.2283859,
  0.05674094, 0.2874711, 0.1880354, 0.2336021, 0.251357, 0.3386045, 0.236253, 
    0.3129759, 0.2706403, 0.303089, 0.3843528, 0.2051879, 0.1661574, 
    0.4202011, 0.2163106, 0.1929996, 0.3119995, 0.3491836, 0.2823747, 
    0.2010818, 0.1955265, 0.3002181, 0.154675, 0.167272, 0.2017074, 
    0.1332841, 0.07573282, 0.1905966, 0.1289237,
  0.1954412, 0.1442946, 0.1892786, 0.165239, 0.135932, 0.1694553, 0.2415511, 
    0.10716, 0.1500896, 0.3440446, 0.2582147, 0.2075275, 0.1645522, 
    0.1422429, 0.08827759, 0.1736182, 0.1038783, 0.1582562, 0.1520793, 
    0.2102447, 0.2229626, 0.2405427, 0.1868732, 0.2004409, 0.2193026, 
    0.3861728, 0.1879952, 0.1258356, 0.1373565,
  0.1597672, 0.1418909, 0.1057136, 0.1554676, 0.1075062, 0.1821259, 
    0.1605244, 0.1568147, 0.2078207, 0.3213772, 0.2529563, 0.2180288, 
    0.2333686, 0.1974421, 0.1712029, 0.1303915, 0.2285545, 0.1316554, 
    0.06245633, 0.05022237, 0.1060387, 0.1574076, 0.1920284, 0.1553711, 
    0.1775427, 0.1228786, 0.1891775, 0.237062, 0.2107294,
  0.1991826, 0.194491, 0.1897993, 0.1851077, 0.180416, 0.1757244, 0.1710328, 
    0.1959819, 0.1983268, 0.2006717, 0.2030167, 0.2053616, 0.2077066, 
    0.2100515, 0.1854349, 0.1947977, 0.2041605, 0.2135233, 0.2228862, 
    0.232249, 0.2416118, 0.2591813, 0.2521651, 0.245149, 0.2381329, 
    0.2311168, 0.2241007, 0.2170846, 0.2029359,
  0.1594303, 0.1140424, 0.1008866, 0.03021031, 0.009492382, 0.004910913, 
    0.01142546, 0.02548126, 0.03118298, 0.05873131, 0.08885769, 0.1134158, 
    0.1396396, 0.1686895, 0.05000271, 0.08009611, 0.1300439, 0.1672089, 
    0.2023309, 0.2429646, 0.3728593, 0.6104698, 0.6150094, 0.5363204, 
    0.3097994, 0.2281991, 0.2193583, 0.235992, 0.2369496,
  0.06282118, 0.1145125, 0.2729256, 0.3433982, 0.2197345, 0.1163107, 
    0.2216281, 0.2475895, 0.2891015, 0.4052854, 0.3682333, 0.2668216, 
    0.211631, 0.1478919, 0.306365, 0.2781772, 0.232546, 0.288449, 0.3268593, 
    0.2362257, 0.2850227, 0.340879, 0.355047, 0.5057802, 0.3280547, 
    0.2426758, 0.2859454, 0.2401789, 0.280797,
  0.3011336, 0.3075865, 0.331085, 0.2974639, 0.2761061, 0.2421764, 0.2417708, 
    0.263348, 0.3916111, 0.3229603, 0.3443504, 0.3123663, 0.2867216, 
    0.3027268, 0.2562829, 0.2613866, 0.2701015, 0.3033372, 0.4038928, 
    0.3249464, 0.3307957, 0.305791, 0.2695676, 0.2741529, 0.2321725, 
    0.2332273, 0.2508874, 0.3576819, 0.3000737,
  0.2609001, 0.2195165, 0.2801003, 0.2471233, 0.2627111, 0.2132462, 0.195912, 
    0.2775002, 0.2768573, 0.2816905, 0.3265103, 0.2488522, 0.1643769, 
    0.1118399, 0.1682681, 0.1283194, 0.1434816, 0.2005498, 0.2459582, 
    0.2059751, 0.247761, 0.1786476, 0.1806613, 0.1446685, 0.1063102, 
    0.1845514, 0.1536456, 0.1544186, 0.2539786,
  0.2021204, 0.1343764, 0.1376117, 0.1362081, 0.1508943, 0.09756353, 
    0.08310208, 0.09687328, 0.1477484, 0.1326895, 0.1254233, 0.1043375, 
    0.07549269, 0.08673542, 0.1594925, 0.1321299, 0.1113941, 0.1355303, 
    0.1275648, 0.146771, 0.1293481, 0.2279298, 0.163929, 0.164808, 0.1843474, 
    0.1370762, 0.1348967, 0.1513552, 0.1378723,
  0.01796847, 0.0112662, 0.05936619, 0.02704438, 0.05540311, 0.1001955, 
    0.02103789, 0.03817573, 0.03065649, 0.03643451, 0.003930756, 0.006120203, 
    0.07389902, 0.0825736, 0.1061977, 0.1547063, 0.1456771, 0.1073059, 
    0.1218056, 0.1506382, 0.1390526, 0.1068981, 0.03872497, 0.009819678, 
    0.06856255, 0.09242921, 0.08041787, 0.07532655, 0.03907847,
  3.173174e-06, 0.0003888113, 0.04555835, 0.02209118, 0.1111835, 0.1532176, 
    0.06154025, 0.03575796, 0.006628092, 0.001910919, 0.01044, -3.006054e-06, 
    0.009167183, 0.1359733, 0.02686677, 0.05467006, 0.02213308, 0.05327369, 
    0.08867011, 0.06915545, 0.0551129, 0.01238558, 3.337179e-07, 
    4.541808e-06, 0.07027201, 0.009434601, 0.06461677, 0.01792071, 0.005256949,
  0.003404629, 0.04166337, 0.007605449, 0.1059578, 0.05747826, 0.04967988, 
    0.03602933, 0.1310234, 0.1062749, 0.04864862, 0.1163424, 0.05628644, 
    0.06650939, 0.0385186, 0.0218592, 0.02177211, 0.03005867, 0.01503154, 
    0.001838491, 0.0008688156, 0.0001141716, 3.560768e-07, 9.434062e-06, 
    0.06943398, 0.0255572, 0.03842189, 0.02471367, 0.0003513514, 8.915061e-07,
  0.004746611, 0.1541633, 0.1142781, 0.06622127, 0.009913998, 0.08685368, 
    0.05141455, 0.01358439, 0.02809922, 0.1154566, 0.06606995, 0.02203883, 
    0.01918666, 0.02009861, 0.05784459, 0.03226231, 0.02579129, 0.02550677, 
    0.01829902, 0.003934128, 0.003243449, 0.0009823637, 0.01826782, 
    0.2514719, 0.1358699, 0.02846951, 0.06034442, 0.03769805, 0.01033684,
  0.003186029, 0.00236398, 0.001128629, 0.0786965, 0.004641421, 0.001977803, 
    0.007452784, 0.008177675, 0.0444643, 0.04564646, 0.1546815, 0.03526554, 
    0.04872171, 0.05062232, 0.02637558, 0.05383831, 0.02529773, 0.0251651, 
    0.03048171, 0.01535538, 0.009651556, 0.09156126, 0.1405566, 0.07274535, 
    0.02006061, 0.03970471, 0.01724536, 0.0004417731, 0.01831611,
  2.215777e-06, 2.531108e-08, 3.087713e-08, 8.430328e-07, 2.249967e-09, 
    7.135417e-11, 0.000463489, 5.45493e-05, 0.1519629, 0.1364487, 0.09206297, 
    0.0203511, 0.04165758, 0.02910221, 0.03970813, 0.03918423, 0.01878084, 
    0.001808231, 1.132016e-05, 1.980415e-06, 9.767384e-07, 0.02422156, 
    0.04139594, 0.08550606, 0.01816633, 0.01683409, 0.005774881, 
    1.370547e-06, -1.716695e-06,
  -5.536094e-06, 4.69172e-07, 3.224378e-06, 0.006158354, 0.02177416, 
    7.809939e-07, -0.000258407, 0.06712343, 0.3026582, 0.1237694, 0.08801129, 
    0.0984733, 0.1933519, 0.06865271, 0.01223304, 0.0482797, 0.1173595, 
    0.04045089, 8.764405e-07, 4.284317e-07, 6.086105e-05, 0.01687342, 
    0.01156697, 0.05904306, 0.1232969, 0.02512495, 0.04159413, 0.0123184, 
    0.005848292,
  0.06946044, 0.03264136, 0.05063752, 0.1630712, 0.02897506, 0.001789558, 
    0.08741938, 0.01908988, 0.001714661, 0.06634269, 0.1383394, 0.07694099, 
    0.1237524, 0.1849326, 0.1261602, 0.09806406, 0.1368885, 0.138553, 
    0.0662219, 0.03514871, 0.02048803, 0.06235409, 0.1850129, 0.1111897, 
    0.1821459, 0.1181517, 0.1390469, 0.1270734, 0.1869265,
  0.1826557, 0.1162054, 0.1780659, 0.1342889, 0.07321981, 0.07204355, 
    0.0880848, 0.21436, 0.145773, 0.1021969, 0.222097, 0.2847692, 0.1940897, 
    0.1485555, 0.1886113, 0.1996643, 0.2701805, 0.2188074, 0.1876936, 
    0.130816, 0.0582846, 0.1025287, 0.1802877, 0.3517552, 0.2380668, 
    0.1712719, 0.1801738, 0.1214723, 0.2755312,
  0.1339575, 0.3303831, 0.2265263, 0.2480901, 0.279877, 0.345153, 0.2305102, 
    0.2786452, 0.2634373, 0.3030089, 0.3617191, 0.2210265, 0.1845484, 
    0.4588523, 0.2226992, 0.1958809, 0.3257344, 0.3501487, 0.2804028, 
    0.2169179, 0.1798312, 0.2879159, 0.1504115, 0.1668309, 0.1856666, 
    0.1152646, 0.1035266, 0.2335105, 0.191348,
  0.23234, 0.176973, 0.197189, 0.1793984, 0.1199929, 0.181189, 0.259149, 
    0.1055823, 0.1619903, 0.3253754, 0.2389492, 0.2140174, 0.1155775, 
    0.1638867, 0.06230221, 0.1186263, 0.1161575, 0.1380645, 0.201852, 
    0.2330237, 0.2084392, 0.2134123, 0.1600992, 0.2677835, 0.1902917, 
    0.4062153, 0.187991, 0.09540815, 0.1342764,
  0.09632328, 0.1105869, 0.1368313, 0.1314438, 0.0771875, 0.1404937, 
    0.147759, 0.1232346, 0.179962, 0.1928425, 0.187749, 0.1989848, 0.2245616, 
    0.165278, 0.0767331, 0.0596224, 0.1517472, 0.07045157, 0.03429926, 
    0.07214274, 0.123297, 0.1261947, 0.1837899, 0.1759045, 0.2263304, 
    0.146676, 0.187779, 0.236917, 0.2265453,
  0.2526399, 0.2478842, 0.2431285, 0.2383728, 0.2336172, 0.2288615, 
    0.2241058, 0.2563362, 0.2624614, 0.2685865, 0.2747117, 0.2808369, 
    0.2869621, 0.2930873, 0.2893992, 0.2989568, 0.3085145, 0.3180721, 
    0.3276297, 0.3371873, 0.3467449, 0.3280882, 0.3171611, 0.3062339, 
    0.2953068, 0.2843797, 0.2734526, 0.2625255, 0.2564445,
  0.1593583, 0.1334233, 0.1051469, 0.07949477, 0.016767, 0.01987735, 
    0.02550735, 0.03446132, 0.03578749, 0.08448654, 0.1319829, 0.1414817, 
    0.155451, 0.1571825, 0.1328874, 0.08465864, 0.1284447, 0.1776448, 
    0.2164192, 0.2702801, 0.4120223, 0.6825855, 0.6307462, 0.4849201, 
    0.2814735, 0.2319893, 0.2120356, 0.2524622, 0.2341119,
  0.04605062, 0.09090989, 0.2506837, 0.3587019, 0.2440525, 0.1373037, 
    0.2233845, 0.2877604, 0.3589595, 0.4510436, 0.3908717, 0.2709751, 
    0.1958515, 0.203005, 0.3237376, 0.30064, 0.2584348, 0.2566392, 0.2952121, 
    0.2069112, 0.2681154, 0.3095885, 0.3144667, 0.502492, 0.3033039, 
    0.2626847, 0.3234566, 0.2317686, 0.2574275,
  0.3118011, 0.311539, 0.3245971, 0.3046126, 0.3022108, 0.2379624, 0.1800374, 
    0.2715597, 0.3732983, 0.3292135, 0.3353773, 0.3080349, 0.2810146, 
    0.3214111, 0.2985631, 0.2643371, 0.2793736, 0.2867754, 0.3867643, 
    0.3215569, 0.3226064, 0.3192513, 0.2962435, 0.2580801, 0.2291511, 
    0.2105228, 0.2449995, 0.3276245, 0.3017522,
  0.2542115, 0.2469324, 0.2665551, 0.2490795, 0.2564632, 0.208667, 0.2138212, 
    0.2950743, 0.2689894, 0.2942553, 0.3339638, 0.2367511, 0.1638501, 
    0.1136531, 0.1960593, 0.1351673, 0.1734466, 0.2221975, 0.2925344, 
    0.2050198, 0.2746207, 0.2039758, 0.2000991, 0.1537315, 0.1242701, 
    0.1989385, 0.1546472, 0.1867313, 0.2428007,
  0.2294678, 0.1443079, 0.1509055, 0.1204654, 0.1721433, 0.1166714, 
    0.1051849, 0.1070649, 0.1698951, 0.1816979, 0.1501466, 0.1293098, 
    0.08660778, 0.09922009, 0.1645231, 0.1759643, 0.1382434, 0.1699234, 
    0.1444209, 0.1592427, 0.1452104, 0.2285836, 0.1762391, 0.177325, 
    0.2121634, 0.1609459, 0.1461789, 0.1751436, 0.1521046,
  0.04181885, 0.0195769, 0.05644449, 0.04298821, 0.06622026, 0.1202605, 
    0.04361121, 0.05324512, 0.06755509, 0.05243639, 0.01897332, 0.002750773, 
    0.05891693, 0.09345173, 0.1095009, 0.1396505, 0.1397247, 0.1124178, 
    0.13069, 0.1352828, 0.1242286, 0.1134445, 0.06275698, 0.01229112, 
    0.07183474, 0.1019182, 0.09813272, 0.1018463, 0.04689069,
  -3.184622e-05, -0.0001085624, 0.05187187, 0.02475797, 0.08848916, 
    0.1319698, 0.06059367, 0.05119429, 0.01828036, 0.03312265, 0.001876734, 
    -2.385321e-05, 0.01255356, 0.1172315, 0.02204104, 0.06554753, 0.03004405, 
    0.05648443, 0.09759684, 0.07152421, 0.05419886, 0.0592019, 0.0005312311, 
    1.219706e-05, 0.07690046, 0.01373441, 0.06044197, 0.04907462, 0.01535664,
  0.000120528, 0.03740407, 0.01429543, 0.1078479, 0.05641159, 0.05071186, 
    0.035032, 0.131473, 0.1037813, 0.04794594, 0.1395213, 0.06925996, 
    0.08886281, 0.0386798, 0.02430794, 0.02132705, 0.02631659, 0.01703255, 
    0.008654685, 0.002658293, 0.001166472, 3.496744e-05, 1.866591e-06, 
    0.06970698, 0.02919954, 0.04781567, 0.03523823, 0.001871755, 2.665479e-05,
  0.003600663, 0.1410948, 0.09994068, 0.06912223, 0.01041398, 0.08158454, 
    0.04516045, 0.01477685, 0.03592596, 0.1222221, 0.05804557, 0.02080283, 
    0.01808147, 0.0209279, 0.05129497, 0.02983247, 0.03433627, 0.03037216, 
    0.0233235, 0.009386851, 0.001940434, 0.002250238, 0.01029564, 0.2683341, 
    0.1415692, 0.0239469, 0.05415787, 0.04058836, 0.01117979,
  0.001989461, 0.0008954684, 0.0003350799, 0.04498681, 0.003863472, 
    0.002925623, 0.0153897, 0.007231393, 0.03579797, 0.03579486, 0.1205067, 
    0.03260785, 0.03955547, 0.04386944, 0.02796884, 0.05134071, 0.03256619, 
    0.0338413, 0.04193816, 0.01768955, 0.01066255, 0.08451067, 0.1474544, 
    0.08374697, 0.02534621, 0.04202806, 0.0223328, 1.84452e-05, 0.01487421,
  9.529078e-07, 2.135173e-08, 1.545164e-08, 1.741924e-07, 2.22734e-09, 
    1.228666e-10, 0.000126285, 2.152356e-05, 0.1589648, 0.1541276, 
    0.08041326, 0.02342837, 0.04141476, 0.03340302, 0.0381705, 0.0373325, 
    0.01976193, 0.01445733, 7.929734e-05, 1.865239e-06, 6.631672e-07, 
    0.04095808, 0.04467435, 0.06971756, 0.01634638, 0.01155331, 0.004750224, 
    4.355342e-07, 5.253279e-07,
  7.497115e-07, 3.306369e-07, 1.429533e-06, 0.00362556, 0.01116271, 
    4.007961e-07, -0.0001194166, 0.05085988, 0.2872894, 0.1285602, 
    0.06737726, 0.138547, 0.1761411, 0.04948106, 0.02378369, 0.05701073, 
    0.1249588, 0.06520376, 0.0001517775, 5.32506e-07, 3.376707e-06, 0.018473, 
    0.01783279, 0.05427814, 0.1526537, 0.03239952, 0.04321782, 0.01087483, 
    0.009875601,
  0.05837994, 0.0298856, 0.04158796, 0.1739084, 0.01664864, 0.001127041, 
    0.08415391, 0.01811866, 0.002850163, 0.05430445, 0.1356439, 0.07922733, 
    0.1326266, 0.2013453, 0.1379827, 0.09917109, 0.1273364, 0.1665209, 
    0.06846857, 0.03060874, 0.01935674, 0.05705929, 0.1757234, 0.1093402, 
    0.1549105, 0.1129603, 0.1170664, 0.1294036, 0.1904759,
  0.2130097, 0.1239622, 0.1934535, 0.1518549, 0.06083219, 0.05272139, 
    0.0932222, 0.2065035, 0.1226776, 0.09665662, 0.1959845, 0.2948504, 
    0.1807232, 0.1540864, 0.194846, 0.1907166, 0.2472043, 0.2619106, 
    0.1831189, 0.1356874, 0.05189657, 0.09308048, 0.1976637, 0.3558441, 
    0.2530393, 0.1613569, 0.2485398, 0.1691862, 0.2847156,
  0.1819606, 0.2977311, 0.1739749, 0.2649187, 0.2820536, 0.3722999, 
    0.2895195, 0.2645146, 0.2336716, 0.3079402, 0.2670745, 0.2281706, 
    0.1902145, 0.4338934, 0.234526, 0.1870456, 0.3000404, 0.3666525, 
    0.2600496, 0.177692, 0.175609, 0.2357385, 0.173544, 0.2077013, 0.1705567, 
    0.1170067, 0.1126534, 0.3004212, 0.2372127,
  0.2113637, 0.2034959, 0.1803895, 0.2800669, 0.1080481, 0.191133, 0.2990382, 
    0.1516723, 0.1466184, 0.2310036, 0.1832373, 0.2005282, 0.09657475, 
    0.1320698, 0.05608945, 0.06116167, 0.1084027, 0.112655, 0.1880941, 
    0.1751356, 0.217711, 0.2455177, 0.176473, 0.1961167, 0.1706995, 
    0.4368883, 0.1880744, 0.08197752, 0.09620734,
  0.0813864, 0.05609416, 0.09874828, 0.08979376, 0.08289022, 0.1460046, 
    0.1594747, 0.1263265, 0.1585576, 0.1483863, 0.1531078, 0.1567526, 
    0.1675641, 0.1552538, 0.06822912, 0.05992391, 0.1190495, 0.03940983, 
    0.006449098, 0.03990082, 0.0393192, 0.1117474, 0.1738117, 0.1528241, 
    0.1922996, 0.1799386, 0.2128799, 0.2704831, 0.2197547,
  0.278973, 0.2743315, 0.26969, 0.2650486, 0.2604071, 0.2557657, 0.2511242, 
    0.2840764, 0.2940463, 0.3040162, 0.313986, 0.3239559, 0.3339258, 
    0.3438956, 0.3644211, 0.3728558, 0.3812906, 0.3897254, 0.3981601, 
    0.4065949, 0.4150296, 0.3754163, 0.3616531, 0.3478899, 0.3341267, 
    0.3203636, 0.3066004, 0.2928372, 0.2826861,
  0.1681137, 0.1527701, 0.1128125, 0.105034, 0.01905426, 0.0392589, 
    0.06009351, 0.06785324, 0.06100178, 0.1241634, 0.1678603, 0.157101, 
    0.2137515, 0.141112, 0.1711013, 0.09613691, 0.1614034, 0.1794933, 
    0.2210526, 0.2558592, 0.4839915, 0.6962254, 0.6435772, 0.4566533, 
    0.2821283, 0.2267045, 0.228861, 0.2257662, 0.2327989,
  0.03803239, 0.1165129, 0.240448, 0.3054781, 0.2570714, 0.1687815, 
    0.2141286, 0.3225294, 0.3708172, 0.454344, 0.4010299, 0.2700103, 
    0.195763, 0.1995315, 0.3137888, 0.309466, 0.2580167, 0.3060797, 
    0.2760691, 0.2590805, 0.2809076, 0.305871, 0.3187105, 0.5047352, 
    0.2568328, 0.2636589, 0.2971547, 0.2509857, 0.2448184,
  0.4160369, 0.3968789, 0.3720634, 0.3308947, 0.313697, 0.2745341, 0.27148, 
    0.3209946, 0.4056938, 0.3643762, 0.3369929, 0.3551448, 0.3318755, 
    0.386975, 0.2972906, 0.3029061, 0.3119473, 0.3240139, 0.3730806, 
    0.3467394, 0.3395638, 0.3464043, 0.3180622, 0.2885846, 0.2577447, 
    0.2502517, 0.2646066, 0.3365036, 0.3410998,
  0.2477888, 0.2766267, 0.2760271, 0.2551416, 0.294558, 0.2385803, 0.2729202, 
    0.309898, 0.2844764, 0.3262259, 0.3648848, 0.27285, 0.1846092, 0.1338453, 
    0.1871567, 0.1428137, 0.2283571, 0.2745694, 0.3572675, 0.2784893, 
    0.2736335, 0.2122695, 0.2223805, 0.156953, 0.1594875, 0.2194351, 
    0.168991, 0.2175764, 0.2674294,
  0.2333584, 0.1663011, 0.1640983, 0.1327533, 0.1799592, 0.1315446, 
    0.1308507, 0.1386404, 0.2111054, 0.2026654, 0.154039, 0.1480499, 
    0.1380444, 0.1181683, 0.1966189, 0.1781178, 0.1759401, 0.2041028, 
    0.180489, 0.1898883, 0.1440752, 0.2486163, 0.1878632, 0.2034201, 
    0.2118907, 0.1809377, 0.153378, 0.1955943, 0.1813528,
  0.08833093, 0.03974651, 0.03621383, 0.06117001, 0.0675592, 0.103959, 
    0.06100376, 0.08678123, 0.0874367, 0.07336033, 0.007641711, 0.003200342, 
    0.04268466, 0.1093662, 0.09884258, 0.1191147, 0.1465565, 0.138658, 
    0.1515085, 0.1375032, 0.1145871, 0.1022021, 0.07392567, 0.01243985, 
    0.05439245, 0.1378129, 0.1030863, 0.1160967, 0.09923492,
  0.001966119, -1.320552e-05, 0.01582898, 0.03094066, 0.08203769, 0.1186144, 
    0.0568821, 0.07022866, 0.05682182, 0.04052907, 0.0001079009, 
    -1.749426e-06, 0.05209703, 0.1147644, 0.0255415, 0.07962219, 0.04780659, 
    0.0526496, 0.1061944, 0.05708492, 0.1032013, 0.06396627, 0.02430035, 
    4.927085e-05, 0.09633005, 0.0213229, 0.04769393, 0.05995079, 0.04243783,
  3.01999e-05, 0.0364567, 0.01241491, 0.1070767, 0.053214, 0.04409397, 
    0.03322303, 0.1023453, 0.09114081, 0.04841, 0.12976, 0.08546361, 
    0.1008218, 0.03277383, 0.02409924, 0.02259159, 0.02388287, 0.01700374, 
    0.009803958, 0.007723365, 0.009674736, 0.002449449, 9.946993e-07, 
    0.06307141, 0.03240493, 0.009794604, 0.04598902, 0.008891344, 0.00115873,
  0.007947085, 0.1254405, 0.08312172, 0.05979429, 0.01296951, 0.06800975, 
    0.03808982, 0.01633848, 0.0381863, 0.1358105, 0.04692818, 0.01872946, 
    0.01706366, 0.02031083, 0.03808268, 0.02689059, 0.03209269, 0.02402853, 
    0.0235859, 0.01301616, 0.002874441, 0.001998204, 0.005159751, 0.2884021, 
    0.1414745, 0.02102364, 0.04319636, 0.03751409, 0.01568111,
  0.001111553, 0.0003897595, 0.0001035599, 0.02729103, 0.003371505, 
    0.006418135, 0.02890416, 0.009909407, 0.02854582, 0.03085674, 0.09320168, 
    0.03007314, 0.03023063, 0.03822408, 0.02928938, 0.05099, 0.04438018, 
    0.04065294, 0.05022913, 0.02072969, 0.01162463, 0.07258702, 0.1434231, 
    0.09050032, 0.03696859, 0.05006619, 0.03157375, 0.001083052, 0.01318163,
  5.842381e-07, 2.089587e-08, 7.913505e-09, 5.485145e-08, 2.960681e-09, 
    9.355992e-11, 5.171389e-05, 8.8117e-05, 0.1641683, 0.1651008, 0.0665259, 
    0.04710348, 0.03648249, 0.02787207, 0.03367507, 0.03775454, 0.02157282, 
    0.02313374, 0.001337774, 1.091037e-06, 4.935634e-07, 0.0496111, 
    0.04010034, 0.0552762, 0.01701478, 0.02455549, 0.01363765, 1.041465e-07, 
    5.050928e-07,
  1.587891e-07, 2.601519e-07, 5.729993e-07, 0.002071241, 0.005352465, 
    2.037364e-07, -5.403096e-05, 0.03711283, 0.2848315, 0.1246946, 
    0.07203417, 0.1605458, 0.1672067, 0.03970419, 0.02866795, 0.07463371, 
    0.1331696, 0.08560763, 0.008088603, 8.42879e-07, 1.732267e-05, 
    0.04165618, 0.01660425, 0.1046683, 0.1542578, 0.04788297, 0.04829507, 
    0.02461708, 0.009807137,
  0.04365544, 0.02344788, 0.02313439, 0.1777846, 0.01129822, 0.0001906599, 
    0.08576936, 0.01135083, 0.0009043969, 0.05134824, 0.1314135, 0.08563781, 
    0.1463077, 0.2223576, 0.1510262, 0.140736, 0.1490126, 0.2104121, 
    0.08661504, 0.03391911, 0.01811904, 0.0680511, 0.1780565, 0.08346125, 
    0.1841951, 0.1279794, 0.1370728, 0.1552835, 0.187832,
  0.2039778, 0.1607942, 0.275334, 0.1574658, 0.04644806, 0.03317508, 
    0.07592514, 0.2145029, 0.1026822, 0.09209018, 0.1832839, 0.2690838, 
    0.1777528, 0.1706183, 0.2125334, 0.2303525, 0.3138593, 0.2811732, 
    0.2171226, 0.1610989, 0.04829925, 0.1028698, 0.2388593, 0.3877334, 
    0.2938385, 0.1479079, 0.3064999, 0.1937061, 0.2826873,
  0.1662814, 0.2939409, 0.1411415, 0.2269412, 0.2523648, 0.3349677, 
    0.2464499, 0.2478045, 0.2255872, 0.3228652, 0.2389561, 0.2233972, 
    0.2050865, 0.4015935, 0.2881748, 0.2053341, 0.3370517, 0.3702698, 
    0.2812196, 0.1416331, 0.1399056, 0.2319198, 0.2155913, 0.2214126, 
    0.1810755, 0.1292563, 0.227166, 0.3096315, 0.2141355,
  0.2594394, 0.2370588, 0.2428173, 0.2738508, 0.1858694, 0.2254987, 
    0.2552524, 0.2062439, 0.1569328, 0.2014722, 0.1989549, 0.2142301, 
    0.07701291, 0.1284449, 0.06850816, 0.07015065, 0.05415403, 0.1254342, 
    0.1525066, 0.1420019, 0.2452035, 0.2266444, 0.1713083, 0.1554844, 
    0.179656, 0.4760479, 0.1979059, 0.0765181, 0.146355,
  0.1048959, 0.06971609, 0.129004, 0.1234931, 0.08102348, 0.1563299, 
    0.1646207, 0.1457788, 0.2875107, 0.1791912, 0.1440326, 0.183274, 
    0.1479615, 0.126241, 0.05154372, 0.04794749, 0.09767392, 0.08400094, 
    0.07839107, 0.04508244, 0.07010765, 0.123802, 0.17521, 0.1472496, 
    0.1827487, 0.2371278, 0.2492499, 0.2654522, 0.2437388,
  0.3066899, 0.3023382, 0.2979865, 0.2936349, 0.2892832, 0.2849315, 
    0.2805799, 0.3092391, 0.3224877, 0.3357362, 0.3489847, 0.3622333, 
    0.3754818, 0.3887303, 0.41149, 0.4165334, 0.4215769, 0.4266203, 
    0.4316638, 0.4367072, 0.4417506, 0.3859322, 0.3719919, 0.3580516, 
    0.3441113, 0.330171, 0.3162307, 0.3022904, 0.3101712,
  0.1790444, 0.1725224, 0.1302841, 0.116925, 0.0183444, 0.06774948, 
    0.09637962, 0.09734163, 0.07077875, 0.1566899, 0.1901857, 0.1764248, 
    0.2235188, 0.1167904, 0.1607812, 0.1310192, 0.1244428, 0.1647488, 
    0.2440661, 0.2796797, 0.53462, 0.7289295, 0.6837897, 0.4070445, 
    0.2989067, 0.2088813, 0.260998, 0.2137885, 0.2278883,
  0.04643273, 0.1533263, 0.2204435, 0.2657841, 0.2594498, 0.1795694, 
    0.2227685, 0.3450654, 0.3646201, 0.4644925, 0.4006643, 0.2589725, 
    0.2020595, 0.1867748, 0.3309787, 0.3106043, 0.2908169, 0.2949808, 
    0.3081867, 0.2789669, 0.2857158, 0.3230844, 0.3356795, 0.5602463, 
    0.2368504, 0.2406265, 0.3141424, 0.2941094, 0.2082174,
  0.4873434, 0.4331864, 0.3272497, 0.3091755, 0.3352357, 0.3369841, 
    0.3967032, 0.4049603, 0.4880725, 0.4192486, 0.334832, 0.4274594, 
    0.3853872, 0.4502995, 0.3203357, 0.3344026, 0.353674, 0.3528342, 
    0.3617678, 0.3592179, 0.3142884, 0.3045233, 0.3352491, 0.3428947, 
    0.3009496, 0.3155425, 0.3497067, 0.3780572, 0.4014911,
  0.2700011, 0.2356819, 0.2768289, 0.282633, 0.3272515, 0.285592, 0.3026621, 
    0.3117084, 0.3239851, 0.3131915, 0.3521536, 0.3139556, 0.2019043, 
    0.1952212, 0.2549744, 0.1964833, 0.2779503, 0.3010131, 0.3862286, 
    0.3300792, 0.2469143, 0.2188692, 0.239481, 0.178806, 0.2174788, 
    0.3107461, 0.2700688, 0.2680965, 0.285675,
  0.2775358, 0.1796576, 0.1432526, 0.1510658, 0.1848133, 0.1245017, 
    0.1580906, 0.1700979, 0.2417373, 0.1963326, 0.1104153, 0.116344, 
    0.1451628, 0.1312328, 0.2047454, 0.1731064, 0.1907072, 0.2415506, 
    0.2209071, 0.2417079, 0.2081662, 0.3103486, 0.1913567, 0.2193628, 
    0.1856543, 0.163587, 0.1510566, 0.1931741, 0.195871,
  0.1613993, 0.05082707, 0.02367699, 0.09004394, 0.09766032, 0.1014215, 
    0.08705152, 0.1322347, 0.1320692, 0.07874479, 0.0007441205, 0.000669287, 
    0.03972051, 0.1044148, 0.1187992, 0.1104633, 0.1591802, 0.1472081, 
    0.1643124, 0.1684058, 0.1054666, 0.102056, 0.08638259, 0.01416773, 
    0.06388944, 0.1244691, 0.1169008, 0.09036506, 0.1021605,
  0.07085037, 2.68369e-07, 0.01041776, 0.05586689, 0.08931768, 0.1061565, 
    0.07286961, 0.0705279, 0.05843319, 0.0157359, 2.15059e-05, -6.077018e-08, 
    0.1001141, 0.1513649, 0.03373692, 0.09105743, 0.05094989, 0.05012522, 
    0.09853178, 0.05707453, 0.1120349, 0.07386725, 0.09093089, 0.0001405074, 
    0.1045658, 0.03919829, 0.04957987, 0.06012952, 0.08220301,
  5.595065e-05, 0.04837811, 0.04715314, 0.1114281, 0.05545544, 0.04064135, 
    0.03470049, 0.09212789, 0.07452622, 0.06451702, 0.1283823, 0.09428254, 
    0.1041345, 0.02819557, 0.02716797, 0.0266802, 0.02582688, 0.02086378, 
    0.01387465, 0.01379625, 0.02284519, 0.02498614, 0.0005378277, 0.06517202, 
    0.0323695, 0.004548503, 0.05799241, 0.032967, 0.01806895,
  0.01443763, 0.1106967, 0.06210829, 0.04732795, 0.0176256, 0.05366249, 
    0.03343689, 0.02203448, 0.04176956, 0.1451713, 0.04451224, 0.01723262, 
    0.01920018, 0.02216874, 0.03344314, 0.02671075, 0.02811255, 0.02066447, 
    0.01995826, 0.01776406, 0.007969538, 0.001556104, 0.003656755, 0.2886486, 
    0.1378307, 0.01949674, 0.03784118, 0.03160535, 0.02216722,
  0.0005292469, 0.0001752186, 2.371767e-05, 0.01762672, 0.01094547, 
    0.01628564, 0.04386722, 0.01887763, 0.01972797, 0.03057434, 0.07075468, 
    0.0276375, 0.02500565, 0.03501159, 0.03310948, 0.04702391, 0.04995754, 
    0.05936017, 0.06312532, 0.02631669, 0.01532379, 0.06509135, 0.1418233, 
    0.08249707, 0.03651252, 0.05742952, 0.03881614, 0.001811131, 0.01054739,
  3.844529e-07, 2.061282e-08, 4.342197e-09, -2.683564e-07, 3.214554e-09, 
    -1.743187e-10, 8.588292e-06, 0.0005635023, 0.1761804, 0.159056, 
    0.0496254, 0.06723142, 0.03609729, 0.03032153, 0.04051875, 0.04435993, 
    0.03088322, 0.04515207, 0.02054894, 4.405587e-06, 4.238998e-07, 
    0.05608865, 0.03933052, 0.04569053, 0.02838404, 0.03826538, 0.04962066, 
    -9.023143e-06, 2.955599e-07,
  -4.505787e-08, 2.178916e-07, -4.857063e-07, 0.001389043, 0.002638086, 
    1.206347e-07, -1.978821e-05, 0.02349531, 0.303644, 0.1215635, 0.06751155, 
    0.1742272, 0.1966378, 0.0458217, 0.05368535, 0.1180936, 0.1734198, 
    0.1051999, 0.04663853, 5.042734e-07, 1.812769e-06, 0.04048986, 
    0.03533994, 0.1247987, 0.1629971, 0.05727034, 0.07992736, 0.09362792, 
    0.009660338,
  0.03013755, 0.01630302, 0.01139958, 0.1609877, 0.004715282, -4.323928e-05, 
    0.09427833, 0.006822168, -0.0001412683, 0.04365029, 0.1345419, 
    0.08507488, 0.1740542, 0.2616449, 0.1767831, 0.2057367, 0.2860078, 
    0.3808401, 0.1439968, 0.03876854, 0.01419207, 0.06512999, 0.1807106, 
    0.08518427, 0.2036795, 0.1724086, 0.1617032, 0.172614, 0.2108298,
  0.161783, 0.1728901, 0.2219933, 0.1205111, 0.04085069, 0.02033352, 
    0.05110572, 0.210994, 0.08321047, 0.09191713, 0.1632797, 0.2681557, 
    0.1742041, 0.1736702, 0.2294583, 0.3168177, 0.325434, 0.3718698, 
    0.2636335, 0.14512, 0.04422562, 0.1190389, 0.2120592, 0.3925348, 
    0.3107321, 0.2073816, 0.3396713, 0.240189, 0.3204223,
  0.1509332, 0.1720961, 0.1248387, 0.245462, 0.2239008, 0.2909138, 0.209183, 
    0.2078204, 0.2193693, 0.2370222, 0.2212162, 0.1877064, 0.1903518, 
    0.4061565, 0.3080207, 0.1901709, 0.3745226, 0.3348602, 0.2429851, 
    0.1266715, 0.09986906, 0.260326, 0.2178927, 0.2114651, 0.1821104, 
    0.1797407, 0.2501848, 0.327176, 0.2279771,
  0.3813705, 0.2023311, 0.2390854, 0.2956517, 0.1867709, 0.2327451, 
    0.3001319, 0.1566363, 0.1621318, 0.1574509, 0.1780859, 0.1920795, 
    0.07523958, 0.1651003, 0.05676914, 0.1044659, 0.04290807, 0.1444336, 
    0.1270643, 0.117173, 0.2823267, 0.216391, 0.1660536, 0.1578627, 0.275905, 
    0.5020798, 0.1893432, 0.09768108, 0.2701889,
  0.173151, 0.0965192, 0.08104584, 0.1318987, 0.06820296, 0.1790808, 
    0.190722, 0.2073226, 0.3144346, 0.2449294, 0.1951177, 0.1971627, 
    0.1755634, 0.1201611, 0.05701687, 0.0689712, 0.1390268, 0.0569815, 
    0.05943899, 0.03466944, 0.08467956, 0.1270684, 0.1459209, 0.1692166, 
    0.1637444, 0.2348266, 0.2409315, 0.3057664, 0.2698415,
  0.3144235, 0.3095978, 0.304772, 0.2999463, 0.2951206, 0.2902948, 0.2854691, 
    0.3058111, 0.3195759, 0.3333407, 0.3471055, 0.3608703, 0.3746351, 
    0.3883999, 0.406537, 0.4111666, 0.4157962, 0.4204258, 0.4250553, 
    0.4296849, 0.4343145, 0.41372, 0.4001514, 0.3865827, 0.3730141, 
    0.3594455, 0.3458769, 0.3323082, 0.3182841,
  0.1805746, 0.1941278, 0.1363114, 0.1254708, 0.01351645, 0.1260149, 
    0.1474364, 0.1311098, 0.07618558, 0.1631058, 0.2036866, 0.1794853, 
    0.2221662, 0.09168491, 0.1705098, 0.1781995, 0.1245294, 0.1307891, 
    0.2171772, 0.312354, 0.5849167, 0.7730079, 0.6874352, 0.3802862, 
    0.283441, 0.2249644, 0.2794218, 0.2149446, 0.2372122,
  0.08703309, 0.1289369, 0.2130687, 0.2349426, 0.2721745, 0.2003336, 
    0.2021661, 0.3642727, 0.3500337, 0.4621046, 0.4047223, 0.2432486, 
    0.1986547, 0.176031, 0.3351901, 0.3112958, 0.2723292, 0.3281341, 
    0.3732488, 0.2518126, 0.3035908, 0.325852, 0.3741555, 0.6054094, 
    0.2278891, 0.2796535, 0.4667354, 0.3328025, 0.2535752,
  0.4892083, 0.3986671, 0.2788211, 0.3210608, 0.3580647, 0.3846777, 
    0.5279611, 0.4563786, 0.5123223, 0.3872623, 0.4168858, 0.4091213, 
    0.4130905, 0.4154964, 0.3670679, 0.405341, 0.4429797, 0.4031399, 
    0.3692346, 0.3325118, 0.287643, 0.2775759, 0.3508451, 0.3874884, 
    0.3592454, 0.4294335, 0.3894387, 0.4666159, 0.4891205,
  0.2425022, 0.2244884, 0.2524352, 0.2912377, 0.349473, 0.3369293, 0.3268642, 
    0.3593022, 0.3268989, 0.3105941, 0.3198708, 0.3711182, 0.2300963, 
    0.2504244, 0.3081398, 0.2606935, 0.2985786, 0.2910819, 0.3223796, 
    0.2748936, 0.2222328, 0.2219699, 0.3268429, 0.199914, 0.2589795, 
    0.3978066, 0.3222159, 0.3211462, 0.2670524,
  0.2818208, 0.1706178, 0.0977825, 0.1433287, 0.1610157, 0.1478948, 
    0.1535176, 0.2199979, 0.3224622, 0.234827, 0.1068553, 0.1067851, 
    0.1434489, 0.1693199, 0.2354473, 0.1713088, 0.3024171, 0.304401, 
    0.3079073, 0.2172532, 0.279026, 0.3642021, 0.2597137, 0.2562757, 
    0.1456574, 0.1354083, 0.1423329, 0.1879, 0.1841906,
  0.1742577, 0.03054965, 0.01655928, 0.07271463, 0.1154426, 0.09704503, 
    0.1014952, 0.155482, 0.160384, 0.07024602, 0.001225044, 8.153501e-05, 
    0.03389037, 0.07548659, 0.09350084, 0.1151826, 0.1700776, 0.1477072, 
    0.180298, 0.2027758, 0.1320546, 0.1728756, 0.1660098, 0.0121729, 
    0.0856178, 0.07441068, 0.08201905, 0.129415, 0.1378219,
  0.234504, -8.658147e-05, 0.004450456, 0.08408593, 0.09163091, 0.09721913, 
    0.06684601, 0.09225632, 0.06743807, 0.008247705, 2.876192e-06, 
    1.450856e-08, 0.04948865, 0.1345575, 0.04218174, 0.08553398, 0.09415004, 
    0.06183917, 0.0998643, 0.0646648, 0.08735665, 0.1555205, 0.1841241, 
    0.0004215642, 0.154661, 0.08349457, 0.06166665, 0.07805035, 0.1090234,
  0.008208604, 0.05599467, 0.01776777, 0.147042, 0.05449569, 0.04963886, 
    0.04916046, 0.1202182, 0.09537286, 0.06941372, 0.1295271, 0.10837, 
    0.1058766, 0.03264566, 0.03699496, 0.04872126, 0.04120117, 0.05294307, 
    0.04711531, 0.05731023, 0.07622548, 0.1165936, 0.009295451, 0.07951991, 
    0.0435083, 0.001666341, 0.07478276, 0.09359424, 0.1195042,
  0.02811637, 0.09448081, 0.04291252, 0.03629757, 0.02486173, 0.05161553, 
    0.05149769, 0.04149716, 0.03900976, 0.1454399, 0.0470174, 0.0202088, 
    0.02421681, 0.02784705, 0.03237242, 0.02930139, 0.02417282, 0.02155463, 
    0.02407169, 0.01435824, 0.01528158, 0.0164464, 0.002442261, 0.2718385, 
    0.1242969, 0.02474494, 0.03839355, 0.03541915, 0.02918796,
  0.0003168314, 6.787818e-05, 5.278768e-06, 0.01294036, 0.007476317, 
    0.03286453, 0.05533969, 0.05457356, 0.01574505, 0.04248093, 0.05781082, 
    0.0304406, 0.02500484, 0.03767154, 0.04221429, 0.0488275, 0.04822651, 
    0.09408749, 0.09421585, 0.04498725, 0.0421937, 0.07463231, 0.1352394, 
    0.065763, 0.04034487, 0.06304052, 0.05927502, 0.004959987, 0.007689368,
  2.927746e-07, 2.15061e-08, 2.595769e-09, -5.07823e-07, 3.237392e-09, 
    -5.692981e-08, -6.381236e-06, 0.006580055, 0.1798476, 0.1469929, 
    0.06529584, 0.07289504, 0.04186314, 0.04731036, 0.05661768, 0.05923035, 
    0.06303146, 0.1425369, 0.1060288, 0.001786094, 3.827603e-07, 0.0629054, 
    0.03832147, 0.04288162, 0.05000427, 0.06250235, 0.1152823, 0.01079803, 
    1.831493e-07,
  -1.292707e-07, 1.903694e-07, -6.787615e-05, 0.0008416352, 0.001589869, 
    9.190504e-08, -6.291681e-06, 0.01151998, 0.3142776, 0.0978433, 
    0.08805707, 0.2096205, 0.2414551, 0.04579774, 0.1123674, 0.2409084, 
    0.1992536, 0.1561909, 0.0859129, 0.0009998288, -0.0001807514, 0.04136392, 
    0.01895091, 0.1777052, 0.1787514, 0.0823563, 0.09123563, 0.1619398, 
    0.007665879,
  0.02294715, 0.009113625, 0.008102486, 0.1533842, 0.003244047, 
    -1.526336e-05, 0.1031934, 0.007857935, -0.0002446781, 0.03887774, 
    0.1282201, 0.08541588, 0.1802494, 0.2865298, 0.2288148, 0.3316563, 
    0.3849426, 0.4594947, 0.2411805, 0.0366021, 0.01181738, 0.06055509, 
    0.1711162, 0.08195326, 0.2204126, 0.2133839, 0.1828578, 0.1603204, 
    0.2533688,
  0.1340958, 0.1365891, 0.1807211, 0.1012104, 0.03925744, 0.01219939, 
    0.04099616, 0.1915222, 0.07660357, 0.09419584, 0.1616807, 0.2803382, 
    0.1901843, 0.1974784, 0.2569518, 0.4208072, 0.4506018, 0.3780877, 
    0.2990126, 0.1283475, 0.04538281, 0.08272456, 0.1790703, 0.3674934, 
    0.3263035, 0.3495407, 0.3745651, 0.2127834, 0.3129246,
  0.1574889, 0.1215502, 0.1355279, 0.2096434, 0.2136568, 0.2912208, 
    0.1855025, 0.1679319, 0.2172485, 0.1759014, 0.190461, 0.1427847, 
    0.1711527, 0.3476928, 0.4471722, 0.2862107, 0.3024362, 0.3161888, 
    0.2259425, 0.1047614, 0.09100446, 0.258953, 0.2123574, 0.2222326, 
    0.2095413, 0.2163693, 0.3861443, 0.4139851, 0.2707185,
  0.4128941, 0.272904, 0.2544084, 0.3562428, 0.295149, 0.25092, 0.2802059, 
    0.1336472, 0.2482851, 0.2308791, 0.1528658, 0.1757182, 0.1329809, 
    0.164341, 0.1009733, 0.1502324, 0.08943557, 0.1704117, 0.1118151, 
    0.1332263, 0.3110158, 0.2696413, 0.2635795, 0.1736783, 0.3743016, 
    0.5306205, 0.1957848, 0.1793301, 0.4219645,
  0.1883478, 0.1758038, 0.1288037, 0.1151984, 0.09804959, 0.2000635, 0.22343, 
    0.2849287, 0.3422056, 0.3159305, 0.323916, 0.3251829, 0.3193758, 
    0.2145032, 0.1346687, 0.1353925, 0.1652008, 0.09888824, 0.1433677, 
    0.09617128, 0.07948809, 0.1077418, 0.1678521, 0.1756065, 0.2223858, 
    0.2491056, 0.2234369, 0.3312043, 0.2794315,
  0.3212804, 0.3160094, 0.3107384, 0.3054675, 0.3001965, 0.2949255, 
    0.2896545, 0.3035257, 0.3169185, 0.3303114, 0.3437043, 0.3570971, 
    0.37049, 0.3838829, 0.4010076, 0.4050877, 0.4091679, 0.413248, 0.4173282, 
    0.4214084, 0.4254885, 0.4179294, 0.4057274, 0.3935253, 0.3813233, 
    0.3691213, 0.3569192, 0.3447172, 0.3254972,
  0.2010247, 0.2315549, 0.1396693, 0.1241032, 0.01901592, 0.1524998, 
    0.1773295, 0.1507539, 0.08067114, 0.1502128, 0.1988718, 0.1900901, 
    0.2235455, 0.05940509, 0.1304217, 0.1638705, 0.1459651, 0.1205304, 
    0.2088829, 0.3734487, 0.6319129, 0.7811663, 0.6739208, 0.3680566, 
    0.2607687, 0.2578195, 0.2833724, 0.2322657, 0.2688136,
  0.06841882, 0.129143, 0.2118963, 0.1695865, 0.2710347, 0.202276, 0.164805, 
    0.3681852, 0.3417673, 0.4407715, 0.3961805, 0.228804, 0.1824288, 
    0.1767235, 0.3436388, 0.3570126, 0.2914709, 0.3677882, 0.3570381, 
    0.2383203, 0.3114976, 0.3081219, 0.3954909, 0.5991884, 0.2252618, 
    0.3298062, 0.508747, 0.3943443, 0.2664244,
  0.3549891, 0.3280002, 0.2436355, 0.3317367, 0.3304114, 0.2981633, 
    0.4425052, 0.406135, 0.4181088, 0.3169745, 0.4112015, 0.3816583, 
    0.4352312, 0.3880345, 0.3693916, 0.3967994, 0.4473672, 0.4063198, 
    0.4033758, 0.2746817, 0.3290944, 0.2909718, 0.3732127, 0.3649834, 
    0.4441653, 0.4611649, 0.4213198, 0.4338757, 0.4139396,
  0.250543, 0.2304456, 0.2613001, 0.2954345, 0.367606, 0.3048298, 0.3267047, 
    0.3584901, 0.3132337, 0.2924628, 0.3388545, 0.3955474, 0.2753907, 
    0.2082924, 0.3232732, 0.297264, 0.2803519, 0.3419591, 0.2872132, 
    0.2009604, 0.1842361, 0.2228346, 0.3134286, 0.2029149, 0.2393862, 
    0.3194807, 0.290044, 0.2704867, 0.2684567,
  0.2247194, 0.1875794, 0.07572054, 0.1475096, 0.1558228, 0.1490842, 
    0.170464, 0.2170122, 0.2861104, 0.1701476, 0.09881437, 0.07565016, 
    0.05105851, 0.2095979, 0.3226726, 0.2014482, 0.2725358, 0.3273373, 
    0.1788056, 0.1567979, 0.2156023, 0.3107828, 0.2129544, 0.2809737, 
    0.1265734, 0.1232538, 0.1352213, 0.1855019, 0.2273053,
  0.2374427, 0.03514343, 0.0239867, 0.08900004, 0.0725442, 0.0991604, 
    0.05885416, 0.1736148, 0.1315133, 0.02850177, 0.002744732, 7.137676e-06, 
    0.02712557, 0.05069166, 0.06968623, 0.087849, 0.1546409, 0.1207169, 
    0.1853609, 0.192536, 0.195061, 0.1801013, 0.2916597, 0.0167002, 
    0.06572299, 0.08052159, 0.05981874, 0.1601443, 0.1250763,
  0.2343166, -0.0001899043, 0.004579179, 0.06344982, 0.048984, 0.06651097, 
    0.04125345, 0.04729985, 0.06799787, 0.008194805, 1.130741e-06, 
    9.379424e-09, 0.02665844, 0.1216787, 0.1070236, 0.1025617, 0.1216757, 
    0.08824594, 0.1149782, 0.06184265, 0.08752023, 0.1239617, 0.3319914, 
    0.0005629167, 0.09969541, 0.0816649, 0.1500084, 0.06056118, 0.1408395,
  0.1267903, 0.05657006, 0.002322547, 0.1369297, 0.0688733, 0.0583258, 
    0.05250717, 0.1097532, 0.07976713, 0.06065389, 0.09141485, 0.08629893, 
    0.1120154, 0.0419566, 0.03884731, 0.06247473, 0.0402538, 0.04782702, 
    0.04371873, 0.04733745, 0.1659789, 0.3000158, 0.2443164, 0.0683452, 
    0.01474224, 0.0004068043, 0.1063574, 0.08736296, 0.2319618,
  0.09262013, 0.06828365, 0.02547175, 0.04454699, 0.1514438, 0.08855471, 
    0.15142, 0.1336591, 0.029611, 0.1403596, 0.04642602, 0.07962923, 
    0.05742854, 0.07037102, 0.06529308, 0.04275697, 0.02885241, 0.02614347, 
    0.03436296, 0.01747599, 0.04786751, 0.04266192, 0.004166536, 0.2080389, 
    0.07614687, 0.02898552, 0.05531997, 0.07682075, 0.09226956,
  0.0001628006, 1.560387e-05, -1.605222e-06, 0.009559136, 0.006351098, 
    0.3031073, 0.05598405, 0.08803133, 0.029518, 0.04915964, 0.06681701, 
    0.03545596, 0.03032715, 0.04936253, 0.05075175, 0.06157519, 0.05603416, 
    0.1361902, 0.1242836, 0.151865, 0.2108387, 0.09694023, 0.1351808, 
    0.05267182, 0.04577315, 0.0936726, 0.2946393, 0.007646503, 0.004898191,
  2.347588e-07, 2.248812e-08, 1.95839e-09, -8.53044e-07, 3.287514e-09, 
    -2.26852e-06, -2.924027e-05, 0.01856679, 0.1551742, 0.1764685, 
    0.08430399, 0.0612659, 0.05072055, 0.04964391, 0.03114265, 0.0431669, 
    0.1376402, 0.1668689, 0.3712745, 0.06988613, -1.428183e-06, 0.08978321, 
    0.05099811, 0.04957953, 0.07989474, 0.1204592, 0.1753314, 0.04637403, 
    1.350817e-07,
  -8.63547e-07, 1.721028e-07, 7.361753e-06, 0.0002727354, 0.001047654, 
    8.147808e-08, -2.815468e-06, 0.004192865, 0.3303767, 0.08764686, 
    0.1165145, 0.2195849, 0.2833418, 0.1368428, 0.226681, 0.2724529, 
    0.185597, 0.2630953, 0.2117182, 0.009663267, -0.000243691, 0.04658652, 
    0.006596856, 0.1311679, 0.1985276, 0.1708146, 0.1602131, 0.220625, 
    0.01253058,
  0.01722733, 0.006116628, 0.005629018, 0.1578714, 0.00866487, -7.777396e-07, 
    0.1097028, 0.007890194, -0.000133164, 0.03451982, 0.1211114, 0.06771139, 
    0.1714199, 0.3122611, 0.3435823, 0.3443792, 0.3462933, 0.4251594, 
    0.3629169, 0.03246215, 0.01040324, 0.0532909, 0.1427195, 0.07954545, 
    0.220189, 0.2631383, 0.153546, 0.1662333, 0.242353,
  0.1193105, 0.1523031, 0.1541469, 0.09543699, 0.03552543, 0.007870222, 
    0.03174955, 0.178935, 0.06330388, 0.08732788, 0.1467787, 0.2795924, 
    0.2336609, 0.2409087, 0.307198, 0.4597616, 0.4256659, 0.3320585, 
    0.2674561, 0.1387315, 0.03172896, 0.06087462, 0.1667434, 0.3537283, 
    0.3167191, 0.4246152, 0.3764142, 0.241061, 0.3077896,
  0.1256476, 0.0828938, 0.1241826, 0.1934166, 0.2087887, 0.2606294, 
    0.1856211, 0.1623907, 0.1994624, 0.1652646, 0.1636023, 0.1350494, 
    0.1595201, 0.3021957, 0.531504, 0.3483034, 0.2739815, 0.3087792, 
    0.2508202, 0.09377085, 0.06892594, 0.2431002, 0.2103932, 0.2213662, 
    0.2509789, 0.2069681, 0.5381071, 0.5199515, 0.2395947,
  0.3417954, 0.1950646, 0.2046641, 0.3089162, 0.2421005, 0.3138703, 
    0.2085479, 0.1804501, 0.1638952, 0.1505598, 0.1386149, 0.1429246, 
    0.192398, 0.2712127, 0.1946146, 0.2294888, 0.09286457, 0.1777483, 
    0.1144526, 0.1727622, 0.3039331, 0.2863586, 0.2872214, 0.2561699, 
    0.4920919, 0.5417914, 0.1813338, 0.1824398, 0.5019071,
  0.225618, 0.1543982, 0.1629142, 0.1194048, 0.1845006, 0.259911, 0.2990112, 
    0.3226554, 0.4074967, 0.3663941, 0.3062594, 0.262679, 0.3155276, 
    0.3391806, 0.2420251, 0.2032884, 0.2043212, 0.1540281, 0.1949091, 
    0.08578948, 0.04955891, 0.119592, 0.1544049, 0.2512657, 0.2277005, 
    0.2570988, 0.2177388, 0.3182596, 0.2719716,
  0.3120373, 0.3075071, 0.302977, 0.2984469, 0.2939168, 0.2893867, 0.2848566, 
    0.2919678, 0.3044602, 0.3169526, 0.3294449, 0.3419373, 0.3544297, 
    0.3669221, 0.3917019, 0.3946968, 0.3976917, 0.4006866, 0.4036815, 
    0.4066764, 0.4096712, 0.3968136, 0.3858565, 0.3748993, 0.3639421, 
    0.352985, 0.3420278, 0.3310707, 0.3156613,
  0.2171474, 0.2365611, 0.1592418, 0.1233369, 0.03833907, 0.1535984, 
    0.1906606, 0.1638373, 0.06394526, 0.1274801, 0.2027296, 0.2214209, 
    0.2571273, 0.02659024, 0.08778723, 0.1757747, 0.1695191, 0.1516994, 
    0.2203344, 0.4201911, 0.6570822, 0.7899641, 0.6637469, 0.3962124, 
    0.2811816, 0.2747826, 0.2560028, 0.2455269, 0.278085,
  0.03163544, 0.07029906, 0.1884235, 0.1331108, 0.2634246, 0.1905727, 
    0.112961, 0.3518736, 0.3235012, 0.4372184, 0.3779599, 0.2120106, 
    0.1721211, 0.1840351, 0.3470306, 0.4033716, 0.3349462, 0.3679955, 
    0.3486058, 0.2226165, 0.3102324, 0.3449318, 0.3845943, 0.6217342, 
    0.2138228, 0.393627, 0.4786715, 0.4730825, 0.2767802,
  0.3052366, 0.2816491, 0.2001843, 0.284603, 0.3105461, 0.2486123, 0.3127972, 
    0.3035493, 0.313981, 0.2549161, 0.3370165, 0.3672255, 0.4376641, 
    0.4264782, 0.3830964, 0.4153284, 0.400689, 0.3903644, 0.4022058, 
    0.2228845, 0.3170142, 0.3102287, 0.3644386, 0.3411312, 0.4479226, 
    0.4292046, 0.3844987, 0.3605227, 0.3324029,
  0.2493056, 0.2310275, 0.2660407, 0.2748626, 0.338687, 0.3227144, 0.3575439, 
    0.3713855, 0.3031822, 0.2818814, 0.2911852, 0.3570093, 0.2695681, 
    0.3230633, 0.3329047, 0.2644638, 0.2775573, 0.3102432, 0.2301726, 
    0.1634951, 0.1293322, 0.1931348, 0.2968273, 0.2093048, 0.2118149, 
    0.2727113, 0.2400091, 0.2299442, 0.3015671,
  0.1986499, 0.1348105, 0.03794435, 0.1349303, 0.1459805, 0.156494, 
    0.2268242, 0.2078649, 0.2454361, 0.1211772, 0.04762603, 0.02991207, 
    0.02004181, 0.165262, 0.3962355, 0.1701918, 0.171174, 0.2142281, 
    0.116553, 0.1260129, 0.1768898, 0.2774009, 0.2199213, 0.2961514, 
    0.09257451, 0.0999407, 0.1452043, 0.1527954, 0.2273498,
  0.1503913, 0.06658001, 0.02207218, 0.03537336, 0.03630448, 0.1139415, 
    0.03356005, 0.07598677, 0.05824401, 0.01493345, 0.002133685, 
    -7.440116e-08, 0.02469925, 0.02973959, 0.06124688, 0.08272196, 0.1569785, 
    0.128358, 0.144126, 0.1571321, 0.1807132, 0.09793363, 0.146738, 
    0.01339014, 0.06831352, 0.04580885, 0.04099334, 0.1011897, 0.1224677,
  0.1636432, -0.001088498, 0.004692154, 0.01657729, 0.02096551, 0.04181091, 
    0.01531927, 0.01854421, 0.02972375, 0.002611665, 5.779259e-07, 
    7.787424e-09, 0.01331231, 0.09179998, 0.09656707, 0.1271911, 0.07879911, 
    0.05137724, 0.05427037, 0.01519065, 0.04275519, 0.04347581, 0.2561856, 
    0.002221634, 0.07763748, 0.06173945, 0.03282697, 0.02620838, 0.1996266,
  0.3179357, 0.04775686, -0.0002237784, 0.086271, 0.03039556, 0.09271761, 
    0.028418, 0.06123306, 0.03419269, 0.08386869, 0.06118799, 0.02601388, 
    0.07689594, 0.03377553, 0.01611002, 0.02324209, 0.01136511, 0.009846019, 
    0.007457563, 0.00917756, 0.05197084, 0.1125278, 0.4330544, 0.04033421, 
    0.002845951, 0.0001095442, 0.0239458, 0.02298055, 0.08388957,
  0.1916502, 0.04370994, 0.01497224, 0.05615185, 0.06667091, 0.04107427, 
    0.06044156, 0.03943278, 0.04056111, 0.1042913, 0.04488969, 0.1192913, 
    0.02360735, 0.03366731, 0.04396028, 0.03715915, 0.02958351, 0.03049647, 
    0.01698189, 0.01621822, 0.04629244, 0.1657957, 0.1038544, 0.1665799, 
    0.04253555, 0.02410814, 0.0749869, 0.1063809, 0.07287574,
  3.322727e-05, 1.14675e-06, -1.549619e-06, 0.005194147, 0.0101089, 
    0.04880461, 0.0713985, 0.01973611, 0.00908212, 0.01922231, 0.06824679, 
    0.02997985, 0.02765534, 0.03459773, 0.02817982, 0.04578968, 0.04041274, 
    0.08940495, 0.0828581, 0.1633495, 0.0829936, 0.05504189, 0.1494963, 
    0.04864033, 0.02119615, 0.04085334, 0.1585608, 0.06867526, 0.0007605659,
  1.916952e-07, 2.336371e-08, 1.683484e-09, -4.401571e-07, 3.290772e-09, 
    -0.0004834304, 8.669846e-05, 0.09109104, 0.1132495, 0.2017864, 
    0.09171809, 0.0562967, 0.02058163, 0.01197969, 0.00767201, 0.03423123, 
    0.07412528, 0.05483451, 0.3812903, 0.2182425, -0.0006758419, 0.07371797, 
    0.02449833, 0.03234641, 0.06437473, 0.0721501, 0.1701688, 0.05449327, 
    1.163083e-07,
  -1.432725e-06, 1.606831e-07, 6.738102e-06, -3.908148e-06, 0.001219347, 
    7.74393e-08, -1.463326e-06, 0.0009039332, 0.3345886, 0.0758673, 
    0.1109491, 0.2485396, 0.3151018, 0.1228182, 0.304923, 0.2312652, 
    0.1578037, 0.2307941, 0.2667748, 0.177746, 0.002259226, 0.04817677, 
    0.009790156, 0.1726496, 0.2062884, 0.1432309, 0.1560907, 0.184397, 
    0.01827318,
  0.0151161, 0.003691095, 0.007271881, 0.1773134, 0.03454366, 9.309788e-08, 
    0.1121454, 0.005190357, -9.132038e-05, 0.02907625, 0.1178714, 0.05521427, 
    0.1680062, 0.358008, 0.4350896, 0.3835744, 0.2920212, 0.3594266, 
    0.3143749, 0.04099926, 0.009075544, 0.05177164, 0.110879, 0.07972333, 
    0.22095, 0.2523643, 0.1501658, 0.1518819, 0.2439279,
  0.1077493, 0.124987, 0.1344344, 0.08349137, 0.03108775, 0.008089408, 
    0.02557091, 0.1634474, 0.04800748, 0.08044697, 0.1259429, 0.2872891, 
    0.2376582, 0.2932863, 0.3847969, 0.4304728, 0.4223141, 0.3042677, 
    0.2150218, 0.1574559, 0.01670737, 0.04073861, 0.1441942, 0.326877, 
    0.2739615, 0.357146, 0.334865, 0.1861569, 0.255882,
  0.07278764, 0.05519641, 0.1050243, 0.1680351, 0.191424, 0.2366421, 
    0.1676947, 0.1411452, 0.1869892, 0.1479684, 0.1398804, 0.1061005, 
    0.1368143, 0.2846435, 0.4892299, 0.4804414, 0.2472641, 0.2806557, 
    0.1903941, 0.08516574, 0.06074262, 0.2147988, 0.1739939, 0.2713903, 
    0.3983553, 0.1877565, 0.4689057, 0.3910667, 0.1456688,
  0.1807375, 0.08540801, 0.1315375, 0.2058409, 0.2255912, 0.2499792, 
    0.1499693, 0.1138188, 0.09452859, 0.107487, 0.1496222, 0.152513, 
    0.1375285, 0.2776501, 0.1940638, 0.2577032, 0.1874788, 0.1757028, 
    0.1594899, 0.1950737, 0.2878835, 0.2977718, 0.2622921, 0.3139562, 
    0.4891007, 0.5188257, 0.1820774, 0.1762439, 0.4157243,
  0.2884715, 0.2860944, 0.208862, 0.2028268, 0.2104317, 0.3139369, 0.3791694, 
    0.4150592, 0.5051602, 0.4355598, 0.3429404, 0.263422, 0.3015032, 
    0.3325827, 0.2626412, 0.2377545, 0.230609, 0.1631173, 0.1437503, 
    0.185828, 0.06739199, 0.1493883, 0.2268974, 0.3507177, 0.2148894, 
    0.2231021, 0.2245708, 0.3151672, 0.20666,
  0.282757, 0.2802002, 0.2776433, 0.2750864, 0.2725295, 0.2699726, 0.2674157, 
    0.2478777, 0.2594422, 0.2710066, 0.282571, 0.2941354, 0.3056998, 
    0.3172642, 0.3494699, 0.3501736, 0.3508773, 0.3515809, 0.3522846, 
    0.3529883, 0.3536919, 0.3346953, 0.3249841, 0.3152729, 0.3055618, 
    0.2958506, 0.2861394, 0.2764282, 0.2848026,
  0.2394395, 0.2503728, 0.1452226, 0.1208883, 0.03435416, 0.1311467, 
    0.1785654, 0.1534144, 0.02985204, 0.07998218, 0.1355781, 0.2124978, 
    0.3283087, 0.006375905, 0.07400536, 0.1921663, 0.2317126, 0.2005033, 
    0.2286572, 0.4513813, 0.6502671, 0.79656, 0.6478051, 0.4019377, 
    0.3053839, 0.2861891, 0.2471689, 0.2595843, 0.2729241,
  0.02109896, 0.03029978, 0.1484697, 0.09825139, 0.2474844, 0.1835824, 
    0.0654057, 0.3191503, 0.3045383, 0.4356179, 0.3533929, 0.1996065, 
    0.1621807, 0.1663687, 0.3533553, 0.4288643, 0.3527945, 0.426578, 
    0.3371934, 0.2163545, 0.2915292, 0.3880284, 0.4294731, 0.6585056, 
    0.2007092, 0.4306502, 0.5485781, 0.465423, 0.2655028,
  0.2727211, 0.2514046, 0.1767678, 0.2114291, 0.2780392, 0.2220569, 
    0.2139473, 0.2177004, 0.2342459, 0.2095474, 0.2692956, 0.318927, 
    0.4227495, 0.4388623, 0.3866581, 0.4456644, 0.3674117, 0.3656423, 
    0.3711343, 0.20612, 0.2521825, 0.3062207, 0.3319159, 0.27893, 0.3793291, 
    0.3891953, 0.3583003, 0.3287793, 0.3110507,
  0.2439546, 0.2382029, 0.2641388, 0.2646503, 0.3378642, 0.3334506, 
    0.3708876, 0.3540739, 0.3191054, 0.2603996, 0.2535969, 0.3165783, 
    0.2223216, 0.2950445, 0.338012, 0.2331004, 0.2483631, 0.270004, 
    0.1974526, 0.1540536, 0.111428, 0.1761064, 0.2650986, 0.1989719, 
    0.1718433, 0.25122, 0.2028731, 0.2143158, 0.2944027,
  0.1860823, 0.08388569, 0.01705901, 0.1177646, 0.1210301, 0.1313017, 
    0.2106992, 0.1499975, 0.1885567, 0.08412204, 0.01838109, 0.01178712, 
    0.008274576, 0.09896306, 0.3877214, 0.1177808, 0.1301499, 0.152206, 
    0.09300923, 0.1002016, 0.1439308, 0.2539237, 0.1647161, 0.3079834, 
    0.1112697, 0.1216914, 0.1246495, 0.1370953, 0.2169057,
  0.06333015, 0.04546362, 0.01633716, 0.01091673, 0.01919559, 0.06999016, 
    0.01466804, 0.05275905, 0.02891641, 0.006657457, 0.0006541515, 
    -2.433822e-06, 0.02405831, 0.02277796, 0.04662416, 0.06419244, 0.1799994, 
    0.08751319, 0.08479124, 0.1195365, 0.0771643, 0.06473126, 0.07284415, 
    0.01548295, 0.04894537, 0.0302953, 0.03302567, 0.0570356, 0.04044466,
  0.09474956, -0.0002545219, 0.004428761, 0.004146642, 0.01098896, 
    0.02174192, 0.002094478, 0.007746889, 0.006807489, 0.0001225894, 
    5.747775e-06, 6.903852e-09, 0.00143302, 0.06839919, 0.04941778, 
    0.09540121, 0.03859362, 0.02189353, 0.02667454, 0.001781417, 0.01517047, 
    0.009781378, 0.1003487, 0.007083529, 0.0597958, 0.06419474, 0.008584525, 
    0.006600303, 0.07358177,
  0.1676365, 0.0399648, -8.953572e-05, 0.07382389, 0.009184699, 0.02517586, 
    0.006512338, 0.03533911, 0.007187576, 0.01257087, 0.04698368, 
    0.004144921, 0.04713879, 0.006703163, 0.00225452, 0.003249416, 
    0.000968312, 0.00102442, 0.0007183973, 0.001301883, 0.01447414, 
    0.03646554, 0.2068213, 0.02267389, 0.0008384588, 3.891988e-05, 
    -0.001553971, 0.004619072, 0.0264178,
  0.06246737, 0.02899079, 0.01710444, 0.05174673, 0.01021129, 0.02393404, 
    0.02182966, 0.008348959, 0.06278386, 0.06844379, 0.03347383, 0.01952272, 
    0.004185266, 0.005108827, 0.02535108, 0.006219112, 0.01154073, 
    0.01159023, 0.001811903, 0.008233734, 0.01461897, 0.08714227, 0.4333816, 
    0.1380899, 0.02841293, 0.006316903, 0.02022257, 0.01948298, 0.02473985,
  0.0001046426, -5.649143e-07, -5.679923e-07, 0.002913859, 0.01631149, 
    0.01408351, 0.04648916, 0.01034098, 0.002529045, 0.004289817, 0.04300777, 
    0.01593794, 0.01108061, 0.008325101, 0.006810344, 0.01561207, 0.01924758, 
    0.03543783, 0.03247309, 0.04305716, 0.02141552, 0.0299505, 0.1827832, 
    0.04044057, 0.00461109, 0.01443896, 0.0420311, 0.09335072, 3.21897e-05,
  1.529753e-07, 2.358021e-08, 1.487739e-09, -1.667938e-07, 3.23778e-09, 
    0.001041677, -6.21902e-05, 0.08137283, 0.08382452, 0.1442723, 0.02232419, 
    0.0190057, 0.005071923, 0.00139582, 0.001006987, 0.01341959, 0.02023606, 
    0.01417786, 0.1809165, 0.2233211, 0.0002508696, 0.07016596, 0.009957052, 
    0.01911134, 0.01583724, 0.08046013, 0.05438655, 0.01952705, 1.075736e-07,
  -8.163527e-07, 1.551678e-07, -6.560177e-07, 1.757917e-05, 0.001381364, 
    7.500143e-08, -9.171728e-07, -0.001211312, 0.3284216, 0.07271194, 
    0.09869927, 0.2616798, 0.2822409, 0.1412683, 0.2055231, 0.2212664, 
    0.154097, 0.1212327, 0.1879813, 0.2116551, 0.001919498, 0.04125495, 
    0.01179457, 0.1430955, 0.1641232, 0.08485006, 0.0964898, 0.08101345, 
    0.02130217,
  0.01171716, 0.001584154, 0.007894211, 0.1700111, 0.04744743, 1.446397e-07, 
    0.1104369, 0.00336818, -7.287897e-05, 0.02361607, 0.1311711, 0.05325268, 
    0.1663216, 0.3988569, 0.4346838, 0.294331, 0.2726794, 0.3270665, 
    0.2745598, 0.0476237, 0.00777918, 0.04117148, 0.08809583, 0.08585943, 
    0.1812157, 0.2217766, 0.1470116, 0.1295759, 0.2168023,
  0.1277243, 0.08418818, 0.1114039, 0.07165644, 0.02441825, 0.008667115, 
    0.01813336, 0.1518147, 0.04359372, 0.06977437, 0.1081271, 0.27958, 
    0.2742565, 0.3376928, 0.4112836, 0.4270836, 0.4148806, 0.2735596, 
    0.1759617, 0.1595076, 0.008459693, 0.02467231, 0.1309929, 0.3031985, 
    0.2616771, 0.3210104, 0.2757023, 0.1300843, 0.2152454,
  0.0421848, 0.04278913, 0.08923511, 0.1445605, 0.1794805, 0.2154173, 
    0.1458852, 0.1138429, 0.1720826, 0.1384155, 0.1205646, 0.08235865, 
    0.1234805, 0.2577497, 0.4286387, 0.4624675, 0.2127059, 0.2474849, 
    0.1533893, 0.0750206, 0.05848144, 0.1873124, 0.1905546, 0.2639963, 
    0.4952025, 0.1967681, 0.3729781, 0.310566, 0.09511669,
  0.114158, 0.03921889, 0.082592, 0.1555068, 0.1748289, 0.2328529, 0.1200211, 
    0.08047429, 0.04652076, 0.06413411, 0.1169787, 0.1282265, 0.09320134, 
    0.193363, 0.1389364, 0.2352336, 0.1906363, 0.1715651, 0.2004487, 
    0.2086486, 0.3779642, 0.4037531, 0.2645577, 0.412187, 0.4854546, 
    0.4809496, 0.1716045, 0.16867, 0.2995016,
  0.2584296, 0.2758379, 0.2126794, 0.1627491, 0.2296827, 0.3813017, 
    0.3753757, 0.4296948, 0.5162884, 0.4599165, 0.370567, 0.3903687, 
    0.3413943, 0.327112, 0.3295338, 0.2918783, 0.2954059, 0.2589501, 
    0.1504832, 0.1801454, 0.1406667, 0.1579864, 0.2055213, 0.3170291, 
    0.1824482, 0.1903796, 0.1954913, 0.3022633, 0.2592049,
  0.2543121, 0.248078, 0.2418438, 0.2356097, 0.2293755, 0.2231413, 0.2169072, 
    0.1703532, 0.1808871, 0.191421, 0.201955, 0.2124889, 0.2230228, 
    0.2335567, 0.2855418, 0.2890391, 0.2925364, 0.2960337, 0.299531, 
    0.3030283, 0.3065256, 0.3110784, 0.3032813, 0.2954843, 0.2876872, 
    0.2798901, 0.2720931, 0.264296, 0.2592995,
  0.2536327, 0.2485329, 0.1009383, 0.1052316, 0.02415731, 0.1045539, 
    0.1317655, 0.1564837, 0.004907423, 0.04918046, 0.0949548, 0.189347, 
    0.3653443, 0.0001194957, 0.1321923, 0.2354062, 0.3291658, 0.2825424, 
    0.2243505, 0.4607776, 0.6360319, 0.7878951, 0.6151549, 0.3915718, 
    0.39087, 0.317479, 0.2389863, 0.2275548, 0.2412649,
  0.0285067, 0.01522458, 0.1087604, 0.06619323, 0.2198193, 0.17441, 
    0.02347141, 0.2746461, 0.2917802, 0.4082065, 0.3190922, 0.2029514, 
    0.1504686, 0.147102, 0.3677644, 0.4399565, 0.3935366, 0.4572607, 
    0.3136688, 0.2262937, 0.2978528, 0.3891908, 0.4264582, 0.6803463, 
    0.1982981, 0.5160803, 0.562979, 0.5018205, 0.2690532,
  0.2178412, 0.2244066, 0.151532, 0.1628232, 0.2155884, 0.171346, 0.1536064, 
    0.1632747, 0.1704498, 0.1642591, 0.212037, 0.2708466, 0.3997448, 
    0.4185431, 0.3373202, 0.4114494, 0.3244625, 0.338558, 0.3167988, 
    0.1754116, 0.2051386, 0.2766173, 0.2726788, 0.2297135, 0.3329603, 
    0.344375, 0.3002177, 0.2852979, 0.2687694,
  0.2383305, 0.2353294, 0.237441, 0.2347031, 0.3293256, 0.3286679, 0.3541003, 
    0.3157881, 0.268137, 0.2254309, 0.2056512, 0.2471392, 0.1567182, 
    0.2079777, 0.3086608, 0.1988217, 0.1772869, 0.2333164, 0.1615131, 
    0.1356572, 0.1021842, 0.1645586, 0.2315232, 0.1757971, 0.1391475, 
    0.1791123, 0.1635479, 0.1866197, 0.2693828,
  0.1708447, 0.05376191, 0.007166047, 0.08495875, 0.08885518, 0.08668866, 
    0.1476536, 0.1004074, 0.1167601, 0.05574477, 0.009040592, 0.004889166, 
    0.00403987, 0.05255701, 0.3627769, 0.07700305, 0.1053314, 0.1327657, 
    0.07052627, 0.07667801, 0.114865, 0.2124089, 0.1063879, 0.2953676, 
    0.08724498, 0.08917842, 0.09738763, 0.1128431, 0.194541,
  0.02634037, 0.01734164, 0.02329878, 0.00430335, 0.01000795, 0.02714799, 
    0.007155368, 0.02114408, 0.01791359, 0.003186838, 0.0002956114, 
    -2.758109e-06, 0.02224707, 0.01385076, 0.03273509, 0.04366335, 0.136157, 
    0.05133621, 0.05073044, 0.07822862, 0.04008091, 0.03965161, 0.04396776, 
    0.01539373, 0.04041986, 0.02177745, 0.02151483, 0.03072878, 0.01694015,
  0.03615839, 0.0005438847, 0.00348234, 0.001845777, 0.003339549, 
    0.008009792, 0.000186388, 0.003230268, 0.001928337, 3.335948e-05, 
    0.0001606726, 6.610696e-09, 0.0005909709, 0.03443353, 0.009252303, 
    0.01794786, 0.01002704, 0.008769465, 0.01312189, 0.0004450196, 
    0.006235151, 0.003122489, 0.03923976, 0.01227509, 0.04950979, 0.06577117, 
    0.002725047, 0.001064988, 0.02423269,
  0.06912838, 0.04289612, 0.0001331775, 0.06690108, 0.002117029, 0.007166298, 
    0.0006377273, 0.01063158, 0.001696371, 0.0004069504, 0.03880765, 
    0.0004824174, 0.02041632, 0.0006953306, 6.004276e-05, 0.0008458591, 
    9.73698e-05, 0.0003361517, 0.0002575104, 0.0005602656, 0.005690837, 
    0.01223378, 0.08773439, 0.007535828, 0.0002239926, 1.345938e-05, 
    -0.001278957, 0.001564305, 0.01016598,
  0.01633405, 0.02203628, 0.02166108, 0.04540537, 0.002304869, 0.01312032, 
    0.01393493, 0.002566732, 0.06655139, 0.0502474, 0.01314756, 0.007742481, 
    0.0004333257, 0.001049094, 0.01192412, 0.0007382716, 0.001193877, 
    0.0008691165, 0.0001584325, 8.424603e-05, 0.001629355, 0.01800888, 
    0.3085324, 0.1244184, 0.02409172, 0.0004512959, 0.003751478, 0.006523528, 
    0.00334801,
  8.409032e-05, -2.497761e-06, -1.486557e-07, 0.003188423, 0.006677777, 
    0.006538349, 0.01206639, 0.001745403, 0.0004153362, 0.00102833, 
    0.02194178, 0.003292503, 0.001650883, 0.0007378064, 0.0003750526, 
    0.003428384, 0.004508245, 0.01113528, 0.00920643, 0.01352878, 0.00882371, 
    0.01269152, 0.2176093, 0.02931667, 0.0004689718, 0.005445641, 0.01256005, 
    0.02794667, -0.0001897557,
  1.325729e-07, 2.339585e-08, 1.359159e-09, 6.335023e-09, 3.166692e-09, 
    1.45933e-05, -0.0002242337, 0.02482072, 0.07089984, 0.06391056, 
    0.005292994, 0.004226915, 0.00107215, 0.0001131634, 2.417133e-05, 
    0.003521482, 0.00678293, 0.005003612, 0.07872389, 0.1268793, 9.41682e-05, 
    0.05867908, 0.004232454, 0.005147463, 0.003455029, 0.02885041, 
    0.02066468, 0.006017949, 1.025064e-07,
  -1.044916e-07, 1.511419e-07, -1.091292e-06, 0.0001222078, 0.001361724, 
    7.35881e-08, -6.860052e-07, -4.474385e-05, 0.3060836, 0.0723802, 
    0.1028114, 0.223018, 0.2346807, 0.1223742, 0.1118552, 0.1797547, 
    0.1050793, 0.04992129, 0.080898, 0.125286, 0.0013594, 0.03237424, 
    0.004049329, 0.1052615, 0.1348975, 0.03966207, 0.04990344, 0.02923854, 
    0.02136699,
  0.007911599, 0.0007564098, 0.006331468, 0.1636926, 0.02039763, 
    1.456293e-07, 0.1000563, 0.002237447, -6.717718e-05, 0.01907022, 
    0.151116, 0.05495595, 0.1527701, 0.4021794, 0.4180212, 0.2362471, 
    0.2278057, 0.3107045, 0.2087292, 0.04510563, 0.00522235, 0.03955702, 
    0.06796859, 0.0813008, 0.1268943, 0.1844805, 0.1167654, 0.09685937, 
    0.1883346,
  0.09780587, 0.06624976, 0.09056414, 0.0603539, 0.01798295, 0.01204464, 
    0.01319108, 0.1364078, 0.0418083, 0.05753602, 0.0934716, 0.2589244, 
    0.2812855, 0.3431139, 0.377664, 0.3616333, 0.3824103, 0.2345469, 
    0.1602295, 0.1402987, 0.005828125, 0.01654037, 0.1131789, 0.2815815, 
    0.224795, 0.283919, 0.211715, 0.08684478, 0.1706089,
  0.02434273, 0.0318368, 0.07367985, 0.1239145, 0.16106, 0.1896744, 
    0.1321317, 0.09805476, 0.152537, 0.1259778, 0.1094718, 0.06743125, 
    0.1035098, 0.2299974, 0.38216, 0.4097909, 0.1815816, 0.2054237, 
    0.1486605, 0.07329909, 0.05744776, 0.1423914, 0.2017613, 0.2401204, 
    0.4062356, 0.1974218, 0.292941, 0.2922408, 0.05747677,
  0.08568473, 0.02338994, 0.0639092, 0.1233041, 0.1189277, 0.2182116, 
    0.1092494, 0.05277583, 0.02885831, 0.0337933, 0.08772572, 0.08799052, 
    0.08301821, 0.1539822, 0.1268689, 0.2173561, 0.1558389, 0.1618451, 
    0.2616208, 0.2133853, 0.4790657, 0.4588087, 0.2370151, 0.4206994, 
    0.5234381, 0.4026824, 0.144665, 0.1478141, 0.2529812,
  0.1956655, 0.2272109, 0.2521561, 0.2709903, 0.3173774, 0.4737029, 
    0.4818095, 0.4514453, 0.4989118, 0.417496, 0.3868387, 0.4158273, 
    0.3922449, 0.3771964, 0.3298087, 0.3024827, 0.3169705, 0.2495606, 
    0.1715064, 0.1780632, 0.1559649, 0.1749954, 0.1636226, 0.289629, 
    0.157689, 0.1765214, 0.1727138, 0.3092778, 0.2788908,
  0.1638406, 0.1553347, 0.1468288, 0.138323, 0.1298171, 0.1213112, 0.1128054, 
    0.1095106, 0.1161759, 0.1228412, 0.1295066, 0.1361719, 0.1428372, 
    0.1495025, 0.1823685, 0.1919615, 0.2015545, 0.2111475, 0.2207405, 
    0.2303336, 0.2399266, 0.2685409, 0.2607884, 0.2530359, 0.2452834, 
    0.237531, 0.2297785, 0.222026, 0.1706453,
  0.2580993, 0.2101724, 0.06701225, 0.08211489, 0.0339504, 0.03264625, 
    0.03220872, 0.05962793, 0.0007310432, 0.005323499, 0.03187731, 0.1938429, 
    0.3675962, -0.006927306, 0.2247294, 0.3240417, 0.3817052, 0.3012386, 
    0.2348743, 0.422128, 0.5949492, 0.7883973, 0.5626062, 0.3730182, 
    0.4110588, 0.3879938, 0.2277987, 0.1762101, 0.2197157,
  0.03681203, 0.009942585, 0.08133455, 0.05280655, 0.1991694, 0.1546383, 
    0.008801241, 0.2259315, 0.2358198, 0.3314549, 0.2671757, 0.2044473, 
    0.1343951, 0.128002, 0.3634707, 0.4758981, 0.3958288, 0.4392937, 
    0.277483, 0.2058471, 0.2894746, 0.3668457, 0.3843114, 0.6525793, 
    0.1919249, 0.5900417, 0.5570457, 0.4780649, 0.272837,
  0.1620376, 0.1880647, 0.1149989, 0.1214878, 0.1630548, 0.1266086, 
    0.1152771, 0.1209734, 0.1252009, 0.1231642, 0.1631452, 0.2160679, 
    0.3577897, 0.3750195, 0.2825567, 0.3256491, 0.2636779, 0.276513, 
    0.255719, 0.130817, 0.1653185, 0.2193527, 0.2113893, 0.176339, 0.2802149, 
    0.2904598, 0.2348731, 0.2277811, 0.2012072,
  0.2276067, 0.2108407, 0.1990583, 0.1952246, 0.2823456, 0.299566, 0.3202649, 
    0.2557903, 0.1995894, 0.1696721, 0.1464061, 0.164491, 0.1028154, 
    0.1378781, 0.2664072, 0.1500795, 0.1207312, 0.1790684, 0.1263267, 
    0.1058122, 0.08399761, 0.1430707, 0.1807621, 0.1566058, 0.1190183, 
    0.1314268, 0.12964, 0.1488814, 0.2391286,
  0.1452493, 0.03398035, 0.003885311, 0.05590272, 0.05437505, 0.05822928, 
    0.09270885, 0.06420065, 0.07116874, 0.03621556, 0.004661489, 0.002417386, 
    0.002278506, 0.02851044, 0.3239825, 0.05255752, 0.07315862, 0.1009519, 
    0.05318319, 0.05140839, 0.08217301, 0.1664597, 0.07292305, 0.286987, 
    0.06298076, 0.03710967, 0.06641325, 0.08014645, 0.1570086,
  0.01541082, 0.007774055, 0.02280768, 0.002510562, 0.004013747, 0.01077157, 
    0.003464273, 0.01166304, 0.01161317, 0.001660642, 0.0002974863, 
    -6.068295e-06, 0.01786231, 0.004026229, 0.0206669, 0.02469395, 
    0.07774726, 0.02920256, 0.03293661, 0.0403943, 0.01860333, 0.02641419, 
    0.02437361, 0.01414263, 0.03810553, 0.01446058, 0.01131617, 0.01321006, 
    0.00772501,
  0.01964627, 0.0004623572, 0.001855105, 0.001104144, 0.0008199607, 
    0.002309481, 5.030574e-05, 0.0003336146, 0.001160044, 3.109063e-05, 
    0.0003526457, 6.42136e-09, 0.0003481522, 0.0147109, 0.002099311, 
    0.006690449, 0.003085149, 0.003462877, 0.005754753, 0.0002363678, 
    0.002891819, 0.001556715, 0.02052972, 0.005714579, 0.03814337, 
    0.06034946, 0.001323144, 0.0004077475, 0.01151419,
  0.03479949, 0.03664548, -0.0002419075, 0.0436068, 0.0004152599, 
    0.002829097, 0.0001551208, 0.001596682, 0.0005065367, -0.001108544, 
    0.0278969, 0.0002623356, 0.005370775, 3.398083e-05, -7.210529e-06, 
    0.000405466, 4.992179e-05, 0.0001909967, 0.0001358303, 0.0003093646, 
    0.003026729, 0.00584741, 0.04543072, 0.003670393, 0.0001263617, 
    7.499478e-06, -0.00059776, 0.0007902096, 0.00504218,
  0.007698852, 0.04936659, 0.02469374, 0.03172317, 0.001121947, 0.006218724, 
    0.007849632, 0.001261561, 0.05250692, 0.04070792, 0.006299049, 
    0.004479707, 0.0001425924, 0.0005364177, 0.006183691, 0.0002259687, 
    0.0002249455, 0.0001580374, 7.573897e-05, 1.569062e-05, 0.0004509417, 
    0.005557448, 0.1418665, 0.1246249, 0.02209091, 6.083728e-05, 0.001071252, 
    0.003910326, 0.001443993,
  3.922347e-05, -1.583416e-06, -4.173163e-08, 0.004700556, 0.003678271, 
    0.003822371, 0.002329694, 0.0007934088, -0.0003724341, 0.0003334768, 
    0.008827124, 0.001227344, 0.0001110878, 3.072804e-05, 2.62321e-05, 
    0.0007097144, 0.0006798746, 0.003300063, 0.002237807, 0.006564674, 
    0.004901703, 0.005660895, 0.2029491, 0.02698365, 2.342527e-05, 
    0.001635941, 0.005869755, 0.01145319, -0.0004773399,
  1.265401e-07, 2.308446e-08, 1.282599e-09, 5.119182e-09, 3.089083e-09, 
    -3.157286e-05, -0.0002886193, 0.005005967, 0.05337167, 0.02802557, 
    0.002063516, 0.001083981, 0.0002221345, 5.689558e-05, 7.495246e-06, 
    0.0009000744, 0.002134322, 0.002616446, 0.04115038, 0.0818845, 
    3.438401e-07, 0.05005096, 0.001227506, -0.0002949, 0.001612556, 
    0.01327708, 0.01052041, 0.00317016, 9.969177e-08,
  3.563747e-08, 1.488692e-07, -9.020785e-07, -8.955957e-06, 0.0009530124, 
    7.222535e-08, -5.777391e-07, 0.002085695, 0.2833847, 0.05683515, 
    0.1087579, 0.1892736, 0.1687546, 0.0880754, 0.07036289, 0.12542, 
    0.06541492, 0.02288581, 0.04532949, 0.07296985, 0.0008444187, 0.02426773, 
    0.00153511, 0.06001354, 0.113849, 0.01555752, 0.03294864, 0.01366855, 
    0.01736088,
  0.006320807, 0.001468408, 0.004222246, 0.1509703, 0.01087508, 1.414341e-07, 
    0.08851501, 0.001363349, -6.431388e-05, 0.01301495, 0.1434441, 0.0595527, 
    0.1414755, 0.3870035, 0.3701026, 0.1765843, 0.1572292, 0.2710754, 
    0.1639507, 0.0417864, 0.003588356, 0.03126973, 0.04965092, 0.06900308, 
    0.08236884, 0.128713, 0.07618061, 0.06509542, 0.138768,
  0.06095287, 0.0521801, 0.07176408, 0.05001054, 0.01139596, 0.0080835, 
    0.01028021, 0.1203924, 0.03524261, 0.04705171, 0.07620537, 0.2346634, 
    0.2499969, 0.3006776, 0.3341929, 0.2949102, 0.3097048, 0.1903523, 
    0.1647347, 0.1177227, 0.003726385, 0.01194316, 0.0936879, 0.2559152, 
    0.1864174, 0.2410189, 0.1520203, 0.04593261, 0.1183678,
  0.01641677, 0.02336658, 0.06247227, 0.1058169, 0.1370007, 0.1623052, 
    0.1159658, 0.08493657, 0.1325485, 0.1085353, 0.1003293, 0.05018615, 
    0.08089815, 0.1853692, 0.3345393, 0.3717134, 0.1481238, 0.1639979, 
    0.1335429, 0.06778856, 0.05106224, 0.1008208, 0.2203391, 0.2408307, 
    0.3405642, 0.157142, 0.2395598, 0.2553895, 0.03337825,
  0.06181215, 0.01436411, 0.05268507, 0.09681949, 0.09916729, 0.192709, 
    0.09176484, 0.03541107, 0.02191652, 0.02639264, 0.06099053, 0.0563903, 
    0.07846791, 0.1343286, 0.1071931, 0.206654, 0.1367199, 0.1495811, 
    0.2645876, 0.1985249, 0.4358059, 0.4299834, 0.189718, 0.3840693, 
    0.4549818, 0.3380386, 0.1318906, 0.1237828, 0.2173869,
  0.1578325, 0.2015494, 0.3239189, 0.3027522, 0.3188198, 0.4123059, 0.466344, 
    0.4179686, 0.4291017, 0.3935642, 0.3893108, 0.390998, 0.3861986, 
    0.3811787, 0.2647535, 0.2897528, 0.3086131, 0.2298405, 0.1604416, 
    0.1720074, 0.1743077, 0.1852224, 0.1141347, 0.2471058, 0.1366914, 
    0.1317144, 0.1456202, 0.2947589, 0.2305744,
  0.1325901, 0.124773, 0.1169559, 0.1091389, 0.1013218, 0.09350474, 
    0.08568767, 0.0542624, 0.05990139, 0.06554039, 0.07117938, 0.07681837, 
    0.08245736, 0.08809636, 0.1333268, 0.1432252, 0.1531236, 0.163022, 
    0.1729204, 0.1828188, 0.1927172, 0.1966792, 0.1889589, 0.1812386, 
    0.1735183, 0.1657979, 0.1580776, 0.1503573, 0.1388437,
  0.2852113, 0.1308956, 0.07156186, 0.02541386, 0.0009953415, 0.006397747, 
    0.004488195, 0.008926769, 0.02721231, 0.03690285, 0.02204792, 0.1485681, 
    0.3075838, -0.008937417, 0.3374715, 0.3815563, 0.3294517, 0.2710194, 
    0.2136659, 0.389128, 0.572473, 0.790086, 0.5015061, 0.3106304, 0.3914497, 
    0.4427109, 0.2149354, 0.1413639, 0.1942936,
  0.04918265, 0.005476454, 0.06532447, 0.04267117, 0.1823372, 0.1301953, 
    0.003988433, 0.1517419, 0.1963763, 0.2509579, 0.2096426, 0.2253164, 
    0.1215599, 0.1207938, 0.3650925, 0.4304262, 0.3831678, 0.3759368, 
    0.2284965, 0.1790684, 0.2600604, 0.313851, 0.3418661, 0.5896098, 
    0.2154624, 0.5939749, 0.4887188, 0.4045994, 0.2595081,
  0.1136773, 0.1362136, 0.08380835, 0.08227946, 0.1162758, 0.08944529, 
    0.08480729, 0.09214158, 0.09175424, 0.08438606, 0.1263838, 0.172191, 
    0.307353, 0.2991408, 0.2079579, 0.2304757, 0.2019874, 0.2115254, 
    0.1989053, 0.09812687, 0.1264607, 0.15631, 0.1501958, 0.12053, 0.2116381, 
    0.2284902, 0.1760929, 0.1716933, 0.1348985,
  0.1914558, 0.1816129, 0.1598892, 0.1510088, 0.2328009, 0.2499446, 
    0.2738224, 0.1962257, 0.1398211, 0.1199237, 0.1001899, 0.1053031, 
    0.06685913, 0.08476712, 0.2179183, 0.1082746, 0.08280848, 0.123404, 
    0.08022647, 0.07539909, 0.05733382, 0.1006463, 0.1327751, 0.1402563, 
    0.0988967, 0.09450704, 0.09397313, 0.1153053, 0.2062355,
  0.1044697, 0.02082211, 0.002264905, 0.03129955, 0.02802043, 0.03528858, 
    0.05500088, 0.03637223, 0.04105334, 0.02491825, 0.002604116, 0.001462352, 
    0.001640042, 0.01638533, 0.2911485, 0.0337536, 0.04927573, 0.06460695, 
    0.03483665, 0.03205595, 0.04340676, 0.1230447, 0.04388541, 0.2709185, 
    0.04452411, 0.01848708, 0.03994641, 0.04705219, 0.1177217,
  0.009198482, 0.004905369, 0.02121185, 0.001518294, 0.001906092, 
    0.005228632, 0.001809995, 0.007383402, 0.008726021, 0.001081725, 
    5.637591e-05, -6.133025e-06, 0.01301574, 0.001382969, 0.01130738, 
    0.01332084, 0.04650261, 0.01463489, 0.02051153, 0.01898976, 0.009004519, 
    0.01507473, 0.0141745, 0.01175285, 0.03720878, 0.007823843, 0.005029289, 
    0.006695408, 0.004540413,
  0.01298594, 6.64803e-05, 0.0006946428, 0.0007626406, -0.0006065577, 
    0.0007285164, 2.336262e-05, 0.0001541384, 0.0008222779, 3.129822e-05, 
    0.0001881951, 6.369007e-09, 0.00023876, 0.007079502, 0.001137738, 
    0.003583099, 0.001481883, 0.00152499, 0.002568982, 0.0001579292, 
    0.001553264, 0.0009646083, 0.01313885, 0.003616437, 0.02792293, 
    0.0614486, 0.0008837288, 0.0002482787, 0.007171214,
  0.02170014, 0.02743985, -0.0004336254, 0.02575665, 0.0001378406, 
    0.001603798, 9.157502e-05, 0.0003762691, 0.0002657385, -0.0006766063, 
    0.01776599, 0.0001655831, 0.0003669978, 1.063755e-05, -4.309185e-06, 
    0.0002442385, 3.258839e-05, 0.0001284096, 8.643721e-05, 0.000201296, 
    0.001952854, 0.003555049, 0.02890087, 0.006580174, 0.0003857531, 
    4.286004e-06, -0.0002473744, 0.0004892964, 0.003171775,
  0.004717178, 0.06838027, 0.01964265, 0.02295541, 0.0006892869, 0.002663333, 
    0.003998753, 0.0008051487, 0.03898832, 0.039002, 0.002790549, 
    0.002241066, 7.574332e-05, 0.0003415986, 0.003142197, 0.0001287725, 
    8.025078e-05, 6.16975e-05, 4.600607e-05, 8.227737e-06, 0.0002475778, 
    0.003155773, 0.08351849, 0.1041435, 0.02117013, 3.852386e-05, 
    0.0006379028, 0.001651442, 0.0009005493,
  2.624888e-05, -7.474026e-07, -9.524462e-09, 0.004717723, 0.001854114, 
    0.002576384, -0.001171628, 0.0005163956, -0.0002528224, 0.0001412096, 
    0.003494452, 0.0006566981, 4.218631e-05, 3.21295e-05, 2.382602e-05, 
    0.000250923, 0.0002195249, 0.001389318, 0.001074033, 0.004256667, 
    0.003296071, 0.002543398, 0.1736259, 0.03045183, 1.355005e-05, 
    0.0006649586, 0.003523271, 0.006918352, -0.0004466733,
  1.270508e-07, 2.252137e-08, 1.252563e-09, 2.190917e-09, 3.04125e-09, 
    -2.027378e-05, -0.000188601, 0.002259698, 0.03958104, 0.009343683, 
    0.0009920644, 0.0004516015, 9.116411e-05, 3.554392e-05, 3.618979e-06, 
    0.0005062146, 0.001210972, 0.00167249, 0.02622835, 0.0596962, 
    -2.502801e-06, 0.0423809, 0.0003623828, -0.001358726, 0.0009984197, 
    0.00810009, 0.00660661, 0.001997641, 9.860165e-08,
  6.118371e-08, 1.484649e-07, -3.383828e-07, -2.884846e-05, 0.0007345834, 
    7.356662e-08, -5.506249e-07, 0.003521717, 0.2542062, 0.0344309, 
    0.09081834, 0.1360926, 0.1142316, 0.04816996, 0.047604, 0.08464387, 
    0.03577947, 0.01152063, 0.02956585, 0.04845989, 0.0005498509, 0.01730072, 
    0.0005061487, 0.03190872, 0.0702191, 0.007583763, 0.02198069, 
    0.006749153, 0.01630249,
  0.003959327, 0.0004151519, 0.002590481, 0.1320962, 0.007451692, 
    1.387021e-07, 0.07627046, 0.0009472911, -5.700974e-05, 0.008559639, 
    0.1252543, 0.06977036, 0.1342897, 0.3494721, 0.2901928, 0.1243443, 
    0.1031711, 0.2164223, 0.1326563, 0.03628729, 0.002681899, 0.02051153, 
    0.03486504, 0.05522347, 0.05193541, 0.0741557, 0.04477844, 0.03641916, 
    0.09217338,
  0.03551925, 0.04219207, 0.05122621, 0.04219643, 0.007355614, 0.004318891, 
    0.008538065, 0.1069797, 0.03038172, 0.03750005, 0.06225463, 0.2095837, 
    0.2283288, 0.2449562, 0.2800696, 0.2400499, 0.2271309, 0.1288223, 
    0.1401648, 0.09929539, 0.001616205, 0.01098025, 0.07417698, 0.2240212, 
    0.1461348, 0.1936503, 0.09561685, 0.02480553, 0.07247338,
  0.01009819, 0.01596223, 0.05279411, 0.08286401, 0.1113981, 0.1327646, 
    0.09601571, 0.06924487, 0.1145631, 0.08986791, 0.09206562, 0.03818716, 
    0.065685, 0.1362773, 0.2628166, 0.3150172, 0.1233201, 0.1328351, 
    0.115266, 0.06201738, 0.04232757, 0.07861277, 0.2436921, 0.2428189, 
    0.2682407, 0.1421486, 0.1833935, 0.1774834, 0.0212436,
  0.04363925, 0.0100828, 0.04755254, 0.08109758, 0.08013846, 0.1484967, 
    0.07815379, 0.02614827, 0.02285199, 0.02572699, 0.04554005, 0.04137082, 
    0.07963806, 0.1136282, 0.0833851, 0.1735461, 0.1173869, 0.137423, 
    0.2620957, 0.2130172, 0.3832978, 0.3652755, 0.1514679, 0.3356613, 
    0.3662146, 0.2910409, 0.1342566, 0.1109299, 0.1871722,
  0.1475583, 0.1794603, 0.2387412, 0.2734975, 0.2372502, 0.325006, 0.3653078, 
    0.3424092, 0.3648969, 0.3418535, 0.3173668, 0.3386565, 0.3031538, 
    0.3035103, 0.207757, 0.2494219, 0.2668542, 0.2044027, 0.1462772, 
    0.1542224, 0.1782732, 0.177158, 0.08538361, 0.217026, 0.113428, 
    0.1032909, 0.118667, 0.2680497, 0.1829453,
  0.1097378, 0.1046833, 0.0996289, 0.09457447, 0.08952003, 0.08446559, 
    0.07941116, 0.07414467, 0.07781326, 0.08148185, 0.08515044, 0.08881903, 
    0.09248763, 0.09615622, 0.1018885, 0.1096976, 0.1175066, 0.1253157, 
    0.1331247, 0.1409338, 0.1487428, 0.1564144, 0.1499912, 0.143568, 
    0.1371448, 0.1307216, 0.1242984, 0.1178752, 0.1137813,
  0.3703603, 0.09421147, 0.05608642, 0.006970232, 0.00135098, 0.007220123, 
    0.005599548, 0.003772465, 0.002122047, 0.02557866, 0.03189069, 
    0.08869485, 0.2597118, -0.007794089, 0.4454839, 0.3823479, 0.3087469, 
    0.2424894, 0.1694117, 0.4426927, 0.5455712, 0.7893414, 0.4541293, 
    0.26928, 0.3611453, 0.4603051, 0.2172244, 0.1316446, 0.1788244,
  0.05983742, 0.008220697, 0.05168947, 0.03549312, 0.1650369, 0.1126771, 
    0.00209055, 0.1191334, 0.17487, 0.1864996, 0.1943059, 0.2321011, 
    0.1103941, 0.1174604, 0.3687629, 0.3942964, 0.3630112, 0.3274006, 
    0.2019243, 0.1608799, 0.2483139, 0.2809708, 0.3077339, 0.5139805, 
    0.2389031, 0.5311374, 0.4106434, 0.3312194, 0.2404081,
  0.08770049, 0.1040131, 0.06672448, 0.06228759, 0.0893158, 0.07179875, 
    0.06750318, 0.07106172, 0.07024379, 0.06185402, 0.1028775, 0.1452271, 
    0.2653589, 0.2461613, 0.1590948, 0.1751191, 0.1608948, 0.1732761, 
    0.1587145, 0.07818501, 0.09874749, 0.1175944, 0.1165553, 0.08681854, 
    0.1647489, 0.1905297, 0.1453267, 0.1334281, 0.1021705,
  0.1614755, 0.157835, 0.1390568, 0.1266823, 0.1986536, 0.2216027, 0.2451625, 
    0.1562727, 0.1043136, 0.08975358, 0.07055236, 0.07285804, 0.04423448, 
    0.05602214, 0.1836082, 0.07898594, 0.06097723, 0.08089127, 0.05384718, 
    0.05497746, 0.03796179, 0.07496086, 0.1018427, 0.1426897, 0.07598309, 
    0.06873981, 0.07105448, 0.09292293, 0.1801555,
  0.06931009, 0.01140139, 0.001550227, 0.01659302, 0.01591841, 0.01934731, 
    0.03464871, 0.0225011, 0.02521251, 0.01673749, 0.001913824, 0.001047673, 
    0.001330166, 0.009668605, 0.2611956, 0.02088165, 0.03344049, 0.04462676, 
    0.02129877, 0.02057674, 0.02411349, 0.08616337, 0.02700902, 0.2535281, 
    0.03266023, 0.0093592, 0.02434029, 0.02683265, 0.08413611,
  0.006258318, 0.003638817, 0.02041392, 0.001140015, 0.001302488, 
    0.003383663, 0.0009321431, 0.005196261, 0.006227472, 0.0008242704, 
    2.57232e-05, -4.371177e-06, 0.01385513, 0.0007686288, 0.00525745, 
    0.0057353, 0.02864206, 0.007741562, 0.01287034, 0.01054306, 0.005008319, 
    0.008075719, 0.009873771, 0.01033289, 0.0327014, 0.004090811, 
    0.002187561, 0.003930074, 0.003286037,
  0.009689844, -5.258697e-05, 0.0001681739, 0.0005753127, -0.0008734284, 
    0.0003803525, 1.437887e-05, 0.0001084607, 0.0006338001, 2.683698e-05, 
    8.264266e-05, 6.362576e-09, 0.0001827737, 0.003785764, 0.00079087, 
    0.002445193, 0.001007081, 0.0007831192, 0.00120129, 0.0001183122, 
    0.001004235, 0.0006912563, 0.009606181, 0.002628636, 0.0237602, 
    0.06046572, 0.000638603, 0.0001778308, 0.005173541,
  0.01547081, 0.0167418, -0.0002832834, 0.01787611, 7.874982e-05, 
    0.001132915, 6.279745e-05, 0.0001881363, 0.0001943633, -0.0004385907, 
    0.01229314, 0.0001217152, -0.0003530231, 1.169392e-05, -3.146495e-06, 
    0.0001715016, 2.469999e-05, 9.704407e-05, 6.320807e-05, 0.0001490366, 
    0.001438563, 0.002525006, 0.02107329, 0.01389427, 0.0009224244, 
    1.91253e-05, -9.987644e-05, 0.0003516416, 0.002319432,
  0.003358836, 0.06972004, 0.01440391, 0.01684837, 0.000492979, 0.001128732, 
    0.00223535, 0.000590189, 0.03017911, 0.04670194, 0.00130503, 0.001287002, 
    4.973464e-05, 0.0002488534, 0.00161405, 9.161331e-05, 5.395259e-05, 
    3.600131e-05, 3.293196e-05, 5.93694e-06, 0.0001677367, 0.00216536, 
    0.05894665, 0.06872129, 0.01756341, 3.087119e-05, 0.0004657302, 
    0.0008797162, 0.0006589348,
  0.0001374026, -3.394716e-07, 1.852856e-08, 0.003064155, 0.0009762871, 
    0.001934758, -0.001323288, 0.0003697031, -0.0001441484, 9.857582e-05, 
    0.00186401, 0.0003103657, 2.941652e-05, 3.326095e-05, 2.042744e-05, 
    0.0001545798, 0.0001095924, 0.0008025797, 0.0007172805, 0.003138183, 
    0.00248036, 0.001311496, 0.1585271, 0.0365505, 7.620032e-06, 0.000356506, 
    0.002490828, 0.004926202, 0.0005377528,
  1.289704e-07, 2.165753e-08, 1.227801e-09, -5.979897e-10, 3.021843e-09, 
    -1.448136e-05, -0.000125659, 0.001461912, 0.03952584, 0.004797843, 
    0.0006710378, 0.0002763699, 5.180991e-05, 2.585855e-05, 2.570343e-06, 
    0.0003570193, 0.0009217464, 0.001222254, 0.01907557, 0.04717182, 
    -3.410423e-06, 0.03512725, 0.0001796192, -0.001530686, 0.000710891, 
    0.005848766, 0.004773733, 0.001450201, 9.847781e-08,
  6.699531e-08, 1.496576e-07, -2.500514e-07, -2.20326e-05, 0.0005827478, 
    7.059183e-08, -1.166881e-06, 0.00469423, 0.2367903, 0.01977911, 
    0.06930829, 0.08144312, 0.07675772, 0.03194354, 0.03286892, 0.05595405, 
    0.02065812, 0.007591485, 0.02203356, 0.0360221, 0.0003936167, 0.01242032, 
    0.0007020999, 0.01777773, 0.03487393, 0.004807283, 0.01458594, 
    0.00412243, 0.01219353,
  0.001762975, 0.0001433518, 0.001845121, 0.1183969, 0.005792318, 
    1.358659e-07, 0.06673036, 0.0007583487, -5.215345e-05, 0.005929676, 
    0.107511, 0.07109597, 0.1241893, 0.3004299, 0.2185737, 0.08959582, 
    0.06999453, 0.156432, 0.09450039, 0.03626101, 0.002594173, 0.01505212, 
    0.02310226, 0.0449038, 0.03763876, 0.04483433, 0.02760712, 0.02096933, 
    0.06388313,
  0.02381445, 0.03289269, 0.03575135, 0.03442872, 0.005237341, 0.002806247, 
    0.007387984, 0.09714399, 0.02854561, 0.03208062, 0.05191758, 0.1945557, 
    0.1808701, 0.1985892, 0.2299038, 0.1982798, 0.1613922, 0.08862659, 
    0.1055197, 0.08759195, 0.001408839, 0.009448572, 0.05986502, 0.1980049, 
    0.1169911, 0.1486405, 0.06162329, 0.01555267, 0.04811344,
  0.006405818, 0.0116402, 0.04421891, 0.07042821, 0.09605863, 0.1106884, 
    0.08313151, 0.06044285, 0.1043703, 0.07832855, 0.08162002, 0.02960993, 
    0.05671808, 0.1157299, 0.2075062, 0.2657409, 0.1040054, 0.1121237, 
    0.1067863, 0.05518108, 0.03980977, 0.07417513, 0.2244481, 0.2401791, 
    0.2071726, 0.1244473, 0.1343282, 0.1123455, 0.01429533,
  0.03105446, 0.008228135, 0.04499611, 0.06613547, 0.0743629, 0.1229466, 
    0.07661133, 0.03541826, 0.03545632, 0.03104549, 0.04001373, 0.03684749, 
    0.09174085, 0.1037258, 0.07922582, 0.1652607, 0.131092, 0.1263268, 
    0.2362257, 0.202857, 0.3389642, 0.3130053, 0.1389115, 0.3003405, 
    0.3196017, 0.2472085, 0.1560706, 0.1018499, 0.1609401,
  0.123186, 0.1570685, 0.1882002, 0.1817263, 0.1730318, 0.2294533, 0.2420376, 
    0.2280748, 0.286613, 0.2657239, 0.2289864, 0.2684371, 0.2208188, 
    0.2058373, 0.1665686, 0.2165776, 0.180311, 0.1642437, 0.1308276, 
    0.1222314, 0.1559462, 0.1637257, 0.07200851, 0.1980266, 0.0970061, 
    0.08392487, 0.1047132, 0.2496302, 0.1684233,
  0.1035665, 0.09938545, 0.0952044, 0.09102335, 0.0868423, 0.08266126, 
    0.07848021, 0.07010201, 0.07290033, 0.07569864, 0.07849696, 0.08129528, 
    0.0840936, 0.08689192, 0.0954553, 0.1024744, 0.1094934, 0.1165125, 
    0.1235316, 0.1305507, 0.1375698, 0.1421279, 0.1364916, 0.1308552, 
    0.1252189, 0.1195825, 0.1139462, 0.1083098, 0.1069113,
  0.30685, 0.0655206, 0.03910422, 0.0053244, 0.0009206465, 0.006235758, 
    0.005546478, 0.003924155, 0.001449674, 0.01693803, 0.02236959, 
    0.08218847, 0.2383142, -0.006666271, 0.5643011, 0.3771947, 0.2466092, 
    0.2463768, 0.1677826, 0.4685898, 0.5154152, 0.7649462, 0.4368799, 
    0.2628313, 0.337417, 0.460489, 0.2234803, 0.1263617, 0.1924764,
  0.06386926, 0.02470638, 0.04860178, 0.03232714, 0.1672942, 0.09239901, 
    0.001444773, 0.1097582, 0.1663353, 0.1740729, 0.17464, 0.2310057, 
    0.1086722, 0.1154978, 0.3638074, 0.3858128, 0.3587729, 0.3013169, 
    0.1871172, 0.1431997, 0.2278996, 0.2770616, 0.2950133, 0.4700288, 
    0.2424559, 0.4821455, 0.3558314, 0.289615, 0.2209075,
  0.07462894, 0.08861214, 0.05801131, 0.05282987, 0.07617709, 0.0637639, 
    0.05932838, 0.05967683, 0.05765001, 0.05134673, 0.08972823, 0.1295668, 
    0.2308005, 0.2125605, 0.1358311, 0.1496765, 0.1409735, 0.1557932, 
    0.1373537, 0.06851607, 0.08247849, 0.09691808, 0.0976396, 0.071311, 
    0.1416444, 0.17212, 0.130555, 0.112682, 0.08676675,
  0.1392943, 0.1369625, 0.1223512, 0.1100291, 0.1752302, 0.1891829, 
    0.2136957, 0.1313696, 0.08868778, 0.07489965, 0.05692262, 0.05722606, 
    0.03387496, 0.0428962, 0.1446386, 0.05978199, 0.0491685, 0.05660203, 
    0.04107695, 0.04524978, 0.02928856, 0.05877272, 0.08154061, 0.1700152, 
    0.05616622, 0.05339836, 0.059839, 0.07783309, 0.152204,
  0.05345255, 0.007937199, 0.001247062, 0.01080685, 0.01112201, 0.01345044, 
    0.02598567, 0.01587393, 0.01832508, 0.01143934, 0.001627219, 
    0.0008752822, 0.001166038, 0.007290104, 0.2729458, 0.01355902, 
    0.02211992, 0.03362512, 0.01363168, 0.01379635, 0.01570906, 0.05694488, 
    0.0186705, 0.2660232, 0.02589807, 0.005829629, 0.01513249, 0.01762617, 
    0.06226692,
  0.004953525, 0.003011797, 0.02660869, 0.0009639825, 0.001088564, 
    0.002608678, 0.0007140283, 0.004158251, 0.004595378, 0.0006717346, 
    1.798139e-05, -2.498084e-06, 0.0169541, 0.0005732112, 0.002877181, 
    0.003235187, 0.01614274, 0.005034645, 0.008599746, 0.006490083, 
    0.003576192, 0.005237118, 0.007839263, 0.009802558, 0.04473928, 
    0.002566162, 0.001327112, 0.00289102, 0.00271169,
  0.008085565, -8.441433e-05, -9.197032e-05, 0.0004830965, -0.0009860601, 
    0.0002777331, 1.137594e-05, 8.968321e-05, 0.0003418127, 2.384521e-05, 
    6.029238e-05, 6.3794e-09, 0.0001548956, 0.002429387, 0.0006356593, 
    0.001881082, 0.0007660023, 0.0005611492, 0.0007723792, 9.777937e-05, 
    0.0007624302, 0.0005614584, 0.007908085, 0.002137732, 0.05071891, 
    0.06576473, 0.000525997, 0.0001443204, 0.004222802,
  0.01248937, 0.008802988, -0.0003990251, 0.0205781, 5.868084e-05, 
    0.000900495, 5.158411e-05, 0.0001453114, 0.0001632164, -0.0004044362, 
    0.009672146, 0.0001031303, -0.0003793439, 1.266368e-05, -2.214933e-06, 
    0.0001385779, 2.112672e-05, 9.323236e-05, 5.30254e-05, 0.0001250707, 
    0.001195501, 0.002064785, 0.01727136, 0.04712318, 0.02291454, 
    0.0004721858, -7.021453e-05, 0.0002910694, 0.001928417,
  0.002710064, 0.1044819, 0.01892047, 0.01838203, 0.000395153, 0.0006722822, 
    0.001484427, 0.0004843838, 0.03726077, 0.09777156, 0.0008520679, 
    0.0008973706, 3.817444e-05, 0.0002025675, 0.001015755, 7.483097e-05, 
    4.286767e-05, 2.68453e-05, 2.720827e-05, 5.570438e-06, 0.0001349917, 
    0.001759342, 0.04655586, 0.06553572, 0.06238104, 2.557475e-05, 
    0.000380246, 0.0006221178, 0.0005430904,
  0.004470002, -9.294237e-07, -1.109425e-06, 0.002662752, 0.0006842598, 
    0.00160466, -0.002913975, 0.0003027029, -0.001643621, 8.453508e-05, 
    0.001345163, 0.0002089863, 2.690364e-05, 2.925442e-05, 1.789523e-05, 
    0.0001170155, 8.478478e-05, 0.0006403975, 0.0005865248, 0.002572138, 
    0.002056817, 0.0008596131, 0.2345557, 0.05560306, 5.281031e-06, 
    0.0002711971, 0.002029133, 0.003957922, 0.02466694,
  1.295441e-07, 2.120022e-08, 1.235602e-09, -7.413451e-10, 3.041096e-09, 
    -1.140076e-05, -9.228406e-05, 0.0009467413, 0.07755069, 0.002845016, 
    0.0005429136, 0.0002100326, 3.901344e-05, 2.173684e-05, 2.220423e-06, 
    0.0002903629, 0.0007843837, 0.001020379, 0.01565976, 0.04045416, 
    -3.602993e-06, 0.03232295, 0.0001299131, -0.001722356, 0.0005774659, 
    0.004742151, 0.003907837, 0.001205828, 9.896686e-08,
  7.00773e-08, 1.513919e-07, -2.04047e-07, -1.426059e-05, 0.0004914041, 
    7.231225e-08, -2.280106e-06, 0.00650484, 0.2503097, 0.02516378, 
    0.05182718, 0.04764972, 0.05107159, 0.0209721, 0.02503416, 0.03343171, 
    0.01349474, 0.005535996, 0.018209, 0.02943882, 0.0003003847, 0.01590059, 
    0.006296007, 0.0113169, 0.01815316, 0.003464446, 0.01027373, 0.003099176, 
    0.009362955,
  0.001109836, -6.011539e-05, 0.001594406, 0.1145927, 0.00491426, 
    1.345931e-07, 0.06080841, 0.0006602286, -4.790282e-05, 0.004595545, 
    0.1018433, 0.05824548, 0.1006528, 0.2219794, 0.1763107, 0.07226302, 
    0.05271459, 0.1157562, 0.07151202, 0.04081344, 0.003280072, 0.01172391, 
    0.01703757, 0.03324109, 0.0307874, 0.03088857, 0.01908221, 0.01438921, 
    0.04770008,
  0.01721506, 0.02891466, 0.02921794, 0.03116667, 0.004153071, 0.002232981, 
    0.006841626, 0.09389102, 0.03230577, 0.03335361, 0.06159069, 0.1983889, 
    0.1402705, 0.1660609, 0.1864891, 0.1710531, 0.1280437, 0.06620771, 
    0.08567147, 0.08868612, 0.00093128, 0.01014533, 0.06667602, 0.2171396, 
    0.1053406, 0.1194176, 0.04566871, 0.01143728, 0.03067236,
  0.004908656, 0.01189778, 0.039706, 0.07258524, 0.1024926, 0.1197563, 
    0.082013, 0.08295342, 0.1145806, 0.08497965, 0.08772034, 0.02978275, 
    0.0776788, 0.1189004, 0.175211, 0.2319213, 0.1060914, 0.103715, 
    0.1286728, 0.05377972, 0.0443635, 0.09798502, 0.2028342, 0.2439729, 
    0.1783019, 0.1064972, 0.1052992, 0.08443335, 0.01108373,
  0.02509598, 0.007494209, 0.04830093, 0.05728787, 0.09573448, 0.1159503, 
    0.09656008, 0.07047655, 0.06839379, 0.05948175, 0.06542138, 0.04337864, 
    0.1255037, 0.09244807, 0.08951169, 0.1528498, 0.1745559, 0.132455, 
    0.2317663, 0.176143, 0.3132985, 0.2766394, 0.1599356, 0.284878, 
    0.2869883, 0.2180579, 0.2044016, 0.1058659, 0.1388142,
  0.1348878, 0.1391018, 0.1561866, 0.1358555, 0.1363049, 0.1952482, 
    0.1961462, 0.169794, 0.2114407, 0.2137058, 0.1849761, 0.2174565, 
    0.1813359, 0.1726138, 0.1458755, 0.1909464, 0.1422631, 0.1416548, 
    0.1182652, 0.1068142, 0.1332764, 0.1508678, 0.06776903, 0.1854817, 
    0.08864737, 0.07366861, 0.09623438, 0.2323913, 0.1899768,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -6.342386e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0004205892, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001735706, 0.0008495311, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -5.96966e-07, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, -3.245306e-05, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 5.442294e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 6.860822e-06, 0, 0, 0, 0, -7.087373e-06, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, -1.618534e-05, 0.0127431, 0.001716627, 0, 0, 0, 
    0, 0, 0, 5.788525e-05, 0, 0, -2.9914e-05, 0, 0, 0, 0, 0.00138384, 0, 0,
  0, 0, 0, 0, 0, 0, 1.871917e-06, 0, 0, 2.340706e-05, 0, 0.0001482248, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, -0.000102098, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0.0005231446, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, -2.136875e-06, 0, -8.581025e-06, 0, -5.150179e-05, 0, 
    0.0006879269, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 9.635152e-05, 0, 0, 0, 0, 0, 2.014572e-05, 0, 0, 0, -4.885477e-11, 
    -5.799434e-05, -6.183608e-06, 2.592714e-05, -1.862892e-06, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, -9.563719e-05, 0.01977615, 0.002711005, 
    -8.793252e-11, 0.0003916571, 0, -5.909663e-05, 0, 0, 0.0008393262, 0, 
    0.0001337681, -0.0002842195, 0, 0, 0, -1.249362e-05, 0.002459488, 
    -3.122435e-05, 0.0008750577,
  0, 0, 0, 0, 0, 0, 0.0003772757, 0, 0, 2.118975e-05, 7.258976e-06, 
    0.001670827, 0, 0, 0, 0, 0, 0, 0, 0, 0, -7.402634e-06, 0.0001923707, 0, 
    0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0.0008934474, 0, -1.458893e-05, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8.228584e-05, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.108377e-06, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0.003088254, 0, 0.001738238, 0, -8.014176e-05, 0, 5.350093e-05, 
    -7.338533e-06, 0.006398053, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0.0001586558, 0, 0, 0, 0, 0, 6.149001e-05, 0.0005091438, 0, 0, 
    -3.300753e-05, 0.0008060274, -2.267629e-05, 0.001814428, -9.870305e-06, 
    1.314081e-05, 0, 0, 0, 0, 0, 0, 0.002563418, -1.250827e-05, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, -9.105158e-05, 0.02791714, 0.005643677, 
    0.002311772, 0.0009383481, 2.674919e-05, -0.0001302569, -3.357912e-05, 
    -5.9825e-05, 0.001352314, 0, 0.0004792959, 0.003684592, -0.0001473303, 0, 
    -1.760366e-05, -7.18571e-05, 0.004539766, 0.001684006, 0.002123941,
  0, 0, 0, 0, 0, -9.046737e-06, 0.006766476, 9.166759e-05, 0, 0.002142925, 
    2.215855e-06, 0.01252668, 0, 0, 0, 0, 0, 0, 0, 0, 0, -6.629505e-05, 
    0.002161752, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, -1.208927e-05, 0.002639116, -2.682527e-05, 
    -8.004777e-05, -6.685972e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001523888, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3.883885e-05, -2.37243e-05, -9.224489e-06, -5.040381e-06, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -2.832067e-05, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3.819614e-05, -1.303445e-05, 0, 
    0, 0, 8.517634e-05, -4.764423e-06, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -5.739249e-06, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0.004929956, 0, 0.004203972, -9.157591e-06, 6.515581e-05, 0, 
    0.001225072, 7.995551e-06, 0.01079161, -4.081506e-05, 6.248865e-05, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0.000232029, -7.724318e-06, 0, 0, 0, 0, -8.632636e-05, 0.001190248, 
    -3.430328e-06, 4.967672e-06, -6.265692e-05, 0.001866304, 0.0005319939, 
    0.002399262, -2.670593e-05, 0.0005369198, 0, 0, 0, 0, 0, -6.769491e-09, 
    0.004419196, 2.44691e-05, 0, -1.190027e-05, 0, 0,
  0, 0, 0, 0, 0, 0, 0, -9.718907e-06, -2.098495e-05, 0.001908925, 0.04053114, 
    0.01581791, 0.005097202, 0.001799321, 0.002626441, 0.0005126832, 
    -9.998952e-05, -0.0001510712, 0.001665955, -6.109474e-06, 0.001628999, 
    0.01000831, 0.0001985195, 0, 0.0001991372, -0.0001259967, 0.006381037, 
    0.005728374, 0.004918064,
  0, 0, 0, 0, 0, -8.5694e-05, 0.01342009, 0.0006349557, -1.191379e-05, 
    0.008459889, 0.005848968, 0.03369533, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -0.0001163006, 0.007139314, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, -0.000171121, 0.003475837, -0.0001310593, 0.001828718, 
    0.005148589, -5.606404e-06, 0, 0, 0, -1.124491e-05, 0, 0, 0, 0, 0, 0, 0, 
    -1.650212e-05, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -5.852925e-05, 0, 0.003875511, 0.001286442, 
    0.000157632, 0, 0, 0, 0, 0, 0, 0, 0.004501072, -0.0001344824, 
    -2.478488e-05, -3.543865e-05, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.00147695, 
    0, 9.171361e-05, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, -5.39459e-07, 4.553324e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, -1.664044e-05, 0, 0, 0, 0, 0, -5.915803e-07, 0, 0, 0,
  0, 0, 0, 5.388694e-05, -2.138131e-08, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.005609586, 0.0001502809, 0.0007321388, 0, -4.566528e-06, 0.002684842, 
    -5.959152e-05, 0, 0, 0, 0, 0.0008176622, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -8.301411e-05, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0.007076292, 0, 0.00761475, -0.0001125187, 0.001411524, 0, 
    0.00307385, 0.004403167, 0.01805509, -3.343229e-05, 7.842499e-05, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0.000189598, -9.121188e-05, 0, 0, 0, -2.516755e-05, 0.003809891, 
    0.0026288, 5.408653e-05, 0.0003433039, -3.527563e-05, 0.01325701, 
    0.0007514787, 0.007784039, -4.976762e-05, 0.0006382718, 0, 0, 0, 0, 0, 
    -3.0432e-05, 0.006041469, 0.0003964189, 0, -4.422442e-05, -1.614611e-05, 0,
  4.550006e-05, 0, -2.052753e-06, 0, 0, 0, 0, 0.0003168219, -4.258727e-05, 
    0.00716552, 0.04759589, 0.02872662, 0.01394618, 0.002034001, 0.003607468, 
    0.004855298, -0.0002958344, -0.0004048032, 0.002854814, 0.000411052, 
    0.005889871, 0.01646629, 0.0005007592, 0, 0.001253966, 0.0004082255, 
    0.01419196, 0.01805273, 0.005745899,
  0, 0, 0, 0, 0, 5.007793e-05, 0.01828089, 0.002580869, 5.608329e-05, 
    0.01628827, 0.01242172, 0.05052364, -7.712339e-06, 0, 0, 0, 0, 0, 0, 0, 
    0, 7.739874e-05, 0.01949499, -7.951252e-07, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, -0.0003680171, 0.008842622, 1.959636e-05, 0.00550442, 
    0.02216046, 1.407528e-05, 0, 0, 0.002178964, -3.934198e-05, 0, 0, 0, 0, 
    0, 0, 0, 0.001175315, 0, 0, 0, 0,
  0, 7.926953e-06, -1.225131e-06, 0, 0, 0, 0, 0, 0, 0, 0.0007842796, 
    2.135213e-05, 0.01021238, 0.002965884, 0.003157244, 0, 0, -3.429538e-06, 
    0, 0, 0, -1.944377e-05, 0.01148874, -0.0001002081, 0.000596045, 
    0.0001550104, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -5.581887e-05, 0, 0, 0, 0, 0, 0, 
    -1.644622e-05, 0.004052139, -4.122944e-05, 0.00297813, 0.000272387, 0, 
    -8.983155e-07, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -5.628969e-05, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001044392, 0, 
    0, -2.087003e-05, 0, 0, -1.460748e-05, 0, 0,
  0, 0, 0, 0.0007389534, 0.00348642, 0, -8.595177e-06, 0, 0, 0, 0, 0, 0, 0, 
    0, -6.204338e-06, 0, 0, 0.0005595066, 0.0002048152, 0, 0.001400252, 0, 
    0.0002967578, 0, 8.449581e-05, 0.0005014488, -2.601777e-06, 0,
  0, 0, 0, 0.0006271726, -1.540007e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.01030338, 0.006930005, 0.006394145, 0.0009504541, 0.002426731, 
    0.007055821, 0.004278251, -1.013659e-06, 0, 0, 0, 0.00165942, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0004592294, 0, 0.0001216661, 0, 
    -1.496276e-05, 8.007001e-05, 0, 0, 0, 0.0009289061, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0.01845479, -1.743932e-06, 0.0180289, 8.528664e-05, 
    0.007145399, 0, 0.01148937, 0.009512443, 0.03303483, 0.0004657477, 
    0.0008474598, -3.050296e-06, 0, 0, 0, 0, 0, -2.661367e-05, 0, 0, 0, 0, 0, 
    0, 0,
  0, 0.0001526179, -0.0002148919, 0, 0, 0, -7.248153e-05, 0.01350547, 
    0.003453615, 0.0006208774, 0.001250421, 0.0004165127, 0.03142405, 
    0.008817073, 0.01643229, -9.68601e-05, 0.002444418, -4.481463e-05, 0, 0, 
    4.580924e-05, 0, -7.481487e-05, 0.008223942, 0.001982359, -6.654036e-05, 
    9.629826e-05, 6.273651e-06, -2.374157e-06,
  0.0003081421, -1.254348e-05, -1.447996e-05, 0, 0, -1.338759e-07, 
    0.000152749, 0.001292781, 0.001864904, 0.02320247, 0.05361378, 
    0.06874087, 0.02649796, 0.003925373, 0.004601125, 0.0105444, 0.001601049, 
    0.002587719, 0.01094272, 0.0006039268, 0.01432973, 0.02563039, 
    0.004208031, 0, 0.003898913, 0.00304004, 0.0197973, 0.04306175, 
    0.008407968,
  0, 0, 0, 0, 0, 5.752529e-05, 0.02691546, 0.0102929, 0.00172879, 0.02326381, 
    0.02439347, 0.08780923, 6.043378e-05, 0, 0, 0, 0, 5.138766e-05, 
    0.000199154, 0, 0, 0.00017358, 0.04577704, 0.0005865178, 0, 
    -0.0001841351, -3.903129e-05, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0.0006734097, 0.01453507, 0.005786767, 0.01863952, 
    0.0504946, 1.831283e-06, 0, 0, 0.004023158, 0.0007580776, 0, 
    -3.09637e-06, 0, 0, 0.000259113, -0.000109891, 5.479153e-05, 0.001796678, 
    0, 0, 0, 0,
  -5.75362e-06, 0.001677203, 0.001493719, 0, 0, 0, 0, 0, -1.437184e-05, 
    -8.605529e-05, 0.003002356, 0.00220553, 0.0310705, 0.01722093, 
    0.006260362, 0.004375538, 0, -3.970893e-05, -5.501452e-09, 0, 0, 
    0.0004250941, 0.02243042, 0.007771041, 0.007222893, 0.002088355, 
    -1.315156e-07, -4.082406e-05, 0,
  0, 0, 0, 0, 0, -2.336981e-06, 0, -6.673404e-05, 0, -8.131301e-05, 0, 0, 0, 
    0.00141632, 0, 0, 0, 0, 0, 0, 2.709559e-05, 0.005346594, -0.0001113727, 
    0.006362559, 0.005137847, -8.684088e-06, 0.0004391221, 0.002082202, 0,
  0, 0, 0, -3.300115e-06, 0, 0, 0, 0, 0.0002876816, 0, 0, 0, 0.0007041529, 0, 
    0, 0, 0, 0, 0, 0, -0.0001154909, 0.0001353169, 0, -2.952466e-06, 0, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0004655422, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0.003306726, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2.873056e-05, 0, 
    0.000229267, -2.207311e-05, 0.002491246, 0, 0, 0.0003547674, 0, 0, 
    0.002948097, 0, 0,
  -8.311529e-08, 0, 0, 0.002491426, 0.007231226, -6.873665e-07, 0.00119557, 
    -7.883244e-08, 0, 0, 0, 0, 0, -1.264014e-06, -1.955157e-05, 0.0001966108, 
    5.686746e-05, 8.450326e-05, 0.005310684, 0.004891541, 0, 0.005272687, 
    -4.400329e-05, 0.006179622, 0, 0.0006298061, 0.001662098, -0.0001095988, 0,
  0, 0, 0.0003335686, 0.003167137, -2.350045e-05, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0002723906, 0.01341528, 0.01646138, 0.02154008, 0.005990866, 
    0.02609224, 0.01279805, 0.01190436, -0.0001325414, 0, 0, 0, 0.002588714, 
    -1.991174e-05, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, -3.808932e-06, 0, 0, 0, 0, 0.003492509, 0.00190578, 
    0.002908823, 0.001536379, -0.0002214118, 0.0005592275, 0, 0, 0, 
    0.0004705814, 8.500442e-05, 0, 0, 0, -1.345812e-09, 0,
  0, 1.671202e-08, 0, 0, 0.02780971, -0.0001533986, 0.02234088, 0.002452637, 
    0.0294284, -1.1002e-06, 0.02704689, 0.01576709, 0.06417029, 0.003888267, 
    0.007691212, 0.001383819, -1.849331e-08, 0, 6.932972e-06, 0, 
    -1.542326e-10, 1.491972e-07, -5.144674e-10, -1.295332e-05, -7.735281e-11, 
    0, -2.054949e-11, -6.297374e-10, -3.745728e-09,
  -7.880596e-06, 0.006161877, 0.000801077, -1.390492e-05, 0, -4.44652e-11, 
    0.0003569188, 0.02444117, 0.01312495, 0.01558463, 0.009119751, 0.0109641, 
    0.08829448, 0.03033643, 0.0346685, 0.0005179937, 0.009389621, 
    -0.0002955483, -1.035799e-06, -8.391953e-10, 0.002231243, 0, 0.002628182, 
    0.02086635, 0.01031699, 0.0003624342, 0.0001789286, 0.005622553, 
    0.0002176627,
  0.004167182, 8.152666e-07, 1.785766e-05, 0, 2.066849e-07, 0.0004458389, 
    0.00515473, 0.01525603, 0.01540318, 0.07738879, 0.07603515, 0.1367999, 
    0.06289208, 0.009433031, 0.008193972, 0.02671742, 0.005351183, 
    0.02020069, 0.02548925, 0.001484983, 0.0253873, 0.04384217, 0.03583186, 
    0.0002251897, 0.00824379, 0.004836475, 0.02467627, 0.06955654, 0.01530837,
  -1.12825e-06, 0, 0, 0, -4.7264e-07, 0.001060474, 0.03306356, 0.04315197, 
    0.009848157, 0.03658715, 0.05024693, 0.1095185, 0.002813095, 
    0.0005217324, 0, -4.492783e-06, 0, 0.003715494, 0.004290683, 0, 0, 
    0.009765498, 0.0677853, 0.001114806, -6.000449e-07, 3.317881e-05, 
    -0.0001255269, 0, 0,
  0, 0, 0, 0, 0, -3.257054e-06, -2.467433e-08, 0.004929751, 0.02348801, 
    0.02158666, 0.03969984, 0.06941526, 0.006757203, -5.239583e-05, 
    -2.538102e-06, 0.005461655, 0.002228589, 0.002989724, -6.561504e-05, 0, 
    0, 0.001611872, 0.001263319, 0.003282374, 0.006903736, 0.0007948261, 
    -1.813002e-05, 0, 0,
  -2.301448e-05, 0.007822327, 0.00354265, 0, 0.0006278346, 6.427071e-05, 
    -1.422367e-06, 0, -2.748068e-05, -6.149743e-05, 0.01224002, 0.01477802, 
    0.05343124, 0.03902749, 0.01452115, 0.005804234, 0.0001606958, 
    0.0001898704, 0.0009391427, 0, 0, 0.00361976, 0.03109472, 0.01515671, 
    0.01350334, 0.008592879, 0.001071624, -6.936724e-05, -1.012657e-05,
  -9.26171e-06, -3.587456e-06, 0.001427652, 0, 0, 0.0007291539, -3.08718e-06, 
    -0.0001793988, 0.0002529089, 0.002563156, 0, -1.439928e-07, 
    -6.374122e-05, 0.002685849, 0, -1.669689e-05, -1.036835e-05, 
    -4.111727e-06, 0.001357712, -3.020362e-05, 0.0002547562, 0.007098265, 
    -0.0002443546, 0.01377166, 0.007567353, 0.002869935, 0.01186497, 
    0.004936536, -4.499734e-06,
  0, -7.495282e-06, 0.0001901835, -6.600484e-06, 0, 0, 0, 0, 0.0009155409, 0, 
    0, 0, 0.002510151, 0.0001360113, 0, 0, 0, 0, 0, -1.221832e-05, 
    0.001975713, 0.003885111, -0.0001548387, -1.050076e-05, 0.003770415, 0, 
    -1.027451e-09, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0.003646244, 0, 0, -8.311287e-07, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0002319962, -1.410054e-05, 0, 
    0, -1.462305e-05, 0.002710464, 0.0009877353, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, -8.606718e-06, 0, 0.004059621, 0, 0.0003657958, 0.002992582, 
    0.0005339844, 0.0007471695, 0, 0, -4.439396e-07, 0, 0, 0, 0.0002113712, 
    0, 0.002000639, 0.001425605, 0.004809568, 0, 0.00244278, 0.00201385, 
    -5.057193e-06, 0, 0.00802965, -0.000112029, 0,
  0.0001268675, 0, -3.9926e-06, 0.003344445, 0.01818217, 0.002260836, 
    0.004980458, 0.001662015, 0.0004263667, 2.010066e-11, 0, 0, 0, 
    0.0002027989, 0.00173379, 0.007690436, 0.004903803, 0.01157608, 
    0.01906249, 0.0220357, -2.686466e-05, 0.0143123, 0.001953177, 0.01435665, 
    0.0002981797, 0.003333827, 0.005073978, -0.000125755, -0.0001250809,
  -1.007044e-05, 0, 0.002594604, 0.009376679, -5.923293e-05, -1.859296e-08, 
    -2.861445e-07, 0, 0, 2.98131e-13, 0, -2.946892e-10, 0, 0.0152595, 
    0.02414079, 0.03055121, 0.03914637, 0.01232054, 0.06180831, 0.02808391, 
    0.01585011, 0.0007262874, -1.267012e-07, -1.285511e-07, 0, 0.008345398, 
    0.002103656, -2.726671e-05, -2.602151e-06,
  -1.350591e-09, 0.0003105788, -2.749045e-09, -1.047956e-09, 3.783191e-08, 0, 
    -1.02133e-05, -2.527359e-07, 1.208541e-05, 4.295448e-06, 6.07043e-07, 
    2.044047e-05, 3.076272e-05, 0.008500069, 0.005653163, 0.006662788, 
    0.006837499, -0.0005811537, 0.001930666, -1.7664e-06, 4.416022e-05, 
    -1.536358e-10, 0.0001209179, 0.0009202119, -1.679511e-06, 0, 
    -2.638599e-07, 8.362126e-05, 4.099259e-06,
  0, 1.727331e-05, 0, 0, 0.03926986, 0.002897125, 0.02823302, 0.06915738, 
    0.07968928, 0.0112695, 0.05108818, 0.06832206, 0.1343165, 0.09563308, 
    0.07126717, 0.03323503, 9.178724e-05, -1.924556e-07, 0.008708041, 
    -1.312581e-09, 7.780257e-06, 0.0002993601, 3.793886e-06, 0.002899015, 
    7.816028e-06, 3.884363e-07, 2.756913e-05, 1.479837e-05, 0.0001673562,
  7.70719e-05, 0.01783071, 0.003721381, -2.761473e-05, -3.259599e-05, 
    3.529586e-05, 0.005886411, 0.09880507, 0.05848976, 0.1039483, 0.1778741, 
    0.1892514, 0.3039606, 0.1353647, 0.1555918, 0.08619868, 0.02493398, 
    0.01400549, -1.33983e-05, 9.250546e-05, 0.01550048, 0.0002766717, 
    0.006309839, 0.06032217, 0.0320931, 0.004019174, 0.004040398, 0.03645924, 
    0.01985088,
  0.02371247, 0.005360571, 0.0007364705, -1.151101e-10, -0.0001597704, 
    0.0432931, 0.129024, 0.4277212, 0.4489015, 0.4343813, 0.3750301, 
    0.4019556, 0.3309522, 0.1603617, 0.05291226, 0.104191, 0.07615776, 
    0.06542128, 0.0489361, 0.00940434, 0.04136391, 0.1738704, 0.116255, 
    0.007822154, 0.01551882, 0.006274417, 0.03029992, 0.1487696, 0.045639,
  0.007988797, 0.0002714226, 2.428997e-06, 9.425109e-06, 0.003126353, 
    0.0180767, 0.08317282, 0.2624839, 0.1592309, 0.1169856, 0.2279714, 
    0.2061689, 0.08595649, 0.002442335, 9.394413e-05, 0.003482752, 
    2.847654e-05, 0.008337314, 0.01318232, 0.003671058, 0.0006555862, 
    0.02740134, 0.1175281, 0.004137074, 0.0008178672, 1.711418e-05, 
    -0.0001738268, 0.0003737571, -5.732654e-06,
  0.0007036509, 0.0001407474, 0, -3.138101e-07, 0, -5.224168e-05, 
    8.362073e-05, 0.008599445, 0.05245634, 0.1642812, 0.2308708, 0.2096885, 
    0.1120415, 0.03354474, 0.02652091, 0.02109093, 0.01759507, 0.008788356, 
    0.0007583909, -3.664909e-06, 0, 0.006153514, 0.03933158, 0.01226858, 
    0.01799607, 0.001204595, -0.0002083645, -1.338525e-05, -1.357578e-05,
  -3.452172e-05, 0.01979165, 0.005598112, 0.0001915681, 0.001924436, 
    0.002255924, -1.307169e-06, 0.000173413, 0.006690509, 0.001337408, 
    0.03998613, 0.06660461, 0.1876878, 0.09142508, 0.04355847, 0.02664186, 
    0.01035535, 0.00611462, 0.002714289, -7.944697e-05, 0, 0.005520075, 
    0.03934349, 0.02160859, 0.02393853, 0.02290258, 0.009128776, 
    -0.0001608233, -1.977678e-05,
  0.0005100632, -1.485969e-05, 0.00346215, 0, 0.0004229026, 0.00226481, 
    -0.0001032784, 0.001534507, 0.002097183, 0.006268782, -8.321743e-05, 
    -0.0001286625, 0.0003790341, 0.004471493, 0, 0.001400417, 0.002587883, 
    0.0009788587, 0.004370776, 0.0002372212, 0.007259897, 0.01252455, 
    0.001498483, 0.02130367, 0.008900745, 0.007921005, 0.03204516, 
    0.01546975, 0.0009030799,
  0, 0.002522465, 0.000338312, -2.01915e-05, 0, 0, 1.121127e-06, 0, 
    0.003299381, 0, 0, 0, 0.007220337, 0.001653813, 0, 0, 0.0007268559, 0, 0, 
    -6.084397e-05, 0.009388013, 0.008821693, 0.003929709, -3.13837e-05, 
    0.009897556, -3.95099e-10, -1.643947e-07, 3.469045e-08, -5.350966e-05,
  0, 0, 0, 0, 0, 0, -9.991852e-05, 0.004990603, 0.0001155892, 0, 
    -2.493386e-06, 0, 0, 0, 0, 0, 0, 0, 0, -8.848617e-06, -0.0003754172, 0, 
    0, 0, -3.66024e-06, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0.0002795945, 0, -2.667997e-08, 0, 0, 0.0001834745, 0, 0, 0, 
    0.0004147484, -5.894385e-05, -1.47323e-05, 0, 4.763341e-05, 0.006687426, 
    0.004641651, -3.743762e-05, 0.003516025, -1.795479e-05, 0, 0, 0, 0, 0,
  0, 0.0001115948, -4.13048e-05, -6.1057e-05, 0.005750044, 0, 0.00285358, 
    0.00380232, 0.003676056, 0.004491576, 0.0005630788, 0.000821643, 
    0.0001688857, 0.0006453948, 0.001186606, -5.827006e-05, 0.002216577, 
    0.0003255367, 0.007026977, 0.008975322, 0.007291569, 0.0008236423, 
    0.002388209, 0.005810417, 0.002738518, -6.868705e-05, 0.01730627, 
    0.001309694, 0,
  0.003192643, -0.0003284833, 0.001132612, 0.007413718, 0.02917264, 
    0.006627543, 0.01045096, 0.00574086, 0.004529074, 0.003141974, 
    0.002745022, 0.0006936654, -9.290058e-09, 0.003292526, 0.005489669, 
    0.01856651, 0.01912914, 0.0288251, 0.04215703, 0.0499184, 0.000745651, 
    0.02798558, 0.006290454, 0.02810931, 0.002057939, 0.009425252, 0.0182837, 
    0.0007606498, -0.0003630342,
  0.001458738, 3.552041e-05, 0.004782102, 0.01398467, 0.0004710435, 
    3.865855e-06, -3.278337e-06, 2.463745e-07, -5.401146e-10, 7.844505e-08, 
    3.504554e-07, 3.931636e-07, 1.598046e-07, 0.02543429, 0.03995889, 
    0.05114678, 0.06241038, 0.04291485, 0.1111514, 0.04285365, 0.02114374, 
    0.007729148, 0.0005112113, 0.0009848877, -4.622404e-06, 0.01526347, 
    0.006035028, 0.001179296, 0.005360926,
  0.01261535, 0.002527426, 6.583404e-05, 4.222573e-06, 0.01311191, 
    -0.0001274245, 0.0007923369, -6.308665e-06, -7.458623e-05, 4.396948e-06, 
    4.054695e-07, 7.567754e-06, 1.097727e-05, 0.006229006, 0.02683442, 
    0.04924607, 0.05492585, 0.01788799, 0.03541589, 0.01431727, 0.00171325, 
    7.337755e-06, 0.001183019, 0.004634729, 0.0007440309, 0.0001967874, 
    0.00935286, 0.0009473572, 0.007238322,
  0.001778876, 0.02903, 0.0006385816, 1.007835e-05, 0.07837338, 0.01404612, 
    0.04253325, 0.099601, 0.1036259, 0.004995839, 0.05448538, 0.02701424, 
    0.1186839, 0.07152793, 0.06384861, 0.03290778, 0.003202963, 2.136407e-05, 
    0.02488583, 6.738117e-06, 0.003638608, 0.01436943, 0.0003327884, 
    0.01895235, 0.005706029, 0.0002581017, -6.43176e-05, 0.00957856, 
    0.001619405,
  0.1124661, 0.2513872, 0.2031709, 0.006022041, 0.003304288, 0.03035262, 
    0.1520016, 0.2266472, 0.2565554, 0.4220275, 0.1324892, 0.1579778, 
    0.258105, 0.1114823, 0.126428, 0.04056511, 0.03332976, 0.008629813, 
    7.319717e-06, 4.271385e-05, 0.03870854, 0.00842353, 0.03288149, 
    0.2195572, 0.1080273, 0.04701969, 0.01997223, 0.1176637, 0.1135592,
  0.1865723, 0.1607441, 0.03255184, -2.005835e-06, 0.003006937, 0.1492747, 
    0.1544644, 0.2660594, 0.4068738, 0.300649, 0.3160917, 0.3455839, 0.24922, 
    0.1236099, 0.06314897, 0.1482056, 0.1204807, 0.09229843, 0.08833383, 
    0.01840123, 0.04688742, 0.1632261, 0.268838, 0.08648795, 0.130812, 
    0.0614203, 0.05426033, 0.2261109, 0.2449062,
  0.1347319, 0.006302192, 0.03622152, 0.0001136837, 0.0009521452, 0.01409845, 
    0.08933333, 0.2123475, 0.1082282, 0.0862454, 0.1782006, 0.1711199, 
    0.07629193, 0.0388419, 0.03126312, 0.03653573, 0.009882182, 0.05731938, 
    0.05595719, 0.04532211, 0.002692441, 0.02574701, 0.1722128, 0.2688262, 
    0.09372582, 0.04258615, 0.00919363, 0.03289813, 0.03615063,
  0.01152193, 0.008755733, 0.0001344481, 0.001075652, -5.793123e-05, 
    -1.570429e-05, 0.0002404983, 0.01306743, 0.09906485, 0.1631598, 
    0.3198007, 0.2931187, 0.1988079, 0.1118244, 0.1014896, 0.1324486, 
    0.1385123, 0.05788939, 0.009665049, 0.002864029, -6.043341e-06, 
    0.05121817, 0.176423, 0.1528855, 0.2538772, 0.07671203, 0.003442692, 
    0.00124484, 0.005446648,
  -0.0001632987, 0.05065509, 0.008194869, 0.0001634111, 0.00840139, 
    0.0155189, 0.0004244352, 0.01206439, 0.04605771, 0.004329067, 0.08859683, 
    0.1554267, 0.2724166, 0.1924316, 0.1047851, 0.1260452, 0.1158231, 
    0.07110292, 0.024873, 2.493857e-05, 0.0002588832, 0.008387648, 0.109886, 
    0.05029994, 0.09086069, 0.06829064, 0.03202061, 0.001164199, 0.009517534,
  0.008404773, -6.082006e-05, 0.007275877, -1.10077e-09, 0.0009033771, 
    0.01033481, 0.007074214, 0.004431176, 0.009583702, 0.01391629, 
    0.0005080146, -0.0002642794, 0.003108689, 0.006174814, 0, 0.009393672, 
    0.01250546, 0.04549697, 0.02320373, 0.005151114, 0.02164252, 0.01807951, 
    0.005760388, 0.0263056, 0.0141186, 0.02279107, 0.04899869, 0.03914062, 
    0.02730179,
  1.156587e-05, 0.007969112, 0.004222514, -3.519888e-06, 0, 0, 0.000277463, 
    -5.733477e-07, 0.00409674, -3.943431e-05, -0.0001243784, 0, 0.009404178, 
    0.012288, -2.22203e-05, 0, 0.008964146, 0.0005776116, -7.202905e-05, 
    -0.0001116241, 0.01577451, 0.02047526, 0.007549897, -7.397924e-06, 
    0.01437306, -0.0001037167, 0.0001860301, 0.00567941, 0.0006670949,
  0, 0, 0, 0, 0.002806202, 0, -0.0001454438, 0.007069902, 0.0004275531, 0, 
    0.0004027745, 0, 0, 0, 0, 0, 0.001354775, -2.728105e-05, -2.752629e-06, 
    -4.045519e-05, -0.0004096055, 0, 0, 0, -1.388874e-05, 0.002599014, 0, 
    -1.63527e-05, 3.304146e-06,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -4.173786e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  5.585922e-06, 0, 0, 0, -3.164709e-05, 0.00111933, 0, -1.679368e-05, 
    -9.505521e-05, 0, 0.001884347, 0, 0, -3.570389e-05, 0.001207453, 
    -0.0001191811, 0.002215589, 0, 0.006650737, 0.01334159, 0.01674071, 
    0.008160221, 0.01117061, 0.004997587, 0.0008204951, -3.293133e-05, 0, 0, 0,
  0.001090162, 0.002583069, -4.663257e-05, 0.001378924, 0.01005216, 
    0.001817578, 0.006201194, 0.01066023, 0.01348369, 0.007009314, 
    0.001926356, 0.004948545, 0.004402287, 0.004499108, 0.004040239, 
    0.001301499, 0.01473282, 0.006153876, 0.01937327, 0.02650147, 0.01561362, 
    0.007739463, 0.005420377, 0.007633456, 0.00739293, 0.0007720565, 
    0.02708147, 0.03320373, 0,
  0.00713819, 0.003816654, 0.01043836, 0.02884046, 0.0444847, 0.01298233, 
    0.01634289, 0.02050806, 0.02482372, 0.01577558, 0.006504463, 0.002805443, 
    0.0003892227, 0.02000504, 0.02543343, 0.04149762, 0.02522455, 0.06003674, 
    0.07741646, 0.08580403, 0.01378267, 0.04697545, 0.01946471, 0.05819624, 
    0.006807279, 0.0254298, 0.02765883, 0.007516561, 0.0008816092,
  0.004165291, 0.0003803971, 0.006855312, 0.02721501, 0.009734013, 
    0.01216926, 0.002793737, 9.85514e-06, 4.905499e-05, -4.409362e-09, 
    7.62343e-06, -1.276579e-05, 1.275578e-07, 0.04373617, 0.08334447, 
    0.07800769, 0.09844715, 0.1414711, 0.2542757, 0.1679303, 0.06104694, 
    0.03225234, 0.03860569, 0.06249827, 0.02687944, 0.02294851, 0.01920931, 
    0.005356831, 0.008223495,
  0.0003210188, 5.402767e-05, 6.605525e-05, 2.355124e-06, 0.004308084, 
    -5.205745e-06, 3.482718e-05, 3.52615e-07, -5.512039e-05, 4.032015e-06, 
    1.111324e-07, 7.243916e-06, 8.449789e-06, 0.004848994, 0.02158724, 
    0.04244395, 0.06315165, 0.01594744, 0.08172289, 0.003858181, 
    0.0009137249, -2.226544e-05, 7.620381e-05, 0.0002156619, 0.003375341, 
    0.0003885199, 0.009161881, 3.941304e-05, 0.01194411,
  4.711609e-05, 0.000231625, 2.955837e-05, -1.454893e-06, 0.06252214, 
    0.01645605, 0.03874629, 0.08191212, 0.09269944, 0.001441462, 0.04698718, 
    0.02541631, 0.1068574, 0.05871693, 0.05414484, 0.02359247, 0.00140958, 
    3.955079e-05, 0.005820162, 1.263108e-06, 6.154341e-05, 0.006442201, 
    1.191856e-05, 0.01114619, 0.003656379, 0.00015857, -8.742417e-05, 
    0.0001322933, 0.0001073751,
  0.05508732, 0.2171304, 0.09801549, 0.00147503, 0.001192807, 0.00352326, 
    0.08049212, 0.1416742, 0.2112348, 0.3757579, 0.08023857, 0.1509528, 
    0.2382869, 0.08665477, 0.08634286, 0.02033727, 0.03620288, 0.006848254, 
    1.673772e-05, 7.089343e-06, 0.01636562, 0.003560589, 0.04555893, 
    0.2004044, 0.08998013, 0.02381945, 0.01599853, 0.07091075, 0.03567579,
  0.1535998, 0.1347221, 0.03147807, 0.0002206068, 0.0002331985, 0.08881874, 
    0.1128748, 0.1138394, 0.3656142, 0.2401424, 0.2572434, 0.3124488, 
    0.1928592, 0.07530041, 0.03561659, 0.1005854, 0.07531873, 0.05374024, 
    0.06558467, 0.01544352, 0.03891911, 0.1185336, 0.2423316, 0.06018569, 
    0.07979411, 0.05187455, 0.04505609, 0.1973335, 0.1874998,
  0.1867823, 0.04023645, 0.03833032, 2.081376e-06, 0.001467778, 0.01445258, 
    0.08729549, 0.1890947, 0.0970052, 0.07124856, 0.149335, 0.1580272, 
    0.04936637, 0.03468849, 0.02349327, 0.02502978, 0.04600221, 0.06052507, 
    0.05839339, 0.01657508, 0.0005435912, 0.01712215, 0.1538723, 0.2107979, 
    0.07519013, 0.01423542, 0.007567896, 0.02918735, 0.02693769,
  0.0534234, 0.08798701, 0.003405528, 0.0223567, 0.005256125, 0.002955638, 
    0.0003984298, 0.0201372, 0.1829583, 0.1330055, 0.3104797, 0.2977666, 
    0.1718352, 0.09939157, 0.1176331, 0.1361569, 0.146048, 0.05487221, 
    0.02952123, 0.02197792, 0.007908795, 0.06056353, 0.1335402, 0.1368731, 
    0.2226786, 0.1042968, 0.05674905, 0.009485697, 0.01564952,
  0.04877281, 0.113817, 0.03586112, 0.01483481, 0.0810818, 0.04740452, 
    0.005498201, 0.1552805, 0.1602226, 0.06482735, 0.1296923, 0.1461966, 
    0.3185436, 0.2282164, 0.1346799, 0.215809, 0.2233015, 0.1202036, 
    0.03200528, 0.007176835, 0.00225154, 0.08325379, 0.1080885, 0.07734852, 
    0.2118671, 0.1689848, 0.1173649, 0.04419922, 0.03870511,
  0.03193186, 0.0006721822, 0.01800821, 0.01052403, 0.02944314, 0.01529745, 
    0.01624521, 0.01471592, 0.02397533, 0.0841514, 0.02298126, 0.02953862, 
    0.03218133, 0.03921898, 0.005937476, 0.04851395, 0.07511339, 0.1305901, 
    0.05527492, 0.008979613, 0.02803721, 0.06080648, 0.03432134, 0.04560985, 
    0.06475039, 0.09654479, 0.1117482, 0.1245728, 0.1211061,
  0.006808089, 0.01400334, 0.008702205, -8.735355e-05, 0, 0, 0.005434705, 
    0.0007162537, 0.01038203, -0.0006883137, 0.002042068, -6.356389e-05, 
    0.01528217, 0.02610905, 0.001549236, 0.001345391, 0.04930956, 0.02680088, 
    0.001123864, 0.001643674, 0.03889616, 0.04647384, 0.04128889, 
    0.008646294, 0.01825869, 0.01420472, 0.009460329, 0.03073982, 0.04321992,
  0.0116828, 0.005421649, -4.228627e-06, 3.000434e-05, 0.007615615, 
    -8.256254e-06, 0.001374022, 0.009142007, 0.009120179, 0.003400906, 
    0.0007796742, -2.258175e-09, 1.223194e-05, 0, -3.411124e-07, 
    -2.557788e-06, 0.001375952, 0.02895365, 0.0279832, 0.01642744, 
    0.005852164, -0.0001619994, -8.103561e-05, -3.945686e-05, 2.8617e-05, 
    0.006445555, -1.296565e-06, 0.003332028, 0.01523172,
  -1.059159e-06, -1.514682e-05, 0, 0, 0, 0, 0, 0, 1.375985e-06, 
    -6.142727e-08, 0, -0.0001038772, -3.711751e-05, 0, 0, 6.540414e-06, 
    -6.122973e-06, -3.759442e-10, 0, 0, 7.25051e-09, 3.722413e-05, 0, 0, 0, 
    0, 0, -4.449004e-07, 3.713919e-08,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0.0001010102, 0, 0, 0, 0, 
    -1.963856e-09, 0, 0, 0, 0, 0.00196883, 0.0001834175, 0, 0, 0,
  0.0005702862, 0, 0, -5.291303e-06, -0.0001469931, 0.004376149, 
    -5.448341e-05, -6.088347e-05, -0.0001232959, 0, 0.001919715, 
    -7.267933e-05, -5.854398e-05, -0.000198036, 0.001880201, 0.001277146, 
    0.003616772, 7.779839e-05, 0.02289932, 0.02874309, 0.03187939, 
    0.02550706, 0.02819538, 0.01048723, 0.006990252, 0.001505208, 
    -9.224346e-05, 0.001158877, -8.575911e-05,
  0.005105713, 0.005299082, 0.001795175, 0.004295308, 0.0155296, 0.005269021, 
    0.01502566, 0.02098628, 0.02398873, 0.01979295, 0.006943903, 0.01631348, 
    0.02579478, 0.008110752, 0.008005415, 0.01227594, 0.0409036, 0.04801129, 
    0.05262018, 0.05164524, 0.04829074, 0.02820298, 0.02046502, 0.01579622, 
    0.02675467, 0.02383765, 0.05619503, 0.04813835, 0.002033486,
  0.02070891, 0.02533884, 0.02274549, 0.05257604, 0.06940988, 0.04835572, 
    0.04005709, 0.04265602, 0.06022395, 0.02445492, 0.02241264, 0.01393606, 
    0.004677495, 0.04334556, 0.05329204, 0.04611797, 0.05035037, 0.1111582, 
    0.1457044, 0.1748762, 0.1168069, 0.1172823, 0.06640799, 0.09299095, 
    0.1128521, 0.0732116, 0.07387308, 0.04173462, 0.02260854,
  0.03116034, 0.02527418, 0.01206646, 0.06463557, 0.04321214, 0.02697225, 
    0.01874109, 0.001252906, 0.001163942, 2.186816e-06, 0.003679851, 
    0.005530681, 0.0001142524, 0.05214552, 0.08219355, 0.1022178, 0.1648361, 
    0.1821026, 0.2686297, 0.1898797, 0.06701037, 0.06248323, 0.0428532, 
    0.1001407, 0.02273969, 0.06579577, 0.07868039, 0.06602608, 0.04276326,
  0.0002659604, 1.286684e-05, 0.0002731511, 4.752737e-07, 0.002073525, 
    0.001439423, -5.350135e-07, 2.365071e-06, 0.001764453, 3.133991e-06, 
    1.956705e-07, 1.431371e-05, 1.066345e-05, 0.01023819, 0.02372156, 
    0.04255555, 0.05236753, 0.01866657, 0.03195838, 9.987386e-05, 
    0.0006216975, 9.859136e-06, 4.146355e-06, 2.282577e-05, 0.0004759828, 
    2.968894e-05, 0.01711707, 0.003082587, 0.006866595,
  8.91287e-06, 3.677374e-05, 4.560035e-06, -8.83561e-06, 0.06175059, 
    0.01613028, 0.03576933, 0.06405163, 0.0964166, 0.001781238, 0.04728505, 
    0.03161227, 0.09990326, 0.04613588, 0.04504101, 0.01240025, 0.001799384, 
    4.596966e-05, 5.061868e-05, 7.304207e-08, 1.260047e-06, 4.646738e-05, 
    2.489562e-06, 0.005180851, 3.198013e-05, 5.159843e-05, 2.206007e-05, 
    1.344034e-05, 1.115318e-05,
  0.003613262, 0.1688314, 0.06326327, 0.0006249225, 0.0009610148, 0.00324396, 
    0.0553815, 0.122435, 0.1498565, 0.3307719, 0.061318, 0.1447774, 
    0.2171735, 0.08356362, 0.07388956, 0.01766145, 0.03731701, 0.008242866, 
    1.278805e-05, 9.801627e-06, 0.001287734, 0.0001155781, 0.05367384, 
    0.1415421, 0.06912445, 0.03172967, 0.01880214, 0.0435334, 0.01121533,
  0.1410467, 0.1252946, 0.03542663, -1.020321e-05, 0.0003163698, 0.03674381, 
    0.1012308, 0.06090477, 0.3074912, 0.1954914, 0.2093679, 0.2853579, 
    0.1558798, 0.05258585, 0.03504252, 0.07689587, 0.07199673, 0.03936225, 
    0.06033323, 0.0153831, 0.03513868, 0.1045195, 0.2145784, 0.04730208, 
    0.04875429, 0.03062692, 0.04034062, 0.1706337, 0.1672856,
  0.1956194, 0.05131172, 0.01733596, 2.419146e-05, 0.0004389782, 0.01463306, 
    0.0751988, 0.1861509, 0.08776584, 0.05908133, 0.1150949, 0.1478674, 
    0.03806698, 0.03020168, 0.01735202, 0.02270111, 0.02765036, 0.05710853, 
    0.04648694, 0.001729787, 0.0009237331, 0.01488508, 0.1477403, 0.1815865, 
    0.06740642, 0.003072611, 0.006323232, 0.0224834, 0.0154037,
  0.05212808, 0.08345407, 0.005000169, 0.0202286, 0.004120252, 0.01100073, 
    0.0006220093, 0.0639039, 0.2131152, 0.1106849, 0.2776284, 0.2657566, 
    0.1438961, 0.1087603, 0.1069436, 0.1131998, 0.1018371, 0.04521319, 
    0.03554311, 0.01950961, 0.05868451, 0.0413017, 0.09346204, 0.1147389, 
    0.1888384, 0.08590227, 0.03262119, 0.01996002, 0.01804884,
  0.1207644, 0.141478, 0.03292191, 0.0686403, 0.09609757, 0.05585174, 
    0.01748108, 0.2390161, 0.20047, 0.1425226, 0.1670991, 0.153459, 
    0.3053602, 0.2166035, 0.1106807, 0.2174617, 0.2273129, 0.1046012, 
    0.04334619, 0.02594302, 0.02654338, 0.06931613, 0.09880972, 0.08430801, 
    0.1668696, 0.1525306, 0.1349081, 0.06808694, 0.05574324,
  0.0914187, 0.08512373, 0.1443436, 0.07249753, 0.1077102, 0.1474885, 
    0.0822707, 0.03455779, 0.0848271, 0.1031819, 0.07396543, 0.0965937, 
    0.08576056, 0.08817408, 0.05851953, 0.1166453, 0.2107812, 0.1761187, 
    0.08320061, 0.02721334, 0.1360904, 0.1092655, 0.04509394, 0.06457735, 
    0.1137321, 0.1679939, 0.1592354, 0.1861184, 0.1695845,
  0.09065729, 0.08380876, 0.04506212, 0.05760759, 0.03409013, 0.03316386, 
    0.01531421, 0.07785847, 0.1133285, 0.04966457, 0.05227342, 0.02751161, 
    0.02481207, 0.1120933, 0.05739237, 0.07718838, 0.09913691, 0.07761333, 
    0.007681048, 0.08768038, 0.1272604, 0.1338566, 0.06168557, 0.02060321, 
    0.04893809, 0.03625971, 0.07192253, 0.145029, 0.1015179,
  0.110156, 0.09429009, 0.02872244, 0.02542799, 0.0520897, 0.03170058, 
    0.042892, 0.02710725, 0.07507803, 0.1051072, 0.03322476, 0.04250097, 
    0.02234645, 0.005414866, 0.03075393, 0.04244049, 0.05797301, 0.07646892, 
    0.04290553, 0.0624379, 0.03856834, 0.01893791, 0.007658255, -0.002984221, 
    0.0188463, 0.007738243, -3.818655e-05, 0.02752936, 0.05663665,
  0.02293015, 0.0310355, 0.01709228, 0.009827565, -0.0003190814, 
    -4.704822e-08, 1.185579e-10, -6.543919e-08, -0.001157478, 0.01215752, 
    0.02039496, 0.01882636, 0.0177852, 0.01407803, 0.01050365, 0.007667587, 
    0.0003414606, 0.0001494706, 9.638455e-05, -2.68045e-05, -1.935371e-05, 
    0.001169959, -1.177087e-05, -7.554088e-05, -4.242311e-05, -9.518614e-06, 
    -6.590797e-05, 0.005344666, 0.02096691,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0.005388514, 0.0002488404, 0, 0, 0, 0, 0.002103017, 0, 0, 0, 0, 0, 0, 
    1.167411e-05, 0.000752598, 0.001170566, 9.275444e-06, 0.0009925318, 
    0.004227137, 0.002019051, -0.0001219569, 0.003842399, -9.37087e-06, 
    0.004396854, 0.005343024, 0.004990905, 0.0005616367, 0, 0.0006865768,
  0.02248277, -0.0001449998, 9.112467e-07, 0.001105004, 0.001318394, 
    0.008684347, 0.001863178, 0.00662608, 0.003412616, 0.003265121, 
    0.01017259, 0.004590739, -0.0002005629, -0.0001522605, 0.03207861, 
    0.02571432, 0.007914051, 0.006509601, 0.05363286, 0.06078199, 0.0590885, 
    0.05534103, 0.0401612, 0.0360558, 0.04150859, 0.0235865, 0.009423789, 
    0.009121227, 0.01723322,
  0.03827124, 0.0363978, 0.01218193, 0.01979865, 0.02686875, 0.04540601, 
    0.04266614, 0.06024761, 0.05839815, 0.05681862, 0.03790884, 0.04251191, 
    0.04822895, 0.04591141, 0.07643618, 0.04170986, 0.1205778, 0.09531246, 
    0.09905157, 0.09643802, 0.1071931, 0.06812572, 0.05465187, 0.03624966, 
    0.09533216, 0.1022974, 0.1018512, 0.1269511, 0.0387112,
  0.1170949, 0.08596438, 0.07164593, 0.1290322, 0.1549994, 0.1020418, 
    0.09001268, 0.08557171, 0.117172, 0.06183061, 0.07371951, 0.0487677, 
    0.06025419, 0.1389481, 0.1160019, 0.06964955, 0.10731, 0.1517341, 
    0.1515959, 0.1579878, 0.1422027, 0.1380089, 0.145827, 0.1430318, 
    0.1108026, 0.1269619, 0.1248474, 0.1138805, 0.08556783,
  0.04429546, 0.02610399, 0.02413592, 0.06017282, 0.02277103, 0.0209221, 
    0.02180912, 0.004466805, 0.01373236, -6.136495e-05, 0.02112426, 
    0.01259282, 0.000694968, 0.0409577, 0.09695577, 0.1311706, 0.1714392, 
    0.1668855, 0.2327481, 0.1821701, 0.04168354, 0.05611822, 0.02055697, 
    0.03973785, 0.009404534, 0.05141922, 0.07088378, 0.06034341, 0.03776304,
  -2.001875e-06, -3.433189e-05, 0.004517664, -8.207935e-08, 0.002683976, 
    0.009420238, -7.363131e-09, -3.287006e-06, 0.01454381, 2.177178e-06, 
    2.052684e-07, 0.003361879, -2.918272e-05, 0.0320315, 0.04093784, 
    0.03347398, 0.04475975, 0.0305537, 0.02594256, 3.334578e-06, 
    0.0001949455, 5.315185e-08, 1.546046e-07, 1.913255e-06, 0.0006071291, 
    2.555406e-05, 0.01601452, 0.02451531, 0.002064645,
  5.64259e-06, 9.661668e-06, 5.033808e-06, -2.349478e-06, 0.06625206, 
    0.01830733, 0.03193018, 0.03419355, 0.09073602, 0.001535852, 0.04358364, 
    0.03326977, 0.1070891, 0.03900094, 0.04934941, 0.003080955, 0.001095474, 
    1.243494e-05, 1.183358e-06, 4.370827e-08, 1.481213e-09, 9.094551e-07, 
    8.897355e-07, 0.0005235513, 5.906546e-06, 0.0001201138, 2.397933e-06, 
    2.639751e-05, 2.801681e-06,
  0.0001398373, 0.1280483, 0.0435853, 0.000511152, 0.0006485221, 0.005081995, 
    0.03391267, 0.09868635, 0.1157749, 0.2659983, 0.04552074, 0.1152369, 
    0.1887523, 0.0731564, 0.07285137, 0.008783528, 0.05306963, 0.00737845, 
    1.920323e-06, 8.587963e-07, 3.228322e-05, 7.819944e-05, 0.01563347, 
    0.1026032, 0.05782706, 0.04735063, 0.03610703, 0.031722, 0.003947945,
  0.1301944, 0.1311487, 0.05027713, -4.316795e-05, 0.000484449, 0.01911366, 
    0.09800222, 0.03610542, 0.2559764, 0.1615977, 0.1836552, 0.23822, 
    0.1276551, 0.04985793, 0.0367799, 0.04367221, 0.05798201, 0.02435212, 
    0.06021452, 0.01445616, 0.03154073, 0.08943323, 0.1537128, 0.02784364, 
    0.0308429, 0.01300288, 0.03790675, 0.1591958, 0.1310029,
  0.1653605, 0.03068193, 0.00849915, 4.76786e-05, -5.426307e-06, 0.01980789, 
    0.0781764, 0.1767607, 0.08111952, 0.05397526, 0.1135852, 0.1362303, 
    0.0283864, 0.007621321, 0.01612099, 0.01586895, 0.01258712, 0.02430423, 
    0.03676165, -0.0001994247, 3.897309e-05, 0.009636416, 0.1376213, 
    0.1477778, 0.05136167, 0.006766179, 0.004572568, 0.02536759, 0.014915,
  0.04464709, 0.07829782, 0.005228157, 0.01254721, 0.001008403, 0.01158338, 
    0.002956115, 0.05654716, 0.2122349, 0.09679643, 0.2559979, 0.2545353, 
    0.1300048, 0.1108187, 0.07195496, 0.09544575, 0.08204481, 0.03288116, 
    0.01906627, 0.006141816, 0.04066907, 0.02975885, 0.06409837, 0.09640109, 
    0.1642962, 0.07240252, 0.01384593, 0.03000163, 0.007047029,
  0.1111546, 0.1305049, 0.02915934, 0.06647557, 0.08186548, 0.04643962, 
    0.06118192, 0.2115333, 0.2008708, 0.1307712, 0.1849085, 0.1388498, 
    0.2840937, 0.1978831, 0.1129922, 0.2211158, 0.2151292, 0.08618169, 
    0.03992809, 0.05953864, 0.1103186, 0.05183524, 0.07987897, 0.07683636, 
    0.1344312, 0.145059, 0.1168221, 0.03860321, 0.03857159,
  0.1195464, 0.1418768, 0.1205949, 0.06749682, 0.1111806, 0.13886, 0.0959348, 
    0.07485953, 0.1571509, 0.151423, 0.1307475, 0.1505436, 0.1406198, 
    0.1343497, 0.1342742, 0.2039454, 0.2173072, 0.1827638, 0.09274361, 
    0.06263059, 0.2018702, 0.08673429, 0.05380984, 0.06726892, 0.1314507, 
    0.1750577, 0.1655456, 0.1665144, 0.1429294,
  0.09934576, 0.08626897, 0.09915577, 0.09029377, 0.0608298, 0.06394267, 
    0.1268165, 0.1492592, 0.1450362, 0.0547285, 0.1153568, 0.1625325, 
    0.09855264, 0.1462802, 0.1370998, 0.1500751, 0.1546952, 0.1412072, 
    0.05152118, 0.1036285, 0.1164604, 0.1506837, 0.1116452, 0.07149374, 
    0.1207265, 0.09080957, 0.1599695, 0.1953361, 0.1291697,
  0.1802821, 0.1356646, 0.07324011, 0.08971793, 0.1633156, 0.1721652, 
    0.08835426, 0.1144653, 0.1537761, 0.1414635, 0.1208499, 0.06825762, 
    0.1340683, 0.04480627, 0.0735518, 0.09311931, 0.09919631, 0.1136047, 
    0.1523193, 0.130958, 0.1037576, 0.1002553, 0.0649868, 0.003429664, 
    0.1282872, 0.01156378, 0.003009788, 0.0862187, 0.1212607,
  0.05082738, 0.07193404, 0.07463422, 0.03415451, 0.02118286, 0.04076299, 
    0.03447947, 0.03553987, 0.03779233, 0.0318686, 0.08012123, 0.09143098, 
    0.08578645, 0.07018009, 0.0685948, 0.08851517, 0.1018392, 0.06155612, 
    0.02812288, 0.006727522, 0.006057789, 0.01444374, 0.02746189, 0.02059255, 
    0.009341117, 0.0001835599, -0.0008002076, 0.028948, 0.05240503,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6.289879e-07, -4.357969e-06, 0, 
    -0.0003264332, 0.004044815, 0, 0, 0, 0, 0, -5.798911e-06, 0, 0, 0, 0, 0,
  0.01726402, 0.01077286, 0.003993069, 0, 0, -0.0001657698, 0.01005685, 
    -0.0001421575, 0, 0, -8.253001e-07, -1.865015e-05, -0.0001401213, 
    0.001457015, 0.00654018, 0.009018349, 0.0001946873, 0.004583432, 
    0.007729654, 0.009634611, 0.009916767, 0.0183055, 0.001075574, 
    0.01652222, 0.007943446, 0.008978295, 0.01190633, 0.0131385, 0.006959607,
  0.07276206, 0.04504716, 0.0171495, 0.02446983, 0.00748271, 0.0234285, 
    0.04845848, 0.03688049, 0.06271301, 0.02786165, 0.02222792, 0.02573574, 
    0.019156, 0.0635942, 0.05604484, 0.1176194, 0.1089913, 0.07688005, 
    0.1346827, 0.1606949, 0.09256069, 0.07282727, 0.06936137, 0.07452166, 
    0.1146919, 0.1102002, 0.06177497, 0.05057508, 0.0858698,
  0.09336307, 0.06252874, 0.09776555, 0.09266417, 0.1294846, 0.1170883, 
    0.09522319, 0.1129563, 0.115805, 0.125304, 0.09755582, 0.1262223, 
    0.1153075, 0.2151976, 0.2352136, 0.1630112, 0.192398, 0.1762701, 
    0.1776754, 0.1359952, 0.1449292, 0.09205897, 0.07693392, 0.1018843, 
    0.09889869, 0.1487865, 0.1985341, 0.1851237, 0.06115406,
  0.1494593, 0.1292961, 0.1447746, 0.1746213, 0.1518051, 0.1090722, 
    0.1004415, 0.1043346, 0.1305549, 0.06732123, 0.08495, 0.1009346, 
    0.1242351, 0.216119, 0.1578282, 0.1470549, 0.1484295, 0.1732259, 
    0.1568175, 0.153104, 0.1157178, 0.1504529, 0.1363177, 0.1866804, 
    0.08959077, 0.1185587, 0.1389922, 0.1113152, 0.1054665,
  0.04725476, 0.01893144, 0.05368345, 0.05165236, 0.01981341, 0.01029482, 
    0.00190946, 0.006109336, 0.01729944, 0.001791984, 0.01983033, 0.0111492, 
    0.009151041, 0.03560375, 0.1138485, 0.1510658, 0.1338696, 0.1646902, 
    0.2144831, 0.1627511, 0.04119868, 0.04505031, 0.01066401, 0.02025758, 
    0.005219522, 0.04375952, 0.05450024, 0.0429821, 0.02914346,
  1.532516e-06, -2.625837e-05, 0.004070447, -1.332764e-07, 0.0134092, 
    0.002908082, -1.145148e-06, -0.0001993753, 0.006210504, -1.569815e-06, 
    3.240342e-07, 0.01303648, 0.0006668377, 0.08353554, 0.05067652, 
    0.04206459, 0.03374479, 0.0319417, 0.01879624, 2.305362e-06, 
    0.0001545742, -1.325699e-06, -2.90195e-09, 1.178315e-07, 0.0005238167, 
    8.761723e-06, 0.0134407, 0.03343872, 0.008607888,
  3.663146e-06, 1.507676e-06, 3.744279e-06, -2.785384e-06, 0.07334751, 
    0.01343384, 0.03016534, 0.007815816, 0.07992367, 0.002151356, 0.03653736, 
    0.03567406, 0.1109153, 0.0296144, 0.05106064, 0.00110621, 0.00158554, 
    4.452086e-06, 3.99549e-07, -1.01292e-10, -2.022525e-11, 2.982281e-08, 
    2.784818e-08, 2.217131e-05, 3.24275e-06, 0.000842512, 9.174573e-06, 
    0.0006709904, 9.800896e-07,
  1.518648e-05, 0.09957745, 0.043519, 0.0003600424, 0.0006573495, 
    0.006589895, 0.01921005, 0.07538942, 0.07955442, 0.1692796, 0.02740284, 
    0.06874997, 0.1424911, 0.05851865, 0.05589544, 0.008193331, 0.05939447, 
    0.005546535, 4.246284e-05, -1.755302e-06, 3.441955e-06, 0.004111288, 
    0.01012445, 0.08442352, 0.05539828, 0.0573098, 0.0483976, 0.0312262, 
    0.001559648,
  0.1021329, 0.11659, 0.1080398, 2.139345e-05, 0.0003322782, 0.01130566, 
    0.07521401, 0.02243015, 0.171426, 0.1478416, 0.144399, 0.1984572, 
    0.1055235, 0.04227094, 0.0330357, 0.02245675, 0.04605824, 0.0115958, 
    0.06247137, 0.01004079, 0.03615106, 0.07855155, 0.113123, 0.02271913, 
    0.02098304, 0.008675148, 0.04143557, 0.1527096, 0.1160645,
  0.1104583, 0.02545858, 0.003514652, 6.493189e-05, 1.13358e-06, 0.03181823, 
    0.07575327, 0.1526701, 0.06205827, 0.05188193, 0.1046614, 0.128645, 
    0.01992358, 0.005162753, 0.01056144, 0.0118713, 0.007775359, 0.008337217, 
    0.02159839, -0.0001211767, 4.374429e-05, 0.006948126, 0.1104234, 
    0.1059882, 0.03405406, 0.003888487, 0.00217859, 0.03510627, 0.01389072,
  0.01938283, 0.07551389, 0.004210456, 0.007827437, -0.0003005904, 
    0.009039194, 0.005454896, 0.0500811, 0.2148717, 0.08367137, 0.2373733, 
    0.2387921, 0.1061725, 0.1115284, 0.05512203, 0.09410576, 0.08453125, 
    0.03066062, 0.0110232, 0.000763429, 0.01732798, 0.02129536, 0.04458164, 
    0.071252, 0.1353116, 0.06536678, 0.004655551, 0.02828453, 0.0162905,
  0.08630525, 0.1192331, 0.02029041, 0.03766385, 0.07702439, 0.04145366, 
    0.1205477, 0.1818574, 0.1862535, 0.09926024, 0.1842964, 0.1283143, 
    0.2469002, 0.1886471, 0.1145586, 0.218349, 0.2162746, 0.07564326, 
    0.03909971, 0.06890144, 0.09737378, 0.04457414, 0.07074047, 0.06758383, 
    0.1139976, 0.1474793, 0.1083183, 0.03257237, 0.04777849,
  0.1176058, 0.114772, 0.1086889, 0.05917657, 0.08316603, 0.1102584, 
    0.1255112, 0.1314184, 0.1821919, 0.1517264, 0.139969, 0.1638128, 
    0.1528715, 0.1264449, 0.1281029, 0.2186465, 0.2203749, 0.1622338, 
    0.09574706, 0.07905411, 0.1898912, 0.07711881, 0.07117262, 0.06820371, 
    0.1294935, 0.1789131, 0.1560327, 0.1539387, 0.1216144,
  0.1432797, 0.1048629, 0.08657116, 0.08173802, 0.09349514, 0.1244434, 
    0.144252, 0.1691291, 0.1596456, 0.08612484, 0.122838, 0.2263499, 
    0.1393593, 0.1594022, 0.1317938, 0.1966315, 0.2066885, 0.1696203, 
    0.1247019, 0.1035211, 0.1100675, 0.163613, 0.1513151, 0.154685, 
    0.2002162, 0.1987353, 0.1862402, 0.2013431, 0.1289548,
  0.1743895, 0.1552931, 0.1048978, 0.100396, 0.1706312, 0.244067, 0.1601985, 
    0.1531993, 0.1763761, 0.1428219, 0.1116545, 0.1055932, 0.1366087, 
    0.05785318, 0.09654429, 0.1061624, 0.1202388, 0.1441754, 0.1515233, 
    0.1840575, 0.1114577, 0.1367204, 0.1343068, 0.03922496, 0.1780875, 
    0.05676551, 0.003334317, 0.1368977, 0.1519116,
  0.1181915, 0.122466, 0.1543382, 0.09316704, 0.09162482, 0.133267, 
    0.1262863, 0.1215396, 0.1135339, 0.09046081, 0.1006395, 0.1085885, 
    0.1217828, 0.1388438, 0.1528066, 0.1474564, 0.129863, 0.08927795, 
    0.1479221, 0.1001492, 0.04214706, 0.0402927, 0.04068027, 0.03641704, 
    0.08835989, 0.01380112, 0.02025139, 0.03583, 0.1043887,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9.89617e-07, 0.0006688809, 
    0.0002178159, 0.005537611, 0.007712838, 0, 0, 0, 0, 0, -1.957309e-05, 
    -2.594771e-05, 0, 0, 0, 0,
  0.03265325, 0.02305072, 0.01473975, 0.00209473, 0.0001919719, -0.000546851, 
    0.01752098, 0.0003863471, -0.0004520747, 0, 9.419947e-05, 0.000482185, 
    -0.001223893, 0.03491586, 0.04382594, 0.0410308, 0.03765881, 0.05776461, 
    0.05659393, 0.1121629, 0.03483898, 0.0445908, 0.01938761, 0.02997401, 
    0.08151399, 0.03924094, 0.05711116, 0.03845429, 0.03446017,
  0.1230473, 0.08046714, 0.08020885, 0.08688661, 0.06048223, 0.08219781, 
    0.1195162, 0.1122162, 0.1477682, 0.1191108, 0.1218814, 0.179657, 
    0.1190766, 0.1856908, 0.141366, 0.1939979, 0.2090704, 0.1644571, 
    0.2115343, 0.2246255, 0.1736124, 0.1274466, 0.158146, 0.0994854, 
    0.1844105, 0.1492076, 0.1287311, 0.1340003, 0.1386853,
  0.1038503, 0.08416809, 0.1071772, 0.1358248, 0.1343166, 0.1471753, 
    0.1404796, 0.1749351, 0.1566925, 0.1884167, 0.1499192, 0.1878973, 
    0.1862691, 0.3124834, 0.3127536, 0.1583218, 0.1924594, 0.1815189, 
    0.1972732, 0.1937763, 0.2085466, 0.1192342, 0.1052101, 0.1237043, 
    0.1424175, 0.1653443, 0.2223846, 0.198708, 0.08317311,
  0.1389208, 0.1131772, 0.1431314, 0.1681735, 0.1540536, 0.1036653, 0.101569, 
    0.09396535, 0.1385159, 0.07994322, 0.09333206, 0.140133, 0.1710508, 
    0.2275472, 0.1800874, 0.1495578, 0.1609639, 0.1994257, 0.1672917, 
    0.1461485, 0.106871, 0.158191, 0.1455335, 0.1871753, 0.07339177, 
    0.1140741, 0.1240097, 0.1095178, 0.1140767,
  0.05479776, 0.008186881, 0.04880594, 0.05200053, 0.009171079, 0.005693211, 
    -1.48471e-05, 0.009137046, 0.03884361, 0.005169945, 0.02266892, 
    0.01478934, 0.008427816, 0.03692138, 0.08717353, 0.1300841, 0.1366871, 
    0.1624103, 0.2063912, 0.1628996, 0.04001037, 0.02902312, 0.01344943, 
    0.01602997, 0.006749763, 0.04112561, 0.04102063, 0.04227941, 0.04071533,
  1.537432e-07, 1.033212e-06, 0.001336377, 5.51363e-08, 0.01214608, 
    0.0004718606, -8.255738e-08, 0.000814671, 0.008493805, -3.298227e-06, 
    9.79555e-07, 0.01123235, 0.003875415, 0.08673631, 0.05812938, 0.02515918, 
    0.0242532, 0.03131001, 0.01830396, 4.469928e-06, 6.200603e-05, 
    -1.454645e-06, 0, -1.914386e-09, 0.0004760234, 1.981821e-05, 0.009888906, 
    0.01910519, 0.002702449,
  8.170811e-07, 7.265312e-06, 2.234368e-06, 0.0001190829, 0.08328246, 
    0.01063074, 0.02700814, 0.00767895, 0.0727711, 0.01078015, 0.02969374, 
    0.03226768, 0.1218043, 0.02213674, 0.05795875, 0.0008930884, 0.002187331, 
    7.35519e-05, 8.513607e-08, 0, 0, -9.180219e-10, 5.044859e-08, 
    4.261843e-05, 1.334845e-05, 3.112803e-05, 0.00148743, -0.0001278321, 
    2.816039e-07,
  5.955661e-06, 0.05434646, 0.0424373, 0.000298269, 0.00118527, 0.007963737, 
    0.01479796, 0.07908534, 0.0493889, 0.08945429, 0.02128018, 0.04225498, 
    0.1239216, 0.05287082, 0.04689218, 0.008343407, 0.05951089, 0.004389771, 
    0.0001033513, 0.0007644967, 2.091347e-06, 0.0003770281, 0.006660142, 
    0.08601578, 0.06038091, 0.07627276, 0.07261517, 0.02233644, 0.004764516,
  0.06768543, 0.1032056, 0.1027529, -5.225424e-06, 0.000361029, 0.01032937, 
    0.0539716, 0.01522837, 0.1059936, 0.1215195, 0.1311612, 0.1809467, 
    0.08748922, 0.03060493, 0.03572446, 0.01760604, 0.0449253, 0.005650936, 
    0.06158622, 0.01233154, 0.03499916, 0.06501421, 0.09335653, 0.02018784, 
    0.01901574, 0.01016652, 0.06032397, 0.1420245, 0.09000009,
  0.06040797, 0.02282269, 0.0007371376, 0.0001352441, 3.364119e-05, 
    0.0381461, 0.06148217, 0.1250201, 0.0581774, 0.05990728, 0.122204, 
    0.1231288, 0.01653869, 0.003994081, 0.006346705, 0.02292225, 0.004341504, 
    0.004678908, 0.0008923461, -1.175571e-05, 2.942809e-05, 0.003552543, 
    0.08875847, 0.0766061, 0.01711345, 0.001884511, 0.007761141, 0.04852508, 
    0.01305773,
  0.0206748, 0.0831006, 0.004049034, 0.009736115, -2.702442e-05, 0.006165416, 
    0.006047847, 0.05678421, 0.2298606, 0.07704266, 0.2338956, 0.1981591, 
    0.09346376, 0.1078579, 0.04048507, 0.08188416, 0.07966527, 0.0314407, 
    0.01230926, 3.155805e-06, 0.003134937, 0.01334629, 0.039961, 0.04962397, 
    0.1077121, 0.05505684, 0.001878311, 0.01946004, 0.01949618,
  0.07507586, 0.1191533, 0.01662689, 0.02860693, 0.07271937, 0.03814518, 
    0.1855926, 0.1396652, 0.152426, 0.08135052, 0.1740658, 0.1141594, 
    0.2211575, 0.1788502, 0.09303761, 0.1978666, 0.2070313, 0.06706901, 
    0.04124301, 0.08342231, 0.08199587, 0.03859449, 0.06154136, 0.06281642, 
    0.09698633, 0.1328351, 0.0725863, 0.03685692, 0.02166598,
  0.1242376, 0.1072345, 0.09558179, 0.05536986, 0.06443883, 0.1014022, 
    0.1206305, 0.1138257, 0.1809138, 0.1308801, 0.1525285, 0.1621171, 
    0.1430809, 0.1094554, 0.1000052, 0.2210329, 0.2154507, 0.1627377, 
    0.09411395, 0.09025525, 0.1722005, 0.07698023, 0.07230848, 0.08567259, 
    0.119971, 0.1700972, 0.1579402, 0.1312001, 0.1268492,
  0.1013439, 0.09778086, 0.07695506, 0.07306209, 0.09583418, 0.1819122, 
    0.1524701, 0.1673295, 0.1673434, 0.09007006, 0.1112147, 0.2151327, 
    0.1365451, 0.1404495, 0.1176463, 0.1905246, 0.2047835, 0.1658198, 
    0.09507193, 0.1254442, 0.09552471, 0.1554895, 0.1596481, 0.1957586, 
    0.222701, 0.2159199, 0.1683725, 0.1932295, 0.1341368,
  0.1431782, 0.1390222, 0.11189, 0.09699637, 0.1535895, 0.252477, 0.1609482, 
    0.1496296, 0.1769052, 0.1297823, 0.1006366, 0.09886374, 0.1353364, 
    0.06566183, 0.1201767, 0.1049579, 0.1045764, 0.1264072, 0.1457181, 
    0.1844562, 0.137053, 0.1348565, 0.1248082, 0.08423202, 0.1986729, 
    0.1135242, 0.01215973, 0.1508628, 0.154904,
  0.1685846, 0.228993, 0.2045937, 0.1440876, 0.1572973, 0.2028664, 0.1812755, 
    0.1678766, 0.1516099, 0.1333979, 0.1296436, 0.1422186, 0.1688765, 
    0.1926692, 0.2390325, 0.2218377, 0.182975, 0.1306929, 0.1605162, 
    0.1218705, 0.08868479, 0.1070938, 0.0657304, 0.02904691, 0.08209497, 
    0.06006841, 0.04728036, 0.07154329, 0.1474669,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.003445406, 0.01152084, 0.01486833, 
    0.02531631, 0.01090618, -2.71336e-05, -8.301684e-07, 0, 0, 3.314715e-05, 
    0.02570331, 0.0402228, 0.01339843, 0.02633776, -0.0002422029, 0,
  0.06307335, 0.05470717, 0.03282851, 0.01600177, 0.001496966, 0.004129547, 
    0.04954462, 0.004859745, 0.000186363, -0.0007887905, 0.001702263, 
    0.001469454, 0.02335962, 0.1251536, 0.1389396, 0.1297342, 0.121968, 
    0.1201599, 0.1102684, 0.1631336, 0.09753048, 0.05760276, 0.04504439, 
    0.09715532, 0.1735824, 0.1522968, 0.1763895, 0.2025269, 0.128539,
  0.1634897, 0.1271808, 0.1495266, 0.1323431, 0.1538881, 0.1541451, 
    0.1431375, 0.1671295, 0.2143217, 0.2153378, 0.2267479, 0.2731135, 
    0.223498, 0.2004726, 0.2480952, 0.2464154, 0.2254744, 0.1522332, 
    0.1988806, 0.2492645, 0.1869007, 0.1542403, 0.2459028, 0.1570037, 
    0.2455688, 0.2067017, 0.135283, 0.1656038, 0.1685588,
  0.102926, 0.1077578, 0.1213183, 0.1263205, 0.1329408, 0.1364675, 0.1640854, 
    0.185533, 0.1783732, 0.1987226, 0.161383, 0.1972164, 0.1906848, 
    0.2753345, 0.2428143, 0.09087137, 0.18683, 0.1641552, 0.1929149, 
    0.1937836, 0.2092336, 0.127819, 0.1231362, 0.1246689, 0.1209791, 
    0.1830323, 0.2182572, 0.1897978, 0.08643208,
  0.105095, 0.09680094, 0.1189782, 0.147498, 0.1501439, 0.1019792, 0.1133425, 
    0.1106923, 0.1376719, 0.09859382, 0.1012731, 0.1337823, 0.1491992, 
    0.2043847, 0.1691208, 0.1481665, 0.146393, 0.1840583, 0.1842541, 
    0.1465949, 0.07593814, 0.1591225, 0.1463675, 0.1864179, 0.05883927, 
    0.09820704, 0.1122761, 0.1078029, 0.09497833,
  0.07212247, 0.004689645, 0.03821319, 0.0504353, 0.007892065, 0.005825111, 
    0.002821545, 0.01842432, 0.0493245, 0.005329497, 0.02343545, 0.01987445, 
    0.005042377, 0.03705664, 0.07044744, 0.1125649, 0.1304169, 0.1637669, 
    0.1839756, 0.1478964, 0.03948437, 0.02897457, 0.01794443, 0.01226067, 
    0.003673272, 0.04112634, 0.03771627, 0.03924182, 0.06159989,
  -1.211619e-06, -2.346331e-06, 0.0009823695, 1.868699e-06, 0.01070153, 
    3.347444e-06, -1.588089e-06, 0.001456625, 0.0004321164, 1.129343e-07, 
    6.712132e-07, 0.003250655, 3.843631e-05, 0.085443, 0.05325003, 
    0.02050901, 0.02333678, 0.03513693, 0.01950868, 2.333562e-06, 
    2.170761e-05, 3.008296e-07, -5.718196e-11, 2.442737e-08, 0.00041002, 
    2.246126e-05, 0.00404167, 0.0002319638, 0.0003999395,
  2.186998e-07, 1.649271e-05, 8.189805e-07, 0.0002629876, 0.08732209, 
    0.008894245, 0.02411218, 0.006288819, 0.0611183, 0.01049437, 0.04084556, 
    0.01712101, 0.1396988, 0.02092072, 0.06675714, 0.001754022, 0.001919883, 
    5.662355e-05, 5.17543e-08, 0, 0, -1.754566e-10, 1.275622e-08, 
    2.32224e-05, 2.408182e-05, 9.582068e-05, 0.006272912, -1.131682e-06, 
    9.317653e-09,
  0.0001580172, 0.04629065, 0.04217182, 0.0002627879, 0.002812684, 
    0.007853647, 0.01590165, 0.08483747, 0.04205919, 0.03733449, 0.02250143, 
    0.03798279, 0.1209527, 0.05301608, 0.04731795, 0.008771989, 0.05695407, 
    0.003781212, 0.001361872, 0.0118541, 5.311804e-05, 0.0006746154, 
    0.005816199, 0.08866249, 0.06899658, 0.08532245, 0.1049336, 0.02978269, 
    0.008992235,
  0.03974836, 0.08042535, 0.1086524, 0.0004148274, 0.0006706182, 0.01540725, 
    0.05037033, 0.01699091, 0.0720347, 0.1084516, 0.1151093, 0.1662779, 
    0.08044446, 0.03314339, 0.04069193, 0.01891773, 0.05268009, 0.005847769, 
    0.08023921, 0.01364208, 0.02981816, 0.05607039, 0.07744558, 0.01913261, 
    0.01995472, 0.01306255, 0.04356891, 0.1244959, 0.07145063,
  0.03876619, 0.02701203, -0.0001443569, 0.001240958, 0.0008080635, 
    0.03548919, 0.06154298, 0.09104367, 0.06545308, 0.06567711, 0.1154837, 
    0.1142293, 0.01494066, 0.003748264, 0.005383128, 0.01752948, 0.003562109, 
    0.001325198, 2.413583e-06, 0.0005589232, 6.608437e-05, 0.001522926, 
    0.0703909, 0.05611722, 0.009990524, 0.008274484, 0.04370496, 0.03436989, 
    0.01821163,
  0.01755371, 0.08749969, 0.005748892, 0.0166854, 5.053848e-05, 0.005165936, 
    0.01641026, 0.06155277, 0.2435665, 0.07255507, 0.2503539, 0.1751398, 
    0.09773764, 0.08323117, 0.01958614, 0.07520707, 0.08769362, 0.0345563, 
    0.01291893, -3.244232e-07, 4.163786e-05, 0.009679676, 0.04195091, 
    0.03901079, 0.09544179, 0.05202177, 0.0001646596, 0.001025689, 0.02261055,
  0.06266475, 0.1220756, 0.0166289, 0.02828708, 0.07411244, 0.02933541, 
    0.1799031, 0.09541364, 0.1076965, 0.07163323, 0.1644857, 0.1062625, 
    0.1964841, 0.176132, 0.08084362, 0.1908491, 0.1816813, 0.07498323, 
    0.04341405, 0.0712781, 0.07084673, 0.03802813, 0.059202, 0.05098128, 
    0.09373804, 0.1346051, 0.06767394, 0.04255469, 0.01332173,
  0.1283166, 0.1061642, 0.08274888, 0.05335901, 0.04943317, 0.08763976, 
    0.1235846, 0.1049864, 0.1781069, 0.1191607, 0.1516736, 0.165168, 
    0.1309211, 0.09715256, 0.07720036, 0.2238028, 0.1979362, 0.1631621, 
    0.08876404, 0.0922128, 0.1707629, 0.08356547, 0.08336242, 0.089138, 
    0.1177964, 0.1758484, 0.1623425, 0.1434862, 0.1207866,
  0.1022433, 0.0964143, 0.07239337, 0.06698503, 0.0986561, 0.1924282, 
    0.1483846, 0.1640467, 0.1636086, 0.08159561, 0.1010627, 0.1884425, 
    0.1373553, 0.1323441, 0.1071846, 0.1849858, 0.1944143, 0.1513983, 
    0.09146177, 0.1170212, 0.07647005, 0.1416229, 0.1689426, 0.2180748, 
    0.2116209, 0.228194, 0.1693003, 0.1855343, 0.1188195,
  0.1239211, 0.1265769, 0.1033261, 0.08627187, 0.1397936, 0.2474108, 
    0.1637749, 0.1332802, 0.1650872, 0.1261531, 0.0877359, 0.1169711, 
    0.1368093, 0.06971627, 0.1205892, 0.09983151, 0.09623728, 0.1071597, 
    0.1334972, 0.1721123, 0.1431869, 0.1273527, 0.1316503, 0.09577135, 
    0.1830388, 0.2136936, 0.03463434, 0.1460475, 0.1622424,
  0.1560806, 0.2120504, 0.1856259, 0.1398025, 0.1515471, 0.2047984, 0.180501, 
    0.1745825, 0.1626266, 0.1318872, 0.1196825, 0.1253574, 0.1581398, 
    0.2028466, 0.2703778, 0.2377025, 0.1912772, 0.1366148, 0.1732086, 
    0.1789415, 0.1768474, 0.1995494, 0.1792131, 0.1193561, 0.1431041, 
    0.06596934, 0.07032181, 0.08349146, 0.1421452,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0001671758, 0.02492593, 0.09135735, 
    0.06887701, 0.05747962, 0.04244315, 0.002951661, 8.962218e-05, 
    -1.804367e-05, 0, 0.01156646, 0.2560562, 0.1342958, 0.08777021, 
    0.05960077, -0.00309674, 0,
  0.1437827, 0.1536002, 0.1429747, 0.09062621, 0.001948207, 0.01197828, 
    0.107335, 0.02730913, 0.0001839119, -0.0007752349, 0.02621359, 
    0.01747656, 0.08534966, 0.1654278, 0.1787622, 0.1596148, 0.1824628, 
    0.1864706, 0.1571368, 0.1679743, 0.1107425, 0.1362351, 0.1258023, 
    0.1840709, 0.2739132, 0.2264848, 0.3031073, 0.301161, 0.2535596,
  0.1765273, 0.1414867, 0.2178582, 0.1439554, 0.2006861, 0.2103884, 
    0.1745121, 0.1968539, 0.2626295, 0.2583875, 0.2308328, 0.3064802, 
    0.2195976, 0.192977, 0.263146, 0.26188, 0.2304607, 0.1626458, 0.2013047, 
    0.2460877, 0.199867, 0.1727912, 0.2694, 0.1912962, 0.2620801, 0.2255885, 
    0.1848639, 0.2023117, 0.189571,
  0.1165789, 0.1381526, 0.1357328, 0.1284252, 0.1171804, 0.1411372, 
    0.1628663, 0.2049509, 0.203054, 0.2064199, 0.1652521, 0.1834261, 
    0.1812532, 0.2537907, 0.2394749, 0.06233284, 0.170796, 0.1746301, 
    0.1756686, 0.1744549, 0.1901773, 0.1380824, 0.1199408, 0.1148637, 
    0.1147022, 0.1844676, 0.2140228, 0.1817778, 0.09520507,
  0.09159012, 0.08747903, 0.0949962, 0.1401824, 0.1479104, 0.0912681, 
    0.09887242, 0.09891055, 0.132691, 0.1108394, 0.105266, 0.1309993, 
    0.1334127, 0.1936448, 0.1590241, 0.1284074, 0.1488357, 0.1674801, 
    0.1858795, 0.1597762, 0.07836327, 0.1668099, 0.1525833, 0.1856328, 
    0.06484266, 0.09699924, 0.1223711, 0.09654751, 0.08571856,
  0.07525831, 0.004173472, 0.03506882, 0.05907875, 0.007822558, 0.006002573, 
    0.0124433, 0.02234807, 0.05659309, 0.01308804, 0.02262947, 0.02236779, 
    0.002029797, 0.03883952, 0.06038994, 0.09624278, 0.1278776, 0.1541785, 
    0.1768052, 0.1585, 0.03217398, 0.04566637, 0.0194806, 0.01297543, 
    0.0003803228, 0.04279722, 0.03856445, 0.03388087, 0.06715549,
  0.0001078341, 8.291642e-08, 0.001075178, 0.0001694053, 0.01229334, 
    1.282147e-07, 5.379095e-06, 0.001287828, 5.752347e-06, 1.134934e-07, 
    1.650489e-07, 0.01880413, 0.002907342, 0.08820193, 0.05859248, 0.0182512, 
    0.02233673, 0.04046854, 0.02192343, -1.437971e-06, 5.282125e-05, 
    -9.037695e-07, -3.725643e-10, 5.069673e-08, 0.0004033585, 1.197389e-05, 
    3.206742e-06, 4.807843e-06, 1.319379e-06,
  2.228944e-07, 1.174705e-05, 3.40977e-07, 0.0003286582, 0.07683603, 
    0.01229999, 0.02518428, 0.01320208, 0.05278742, 0.01184634, 0.05557876, 
    0.01191313, 0.1509533, 0.01995542, 0.06760675, 0.002921517, 0.001391728, 
    4.820832e-05, 1.22606e-07, 2.739569e-11, -4.794927e-10, 0, 1.614117e-08, 
    4.008227e-05, 0.0002947471, -2.379016e-05, 0.01875011, -1.648062e-07, 
    9.321984e-10,
  0.004015098, 0.04294081, 0.04242057, 0.001868266, 0.003242227, 0.005453278, 
    0.01655757, 0.0643305, 0.04536206, 0.01688122, 0.0273536, 0.03201867, 
    0.1259053, 0.06430364, 0.0461671, 0.009567757, 0.05884716, 0.0007147187, 
    9.501913e-05, 0.01317594, 0.005534403, 8.190041e-06, 0.01345208, 
    0.09869538, 0.08224447, 0.09922421, 0.1150286, 0.01324357, 0.01035818,
  0.02751408, 0.06079526, 0.1111825, 0.01174142, 0.0009335595, 0.02760527, 
    0.03033566, 0.03282674, 0.06248474, 0.1092897, 0.1029145, 0.1581911, 
    0.08452912, 0.03911651, 0.03548939, 0.03538242, 0.0650187, 0.01535378, 
    0.1040542, 0.0215783, 0.02378993, 0.05547267, 0.07842114, 0.01735069, 
    0.01972037, 0.0148473, 0.04221813, 0.1212146, 0.0663733,
  0.08615381, 0.03507679, -0.00038269, 0.0007125382, 0.000798338, 0.0349033, 
    0.06686441, 0.08691248, 0.06180019, 0.06740208, 0.1351959, 0.1104937, 
    0.01687269, 0.004261422, 0.004463256, 0.01265614, 0.005387404, 
    1.326877e-05, 4.937969e-07, 0.02442529, 0.0003364144, 0.003360556, 
    0.05983039, 0.04703315, 0.008166011, 0.009742998, 0.02279209, 0.02931203, 
    0.01617264,
  0.02078304, 0.08019952, 0.003329814, 0.01337696, -0.0002029503, 0.00330763, 
    0.01567461, 0.06522039, 0.2699941, 0.07972437, 0.2693781, 0.1816637, 
    0.09859498, 0.06419592, 0.02055043, 0.07373981, 0.08347196, 0.02602683, 
    0.01368451, -1.218161e-07, -4.927725e-05, 0.008337268, 0.03346348, 
    0.04019025, 0.08398975, 0.04756021, -0.000665533, 1.254711e-05, 0.02879892,
  0.05190236, 0.1149524, 0.01846522, 0.02899841, 0.07213341, 0.02633503, 
    0.1728912, 0.06221366, 0.06578848, 0.06516019, 0.1653076, 0.09747246, 
    0.1811351, 0.1672206, 0.08011902, 0.1836549, 0.1629627, 0.05687159, 
    0.04040557, 0.06441643, 0.0708099, 0.04950614, 0.05914719, 0.04832803, 
    0.09129356, 0.1405343, 0.0757774, 0.02743661, 0.005632896,
  0.1285491, 0.109252, 0.07871286, 0.0512912, 0.04180343, 0.08488467, 
    0.131186, 0.1000105, 0.1758795, 0.1118911, 0.1632689, 0.1653788, 
    0.1208219, 0.1010634, 0.072244, 0.222872, 0.1934454, 0.1606538, 
    0.09566168, 0.08823664, 0.1770172, 0.08690481, 0.07091872, 0.09864462, 
    0.1186345, 0.2009587, 0.1564944, 0.1332207, 0.09105278,
  0.09886844, 0.09267434, 0.07461149, 0.06899145, 0.09168705, 0.2161436, 
    0.1533184, 0.1537815, 0.1575001, 0.07938024, 0.08836061, 0.1609096, 
    0.1361849, 0.1252409, 0.1095618, 0.1795351, 0.2071616, 0.1498868, 
    0.09612952, 0.09755666, 0.0706132, 0.1254864, 0.1743243, 0.2418008, 
    0.1845831, 0.2464274, 0.1602175, 0.1744758, 0.1212238,
  0.1229796, 0.1133599, 0.09509683, 0.08628271, 0.1410875, 0.2485168, 
    0.1690156, 0.1331592, 0.1570919, 0.1292456, 0.0823146, 0.1092962, 
    0.128843, 0.0788365, 0.1105703, 0.08828551, 0.09457747, 0.1027645, 
    0.1354219, 0.1611021, 0.1362527, 0.1343187, 0.1381613, 0.1168573, 
    0.1744609, 0.3510548, 0.07865889, 0.1463467, 0.1629762,
  0.1447208, 0.2071034, 0.2088847, 0.1405278, 0.1492106, 0.2031971, 
    0.1864486, 0.1853665, 0.1687615, 0.1343189, 0.1129372, 0.1124595, 
    0.1385479, 0.1922632, 0.2693063, 0.2395394, 0.1957734, 0.1395045, 
    0.1509604, 0.2046798, 0.1893916, 0.2269899, 0.2374186, 0.1607191, 
    0.1505595, 0.09937992, 0.1180822, 0.09222175, 0.1263481,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001180089, 0.1387099, 0.1261118, 
    0.1184558, 0.1535679, 0.11859, 0.03684128, 0.01801114, 0.002305011, 
    -2.080873e-06, 0.04951349, 0.3410966, 0.2339803, 0.1842272, 0.1481351, 
    0.03950402, 0,
  0.2001397, 0.2133516, 0.2097097, 0.1649234, 0.004860216, 0.04869833, 
    0.1453346, 0.05143245, 0.0451904, 0.01348285, 0.04211139, 0.03197166, 
    0.144653, 0.177297, 0.2106174, 0.2084023, 0.169562, 0.2017178, 0.1772134, 
    0.2334344, 0.1736716, 0.1986589, 0.1819674, 0.3096199, 0.3398849, 
    0.290286, 0.3420925, 0.3708526, 0.3361712,
  0.1782124, 0.1750817, 0.2478146, 0.2055396, 0.2562045, 0.273686, 0.1780267, 
    0.1882461, 0.2631966, 0.3156897, 0.2237267, 0.2884396, 0.2014162, 
    0.1888217, 0.2317333, 0.2672474, 0.2296981, 0.1468957, 0.1723389, 
    0.2200775, 0.1820833, 0.1986122, 0.301876, 0.2037272, 0.2624546, 
    0.2692548, 0.2030509, 0.2074263, 0.2187216,
  0.120075, 0.1269227, 0.1357409, 0.1398081, 0.1209072, 0.1447166, 0.1570603, 
    0.2221799, 0.2153738, 0.2067759, 0.173878, 0.1740746, 0.2086479, 
    0.2238948, 0.2353588, 0.05316889, 0.1689365, 0.1445747, 0.1755697, 
    0.1748177, 0.1703973, 0.1457056, 0.101071, 0.1024787, 0.1063405, 
    0.1609275, 0.2035098, 0.1752566, 0.09593457,
  0.07138778, 0.09848507, 0.08010408, 0.1493888, 0.1492015, 0.09566632, 
    0.1057635, 0.1188777, 0.1283128, 0.1167272, 0.1220229, 0.1306985, 
    0.1240317, 0.1711842, 0.1570412, 0.1181315, 0.1433178, 0.1744245, 
    0.2044174, 0.1533947, 0.07303204, 0.128619, 0.1323094, 0.1880405, 
    0.05758324, 0.09758011, 0.1216223, 0.0778955, 0.07977398,
  0.0855843, 0.006640422, 0.02884809, 0.05938987, 0.008965693, 0.00696545, 
    0.01930926, 0.03219148, 0.03530875, 0.01071569, 0.0185747, 0.01488859, 
    0.001795797, 0.04358631, 0.06916196, 0.09415534, 0.1184944, 0.1417971, 
    0.1642615, 0.1732158, 0.02681288, 0.04336128, 0.01779699, 0.01162755, 
    -0.0001545159, 0.04779229, 0.03863423, 0.04848451, 0.08521444,
  3.871936e-07, 4.504511e-08, 0.0008745306, 8.980378e-05, 0.009765869, 
    2.44569e-08, 0.0002591834, 0.00345885, 0.0001120195, 1.986189e-07, 
    3.150352e-08, 0.002584332, 0.009986182, 0.08116646, 0.05166321, 
    0.01360771, 0.02248657, 0.04613449, 0.02033728, 3.779872e-06, 
    0.0003499457, -1.782205e-06, -2.010459e-12, 1.271573e-07, 0.0003646095, 
    7.790725e-06, -0.0002442559, 4.024639e-07, 1.473395e-07,
  3.27171e-07, -5.669777e-06, -1.398914e-06, 0.0001598663, 0.06853751, 
    0.0117926, 0.02864934, 0.02501535, 0.04255233, 0.005346451, 0.0601702, 
    0.0178746, 0.15701, 0.02477256, 0.06901479, 0.003077107, 0.001387061, 
    0.0001962731, 5.688352e-07, 6.295838e-09, 3.795516e-10, 4.563398e-10, 
    3.143634e-08, 0.0003923636, 0.0002949642, 1.975968e-05, 0.00279025, 
    1.486056e-08, 8.030796e-08,
  0.04596582, 0.04391585, 0.03802336, 0.006381816, 0.003921936, 0.008380118, 
    0.0235698, 0.06786042, 0.04508895, 0.01182904, 0.03054928, 0.02962447, 
    0.144989, 0.06281731, 0.03888686, 0.01868509, 0.05208053, 0.0006411732, 
    1.418667e-05, 0.02956935, 0.0486365, 0.0002998428, 0.01496599, 0.124171, 
    0.08866403, 0.09760842, 0.1126019, 0.01418717, 0.004932843,
  0.02113304, 0.03680553, 0.06143362, 0.1318857, 0.0009879322, 0.01162707, 
    0.02344151, 0.04994032, 0.07528823, 0.1248496, 0.1152888, 0.1603568, 
    0.08648689, 0.05063474, 0.03767259, 0.04785339, 0.06317316, 0.02628973, 
    0.1175303, 0.02762216, 0.03000524, 0.06629498, 0.08517803, 0.01750599, 
    0.01970713, 0.02013062, 0.04403618, 0.1251264, 0.06909622,
  0.09703626, 0.02040228, 0.000526815, -6.372383e-05, 0.000978122, 
    0.04022309, 0.0581148, 0.1262653, 0.06974362, 0.08156042, 0.1567828, 
    0.125287, 0.02075344, 0.005303605, 0.003781104, 0.01013458, 0.004424295, 
    1.987729e-06, 4.153003e-06, 0.003882887, 0.0004645541, 0.006783982, 
    0.05367081, 0.04633807, 0.008138141, 0.00942067, 0.02853598, 0.03274096, 
    0.02529863,
  0.01604976, 0.05263092, 0.0005303433, 0.006998661, 0.004766599, 
    0.001706081, 0.009454011, 0.06200309, 0.2723009, 0.08029978, 0.2703502, 
    0.188823, 0.09692731, 0.04423804, 0.02456319, 0.08099245, 0.073139, 
    0.02150821, 0.005463976, 5.887299e-07, -0.000350837, 0.006235778, 
    0.03249957, 0.03131254, 0.07658822, 0.04202205, -0.0002995541, 
    1.915823e-05, 0.02218059,
  0.03882596, 0.09488135, 0.02045902, 0.02939214, 0.0749447, 0.02338191, 
    0.1647014, 0.03719584, 0.04001591, 0.06618038, 0.1695091, 0.0804193, 
    0.1686616, 0.1539285, 0.07564542, 0.1817698, 0.1464559, 0.06059549, 
    0.04068372, 0.05542766, 0.07949211, 0.03616099, 0.0708934, 0.04142275, 
    0.08451888, 0.1339706, 0.06282614, 0.02176494, 0.003023418,
  0.1327372, 0.1071532, 0.08684096, 0.05514259, 0.04773521, 0.09478765, 
    0.1448282, 0.09407832, 0.175749, 0.1063983, 0.1673943, 0.1697074, 
    0.1020065, 0.1123391, 0.07980376, 0.2306103, 0.2241039, 0.1487717, 
    0.1072097, 0.09233289, 0.1574777, 0.09314701, 0.06750973, 0.09563875, 
    0.1128986, 0.1795314, 0.1367981, 0.1161199, 0.1038196,
  0.1058563, 0.09425407, 0.07758459, 0.07231293, 0.08298755, 0.224336, 
    0.161986, 0.1480488, 0.1533554, 0.08367991, 0.08509591, 0.1250558, 
    0.139509, 0.1283839, 0.1126117, 0.1936526, 0.2148339, 0.1530938, 
    0.1162711, 0.08005825, 0.07448471, 0.1152934, 0.2050868, 0.2430014, 
    0.1751088, 0.2672622, 0.1940961, 0.156886, 0.09443022,
  0.09287565, 0.0949268, 0.06982812, 0.07630903, 0.1496913, 0.2468675, 
    0.1840038, 0.1298903, 0.1457704, 0.1342229, 0.07433221, 0.105601, 
    0.1513296, 0.08384399, 0.1324695, 0.07230095, 0.09288459, 0.09622028, 
    0.1498825, 0.1448998, 0.1462446, 0.130304, 0.1337671, 0.129518, 
    0.1441739, 0.4185877, 0.2514073, 0.1444856, 0.1617799,
  0.1278685, 0.2240013, 0.2412443, 0.1512187, 0.1460281, 0.2091719, 
    0.1893215, 0.1843222, 0.1803125, 0.1526195, 0.120311, 0.1164253, 
    0.1255094, 0.1908576, 0.2780393, 0.241079, 0.2109676, 0.1412399, 
    0.1274004, 0.2009407, 0.2032662, 0.2396842, 0.2580104, 0.1702489, 
    0.1547034, 0.1446885, 0.1398612, 0.08832178, 0.1124763,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0.0001204821, -3.668194e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, -4.428965e-05, 
    0.00222999, 0.2008225, 0.1764324, 0.1963225, 0.1797941, 0.1862451, 
    0.1324657, 0.04673965, 0.005868625, 0.001671866, 0.1429112, 0.4119538, 
    0.3375588, 0.2205141, 0.2204868, 0.07350474, 0.001181685,
  0.2066622, 0.2631941, 0.2177175, 0.2121623, 0.01532114, 0.1225758, 
    0.2096098, 0.108132, 0.08509007, 0.06505127, 0.08893563, 0.1075616, 
    0.1637887, 0.1800447, 0.2172519, 0.2685436, 0.2224423, 0.2379624, 
    0.1981031, 0.2559933, 0.2314737, 0.3072546, 0.2694827, 0.3737104, 
    0.3490904, 0.2618795, 0.3171606, 0.3709868, 0.362695,
  0.177927, 0.2104667, 0.2823597, 0.2153679, 0.3036214, 0.2890249, 0.1920567, 
    0.1818572, 0.2733188, 0.3365491, 0.2178661, 0.2670187, 0.2192165, 
    0.1955426, 0.2046973, 0.2448026, 0.213287, 0.1427147, 0.1817673, 
    0.2346319, 0.2075679, 0.2650252, 0.3045834, 0.248063, 0.2523471, 
    0.2699877, 0.2188851, 0.2269721, 0.2274712,
  0.1193114, 0.1208015, 0.1407945, 0.1586432, 0.1439808, 0.155642, 0.1420703, 
    0.2237344, 0.2284265, 0.2090585, 0.1660434, 0.16863, 0.1815049, 
    0.2035366, 0.2419906, 0.06879608, 0.1763859, 0.1426191, 0.1914697, 
    0.1565339, 0.1789517, 0.1422596, 0.09832372, 0.09452054, 0.1058651, 
    0.1505598, 0.1812807, 0.1650624, 0.09226005,
  0.06903129, 0.1098116, 0.08998568, 0.1483835, 0.1566818, 0.1033587, 
    0.10525, 0.1175218, 0.1418587, 0.1216373, 0.1359271, 0.1261416, 
    0.1227262, 0.1713228, 0.1611672, 0.1052545, 0.137162, 0.2016598, 
    0.1973557, 0.1369941, 0.07242516, 0.1199277, 0.1291698, 0.1955403, 
    0.05853856, 0.08422367, 0.1075382, 0.08034135, 0.09814645,
  0.07097904, 0.00959245, 0.02252758, 0.06338948, 0.01595027, 0.009647884, 
    0.02458377, 0.02978409, 0.03860816, 0.004839531, 0.01866009, 0.01100237, 
    0.002417614, 0.04547407, 0.0725809, 0.09639858, 0.09909628, 0.1178938, 
    0.1534318, 0.1852171, 0.0221585, 0.04400975, 0.01762822, 0.01230184, 
    0.0005423474, 0.05729344, 0.03614461, 0.04624944, 0.0807504,
  5.486423e-08, 3.303039e-08, 0.0009293883, 2.812573e-05, 0.005808268, 
    5.757455e-08, 0.001956748, 0.01048624, 2.912944e-05, 2.799886e-07, 
    2.342251e-07, 1.347824e-05, 0.01297679, 0.09531676, 0.04750461, 
    0.01496978, 0.01812022, 0.05704643, 0.0173666, 0.0004662772, 0.001452773, 
    -4.581185e-05, 1.622052e-10, 2.62145e-07, 0.0004593536, 9.308043e-06, 
    0.0003992932, 3.402336e-07, 6.838023e-08,
  6.04912e-07, 4.695983e-05, 1.188489e-06, 3.276216e-05, 0.06764203, 
    0.01754928, 0.03229284, 0.02913701, 0.03928488, 0.001917389, 0.0708299, 
    0.01873131, 0.1678169, 0.03410663, 0.06043593, 0.003568907, 0.001788137, 
    0.0003416289, 6.572383e-06, 6.764666e-09, 1.222113e-09, 2.275849e-08, 
    1.235591e-06, 0.0007811998, 0.000439368, 3.588618e-05, 2.968743e-05, 
    -2.972276e-08, 5.664558e-07,
  0.05815379, 0.05949262, 0.03631026, 0.006327282, 0.002277687, 0.01606337, 
    0.0355061, 0.0725093, 0.05276094, 0.01328431, 0.05871852, 0.04445081, 
    0.1801479, 0.06585029, 0.03961798, 0.03072713, 0.05118307, 0.008195694, 
    0.002471086, 0.03507422, 0.00771665, 0.001731372, 0.02633392, 0.1465566, 
    0.0938206, 0.1069233, 0.1047283, 0.0104609, 0.00476779,
  0.01823274, 0.02025918, 0.03094508, 0.326455, 0.0009080045, 0.01061901, 
    0.02849361, 0.05438656, 0.1354861, 0.1702828, 0.1718017, 0.1931262, 
    0.1007668, 0.05747385, 0.05175886, 0.05289984, 0.06103682, 0.04172331, 
    0.1170155, 0.04094392, 0.03637561, 0.08562917, 0.109761, 0.02484654, 
    0.02947354, 0.0291713, 0.05295388, 0.1381205, 0.08964126,
  0.03259435, 0.00835566, 6.415645e-05, -6.549559e-05, -3.497048e-05, 
    0.03967693, 0.05836391, 0.1413177, 0.1084523, 0.09872994, 0.1978786, 
    0.13985, 0.02579317, 0.006486046, 0.004184887, 0.01054699, 0.004112777, 
    1.310945e-06, 5.143377e-05, 0.0003956201, 0.0005722452, 0.006589847, 
    0.06074825, 0.0548997, 0.008833187, 0.008592688, 0.042358, 0.03979766, 
    0.02735636,
  0.003651034, 0.0216229, 0.0003906211, 0.003364978, 0.001248165, 
    4.224294e-05, 0.004401852, 0.06792689, 0.2853985, 0.07797798, 0.2682713, 
    0.2011554, 0.1055984, 0.04499447, 0.03222523, 0.09242105, 0.07489712, 
    0.02439103, 0.005136283, 3.00958e-06, -0.0004498302, 0.006562131, 
    0.03954788, 0.0370867, 0.09672044, 0.0396063, 0.0005251507, 3.695545e-05, 
    0.007243105,
  0.04040931, 0.07829598, 0.02546991, 0.03018646, 0.07087499, 0.01922512, 
    0.16313, 0.02385125, 0.0351437, 0.06319766, 0.1719443, 0.0674924, 
    0.1507205, 0.1459153, 0.06793573, 0.165405, 0.146749, 0.06327925, 
    0.04362953, 0.04700183, 0.08180658, 0.02960556, 0.05848306, 0.03806088, 
    0.08496263, 0.1562094, 0.06066512, 0.02845166, 0.004211102,
  0.1481029, 0.1256201, 0.1110418, 0.05574598, 0.07141262, 0.09481832, 
    0.1499889, 0.08718568, 0.1632446, 0.1009195, 0.1805425, 0.1591083, 
    0.1098079, 0.1301176, 0.09184309, 0.218866, 0.1761789, 0.1312493, 
    0.1131147, 0.1082513, 0.1769743, 0.1098148, 0.07672071, 0.1105609, 
    0.122177, 0.1631595, 0.1279914, 0.1162339, 0.07439539,
  0.1076261, 0.07662917, 0.07553049, 0.07300598, 0.07558189, 0.2288139, 
    0.1546632, 0.1396783, 0.151886, 0.09336711, 0.08747815, 0.1051899, 
    0.1267662, 0.1253811, 0.1194998, 0.2095334, 0.2245733, 0.1598214, 
    0.1070801, 0.07638805, 0.07144535, 0.1081048, 0.2154697, 0.2440543, 
    0.2196266, 0.2986427, 0.190974, 0.1468354, 0.08294196,
  0.1013799, 0.07110579, 0.0910339, 0.1045546, 0.1174055, 0.2207856, 
    0.1969667, 0.1106305, 0.1387505, 0.1472165, 0.08046429, 0.1073852, 
    0.1321047, 0.1321357, 0.1340853, 0.06322084, 0.07320443, 0.09785799, 
    0.1704693, 0.1428152, 0.1501712, 0.1408261, 0.1487306, 0.1337096, 
    0.1168196, 0.4232397, 0.2880867, 0.1616212, 0.1645312,
  0.1165417, 0.213773, 0.2306554, 0.1627724, 0.1281944, 0.1915511, 0.1945241, 
    0.196924, 0.2024447, 0.1718228, 0.1251824, 0.1406616, 0.1387719, 
    0.2240379, 0.3087786, 0.2472241, 0.2068386, 0.1718102, 0.1317695, 
    0.2323897, 0.2142387, 0.2677571, 0.2848909, 0.1781463, 0.1698548, 
    0.1398642, 0.1389582, 0.08752554, 0.1163275,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.752926e-05, -1.752926e-05, 
    -1.752926e-05, -1.752926e-05, -1.752926e-05, -1.752926e-05, 
    -1.752926e-05, 0, 0, 0, 0, 0, 0, 0, 0,
  0.0004958096, 0.0005761356, -2.044862e-05, 0, 0, -3.415105e-06, 
    -1.952542e-05, 0, 0, 0, -4.211217e-05, 0.001487181, 0.01176753, 
    0.2225032, 0.1957116, 0.1850153, 0.1798922, 0.1817148, 0.1576579, 
    0.1681365, 0.06566303, 0.05812815, 0.2153703, 0.4288198, 0.3486374, 
    0.2185599, 0.2204762, 0.1545638, 0.02267076,
  0.2020776, 0.2734941, 0.2146528, 0.2251337, 0.04621755, 0.2079906, 
    0.2539155, 0.2146882, 0.1720566, 0.1324931, 0.1266254, 0.1426684, 
    0.1865584, 0.1854459, 0.2309877, 0.2531192, 0.2135868, 0.2415989, 
    0.2382905, 0.2714102, 0.2404922, 0.3040979, 0.2821372, 0.3814827, 
    0.3417215, 0.2423107, 0.3011125, 0.3656512, 0.3636218,
  0.1959501, 0.2069008, 0.2837651, 0.2299994, 0.284249, 0.3036454, 0.206671, 
    0.1830318, 0.2795833, 0.3734338, 0.2240916, 0.2978054, 0.2003724, 
    0.1944288, 0.2029633, 0.2415845, 0.2096566, 0.1462676, 0.1601038, 
    0.2339292, 0.251317, 0.226889, 0.3056265, 0.2500417, 0.245301, 0.2600145, 
    0.190533, 0.1914828, 0.2117006,
  0.1158002, 0.1197076, 0.1469606, 0.1576542, 0.152288, 0.1451707, 0.1436896, 
    0.2421428, 0.2272004, 0.2047317, 0.1950811, 0.188641, 0.1711482, 
    0.1958588, 0.2180668, 0.08051741, 0.1921035, 0.1374611, 0.1733298, 
    0.1609087, 0.1901998, 0.156798, 0.09718763, 0.09281443, 0.104176, 
    0.1344711, 0.1655986, 0.1354342, 0.09649431,
  0.05894088, 0.1256024, 0.08797003, 0.1533688, 0.1639873, 0.1133785, 
    0.1068627, 0.1176495, 0.1517012, 0.1424004, 0.149188, 0.14023, 0.1101388, 
    0.172862, 0.1530037, 0.1041854, 0.1468033, 0.1699741, 0.1924027, 
    0.1325364, 0.08322566, 0.1340714, 0.1343426, 0.1951724, 0.05522465, 
    0.08172196, 0.1197772, 0.07706008, 0.09143467,
  0.07949762, 0.007915412, 0.02136888, 0.07699173, 0.02410739, 0.01095262, 
    0.02859196, 0.03475469, 0.03825564, 0.002629892, 0.01482135, 0.006757862, 
    0.003920823, 0.04940748, 0.07298727, 0.1051514, 0.0982435, 0.1096165, 
    0.133332, 0.2014422, 0.0218777, 0.04535107, 0.02444213, 0.0100247, 
    0.01397082, 0.06170911, 0.03649731, 0.05042401, 0.0696355,
  2.66273e-08, 2.796002e-08, 0.001215637, 1.978673e-05, 0.004553053, 
    1.37776e-07, 0.008273729, 0.03700374, 2.933469e-06, 2.148943e-07, 
    2.632361e-07, 1.639035e-06, 0.02259975, 0.118816, 0.05080647, 0.01655179, 
    0.01073881, 0.07175555, 0.0196268, 0.001171422, 0.0158471, -6.960583e-05, 
    1.181885e-08, 3.032007e-07, 0.0006707889, 1.795371e-05, 0.002369293, 
    -6.745649e-06, 6.349283e-08,
  1.837579e-06, 0.0001404347, -2.068676e-06, 0.0001936749, 0.0686754, 
    0.02625902, 0.03116798, 0.03469036, 0.04070792, 0.003170482, 0.06610321, 
    0.01796283, 0.1707813, 0.0455281, 0.0571031, 0.003442349, 0.002471386, 
    0.0006172349, 5.603251e-05, 1.268224e-08, -9.234374e-08, 9.055009e-08, 
    4.426826e-06, 0.001403524, 0.0005271069, 5.106835e-05, 0.0001762291, 
    -7.259468e-08, 4.571253e-06,
  0.02949019, 0.09715178, 0.04827567, 0.003218418, 0.001737014, 0.01625245, 
    0.03319284, 0.08320943, 0.05957557, 0.024475, 0.08153155, 0.05401361, 
    0.2015803, 0.07565565, 0.04182545, 0.03460414, 0.05125842, 0.02573282, 
    0.01999755, 0.03924939, 0.001079869, 0.003524975, 0.05019191, 0.1725414, 
    0.1109214, 0.1040036, 0.09942834, 0.01385858, 0.007157018,
  0.0185168, 0.01652752, 0.01822376, 0.3131444, 0.0007978939, 0.008108527, 
    0.04191368, 0.05146429, 0.1696934, 0.1849755, 0.2206306, 0.2275282, 
    0.1117866, 0.0531837, 0.0514243, 0.05480233, 0.05879622, 0.03902834, 
    0.1174189, 0.04012893, 0.0415976, 0.09950244, 0.1307492, 0.03596683, 
    0.03628628, 0.04248306, 0.07788473, 0.1582855, 0.1236536,
  0.004198022, 0.000450271, 1.491827e-05, -1.325651e-05, -5.137204e-06, 
    0.02847383, 0.07334461, 0.1184109, 0.1389534, 0.09900941, 0.204703, 
    0.136432, 0.02785918, 0.005184363, 0.003850431, 0.01220346, 0.005996275, 
    4.220146e-06, 0.0001758001, 1.156507e-05, 0.000126663, 0.007410646, 
    0.0669412, 0.06936779, 0.00782191, 0.004893323, 0.0381918, 0.03769984, 
    0.017746,
  0.0002185446, 0.001641973, 0.0004591382, 0.0003744867, 0.0001897375, 
    2.136821e-05, 0.004167906, 0.09232712, 0.307406, 0.06606743, 0.2555485, 
    0.2136009, 0.1072293, 0.06643976, 0.03228079, 0.08049977, 0.08680217, 
    0.02412405, 0.01054372, 3.35469e-06, -0.0003534426, 0.009069922, 
    0.05259912, 0.04877841, 0.1463281, 0.03781026, 0.003950346, 0.0001861452, 
    0.001509741,
  0.04478791, 0.05201976, 0.0209343, 0.03099991, 0.07339365, 0.008289056, 
    0.1507723, 0.01728329, 0.02316426, 0.06979549, 0.1894858, 0.06308071, 
    0.141414, 0.1426941, 0.08473957, 0.1528462, 0.1544079, 0.06460908, 
    0.04511714, 0.0385257, 0.05039159, 0.02367236, 0.06441151, 0.0478783, 
    0.08075282, 0.1754169, 0.05954415, 0.03596646, 0.003563774,
  0.154132, 0.1582463, 0.114379, 0.07272217, 0.08690884, 0.1035333, 
    0.1287082, 0.07985715, 0.1414467, 0.07659103, 0.1888095, 0.1685022, 
    0.08998054, 0.1248486, 0.1188549, 0.2513812, 0.193072, 0.1503177, 
    0.1393546, 0.1202524, 0.1694068, 0.1017349, 0.08960063, 0.128167, 
    0.1262236, 0.1601862, 0.120964, 0.1358395, 0.06164549,
  0.1208314, 0.08418765, 0.09299384, 0.09949328, 0.07086173, 0.2257079, 
    0.1699812, 0.1328619, 0.1490888, 0.08057901, 0.08745274, 0.0986862, 
    0.1204301, 0.1667055, 0.1437529, 0.2576412, 0.2177339, 0.1802633, 
    0.09373004, 0.06691679, 0.06893095, 0.129409, 0.2292174, 0.2498733, 
    0.2059588, 0.3123951, 0.2032588, 0.1401898, 0.09347879,
  0.108744, 0.04791126, 0.1029241, 0.1122266, 0.1584539, 0.2503728, 
    0.2089134, 0.1179737, 0.1335221, 0.1535965, 0.1059441, 0.1032482, 
    0.1215715, 0.1116462, 0.08850719, 0.05367168, 0.07529048, 0.13141, 
    0.1655145, 0.1314256, 0.1552677, 0.1632769, 0.145974, 0.1322511, 
    0.06522761, 0.4400298, 0.3080158, 0.1719445, 0.1703475,
  0.124277, 0.2008403, 0.2378862, 0.1570603, 0.1702313, 0.236553, 0.2544229, 
    0.2672151, 0.2503372, 0.1987239, 0.1685651, 0.1879618, 0.1763502, 
    0.2494534, 0.3275089, 0.2394776, 0.187035, 0.1382114, 0.09234121, 
    0.2511293, 0.276489, 0.3163438, 0.3333112, 0.1863577, 0.1865728, 
    0.1478551, 0.1311656, 0.09022486, 0.114968,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -6.310168e-05, -6.310168e-05, 
    -6.310168e-05, -6.310168e-05, -6.310168e-05, -6.310168e-05, 
    -6.310168e-05, 0, 0, 0, 0, 0, 0, 0, 0,
  0.02516185, 0.007534817, -0.0003580235, 0, 0, 4.734836e-05, -2.913667e-05, 
    0, 0, 0, 0.001992492, 0.00104598, 0.03017277, 0.2155555, 0.2008607, 
    0.1972815, 0.1917034, 0.1840394, 0.1583435, 0.204354, 0.1306812, 
    0.1796623, 0.2343133, 0.4575968, 0.3627736, 0.1989827, 0.1965649, 
    0.1787165, 0.04871317,
  0.2121019, 0.3093474, 0.2104404, 0.2482786, 0.128748, 0.2779049, 0.2908217, 
    0.2665525, 0.2445004, 0.1929148, 0.192414, 0.1583067, 0.2120279, 
    0.2270793, 0.2684316, 0.2322612, 0.222017, 0.2568046, 0.2472981, 
    0.2689485, 0.2677808, 0.2991648, 0.2677458, 0.3947901, 0.3384871, 
    0.2154824, 0.2934543, 0.3715642, 0.3313905,
  0.2229417, 0.2156661, 0.2763326, 0.2512414, 0.2888012, 0.3542418, 
    0.2448649, 0.1813868, 0.2333651, 0.3602635, 0.2565255, 0.3054613, 
    0.2356727, 0.1922253, 0.2336385, 0.2399117, 0.1900185, 0.1255074, 
    0.1700419, 0.2261792, 0.244163, 0.2169006, 0.3204584, 0.2486539, 
    0.2290115, 0.2321877, 0.2294452, 0.2067549, 0.2595255,
  0.1063002, 0.1252085, 0.1417764, 0.1734135, 0.1827535, 0.1894442, 
    0.1505858, 0.2770484, 0.2254518, 0.2067788, 0.2223254, 0.1857105, 
    0.1836567, 0.1957725, 0.2113011, 0.09098657, 0.2009899, 0.1577396, 
    0.1815499, 0.1527209, 0.1899856, 0.1678235, 0.104232, 0.08546971, 
    0.1101326, 0.1378857, 0.1625388, 0.1384498, 0.1122545,
  0.07516988, 0.1479949, 0.09171463, 0.1478736, 0.182935, 0.1269829, 
    0.1075214, 0.1341212, 0.1440706, 0.1395438, 0.1600894, 0.1350286, 
    0.107827, 0.1761926, 0.1478149, 0.1115322, 0.1487782, 0.1657802, 
    0.190529, 0.1269611, 0.08898354, 0.1357166, 0.1524978, 0.1915319, 
    0.0723936, 0.094308, 0.1183397, 0.08365538, 0.08398344,
  0.09317434, 0.01363921, 0.02247016, 0.09692878, 0.01916719, 0.01975737, 
    0.0290937, 0.03852113, 0.03350562, 0.00148579, 0.01029638, 0.01213272, 
    0.006887258, 0.05572612, 0.0792488, 0.1138385, 0.09874867, 0.1087662, 
    0.1314036, 0.1951094, 0.02559517, 0.04415504, 0.03485648, 0.005350142, 
    0.01695469, 0.07684908, 0.03773015, 0.06037818, 0.07647995,
  2.279063e-08, -1.375484e-08, 0.002425519, 4.845475e-05, 0.01098669, 
    1.316962e-05, 0.007303972, 0.04735485, 8.933729e-07, -1.412831e-06, 
    1.923177e-07, 9.309466e-08, 0.03515844, 0.1364903, 0.05839886, 
    0.01708614, 0.008213542, 0.08154603, 0.02027392, 0.001412289, 0.03544756, 
    9.437681e-05, 3.566792e-08, 2.916988e-07, 0.001677083, 0.0002766342, 
    0.009057119, 0.0001751105, 6.347917e-08,
  4.442115e-05, 7.484729e-05, 9.238687e-07, 0.001380397, 0.07040355, 
    0.02498026, 0.02408204, 0.0379364, 0.03023935, 0.002528938, 0.06247705, 
    0.01261513, 0.1313914, 0.04637841, 0.05832963, 0.005377904, 0.005630253, 
    0.001558007, 0.0001365191, 1.462688e-08, 1.720716e-08, 5.068554e-07, 
    1.140795e-05, 0.00198413, 0.0004330338, 8.383704e-05, 0.0005988647, 
    6.314976e-07, 1.7024e-05,
  0.01856847, 0.1380323, 0.05133098, 0.002054785, 0.00150591, 0.01627216, 
    0.03838846, 0.0757909, 0.04976435, 0.03254519, 0.07956968, 0.02829199, 
    0.1449206, 0.06525162, 0.04084209, 0.03701466, 0.04973295, 0.014529, 
    0.0131317, 0.02279497, 0.001437714, 0.008960743, 0.04943236, 0.2220582, 
    0.12469, 0.08358641, 0.09759337, 0.01564405, 0.0180582,
  0.01131515, 0.009802211, 0.00906902, 0.2046681, 0.001418245, 0.006231688, 
    0.0492936, 0.03308435, 0.07770754, 0.1228717, 0.1383204, 0.1526057, 
    0.08404469, 0.04060713, 0.04264034, 0.04572534, 0.04991955, 0.03894382, 
    0.1272013, 0.03146651, 0.03665824, 0.08079477, 0.1255184, 0.03874725, 
    0.03568553, 0.05574086, 0.0721771, 0.1417891, 0.1336821,
  0.002044281, -2.256464e-05, 8.263039e-06, 1.195619e-07, 2.618605e-07, 
    0.004912624, 0.06432736, 0.04073876, 0.1813714, 0.09452973, 0.1697099, 
    0.1133882, 0.02409313, 0.005625924, 0.005554063, 0.008421451, 
    0.007160849, 4.632896e-06, 4.73138e-05, 1.483988e-06, 3.192484e-06, 
    0.0073436, 0.05316125, 0.06445307, 0.007251314, 0.003814095, 0.02315719, 
    0.02131443, 0.005499698,
  2.258937e-05, 0.0001954621, 1.261632e-05, -1.990876e-05, 5.681538e-06, 
    4.085735e-06, 0.003172125, 0.1023007, 0.3406293, 0.05555102, 0.192939, 
    0.1983417, 0.1027647, 0.06746181, 0.02603422, 0.06946918, 0.09646361, 
    0.01976349, 0.01646586, 1.586433e-06, -0.000161162, 0.01307038, 
    0.05031164, 0.04990481, 0.177975, 0.03872579, 0.005997581, 0.0005988349, 
    0.0013688,
  0.04683994, 0.04080773, 0.01595322, 0.03420212, 0.05343334, 0.006040664, 
    0.1499728, 0.006804817, 0.008748237, 0.06549132, 0.2406929, 0.06466792, 
    0.1464501, 0.1345512, 0.09766264, 0.1875434, 0.1775486, 0.06950222, 
    0.0481644, 0.03883824, 0.0243966, 0.02068939, 0.08587514, 0.06175626, 
    0.08628106, 0.1881148, 0.06798087, 0.04075887, 0.003911041,
  0.151194, 0.163557, 0.140372, 0.1109929, 0.06262077, 0.1214531, 0.1136839, 
    0.08072659, 0.1199432, 0.06702907, 0.2069417, 0.1606131, 0.08817988, 
    0.1279865, 0.1807118, 0.2684084, 0.2125626, 0.1441705, 0.14826, 0.140884, 
    0.1574641, 0.08575172, 0.1107674, 0.1223664, 0.1296681, 0.1475188, 
    0.1210196, 0.1314975, 0.06732371,
  0.1313775, 0.080917, 0.1023399, 0.1103035, 0.1005317, 0.2421215, 0.1773832, 
    0.1455564, 0.1601596, 0.08093248, 0.07949086, 0.1205013, 0.1173498, 
    0.1346417, 0.1605719, 0.2326015, 0.242315, 0.2129169, 0.09001581, 
    0.06751077, 0.08158258, 0.1383986, 0.2328458, 0.2661427, 0.1769591, 
    0.3158741, 0.1975598, 0.1462421, 0.09888811,
  0.08786116, 0.06391685, 0.1061435, 0.1039951, 0.1226996, 0.2267163, 
    0.211962, 0.1134213, 0.1353513, 0.1656432, 0.08293653, 0.1133282, 
    0.156041, 0.1050313, 0.1019365, 0.0381487, 0.07999226, 0.1641991, 
    0.1730732, 0.1500356, 0.1843342, 0.1639621, 0.1856416, 0.1298877, 
    0.05768161, 0.4560735, 0.3274637, 0.1621868, 0.1706939,
  0.1033385, 0.2060614, 0.2562474, 0.1781958, 0.2043191, 0.246637, 0.2217945, 
    0.2363773, 0.2466387, 0.1761163, 0.1312112, 0.1988845, 0.1670427, 
    0.2064844, 0.2966024, 0.2373273, 0.207872, 0.1752915, 0.1510244, 
    0.2461667, 0.3111069, 0.3170692, 0.3528787, 0.2034922, 0.1846027, 
    0.1387732, 0.1147461, 0.1031394, 0.1005044,
  0.001202133, 0.0006541673, 0.0001062011, -0.0004417651, -0.0009897313, 
    -0.001537698, -0.002085664, -0.0003548568, -0.0002345664, -0.0001142759, 
    6.014522e-06, 0.000126305, 0.0002465954, 0.0003668859, -0.005060323, 
    -0.003962633, -0.002864943, -0.001767253, -0.0006695627, 0.0004281274, 
    0.001525818, -0.000157033, -0.0008270474, -0.001497062, -0.002167076, 
    -0.002837091, -0.003507105, -0.004177119, 0.001640506,
  0.0335715, 0.01821303, 0.0004035453, 0, 0, -0.0006981959, 0.0001635972, 0, 
    -6.625994e-08, 0, 0.004852092, 0.01321254, 0.06443733, 0.2140889, 
    0.1774149, 0.2093987, 0.1683237, 0.1777897, 0.1504618, 0.1883638, 
    0.1914034, 0.2831946, 0.2668545, 0.485863, 0.3799132, 0.171566, 
    0.1854274, 0.1827636, 0.1023377,
  0.2209061, 0.3070619, 0.2117909, 0.280881, 0.1936452, 0.3075067, 0.3189157, 
    0.3422411, 0.2944527, 0.2243302, 0.2006484, 0.1468152, 0.2332764, 
    0.2390187, 0.278568, 0.2762131, 0.2604596, 0.3002456, 0.278434, 
    0.2800579, 0.2839279, 0.3074133, 0.2715246, 0.4179284, 0.3383101, 
    0.2217672, 0.3087657, 0.3905103, 0.3359781,
  0.2548275, 0.2236188, 0.2743094, 0.294571, 0.306743, 0.3868317, 0.308104, 
    0.2712364, 0.2561862, 0.4003004, 0.3040524, 0.3273366, 0.2455509, 
    0.1871716, 0.2306457, 0.2328608, 0.2082313, 0.1436557, 0.1755903, 
    0.2631143, 0.2813253, 0.2542205, 0.3090899, 0.2369103, 0.2231779, 
    0.2472602, 0.2382367, 0.2784162, 0.3664259,
  0.1390942, 0.1333797, 0.1587834, 0.1886871, 0.1925608, 0.194185, 0.154982, 
    0.2625347, 0.2510708, 0.2218314, 0.2268834, 0.1899688, 0.1687755, 
    0.1882385, 0.2299929, 0.09970805, 0.1948199, 0.1874729, 0.1951606, 
    0.1572178, 0.1821093, 0.1761275, 0.1089468, 0.09972904, 0.1088255, 
    0.1511342, 0.1598912, 0.1353486, 0.1086429,
  0.09928901, 0.1575099, 0.1141132, 0.1385524, 0.1958288, 0.1301003, 
    0.1316358, 0.1436825, 0.1612318, 0.1429198, 0.1566975, 0.1348547, 
    0.1190956, 0.1848599, 0.1611465, 0.1285715, 0.1630793, 0.171227, 
    0.1809635, 0.1277917, 0.09607153, 0.1232088, 0.142377, 0.18853, 
    0.1099821, 0.1085619, 0.1184254, 0.09779614, 0.08494178,
  0.1098797, 0.02293279, 0.02732026, 0.09259175, 0.03079346, 0.02613368, 
    0.03345479, 0.05075914, 0.02950429, 0.006342174, 0.008932141, 0.01037236, 
    0.006878926, 0.06403105, 0.08444522, 0.1167438, 0.1050457, 0.1179993, 
    0.1244437, 0.2277315, 0.03674332, 0.05306321, 0.05480213, 0.006524746, 
    0.0431235, 0.09022982, 0.04208227, 0.06653729, 0.08384688,
  8.538932e-08, -1.1076e-05, 0.004016584, 0.0002682482, 0.01535375, 
    0.0007774312, 0.007714173, 0.0609917, 0.0001413192, 1.060475e-05, 
    6.632781e-08, 9.602602e-08, 0.04403912, 0.1359381, 0.05930854, 
    0.01702258, 0.00202464, 0.08701174, 0.02207982, 0.007906825, 0.04279957, 
    0.001935144, 6.105208e-08, 2.664831e-07, 0.007781289, 0.001057485, 
    0.01451558, 0.00056107, 6.395414e-08,
  6.464132e-06, 1.994854e-05, 3.323067e-06, 0.005645555, 0.07476113, 
    0.02413637, 0.0194559, 0.04407321, 0.02569674, 0.001803578, 0.0538268, 
    0.01413914, 0.1187814, 0.04153595, 0.06624409, 0.00922008, 0.008869262, 
    0.003386696, 0.0003974674, -1.87509e-06, 1.024473e-08, 5.414094e-07, 
    9.830939e-06, 0.005236808, 0.0004882272, 0.0002212961, 0.0004948733, 
    1.83546e-06, 4.022876e-05,
  0.01024853, 0.09925333, 0.03951254, 0.002215041, 0.001260761, 0.01298578, 
    0.04240586, 0.05709473, 0.04357425, 0.02991215, 0.06985474, 0.01909802, 
    0.1030594, 0.05225942, 0.04368654, 0.03152248, 0.05029679, 0.01582759, 
    0.006293019, 0.002633265, 0.007217659, 0.01536284, 0.03860567, 0.2268745, 
    0.1353242, 0.06653063, 0.1121704, 0.02329723, 0.01214809,
  0.00590877, 0.009455032, 0.01312201, 0.1090737, 0.002730198, 0.004328416, 
    0.05673841, 0.03272494, 0.05414465, 0.09417288, 0.0859849, 0.1140108, 
    0.07422093, 0.03452475, 0.04288019, 0.04868389, 0.0393528, 0.04922496, 
    0.123122, 0.02282867, 0.03934143, 0.07603806, 0.1104845, 0.03938855, 
    0.03830994, 0.07079063, 0.06724621, 0.1094539, 0.08665619,
  0.0007004774, 9.788327e-06, 5.045796e-06, 1.914739e-07, 4.321765e-08, 
    0.0002895999, 0.06195923, 0.02211261, 0.1635992, 0.1051455, 0.1622418, 
    0.0958014, 0.02323094, 0.008114315, 0.00657658, 0.006898602, 0.004860398, 
    2.313883e-06, -3.769617e-06, 3.537078e-07, 5.097785e-07, 0.007649099, 
    0.03721511, 0.03738588, 0.008984564, 0.006450742, 0.009437943, 
    0.00302506, 0.002356508,
  8.384738e-06, 7.353428e-05, 1.045814e-06, 5.442238e-06, 2.197508e-05, 
    7.941579e-07, 0.0005497232, 0.1991603, 0.3807961, 0.05362504, 0.1521357, 
    0.1799276, 0.08913513, 0.04351949, 0.01669316, 0.05032691, 0.1009831, 
    0.0186935, 0.01631401, 1.06189e-06, -2.114545e-05, 0.01186205, 
    0.05585931, 0.04477918, 0.1396526, 0.04018797, 0.01175502, 0.002396021, 
    0.0008216384,
  0.05274194, 0.04220521, 0.01062364, 0.03165753, 0.03575633, 0.008725887, 
    0.1364615, 0.007622909, 0.00652932, 0.04837557, 0.268064, 0.08230641, 
    0.1374737, 0.1308211, 0.1122516, 0.1813833, 0.178705, 0.07587636, 
    0.05921979, 0.03786789, 0.0138276, 0.01468724, 0.08972871, 0.04786702, 
    0.09185882, 0.1883492, 0.0728462, 0.04495976, 0.01665442,
  0.179095, 0.1818191, 0.1691731, 0.1239673, 0.04894432, 0.08898491, 
    0.07342059, 0.07918638, 0.08983365, 0.07983822, 0.2194652, 0.1651789, 
    0.08135268, 0.1311435, 0.2314492, 0.3066662, 0.2488442, 0.1915232, 
    0.139154, 0.1816817, 0.1650135, 0.06519957, 0.1040136, 0.1614922, 
    0.1493936, 0.1574412, 0.1421405, 0.1773458, 0.06901811,
  0.1410996, 0.08923654, 0.1109547, 0.1013949, 0.1087522, 0.2370281, 
    0.1951823, 0.1536043, 0.1642107, 0.09155951, 0.08889531, 0.1671329, 
    0.1238481, 0.1232727, 0.1812914, 0.2418775, 0.2636319, 0.2665946, 
    0.1028271, 0.07753787, 0.1053838, 0.1326019, 0.2306509, 0.2885766, 
    0.1782502, 0.311255, 0.2101187, 0.1419101, 0.1173444,
  0.1388782, 0.0789473, 0.1239323, 0.1104926, 0.1826022, 0.2711857, 
    0.2259983, 0.134345, 0.1509233, 0.1757888, 0.1302241, 0.1029171, 
    0.1468309, 0.1369248, 0.1004458, 0.05914513, 0.1125052, 0.1771188, 
    0.1809836, 0.1347118, 0.1830924, 0.1804711, 0.1844431, 0.12315, 
    0.05190919, 0.4571783, 0.3140958, 0.1865222, 0.1779568,
  0.1308055, 0.2431858, 0.2880507, 0.1781965, 0.1450825, 0.1598923, 0.158405, 
    0.1915661, 0.1660686, 0.1578695, 0.1110278, 0.1622759, 0.1535373, 
    0.1920848, 0.3081253, 0.2677901, 0.2163479, 0.1987448, 0.1350984, 
    0.2469809, 0.3075967, 0.278708, 0.3703818, 0.19641, 0.1946856, 0.13074, 
    0.1088221, 0.1106713, 0.133858,
  0.02846045, 0.02513455, 0.02180865, 0.01848275, 0.01515685, 0.01183094, 
    0.008505044, 0.01211774, 0.0136193, 0.01512086, 0.01662242, 0.01812398, 
    0.01962554, 0.02112709, 0.01536664, 0.02255501, 0.02974338, 0.03693175, 
    0.04412011, 0.05130848, 0.05849685, 0.06026891, 0.05490489, 0.04954086, 
    0.04417684, 0.03881281, 0.03344879, 0.02808476, 0.03112117,
  0.07290995, 0.02468314, 0.009912843, -0.0001942209, -3.607374e-06, 
    -0.0007650542, -0.001872539, -0.001155611, 0.0003058097, 0.0003534213, 
    0.005716602, 0.05486877, 0.1184017, 0.2016234, 0.1630906, 0.2104014, 
    0.1651128, 0.1578602, 0.1475464, 0.1598183, 0.1913778, 0.3416512, 
    0.2986235, 0.5142877, 0.3771623, 0.1482725, 0.1939641, 0.1812471, 
    0.1179804,
  0.2502098, 0.2963357, 0.2382747, 0.2981966, 0.2396655, 0.3155515, 
    0.3225031, 0.4195329, 0.3278838, 0.2227133, 0.2034493, 0.1387134, 
    0.2462542, 0.2405087, 0.3166384, 0.2922728, 0.2653477, 0.2700216, 
    0.2664914, 0.2861641, 0.2634614, 0.2854369, 0.2451598, 0.4074989, 
    0.3576833, 0.1904425, 0.2754555, 0.3990997, 0.3500845,
  0.2865268, 0.2347467, 0.3079888, 0.3476508, 0.3392694, 0.4022874, 
    0.2860516, 0.300279, 0.3248807, 0.4192214, 0.310179, 0.3411432, 
    0.2582991, 0.1871134, 0.2379885, 0.2590356, 0.2248418, 0.1497587, 
    0.228631, 0.3365038, 0.3277708, 0.26873, 0.3266975, 0.2611657, 0.2120394, 
    0.2496376, 0.2301246, 0.2304183, 0.3463225,
  0.1772361, 0.1756002, 0.2140541, 0.2229863, 0.2033544, 0.1945886, 
    0.1654864, 0.2802623, 0.2326893, 0.2613945, 0.211294, 0.1816447, 
    0.1736277, 0.2010576, 0.2308747, 0.1303286, 0.2249919, 0.1697323, 
    0.2177533, 0.1709263, 0.2200706, 0.1789568, 0.1207133, 0.119716, 
    0.1167208, 0.172187, 0.165436, 0.1664158, 0.1135586,
  0.1416499, 0.1870804, 0.1460288, 0.1382625, 0.2355798, 0.1431976, 
    0.1594319, 0.1737022, 0.1803635, 0.1570113, 0.1638912, 0.1507528, 
    0.1335413, 0.2031329, 0.1792393, 0.13993, 0.1890896, 0.1724408, 
    0.1846474, 0.1555036, 0.132918, 0.1263366, 0.1393334, 0.1874969, 
    0.1312272, 0.1355916, 0.1213993, 0.1097257, 0.107894,
  0.1292615, 0.032622, 0.04353419, 0.08598723, 0.05235087, 0.0306603, 
    0.04147521, 0.07299972, 0.0291687, 0.01569707, 0.007864185, 0.01823725, 
    0.01661086, 0.07549474, 0.09197142, 0.1186246, 0.1138519, 0.1290253, 
    0.1156386, 0.2470475, 0.05684907, 0.06856833, 0.06290282, 0.007615882, 
    0.05793208, 0.09803694, 0.04713987, 0.081882, 0.09341779,
  2.408866e-07, -3.312241e-06, 0.02825247, 0.001954111, 0.0296066, 
    0.01126901, 0.0146598, 0.07296845, 0.004526228, 9.526951e-05, 
    1.564171e-08, 0.000173628, 0.04774438, 0.1113984, 0.06875639, 0.01659291, 
    0.002544777, 0.09724113, 0.03562451, 0.03297022, 0.05388166, 0.005388636, 
    -1.089291e-07, 1.61259e-07, 0.02537391, 0.004137087, 0.02347428, 
    0.003174407, -1.284258e-06,
  4.347727e-06, -3.404441e-05, 5.522326e-05, 0.02230233, 0.07425705, 
    0.02854366, 0.02124356, 0.04244918, 0.02303591, 0.002373973, 0.05051536, 
    0.01698427, 0.1218837, 0.0432379, 0.06435546, 0.01904474, 0.01616704, 
    0.006273963, 0.001889748, 0.0001429148, 2.197717e-09, 3.166669e-07, 
    3.361081e-06, 0.006895492, 0.001041829, 0.003209051, 0.01111169, 
    2.170166e-05, 2.518958e-05,
  0.006342549, 0.09728961, 0.04356156, 0.002269929, 0.001230416, 0.0122098, 
    0.0507652, 0.05246048, 0.0424974, 0.03480808, 0.07017206, 0.0143797, 
    0.08935729, 0.04863612, 0.05072391, 0.03637476, 0.05536652, 0.02243987, 
    0.02007294, 0.0003314164, 0.002750689, 0.003229576, 0.0400987, 0.2245903, 
    0.1498902, 0.06213506, 0.1250195, 0.03439464, 0.008545844,
  0.005382496, 0.007486293, 0.008797026, 0.04302385, 0.001001667, 
    0.004923975, 0.07882663, 0.02549646, 0.04173483, 0.08144046, 0.04903096, 
    0.1024487, 0.06512508, 0.03927634, 0.04523084, 0.04559979, 0.04024922, 
    0.07216282, 0.1240734, 0.01210468, 0.05164596, 0.07420775, 0.1016244, 
    0.04103881, 0.0371539, 0.07167434, 0.05798899, 0.09710844, 0.08008774,
  0.0001649583, 6.223833e-06, 3.294102e-06, 1.079004e-07, 2.691716e-08, 
    -8.954803e-05, 0.06829356, 0.01300721, 0.1691836, 0.09963182, 0.148594, 
    0.09268766, 0.02660549, 0.01487771, 0.01091711, 0.01028429, 0.0041353, 
    -2.598287e-08, -2.497209e-06, 1.368847e-07, 6.71196e-07, 0.009852051, 
    0.03170563, 0.04694108, 0.01146028, 0.01436267, 0.0001863321, 
    0.0006894639, 0.001567934,
  5.535823e-06, 4.738423e-05, 5.377355e-07, 3.163211e-06, 8.790277e-06, 
    2.974004e-07, -0.0006019594, 0.2838531, 0.3861737, 0.043818, 0.1349174, 
    0.164108, 0.08483518, 0.03131887, 0.02231368, 0.09066661, 0.08342776, 
    0.02183692, 0.01446372, 7.447876e-07, 8.831564e-07, 0.009758358, 
    0.04938914, 0.03526253, 0.1258664, 0.03632425, 0.02140848, 0.00545363, 
    7.247721e-05,
  0.04390343, 0.0388502, 0.004801845, 0.03111215, 0.01890584, 0.00425625, 
    0.1109277, 0.01092484, 0.006290535, 0.04694549, 0.2850015, 0.1041839, 
    0.1389188, 0.123858, 0.138264, 0.1551603, 0.2054489, 0.07040641, 
    0.07227939, 0.05031531, 0.00959802, 0.01035886, 0.08535133, 0.03968138, 
    0.06170567, 0.1697815, 0.06276696, 0.05327721, 0.01535516,
  0.2586448, 0.210945, 0.1807, 0.1004613, 0.05752286, 0.09672477, 0.06639504, 
    0.0945582, 0.0921038, 0.1319289, 0.2459995, 0.2142876, 0.08745547, 
    0.1737172, 0.2526231, 0.2813179, 0.2671504, 0.2146197, 0.1328051, 
    0.2057124, 0.1293912, 0.06098, 0.103117, 0.1855473, 0.1655978, 0.1510281, 
    0.1374558, 0.167095, 0.07898405,
  0.1479229, 0.1114422, 0.1101282, 0.1195049, 0.1399192, 0.2671849, 
    0.2462267, 0.1766967, 0.1585195, 0.09423602, 0.1061115, 0.2027116, 
    0.1589762, 0.189495, 0.1962729, 0.2563542, 0.3059084, 0.3251645, 
    0.1326445, 0.08023086, 0.1054471, 0.1732045, 0.2125336, 0.3067497, 
    0.2018703, 0.3201773, 0.2584755, 0.1438634, 0.1037783,
  0.1894555, 0.06961953, 0.1422019, 0.1312528, 0.1867671, 0.2587779, 
    0.2443264, 0.1762363, 0.1996271, 0.201808, 0.1359051, 0.1090222, 
    0.1821267, 0.1453452, 0.1759087, 0.09645279, 0.1180213, 0.2012472, 
    0.1804457, 0.1473475, 0.1969738, 0.2057552, 0.2082922, 0.1096748, 
    0.06907322, 0.4280198, 0.3116394, 0.1723735, 0.1866488,
  0.154817, 0.2703875, 0.2811407, 0.1707522, 0.1779952, 0.1711422, 0.1712917, 
    0.2018289, 0.1711118, 0.2046643, 0.1673822, 0.2402926, 0.2515811, 
    0.2838975, 0.3393277, 0.3497975, 0.3325506, 0.3202307, 0.2064466, 
    0.285972, 0.3569647, 0.34001, 0.3892531, 0.2019361, 0.1921927, 0.1418679, 
    0.1245481, 0.1066282, 0.1512447,
  0.07693093, 0.07670315, 0.07647537, 0.07624759, 0.0760198, 0.07579202, 
    0.07556424, 0.1031714, 0.1092391, 0.1153069, 0.1213747, 0.1274425, 
    0.1335102, 0.139578, 0.1248448, 0.1282206, 0.1315965, 0.1349723, 
    0.1383481, 0.1417239, 0.1450998, 0.1248119, 0.1155961, 0.1063802, 
    0.09716443, 0.08794862, 0.0787328, 0.06951699, 0.07711316,
  0.08872149, 0.05468274, 0.02009241, 0.00241976, -0.0006976654, 0.007018178, 
    0.002843042, 0.002573826, 0.001656383, 0.002330404, 0.01770627, 
    0.1013065, 0.1626809, 0.2080076, 0.1530759, 0.1803427, 0.1595632, 
    0.1451481, 0.1457837, 0.1560421, 0.2145406, 0.3608635, 0.3470549, 
    0.5262598, 0.3835413, 0.1277936, 0.2129931, 0.1715576, 0.1491212,
  0.2446735, 0.3246088, 0.2779773, 0.2823255, 0.3215525, 0.3231295, 
    0.3145132, 0.4739742, 0.3520871, 0.2305549, 0.2085349, 0.14756, 
    0.2519139, 0.2581726, 0.2800582, 0.2689335, 0.2437135, 0.2729422, 
    0.2964559, 0.2973328, 0.3014988, 0.2590787, 0.2217548, 0.3935052, 
    0.3507277, 0.1739909, 0.2596515, 0.3966311, 0.3373199,
  0.2755736, 0.2335631, 0.3073275, 0.2968345, 0.2894666, 0.367389, 0.2617307, 
    0.2311551, 0.336654, 0.3669553, 0.272377, 0.3643455, 0.2709654, 
    0.1920409, 0.2626101, 0.2756603, 0.2505274, 0.1775814, 0.2269264, 
    0.3397845, 0.3083058, 0.2945771, 0.3499061, 0.2820757, 0.2112862, 
    0.2589411, 0.2629431, 0.2740384, 0.3173277,
  0.2019835, 0.216666, 0.2635434, 0.2467978, 0.2376501, 0.2002965, 0.1942672, 
    0.2880178, 0.2302782, 0.2867917, 0.2343148, 0.1949445, 0.1756297, 
    0.2003028, 0.2506337, 0.1200008, 0.229178, 0.2396418, 0.2531967, 
    0.2156419, 0.2241117, 0.1884939, 0.1350292, 0.1415821, 0.1017063, 
    0.1655181, 0.1734409, 0.1562663, 0.1090318,
  0.1534102, 0.215626, 0.1646843, 0.1428608, 0.2542071, 0.1992452, 0.1785957, 
    0.1948604, 0.1968043, 0.1758049, 0.1781612, 0.1604815, 0.1452232, 
    0.2208881, 0.2053964, 0.1535344, 0.2164737, 0.1811191, 0.2016577, 
    0.15373, 0.1695882, 0.1580785, 0.1487114, 0.1848103, 0.1405129, 
    0.1410923, 0.1237373, 0.1259059, 0.132847,
  0.1412882, 0.04047035, 0.06296425, 0.08043836, 0.03642521, 0.0423091, 
    0.04688536, 0.07839569, 0.04519345, 0.02928978, 0.007846729, 0.01024108, 
    0.0458839, 0.08886504, 0.1044382, 0.1265386, 0.1245246, 0.1197044, 
    0.1037972, 0.2614054, 0.0799498, 0.07703017, 0.07202944, 0.009001444, 
    0.06593475, 0.114344, 0.06778385, 0.09024806, 0.105103,
  4.971677e-05, 1.023874e-07, 0.01158627, 0.005323161, 0.05193556, 
    0.01921291, 0.02189662, 0.08485428, 0.01109869, 0.0001008243, 
    3.596075e-09, 0.005702284, 0.05158316, 0.09999274, 0.1189161, 0.0249306, 
    0.008419082, 0.09920879, 0.05460213, 0.04201346, 0.09313269, 0.02225165, 
    -9.435757e-06, 2.059089e-07, 0.0300501, 0.01032445, 0.03164957, 
    0.01507718, 0.0001274307,
  1.476567e-06, 0.0002281078, 0.0003627595, 0.06260984, 0.08568388, 
    0.03839481, 0.02713926, 0.04064447, 0.02282574, 0.004806281, 0.05248029, 
    0.04013639, 0.1231333, 0.04706762, 0.06267215, 0.02869882, 0.01814131, 
    0.004431425, 0.004672813, 0.001447585, -1.209224e-06, 1.493559e-07, 
    1.076696e-06, 0.008814631, 0.0194172, 0.1040252, 0.04061628, 0.001612715, 
    8.755237e-06,
  0.00277776, 0.1003211, 0.04968264, 0.009452643, 0.002109363, 0.01326771, 
    0.05592887, 0.04673471, 0.04308846, 0.03924824, 0.06829698, 0.01252487, 
    0.07335664, 0.04329495, 0.05283514, 0.04525772, 0.06473707, 0.03403941, 
    0.02842274, 0.000100515, 0.0018203, 0.003211378, 0.03302942, 0.2081625, 
    0.1606952, 0.04998989, 0.1296911, 0.04237784, 0.007336189,
  0.00656527, 0.005782769, 0.003263507, 0.009120602, 0.0006315637, 
    0.005102214, 0.07983346, 0.02157239, 0.03246456, 0.06095471, 0.03316091, 
    0.08915211, 0.06281794, 0.04663696, 0.05059138, 0.05048312, 0.03711426, 
    0.09735312, 0.1236048, 0.006682565, 0.06318126, 0.07644317, 0.1014899, 
    0.0482643, 0.0403068, 0.07888197, 0.05475452, 0.08439928, 0.08544708,
  1.52798e-05, 3.824678e-06, 1.920374e-06, 3.384436e-08, 2.410036e-08, 
    -2.789481e-06, 0.05807006, 0.01171541, 0.1600818, 0.1144192, 0.1287899, 
    0.09028897, 0.02965278, 0.03032129, 0.02553486, 0.01523371, 0.004657583, 
    0.0005685635, 3.411324e-06, 1.206717e-07, 7.238723e-07, 0.009121113, 
    0.02516395, 0.04553263, 0.01494161, 0.01862059, -3.672068e-05, 
    0.0001083126, 0.0003164616,
  3.966237e-06, 1.987171e-05, 4.184222e-07, 2.085498e-06, 9.651748e-07, 
    9.98615e-08, -0.000595475, 0.22158, 0.3537986, 0.03625606, 0.1301285, 
    0.1484962, 0.08517066, 0.02739147, 0.04494637, 0.08168224, 0.08187187, 
    0.02433375, 0.01264904, 2.226686e-06, 1.130836e-06, 0.005656829, 
    0.05241272, 0.03277305, 0.1013386, 0.03956607, 0.03362558, 0.008011614, 
    7.251198e-06,
  0.03350665, 0.03460297, 0.004105151, 0.03394287, 0.0109685, 0.002071009, 
    0.08536728, 0.008050305, 0.00298908, 0.03907561, 0.3164077, 0.1042076, 
    0.1367417, 0.1187508, 0.1510228, 0.1586606, 0.2132294, 0.06566513, 
    0.07584159, 0.05463297, 0.01011132, 0.01059759, 0.08568309, 0.05150936, 
    0.06718542, 0.1624157, 0.06018531, 0.04723589, 0.0165145,
  0.2240821, 0.2125362, 0.1790354, 0.08290399, 0.06495054, 0.08570675, 
    0.05186297, 0.1161594, 0.1193095, 0.1488107, 0.2529563, 0.2242212, 
    0.08282059, 0.1720519, 0.2045965, 0.3408982, 0.2614203, 0.2127027, 
    0.139424, 0.1939866, 0.1182144, 0.05248313, 0.07965273, 0.2176824, 
    0.1684527, 0.1668342, 0.1327803, 0.1814277, 0.08153977,
  0.1435372, 0.1353988, 0.1196298, 0.1138944, 0.3007391, 0.3174798, 
    0.2421561, 0.1673761, 0.1823009, 0.1059781, 0.1666589, 0.2451382, 
    0.1680853, 0.2055924, 0.2729324, 0.234427, 0.3469614, 0.3419343, 
    0.1346286, 0.09679018, 0.1167741, 0.1815011, 0.2072841, 0.302726, 
    0.1973681, 0.3309772, 0.260976, 0.1721629, 0.1221437,
  0.2704171, 0.1915361, 0.1345443, 0.1423906, 0.2216533, 0.2923558, 
    0.2910518, 0.1809413, 0.1943949, 0.2013782, 0.1811261, 0.1309378, 
    0.2194626, 0.1587467, 0.1376521, 0.0831307, 0.1502707, 0.2220846, 
    0.140948, 0.1446074, 0.202445, 0.2004009, 0.2224592, 0.09715015, 
    0.08120435, 0.4008694, 0.2948115, 0.1723147, 0.2219761,
  0.09060984, 0.2328014, 0.2591974, 0.1907799, 0.1561511, 0.141609, 
    0.1712674, 0.1904096, 0.1970702, 0.2395615, 0.24055, 0.3124381, 
    0.3127162, 0.3519969, 0.349004, 0.347981, 0.2992863, 0.2334139, 
    0.1113352, 0.1753547, 0.3002841, 0.3535245, 0.4371428, 0.2239653, 
    0.2312677, 0.1507586, 0.1333984, 0.1079106, 0.08029781,
  0.1006265, 0.1005999, 0.1005733, 0.1005467, 0.1005201, 0.1004935, 
    0.1004668, 0.1351729, 0.1456369, 0.1561009, 0.1665649, 0.1770289, 
    0.187493, 0.197957, 0.2007695, 0.2013274, 0.2018854, 0.2024433, 
    0.2030012, 0.2035592, 0.2041171, 0.1753349, 0.1643396, 0.1533443, 
    0.1423489, 0.1313536, 0.1203583, 0.1093629, 0.1006478,
  0.1012162, 0.07676516, 0.03771538, 0.01404703, 0.002951419, 0.02663934, 
    0.04057451, 0.03863859, 0.02323557, 0.007313732, 0.05798226, 0.1252359, 
    0.181601, 0.2062911, 0.1511407, 0.133466, 0.1423394, 0.1343613, 
    0.1460302, 0.1429685, 0.2399686, 0.3686879, 0.4133964, 0.5345943, 
    0.3925084, 0.1231253, 0.2214582, 0.1497265, 0.1603406,
  0.2466433, 0.3088153, 0.3070039, 0.298492, 0.3924966, 0.3365572, 0.3288312, 
    0.4659361, 0.3603081, 0.2518253, 0.21673, 0.1582009, 0.2402573, 
    0.2700093, 0.2866013, 0.2557878, 0.2620544, 0.2593197, 0.2880507, 
    0.2655324, 0.296387, 0.3022606, 0.2379123, 0.4105284, 0.3195853, 
    0.2025366, 0.2722627, 0.4126486, 0.3165458,
  0.2183362, 0.2583255, 0.3618321, 0.3016406, 0.3091175, 0.3291619, 
    0.3353376, 0.2433959, 0.319565, 0.3577858, 0.2553977, 0.3451329, 
    0.2625993, 0.279729, 0.2821968, 0.2487735, 0.2432903, 0.1553247, 
    0.1952347, 0.3051057, 0.3044325, 0.2934544, 0.3285593, 0.2965724, 
    0.1881399, 0.2715524, 0.2806962, 0.2878968, 0.2802365,
  0.2319933, 0.2374048, 0.2747565, 0.2778349, 0.2573393, 0.210108, 0.1853994, 
    0.3051668, 0.2452586, 0.282047, 0.2451936, 0.2036854, 0.2360332, 
    0.2046748, 0.2925314, 0.1516253, 0.2391511, 0.3090727, 0.3073425, 
    0.2502367, 0.2132883, 0.1920044, 0.1584484, 0.1422025, 0.1059229, 
    0.155291, 0.1760589, 0.1766683, 0.1500369,
  0.1865926, 0.2389136, 0.1974735, 0.1792744, 0.2603841, 0.2101769, 
    0.1705565, 0.2185276, 0.1889334, 0.2062444, 0.196837, 0.1814215, 
    0.1450061, 0.2348115, 0.2314824, 0.1798526, 0.2362352, 0.1895058, 
    0.2033636, 0.1434501, 0.1896114, 0.1622235, 0.1839217, 0.1968113, 
    0.1544296, 0.1543386, 0.150028, 0.1539476, 0.1480156,
  0.1473609, 0.0558205, 0.07576936, 0.06633598, 0.0282103, 0.05579151, 
    0.05885402, 0.09036554, 0.05428564, 0.03389375, 0.02171298, 0.02093279, 
    0.05151995, 0.09669238, 0.099714, 0.1330641, 0.1209927, 0.1036264, 
    0.099452, 0.2580037, 0.08414787, 0.09121581, 0.0732512, 0.00717626, 
    0.06949808, 0.1155032, 0.08475568, 0.08648514, 0.1098514,
  0.01218202, -2.323427e-06, 0.03129783, 0.005979912, 0.04229461, 0.04896896, 
    0.04111392, 0.08321749, 0.01218557, 0.0003264074, 2.718541e-09, 
    0.001521679, 0.05197594, 0.089604, 0.1573979, 0.02645185, 0.01642098, 
    0.08640467, 0.05303212, 0.0604519, 0.1109263, 0.03686577, -6.565773e-05, 
    2.831559e-07, 0.02118428, 0.03877069, 0.04291647, 0.04490995, 0.008034643,
  1.322628e-06, -7.705453e-05, 0.0009135455, 0.1167229, 0.07809733, 
    0.0582734, 0.03715888, 0.0387552, 0.01905222, 0.01550477, 0.07356995, 
    0.06623444, 0.1121623, 0.04327871, 0.05352064, 0.02992514, 0.02237073, 
    0.006521064, 0.006812545, 0.001699299, 0.0001355426, 3.027741e-07, 
    1.589326e-07, 0.00910764, 0.005893107, 0.03107153, 0.06054838, 
    0.007460785, 1.475977e-05,
  0.001352228, 0.1050503, 0.06091498, 0.01390065, 0.008504323, 0.01718613, 
    0.05556255, 0.03931846, 0.04643618, 0.0459805, 0.07934343, 0.01148858, 
    0.05051025, 0.03608933, 0.04866359, 0.04111689, 0.05936695, 0.04377537, 
    0.02438397, 0.001519013, 0.000520922, 0.002893355, 0.02451414, 0.2015099, 
    0.1648295, 0.03762452, 0.1139989, 0.03630765, 0.00493812,
  0.007240937, 0.003546708, 0.001374342, 0.003517829, 0.0005010164, 
    0.00693452, 0.06994952, 0.0174987, 0.02129262, 0.04894458, 0.02529465, 
    0.07465443, 0.0556726, 0.04880663, 0.05552129, 0.06123624, 0.03766088, 
    0.1045218, 0.1207462, 0.008323351, 0.06314649, 0.07630417, 0.1041759, 
    0.06380359, 0.03852007, 0.08744841, 0.06341166, 0.06361809, 0.0704417,
  2.993632e-06, 2.602533e-06, 1.001669e-06, 1.502744e-08, 1.210901e-08, 
    -1.223823e-07, 0.04523313, 0.01162827, 0.1466658, 0.1141458, 0.1118234, 
    0.08037618, 0.02914927, 0.03397707, 0.04046556, 0.02627808, 0.01290833, 
    0.0060718, 1.5972e-06, 8.844224e-08, 4.758202e-07, 0.009862345, 
    0.02072369, 0.02564586, 0.02610783, 0.0284442, 0.0005444571, 
    1.269862e-06, 5.168179e-05,
  2.462947e-06, 8.109447e-06, 2.44345e-07, 1.607403e-06, 6.949048e-07, 
    6.61486e-08, -0.0003378169, 0.1343383, 0.3589616, 0.03304541, 0.1234815, 
    0.1441076, 0.08089269, 0.02962856, 0.08114189, 0.05943324, 0.118737, 
    0.05040013, 0.009154448, 6.735174e-05, 9.682809e-07, 0.003415291, 
    0.0568145, 0.03280303, 0.07137437, 0.05075242, 0.04350187, 0.008137431, 
    3.081112e-06,
  0.02241307, 0.01418149, 0.002835993, 0.0366034, 0.00422931, 0.0005795287, 
    0.06738119, 0.004878723, 0.0002732234, 0.02968824, 0.3364855, 0.09865326, 
    0.1148715, 0.1268331, 0.121981, 0.1888362, 0.2106134, 0.06436092, 
    0.07452403, 0.05441921, 0.005938642, 0.007980547, 0.07073786, 0.05821782, 
    0.09298379, 0.1671771, 0.06816195, 0.06513951, 0.01914074,
  0.2155372, 0.2245187, 0.1664497, 0.1160849, 0.04881724, 0.04299957, 
    0.04055451, 0.1241308, 0.1157353, 0.1056918, 0.2804084, 0.2458674, 
    0.08226655, 0.1572704, 0.2145819, 0.3686633, 0.2629104, 0.2045128, 
    0.142345, 0.2233387, 0.0913915, 0.0317169, 0.07233556, 0.2248868, 
    0.1688717, 0.1766883, 0.1455059, 0.1708546, 0.110131,
  0.1509987, 0.1131789, 0.1469216, 0.1386394, 0.3268635, 0.3163632, 
    0.2213622, 0.1703547, 0.1847548, 0.1041889, 0.1578306, 0.2203279, 
    0.1752063, 0.2000285, 0.2675405, 0.2512708, 0.350119, 0.350176, 
    0.1299137, 0.09610894, 0.1094659, 0.1516841, 0.1975743, 0.2680072, 
    0.1688307, 0.3454312, 0.2473755, 0.1737922, 0.1201212,
  0.2068923, 0.1275641, 0.1493386, 0.1350463, 0.2296917, 0.3509909, 0.260134, 
    0.1571737, 0.178416, 0.2113638, 0.1812886, 0.1077934, 0.1905397, 
    0.1378775, 0.1255463, 0.056555, 0.1216467, 0.2122322, 0.1113482, 
    0.1558961, 0.2019704, 0.2185202, 0.249228, 0.1201645, 0.08166525, 
    0.422319, 0.3134364, 0.1683574, 0.2624834,
  0.102064, 0.2163989, 0.2421812, 0.160171, 0.142591, 0.1259263, 0.1532827, 
    0.1710414, 0.1543163, 0.1659684, 0.1948809, 0.2087208, 0.1909257, 
    0.2906035, 0.3130494, 0.2642104, 0.2496322, 0.1892753, 0.1190728, 
    0.1367708, 0.2741086, 0.3254513, 0.4073549, 0.2326158, 0.2365949, 
    0.1813108, 0.1749172, 0.08850585, 0.07912882,
  0.1411746, 0.1400149, 0.1388552, 0.1376954, 0.1365357, 0.135376, 0.1342163, 
    0.1941987, 0.2055332, 0.2168677, 0.2282022, 0.2395368, 0.2508713, 
    0.2622058, 0.2521214, 0.2549853, 0.2578491, 0.260713, 0.2635768, 
    0.2664407, 0.2693045, 0.2432896, 0.2302509, 0.2172123, 0.2041736, 
    0.191135, 0.1780964, 0.1650577, 0.1421024,
  0.1092212, 0.09070639, 0.07870397, 0.02773273, 0.01787497, 0.08339926, 
    0.1107565, 0.08251177, 0.02241365, 0.00946724, 0.06504352, 0.1470666, 
    0.200003, 0.2026962, 0.166411, 0.1109839, 0.1178936, 0.129839, 0.1380012, 
    0.1257422, 0.2858934, 0.4065974, 0.4873575, 0.5355578, 0.3658411, 
    0.1354413, 0.2127934, 0.1326614, 0.1675218,
  0.2710937, 0.2656405, 0.2787902, 0.2782664, 0.3994306, 0.3429341, 
    0.3164304, 0.4142591, 0.3485357, 0.247441, 0.2218277, 0.1869578, 
    0.2346906, 0.2448836, 0.315447, 0.2888799, 0.2962092, 0.291939, 
    0.3109673, 0.305021, 0.3430066, 0.305539, 0.2098445, 0.3954052, 
    0.3209946, 0.2019507, 0.3339331, 0.4791216, 0.3443971,
  0.302479, 0.3605816, 0.3592252, 0.3269428, 0.3761897, 0.3285367, 0.3953064, 
    0.3025101, 0.3390278, 0.3981579, 0.3085631, 0.380342, 0.3546444, 
    0.3210849, 0.3242093, 0.3007485, 0.2924479, 0.1920272, 0.2443605, 
    0.3666455, 0.3319618, 0.2895563, 0.3542911, 0.2889443, 0.2126322, 
    0.3311913, 0.2894678, 0.2779846, 0.3322642,
  0.2593494, 0.2548028, 0.2830163, 0.2682206, 0.2557708, 0.2252877, 
    0.1898514, 0.3042519, 0.250047, 0.3192759, 0.2744513, 0.2424165, 
    0.2480038, 0.2911429, 0.3418589, 0.1935817, 0.2445963, 0.339518, 
    0.325541, 0.2454581, 0.2387709, 0.2211685, 0.2076623, 0.1626385, 
    0.1118781, 0.1761422, 0.2133681, 0.2433568, 0.2080569,
  0.3052821, 0.2586192, 0.2131201, 0.2232981, 0.280163, 0.19266, 0.1723624, 
    0.2177331, 0.2017725, 0.2347016, 0.2205039, 0.1933598, 0.1458227, 
    0.2194599, 0.2724293, 0.1796541, 0.2404003, 0.2127133, 0.2487151, 
    0.1941963, 0.1569761, 0.1733766, 0.207745, 0.2107521, 0.174557, 0.19227, 
    0.1857475, 0.203582, 0.1743544,
  0.1621488, 0.06838401, 0.06639074, 0.08372748, 0.04670717, 0.08634572, 
    0.07990663, 0.1180223, 0.06660179, 0.0860123, 0.01587478, 0.04595195, 
    0.01749719, 0.095634, 0.0893966, 0.1292049, 0.1260853, 0.1035402, 
    0.1155618, 0.2579725, 0.115339, 0.1081519, 0.09354674, 0.006340874, 
    0.08881249, 0.1411376, 0.08232448, 0.08325671, 0.124362,
  0.04608097, -2.526381e-05, 0.008430885, 0.006657115, 0.04249624, 
    0.06576001, 0.05109207, 0.1167439, 0.1177025, 0.03016794, 9.220674e-10, 
    4.227217e-05, 0.07857931, 0.09489682, 0.1822698, 0.03365601, 0.02643346, 
    0.09130152, 0.06119338, 0.08279107, 0.1124797, 0.06748136, 0.002179605, 
    1.327193e-07, 0.02567694, 0.04800368, 0.03791972, 0.06631058, 0.1064218,
  2.14121e-06, -4.209827e-05, 0.000882919, 0.1317696, 0.06451847, 0.05209043, 
    0.0406977, 0.04327783, 0.02154747, 0.03830076, 0.1226791, 0.08743446, 
    0.1042355, 0.03851761, 0.04611292, 0.02908428, 0.02187315, 0.007709846, 
    0.01076631, 0.006911473, 0.0005182839, 3.464706e-06, 6.767854e-08, 
    0.01308013, 0.006376951, 0.001339482, 0.05651979, 0.02031998, 0.001193729,
  0.001121528, 0.1077391, 0.06351095, 0.01218861, 0.01841459, 0.02096523, 
    0.04781543, 0.03644064, 0.05052447, 0.06350534, 0.0618602, 0.01150015, 
    0.04004348, 0.0285699, 0.04307491, 0.03088512, 0.04814152, 0.03990341, 
    0.02501092, 0.008121112, 0.001670293, 0.001522099, 0.01222336, 0.1982454, 
    0.162927, 0.03237461, 0.09260339, 0.03301673, 0.003899416,
  0.006880362, 0.001847483, 0.0006287154, 0.0008390447, 0.0003446375, 
    0.01085422, 0.05888547, 0.01432854, 0.0158578, 0.03833803, 0.02349594, 
    0.05994063, 0.04205089, 0.04498189, 0.05876362, 0.06196819, 0.04885351, 
    0.1090483, 0.1234135, 0.01569888, 0.06640267, 0.07835551, 0.1073028, 
    0.06989442, 0.03331866, 0.1027565, 0.09166722, 0.05823788, 0.05442683,
  2.662604e-06, 1.914147e-06, 4.074466e-07, 7.475377e-09, 8.956329e-09, 
    -4.028838e-06, 0.03479863, 0.01144457, 0.1538008, 0.1024474, 0.09311967, 
    0.06664598, 0.02496131, 0.02604347, 0.0346615, 0.02637011, 0.03838083, 
    0.02824184, 0.000741106, 1.864185e-07, 2.215234e-07, 0.0109495, 
    0.02052463, 0.01315174, 0.02327879, 0.04885305, 0.01300875, 5.576154e-07, 
    9.470869e-06,
  1.589342e-06, 4.783845e-06, 9.423765e-08, 1.375478e-06, 6.660098e-07, 
    4.479624e-08, -0.0002527238, 0.08534884, 0.3512244, 0.03061756, 
    0.1138382, 0.1508238, 0.07233246, 0.04224252, 0.09059939, 0.06900142, 
    0.1256141, 0.05664412, 0.02142175, 0.0002197389, 8.120119e-07, 
    0.002653931, 0.06607822, 0.03489432, 0.05103071, 0.05084421, 0.07202725, 
    0.02543347, -0.0001195707,
  0.01419859, 0.00695987, 0.00124973, 0.04218752, 0.001536713, 8.69382e-05, 
    0.05148259, 0.003428527, 3.956744e-05, 0.02277559, 0.3251629, 0.1136517, 
    0.1105758, 0.1248638, 0.149411, 0.2299769, 0.2280158, 0.0684427, 
    0.09732771, 0.06129194, 0.005165494, 0.01077659, 0.05427397, 0.06018566, 
    0.1101162, 0.1793736, 0.1026781, 0.1020326, 0.02937981,
  0.1950214, 0.2342254, 0.1436197, 0.08070779, 0.03893385, 0.02494589, 
    0.03029565, 0.1577837, 0.1139538, 0.07338403, 0.2918619, 0.2490748, 
    0.07856315, 0.1308086, 0.2860025, 0.4157248, 0.3005746, 0.242428, 
    0.1452813, 0.2381307, 0.06975785, 0.01533365, 0.06050495, 0.2018338, 
    0.1614956, 0.1904278, 0.1672169, 0.1689898, 0.1565715,
  0.1706506, 0.1491187, 0.1945345, 0.1370866, 0.2544542, 0.3157022, 
    0.2059332, 0.1526516, 0.1682075, 0.1102854, 0.1524432, 0.2136798, 
    0.1586673, 0.2391992, 0.3130227, 0.3165438, 0.3358034, 0.3821984, 
    0.1335683, 0.06915488, 0.1114899, 0.1529628, 0.1686853, 0.2519587, 
    0.1603337, 0.3157794, 0.2594511, 0.2353816, 0.1204831,
  0.1830175, 0.1043573, 0.1952458, 0.1571316, 0.2388291, 0.3104486, 
    0.2531326, 0.1402693, 0.1779913, 0.2806783, 0.2194106, 0.1456688, 
    0.1651442, 0.129509, 0.1664842, 0.09221508, 0.1628577, 0.1603195, 
    0.1311188, 0.1721964, 0.2110227, 0.20569, 0.2861592, 0.1685493, 
    0.09277325, 0.4516873, 0.3087805, 0.1709342, 0.3197281,
  0.1514169, 0.2351508, 0.2364045, 0.1380837, 0.1327839, 0.1671679, 
    0.1818471, 0.1775774, 0.2252778, 0.2129381, 0.2028772, 0.2002851, 
    0.1926184, 0.2551676, 0.2872095, 0.2642874, 0.2798181, 0.2297857, 
    0.2285078, 0.2326515, 0.3243597, 0.375857, 0.391295, 0.2558005, 
    0.2206164, 0.2391622, 0.1936547, 0.05015972, 0.1094132,
  0.1754344, 0.1767438, 0.1780531, 0.1793625, 0.1806718, 0.1819812, 
    0.1832905, 0.2570783, 0.2706865, 0.2842947, 0.2979029, 0.3115111, 
    0.3251193, 0.3387275, 0.3469419, 0.3465004, 0.3460589, 0.3456174, 
    0.3451759, 0.3447344, 0.3442928, 0.2797535, 0.2652774, 0.2508014, 
    0.2363253, 0.2218493, 0.2073732, 0.1928972, 0.1743869,
  0.1202212, 0.1171027, 0.1233073, 0.04676189, 0.03676148, 0.1375653, 
    0.1773102, 0.1338959, 0.01601792, 0.0407158, 0.07506795, 0.1616465, 
    0.2096689, 0.1990869, 0.1539664, 0.1346174, 0.1172158, 0.144609, 
    0.1543461, 0.1319167, 0.3445749, 0.4342953, 0.5747386, 0.5045014, 
    0.3832673, 0.1792045, 0.1947163, 0.11907, 0.1752697,
  0.2870125, 0.2867038, 0.2492503, 0.2316861, 0.3904304, 0.3419431, 
    0.2938331, 0.396685, 0.3441147, 0.2419353, 0.2206051, 0.1953889, 
    0.2451635, 0.2125976, 0.3609992, 0.2977495, 0.2798744, 0.2757857, 
    0.3083407, 0.3464085, 0.3381769, 0.3051069, 0.2207513, 0.382944, 
    0.347272, 0.2559416, 0.3522089, 0.5018623, 0.3441329,
  0.4280332, 0.3483935, 0.3850695, 0.361621, 0.4147016, 0.3686183, 0.5173806, 
    0.4160855, 0.4590869, 0.4777992, 0.4827805, 0.4938625, 0.4418077, 
    0.3498044, 0.4116452, 0.341676, 0.3419316, 0.2128179, 0.3949105, 
    0.3886579, 0.3008213, 0.2337274, 0.3262614, 0.3359544, 0.3153758, 
    0.3633225, 0.3438409, 0.3332274, 0.3915349,
  0.2777312, 0.2058452, 0.3047207, 0.2643983, 0.2331071, 0.2139741, 
    0.2201418, 0.2802258, 0.2404916, 0.2794128, 0.2926653, 0.3203321, 
    0.2738807, 0.3482152, 0.3565743, 0.2969435, 0.3067522, 0.4086039, 
    0.3445892, 0.2849054, 0.2701415, 0.2369367, 0.2591416, 0.2120692, 
    0.140749, 0.1868661, 0.2276776, 0.3288965, 0.316692,
  0.2739807, 0.2644855, 0.1721157, 0.2352994, 0.2705841, 0.1915907, 
    0.1533729, 0.201795, 0.1904376, 0.2423023, 0.2023938, 0.1721017, 
    0.1373198, 0.1963622, 0.2866565, 0.1853808, 0.2148557, 0.2478977, 
    0.2900874, 0.2278277, 0.170576, 0.1762961, 0.1886767, 0.2262966, 
    0.2497821, 0.1817148, 0.1905454, 0.3152785, 0.230688,
  0.1373896, 0.111538, 0.04282613, 0.07779845, 0.08941615, 0.1460377, 
    0.1285191, 0.1720315, 0.1351933, 0.1193244, 0.01221202, 0.02446853, 
    0.01323393, 0.09972943, 0.1315493, 0.1143604, 0.1134143, 0.104173, 
    0.1278812, 0.2548434, 0.09223001, 0.1370934, 0.1321844, 0.006492281, 
    0.09454633, 0.1486066, 0.1056292, 0.1156677, 0.1222085,
  0.1975163, -0.0002271394, 0.001101093, 0.0280451, 0.050288, 0.0596146, 
    0.05209737, 0.1301909, 0.1226918, 0.02316443, 1.932358e-10, 1.858583e-06, 
    0.1280797, 0.1739364, 0.1818216, 0.05765642, 0.07046562, 0.1035066, 
    0.1011198, 0.07570191, 0.1085517, 0.1074177, 0.01856956, -1.205208e-07, 
    0.04167211, 0.05097091, 0.05883105, 0.1185602, 0.2694218,
  0.000752219, -7.766424e-06, 0.002632213, 0.1060978, 0.05977704, 0.046376, 
    0.04601504, 0.04015036, 0.02557032, 0.05032671, 0.1569149, 0.0836597, 
    0.1056382, 0.03684139, 0.03969742, 0.0310103, 0.03155995, 0.0103546, 
    0.01648104, 0.0315165, 0.01981846, 0.002766526, 5.850841e-07, 0.02390669, 
    0.004775713, 5.321283e-05, 0.06272744, 0.04154821, 0.03051027,
  0.005588041, 0.1201057, 0.05724854, 0.01111997, 0.02689455, 0.02610721, 
    0.04153894, 0.03556102, 0.05590186, 0.08490498, 0.04591071, 0.01500039, 
    0.02788582, 0.02731203, 0.03525855, 0.02380881, 0.03663737, 0.02995332, 
    0.01995293, 0.01170071, 0.01154596, 0.005027262, 0.008303586, 0.1934505, 
    0.1691512, 0.03029059, 0.07720621, 0.03364552, 0.01698361,
  0.006038126, 0.0009733833, 0.0002623209, 0.0001606882, 0.0001895166, 
    0.01530344, 0.05225741, 0.0151321, 0.01227424, 0.02968659, 0.02111696, 
    0.05229031, 0.03432086, 0.03947498, 0.0567401, 0.05714893, 0.05450987, 
    0.1084681, 0.1273657, 0.02696434, 0.07214507, 0.07297612, 0.1205261, 
    0.0588995, 0.02999653, 0.1024085, 0.1031008, 0.0612229, 0.04534917,
  1.982514e-06, 1.610894e-06, 1.956444e-07, 4.833409e-09, 7.99694e-09, 
    -8.320383e-05, 0.02710648, 0.01018141, 0.1583653, 0.09073232, 0.07193093, 
    0.05882496, 0.02757645, 0.02788618, 0.03317046, 0.02581886, 0.03858204, 
    0.09798373, 0.03366971, 0.0003319016, 7.651229e-08, 0.01706431, 
    0.02643781, 0.007903989, 0.03111368, 0.0732341, 0.06116167, 4.353068e-07, 
    7.8304e-06,
  1.029433e-06, 3.296256e-06, 3.663117e-08, 1.193675e-06, 5.895317e-07, 
    3.506098e-08, -0.0001413604, 0.06285068, 0.3738606, 0.0272311, 0.1069636, 
    0.157571, 0.0685464, 0.05306413, 0.1116856, 0.09837825, 0.1559482, 
    0.07844176, 0.08058395, 0.002028157, 5.237781e-07, 0.003218023, 
    0.07561073, 0.03895786, 0.03944386, 0.04912124, 0.09875773, 0.05875241, 
    -0.0002572846,
  0.00754378, 0.005804056, 0.0004525498, 0.04350265, -0.0003279154, 
    7.503083e-07, 0.04421467, 0.00149452, -3.337704e-05, 0.02521843, 
    0.3288833, 0.1442032, 0.1333731, 0.1453347, 0.2303144, 0.2694001, 
    0.250746, 0.0854262, 0.1492507, 0.06395701, 0.005351977, 0.01988062, 
    0.0488103, 0.05921631, 0.11757, 0.206954, 0.132311, 0.1393784, 0.0518401,
  0.2050386, 0.2165931, 0.1341469, 0.02360389, 0.01817903, 0.0141619, 
    0.02471031, 0.1400202, 0.1119155, 0.06039895, 0.2691137, 0.2514014, 
    0.08323883, 0.1402591, 0.3313693, 0.4807033, 0.3695763, 0.2730014, 
    0.1573901, 0.225058, 0.05898852, 0.01122262, 0.04451982, 0.204905, 
    0.1572334, 0.1926017, 0.2255201, 0.2124385, 0.1260276,
  0.1696943, 0.108202, 0.1195317, 0.1109049, 0.22251, 0.2741372, 0.1824868, 
    0.1681498, 0.1369832, 0.09379236, 0.118981, 0.2089963, 0.1529823, 
    0.2280945, 0.3787969, 0.3298752, 0.3136614, 0.4022842, 0.1583976, 
    0.04620135, 0.08516096, 0.1376914, 0.1472545, 0.234865, 0.185648, 
    0.2791171, 0.3236291, 0.3000598, 0.2129809,
  0.2516929, 0.1613613, 0.2551609, 0.23812, 0.277037, 0.2682954, 0.225745, 
    0.1629937, 0.1829391, 0.2485011, 0.2293755, 0.1227954, 0.1430578, 
    0.1445622, 0.2183007, 0.1751359, 0.178477, 0.1791551, 0.1236068, 
    0.2228215, 0.2106605, 0.2422809, 0.2776356, 0.217169, 0.1149281, 
    0.4584281, 0.297426, 0.1642637, 0.3368,
  0.1983068, 0.2722601, 0.2731971, 0.1639696, 0.1621854, 0.2676493, 
    0.2435529, 0.2629583, 0.3902363, 0.3222352, 0.1934635, 0.2507217, 
    0.2146997, 0.236394, 0.3001224, 0.2989334, 0.3328216, 0.3779605, 
    0.2330021, 0.3038103, 0.3801328, 0.4044448, 0.3692864, 0.2734677, 
    0.2496295, 0.2690938, 0.1887988, 0.05480887, 0.1384468,
  0.1895771, 0.1931944, 0.1968118, 0.2004292, 0.2040465, 0.2076639, 
    0.2112812, 0.3061634, 0.3213109, 0.3364584, 0.3516059, 0.3667534, 
    0.3819009, 0.3970484, 0.4062448, 0.40234, 0.3984352, 0.3945305, 
    0.3906257, 0.386721, 0.3828162, 0.2974379, 0.2825778, 0.2677177, 
    0.2528577, 0.2379976, 0.2231375, 0.2082774, 0.1866832,
  0.1233328, 0.1466324, 0.1561703, 0.1040387, 0.05439635, 0.1936619, 
    0.1971588, 0.1842649, 0.01542061, 0.0447925, 0.08180118, 0.1663744, 
    0.2223108, 0.1658676, 0.1545056, 0.1383399, 0.1135853, 0.1472543, 
    0.1505588, 0.1507812, 0.3595549, 0.4428646, 0.6288491, 0.4701809, 
    0.3839136, 0.2076581, 0.1554919, 0.09333852, 0.1763998,
  0.3184813, 0.2730508, 0.2400982, 0.1967756, 0.401685, 0.3244646, 0.2432081, 
    0.370546, 0.3440843, 0.2525832, 0.2320096, 0.2056797, 0.2518054, 
    0.2033353, 0.3471163, 0.3387839, 0.2995722, 0.3325507, 0.3255494, 
    0.3889156, 0.3239138, 0.3094072, 0.2466869, 0.3810586, 0.3482626, 
    0.3100743, 0.3977443, 0.5306737, 0.3464204,
  0.466173, 0.2694372, 0.3599477, 0.3699591, 0.4259132, 0.4254725, 0.5870388, 
    0.4699312, 0.5658818, 0.574136, 0.5516154, 0.5637863, 0.4044585, 
    0.4531085, 0.4349862, 0.3621472, 0.3795705, 0.3459999, 0.4312484, 
    0.3629039, 0.2688828, 0.2013365, 0.3176773, 0.3529356, 0.3343315, 
    0.4367427, 0.4325552, 0.4108693, 0.4329676,
  0.3117671, 0.2554054, 0.3161395, 0.2096618, 0.2288375, 0.1837322, 
    0.1936684, 0.2384467, 0.2736465, 0.2543694, 0.3005933, 0.3062407, 
    0.2563461, 0.3175522, 0.3422074, 0.432045, 0.3549273, 0.4290676, 
    0.4227598, 0.2976428, 0.2811767, 0.2278481, 0.2565499, 0.2450647, 
    0.1572038, 0.2071629, 0.4274181, 0.3663688, 0.3513536,
  0.214088, 0.2052002, 0.1197942, 0.200289, 0.2149525, 0.187144, 0.1663373, 
    0.2446, 0.2194307, 0.2372549, 0.1891727, 0.1756747, 0.1065894, 0.1576232, 
    0.330424, 0.1589472, 0.2222283, 0.246093, 0.259586, 0.1877116, 0.1862306, 
    0.1993392, 0.1979471, 0.2637764, 0.2425952, 0.1791686, 0.2633476, 
    0.3052906, 0.2516251,
  0.1748975, 0.07297578, 0.02846446, 0.111333, 0.1055925, 0.1342067, 
    0.1467968, 0.2241879, 0.1510853, 0.1235142, 0.003442038, 0.0160749, 
    0.0119999, 0.05922586, 0.1386664, 0.06966933, 0.08965421, 0.0862923, 
    0.1440185, 0.2473443, 0.121529, 0.09998025, 0.1142927, 0.008794255, 
    0.1170933, 0.1495635, 0.1059355, 0.1355945, 0.1281262,
  0.223924, -0.0002854905, 0.000384461, 0.03043164, 0.06507545, 0.07630769, 
    0.0763982, 0.108023, 0.1305673, 0.003005354, 3.184341e-11, 1.849253e-07, 
    0.07113855, 0.2160045, 0.189558, 0.07080988, 0.07142654, 0.1531727, 
    0.08628061, 0.07155746, 0.1301252, 0.1854829, 0.1665254, -1.350485e-06, 
    0.04928604, 0.08280417, 0.06782172, 0.1640786, 0.2584664,
  0.05814337, 1.205513e-06, 0.001616329, 0.06920605, 0.05115991, 0.04747675, 
    0.07991516, 0.07225452, 0.0732728, 0.08556, 0.1358107, 0.09435973, 
    0.1167962, 0.04214476, 0.05040117, 0.06529988, 0.04210273, 0.03044422, 
    0.04626177, 0.09657168, 0.1556207, 0.08192345, 8.46136e-06, 0.05958434, 
    0.002778911, 4.71518e-06, 0.1007779, 0.08389072, 0.1595935,
  0.02792997, 0.1032873, 0.03929154, 0.01659733, 0.03989879, 0.06753573, 
    0.04176014, 0.0397035, 0.04697576, 0.1131428, 0.0490353, 0.02156552, 
    0.02647766, 0.03229502, 0.03064029, 0.02335109, 0.02956949, 0.02392318, 
    0.02124609, 0.01283834, 0.0195071, 0.03404154, 0.0004804358, 0.1995936, 
    0.1524743, 0.03316602, 0.06941208, 0.04078226, 0.0311189,
  0.003970796, 0.0006603586, 0.0001135127, -3.555354e-05, 7.395011e-05, 
    0.02609398, 0.04848022, 0.02316153, 0.008561688, 0.02734083, 0.02185177, 
    0.04694572, 0.03429452, 0.03994624, 0.05455539, 0.0526287, 0.05970101, 
    0.1104672, 0.119064, 0.03984181, 0.06711765, 0.06923481, 0.1092252, 
    0.04077207, 0.03380198, 0.0896772, 0.1200991, 0.0784777, 0.03435048,
  1.55721e-06, 1.381501e-06, 9.528726e-08, 4.063731e-09, 8.559712e-09, 
    0.0005323233, 0.01801034, 0.01050286, 0.1608803, 0.08494885, 0.0582513, 
    0.0633945, 0.03831437, 0.04980309, 0.0490309, 0.03407129, 0.03873967, 
    0.1081385, 0.1249971, 0.01723233, -1.450404e-06, 0.02225226, 0.0338443, 
    0.005251042, 0.03838405, 0.07010783, 0.1350603, -9.863817e-06, 
    2.843742e-06,
  7.18709e-07, 2.595732e-06, 2.421145e-08, 1.060533e-06, 5.113734e-07, 
    3.214377e-08, -0.0001149487, 0.06389439, 0.3740218, 0.02471427, 
    0.1187977, 0.1716417, 0.09300122, 0.08745527, 0.1577664, 0.1460164, 
    0.2345075, 0.1128845, 0.2114152, 0.06368183, 2.932398e-07, 0.006374214, 
    0.06567296, 0.04627109, 0.07045022, 0.0849157, 0.1204843, 0.09508041, 
    4.986658e-05,
  0.003173183, 0.004478656, 0.000153463, 0.04756044, -0.0005219112, 
    -4.855524e-05, 0.04082456, 0.0003672866, -4.329887e-05, 0.01014934, 
    0.3382839, 0.1826956, 0.1885314, 0.1985255, 0.3905435, 0.3187854, 
    0.2759439, 0.1179095, 0.2043995, 0.06430683, 0.006543284, 0.02684453, 
    0.02985041, 0.04830127, 0.1321857, 0.2454094, 0.1962402, 0.2542355, 
    0.1098284,
  0.2051683, 0.2166119, 0.1292195, 0.007105665, 0.003276716, 0.01124405, 
    0.03161358, 0.1378499, 0.1062162, 0.0397989, 0.23264, 0.2503788, 
    0.1171106, 0.1823735, 0.4324856, 0.5483959, 0.4145997, 0.2626849, 
    0.1795663, 0.2033272, 0.04077023, 0.009369478, 0.02884881, 0.2199791, 
    0.1564616, 0.1917394, 0.257645, 0.2516139, 0.1222684,
  0.1452028, 0.09120344, 0.09721918, 0.07429387, 0.1888861, 0.2146264, 
    0.1396174, 0.1271389, 0.1220362, 0.05522045, 0.09336276, 0.1682107, 
    0.1377147, 0.2051993, 0.3406709, 0.3113235, 0.3305826, 0.3890631, 
    0.1524703, 0.02626697, 0.05510718, 0.1192875, 0.1383967, 0.2219855, 
    0.2059778, 0.2414545, 0.4195088, 0.361111, 0.1879089,
  0.2334772, 0.2141043, 0.3000036, 0.2766975, 0.2717987, 0.3407617, 
    0.2577049, 0.1496431, 0.1724635, 0.211826, 0.184626, 0.1219342, 
    0.1300534, 0.1529837, 0.2304302, 0.1588347, 0.2027269, 0.2065542, 
    0.09795848, 0.2538162, 0.2411806, 0.2623758, 0.2570246, 0.2475897, 
    0.1800767, 0.400997, 0.293259, 0.1581997, 0.3124628,
  0.2400448, 0.3491526, 0.3464862, 0.2489279, 0.3418907, 0.3778504, 
    0.3836325, 0.2971166, 0.3887495, 0.3624586, 0.3204822, 0.2752138, 
    0.3856125, 0.3367467, 0.3436057, 0.3230545, 0.371794, 0.3871475, 
    0.3003547, 0.3537561, 0.4444357, 0.4123688, 0.3343282, 0.294329, 
    0.3243567, 0.301021, 0.2024637, 0.08610633, 0.1872059,
  0.2042726, 0.2089887, 0.2137048, 0.2184209, 0.223137, 0.2278531, 0.2325692, 
    0.3185329, 0.3334352, 0.3483376, 0.3632399, 0.3781423, 0.3930446, 
    0.407947, 0.4268204, 0.4205335, 0.4142467, 0.4079599, 0.401673, 
    0.3953862, 0.3890994, 0.3006705, 0.2873389, 0.2740072, 0.2606756, 
    0.247344, 0.2340123, 0.2206807, 0.2004997,
  0.1450891, 0.1761244, 0.1915476, 0.1166482, 0.09962692, 0.2305968, 
    0.2204935, 0.201605, 0.01726659, 0.04934052, 0.08890676, 0.1562986, 
    0.2211185, 0.1170043, 0.1485933, 0.1420733, 0.133343, 0.1552688, 
    0.1385108, 0.1529962, 0.3381466, 0.4200128, 0.6154049, 0.4298816, 
    0.3368471, 0.2159481, 0.112617, 0.06235851, 0.1869854,
  0.3174059, 0.2248269, 0.2415239, 0.1334981, 0.3990258, 0.3087982, 
    0.1714106, 0.3613268, 0.3208266, 0.2543066, 0.230451, 0.203542, 
    0.2684447, 0.2099807, 0.3436518, 0.3915813, 0.3584491, 0.3675252, 
    0.3214633, 0.3937016, 0.369044, 0.3522548, 0.2159356, 0.3738192, 
    0.3567988, 0.3283088, 0.4941024, 0.4827293, 0.3643487,
  0.4895643, 0.2253673, 0.2958619, 0.2902144, 0.3367688, 0.3875818, 
    0.4871825, 0.4419692, 0.5101134, 0.5105162, 0.4517374, 0.5435038, 
    0.4018668, 0.4375973, 0.3827883, 0.3545472, 0.3977447, 0.4631857, 
    0.3574792, 0.3083369, 0.2643327, 0.1904029, 0.3116855, 0.3264645, 
    0.3027406, 0.4876173, 0.4872749, 0.4799557, 0.5202631,
  0.3088415, 0.2811044, 0.2733514, 0.1841279, 0.1907855, 0.1675579, 
    0.1787759, 0.1938395, 0.2633543, 0.282593, 0.2402686, 0.2405954, 
    0.2302627, 0.2287504, 0.3495915, 0.2903045, 0.3829444, 0.4730142, 
    0.4312113, 0.284029, 0.3053477, 0.2189036, 0.2099807, 0.2522708, 
    0.1664942, 0.28835, 0.4133879, 0.3159028, 0.2666497,
  0.1635313, 0.1312573, 0.05787729, 0.1291893, 0.183871, 0.1854783, 
    0.2389538, 0.2776407, 0.2551906, 0.2285169, 0.168334, 0.1068903, 
    0.06373022, 0.1531941, 0.4111941, 0.1112256, 0.1863186, 0.2306855, 
    0.233034, 0.1719908, 0.1327433, 0.175156, 0.2690314, 0.3109249, 
    0.1820148, 0.1627591, 0.2613425, 0.2460763, 0.1883861,
  0.1612035, 0.06107927, 0.02183949, 0.08999295, 0.09293447, 0.1012046, 
    0.1093368, 0.1507734, 0.1102788, 0.07356469, 0.0009651756, 0.005824686, 
    0.009688948, 0.03677267, 0.06449484, 0.05075482, 0.07823344, 0.08739199, 
    0.1218368, 0.1765501, 0.1081179, 0.07131578, 0.1494792, 0.02190362, 
    0.0747841, 0.09483475, 0.07633886, 0.1032325, 0.1305972,
  0.2068033, 0.0156721, 0.0001193703, 0.1333451, 0.06231928, 0.02605177, 
    0.03195497, 0.06903691, 0.1152517, 0.0005117728, 8.682186e-12, 
    5.3145e-08, 0.03448028, 0.1427664, 0.1664527, 0.08809139, 0.1353973, 
    0.1245234, 0.07214489, 0.04670828, 0.09984359, 0.1667511, 0.4116165, 
    -9.478748e-06, 0.07361095, 0.05920363, 0.07693344, 0.08471545, 0.1200873,
  0.413608, 0.0002329168, 0.00130339, 0.04768742, 0.05383955, 0.05453653, 
    0.04748639, 0.1145044, 0.04643543, 0.04640877, 0.07073352, 0.0859063, 
    0.1176619, 0.05484899, 0.06050375, 0.09181663, 0.05385135, 0.1072688, 
    0.06586181, 0.09316415, 0.1412075, 0.4287217, -2.207448e-05, 0.06712984, 
    0.0005797757, -9.463674e-06, 0.0677037, 0.04943791, 0.2918147,
  0.08662749, 0.08536089, 0.01629174, 0.02668871, 0.08840051, 0.05356138, 
    0.09074122, 0.0587238, 0.02958165, 0.0984213, 0.08501562, 0.042415, 
    0.06431238, 0.04163706, 0.03102772, 0.03155592, 0.03179407, 0.02265288, 
    0.03664769, 0.02199153, 0.03371001, 0.09272711, 0.004484734, 0.16946, 
    0.1136655, 0.04712974, 0.08569243, 0.1020888, 0.04956338,
  0.00151417, 0.0005166779, 4.586151e-05, -4.892068e-05, 1.892866e-06, 
    0.03049566, 0.04498718, 0.02536967, 0.006289376, 0.02846498, 0.02249063, 
    0.05122688, 0.04215678, 0.04365679, 0.05329107, 0.06246109, 0.06079447, 
    0.1396678, 0.1260495, 0.1574681, 0.09218726, 0.07168576, 0.1028347, 
    0.03787034, 0.06893708, 0.1052881, 0.1679159, 0.08533935, 0.02302661,
  1.30285e-06, 1.26278e-06, 5.816266e-08, 3.207397e-09, 7.644253e-09, 
    0.01257282, 0.01029545, 0.01094524, 0.1203853, 0.08379917, 0.06120386, 
    0.06450508, 0.03239236, 0.04466676, 0.06910662, 0.06424628, 0.06354858, 
    0.1157037, 0.2674213, 0.03125357, -1.523588e-05, 0.0345966, 0.05151088, 
    0.01149116, 0.04544132, 0.06508757, 0.202102, 0.001188375, 2.772578e-06,
  6.011628e-07, 2.214156e-06, 1.630593e-08, 9.599325e-07, 4.396801e-07, 
    3.081114e-08, -3.330942e-05, 0.06819173, 0.360062, 0.02442843, 0.2013924, 
    0.2018251, 0.1018854, 0.1492415, 0.2188293, 0.1413818, 0.2172226, 
    0.1584375, 0.329006, 0.1421091, 1.836424e-07, 0.01436895, 0.04717034, 
    0.06913217, 0.05912196, 0.179619, 0.1190164, 0.2835456, -0.0005488262,
  4.243774e-05, 0.002466794, 8.589526e-05, 0.06269367, -0.0005397452, 
    -1.436368e-05, 0.03375724, 0.0001477525, -5.217087e-05, 0.005152609, 
    0.3238018, 0.195516, 0.2614202, 0.3909091, 0.546818, 0.43811, 0.336513, 
    0.2320387, 0.358743, 0.06361161, 0.00742352, 0.04909019, 0.02568947, 
    0.05499429, 0.1758848, 0.2633992, 0.2606986, 0.4058065, 0.1431155,
  0.1802539, 0.1802862, 0.1225071, 0.001797586, 0.002782901, 0.008027699, 
    0.02991571, 0.1365181, 0.09285787, 0.03184336, 0.1926184, 0.2030029, 
    0.1717845, 0.1802448, 0.3942861, 0.5782016, 0.4288615, 0.2986268, 
    0.2290428, 0.1710161, 0.02992246, 0.007918377, 0.02928952, 0.193519, 
    0.1401453, 0.2307513, 0.291669, 0.3227847, 0.1579901,
  0.1404785, 0.07066515, 0.07886296, 0.05449704, 0.160313, 0.1382383, 
    0.1184644, 0.09731583, 0.103218, 0.04281064, 0.05699576, 0.1433381, 
    0.1267671, 0.1643299, 0.3599657, 0.4460401, 0.3107858, 0.3381003, 
    0.1160732, 0.01403651, 0.02833252, 0.1001102, 0.1260965, 0.204408, 
    0.2166434, 0.2258818, 0.459798, 0.4022327, 0.2680401,
  0.1984624, 0.236152, 0.4026622, 0.3397619, 0.2755157, 0.3503681, 0.2811738, 
    0.1827707, 0.1623302, 0.2155513, 0.1712098, 0.1382321, 0.1295148, 
    0.1384854, 0.2600407, 0.1683193, 0.2321193, 0.2022656, 0.08750501, 
    0.2959944, 0.3137378, 0.3881599, 0.2587497, 0.3377616, 0.1486988, 
    0.4009122, 0.285018, 0.1600893, 0.3253063,
  0.2629067, 0.4518628, 0.4133481, 0.3844329, 0.4877756, 0.4860838, 
    0.4440095, 0.430101, 0.397018, 0.3660693, 0.3966593, 0.37257, 0.3954536, 
    0.3602293, 0.3641214, 0.3767853, 0.443502, 0.3740228, 0.3472761, 
    0.4444765, 0.5256665, 0.4117961, 0.2963001, 0.3734846, 0.3289063, 
    0.3292763, 0.1671381, 0.08454943, 0.1882003,
  0.2365253, 0.2409665, 0.2454076, 0.2498487, 0.2542898, 0.2587309, 0.263172, 
    0.3210989, 0.335615, 0.350131, 0.3646471, 0.3791631, 0.3936791, 
    0.4081952, 0.4305876, 0.4218192, 0.4130507, 0.4042822, 0.3955137, 
    0.3867452, 0.3779767, 0.2961265, 0.2859378, 0.2757492, 0.2655605, 
    0.2553719, 0.2451832, 0.2349945, 0.2329725,
  0.1425191, 0.216225, 0.2149035, 0.1319423, 0.1234646, 0.2520701, 0.2503372, 
    0.2362856, 0.01235223, 0.03784836, 0.09958936, 0.1438767, 0.2275197, 
    0.06242814, 0.165246, 0.1647716, 0.1690755, 0.1526522, 0.1408863, 
    0.1457829, 0.3184812, 0.3775223, 0.5702679, 0.3799106, 0.3069043, 
    0.2066076, 0.0510488, 0.05222273, 0.1857516,
  0.3136883, 0.1873664, 0.2015227, 0.09109654, 0.3524534, 0.2891621, 
    0.1002243, 0.3407575, 0.2991611, 0.2470369, 0.2386637, 0.2064836, 
    0.2648214, 0.2090582, 0.3335532, 0.4163386, 0.4212569, 0.3831561, 
    0.3607973, 0.3742201, 0.4085212, 0.4068922, 0.1982286, 0.3742847, 
    0.3715691, 0.3539522, 0.5697535, 0.493478, 0.4097926,
  0.4596789, 0.2127502, 0.2168516, 0.2433004, 0.2374031, 0.2647251, 
    0.4016847, 0.3463811, 0.4138221, 0.3971537, 0.3924436, 0.4801309, 
    0.3850004, 0.3307905, 0.3780538, 0.3543821, 0.3933227, 0.3603613, 
    0.3241961, 0.2727958, 0.2390094, 0.1578527, 0.2672409, 0.2900213, 
    0.3220839, 0.5060484, 0.5164316, 0.5265386, 0.5731994,
  0.2506828, 0.2382192, 0.2363434, 0.175131, 0.1696527, 0.1665689, 0.1324954, 
    0.1744203, 0.23359, 0.2730083, 0.1960621, 0.211487, 0.1871063, 0.2055237, 
    0.3135247, 0.2020269, 0.3862235, 0.4395498, 0.4232066, 0.2725598, 
    0.2582771, 0.2349623, 0.1947315, 0.2390821, 0.1450771, 0.2841471, 
    0.3958057, 0.3119293, 0.2344883,
  0.1625946, 0.09476592, 0.03414937, 0.08435921, 0.1592041, 0.1741911, 
    0.2307536, 0.2545462, 0.257172, 0.1884587, 0.1367125, 0.07567906, 
    0.02924899, 0.1300809, 0.4413892, 0.09150033, 0.1569488, 0.2119222, 
    0.2145068, 0.1487551, 0.1542537, 0.1354571, 0.1698401, 0.3255528, 
    0.1299109, 0.1080058, 0.1676961, 0.1740463, 0.1226995,
  0.0783092, 0.04651202, 0.01346171, 0.07666533, 0.1023915, 0.07683294, 
    0.04705207, 0.08547018, 0.06834175, 0.01954068, 0.0004239534, 
    0.001080292, 0.01093085, 0.02444397, 0.04510043, 0.0435965, 0.07270437, 
    0.09239078, 0.1285219, 0.1063831, 0.04931955, 0.04204303, 0.1140759, 
    0.03143113, 0.05348444, 0.07117285, 0.03884564, 0.06876664, 0.07974429,
  0.1177385, 0.02290764, -5.921607e-05, 0.1481044, 0.02347482, 0.004701525, 
    0.01561877, 0.06454979, 0.03659328, 0.000198068, 4.154014e-12, 
    1.858114e-09, 0.02039853, 0.09463286, 0.09987865, 0.08863446, 0.1295337, 
    0.1370786, 0.02703501, 0.01225151, 0.04086316, 0.07174651, 0.3065361, 
    -0.0004293736, 0.09930822, 0.03271485, 0.03657905, 0.02753428, 0.03865238,
  0.4400539, 0.01151673, 0.0002375187, 0.06249363, 0.03777923, 0.01913085, 
    0.01802629, 0.06161637, 0.007739777, 0.005706717, 0.03965188, 0.02053737, 
    0.09997868, 0.04874504, 0.03213703, 0.01996038, 0.01388452, 0.02555708, 
    0.0261891, 0.01667498, 0.03487987, 0.1556493, 0.2461243, 0.01565341, 
    3.828399e-05, -1.522672e-06, 0.007760173, 0.007253022, 0.09820744,
  0.3045032, 0.05733247, 0.005843489, 0.03119326, 0.07301395, 0.01923782, 
    0.03300577, 0.03362551, 0.0311394, 0.05431723, 0.02933587, 0.04125408, 
    0.03286541, 0.02069142, 0.03012212, 0.01762534, 0.03592561, 0.02357783, 
    0.01968181, 0.03000787, 0.1076645, 0.229024, 0.0502358, 0.1123275, 
    0.06523939, 0.03487997, 0.04844327, 0.06336948, 0.1029442,
  0.0006553441, 0.0004198973, 1.733169e-05, -1.225679e-05, 3.275033e-06, 
    0.007246761, 0.03933568, 0.006485313, 0.001326546, 0.01867533, 
    0.02129412, 0.06566407, 0.03018823, 0.02191523, 0.0393731, 0.0431634, 
    0.04192278, 0.09680115, 0.08593512, 0.1916117, 0.1608992, 0.1010761, 
    0.1042691, 0.02410243, 0.06746224, 0.08304762, 0.1651274, 0.2194996, 
    0.0153516,
  1.148898e-06, 1.171265e-06, 4.664682e-08, 2.721358e-09, 7.122238e-09, 
    0.2271453, 0.00733381, 0.01002353, 0.103106, 0.08910223, 0.07626494, 
    0.045881, 0.008265074, 0.01050217, 0.04090845, 0.1045187, 0.02487211, 
    0.07403649, 0.2345928, 0.3823929, 0.0007464391, 0.04564857, 0.03488972, 
    0.001536262, 0.01420143, 0.01482817, 0.05846243, 0.2030916, 2.855513e-07,
  5.566455e-07, 1.985932e-06, 1.142725e-08, 8.927707e-07, 3.893518e-07, 
    3.004919e-08, -1.438848e-05, 0.07584102, 0.346031, 0.02583124, 0.2115581, 
    0.2972217, 0.1341246, 0.1772887, 0.2714234, 0.1701304, 0.1894084, 
    0.07954765, 0.2091466, 0.1508465, 1.445042e-07, 0.02302109, 0.04196697, 
    0.09337522, 0.06607276, 0.05564784, 0.05185697, 0.2023013, 0.004286696,
  -0.00109112, 0.001820222, 4.772263e-05, 0.08058947, 0.0008275307, 
    -4.267749e-06, 0.02627195, 3.211505e-05, -4.47981e-05, 0.0018432, 
    0.3019612, 0.2518769, 0.4345347, 0.5916748, 0.5212927, 0.3894653, 
    0.3904971, 0.4526917, 0.3399944, 0.05284125, 0.007700949, 0.04105759, 
    0.01979162, 0.03487311, 0.248184, 0.2678359, 0.209609, 0.3372071, 
    0.1533007,
  0.1688296, 0.1469702, 0.1164184, 0.0001426825, 0.007594326, 0.005423446, 
    0.02313869, 0.1388153, 0.08825514, 0.03654143, 0.1703887, 0.1794745, 
    0.371072, 0.26727, 0.4674626, 0.6368868, 0.4618717, 0.367916, 0.2881167, 
    0.1567788, 0.02357147, 0.01351551, 0.02504628, 0.1746229, 0.133791, 
    0.2452269, 0.3219194, 0.4172354, 0.1539543,
  0.1553987, 0.05652599, 0.0658152, 0.04784576, 0.107131, 0.08246177, 
    0.09064569, 0.06995559, 0.08534595, 0.03369644, 0.03962544, 0.1381865, 
    0.1140185, 0.1322227, 0.3805712, 0.4585578, 0.2854787, 0.3276146, 
    0.1112548, 0.008186348, 0.01894244, 0.0857277, 0.1162489, 0.1988093, 
    0.2769935, 0.2541839, 0.5282601, 0.3977788, 0.2187479,
  0.2817008, 0.3577886, 0.3759144, 0.4327276, 0.2848973, 0.3233947, 
    0.2507725, 0.1759323, 0.1287679, 0.1818368, 0.1472353, 0.1022204, 
    0.0863702, 0.1182221, 0.2529528, 0.1856732, 0.1783013, 0.2275473, 
    0.1906856, 0.2792397, 0.4704728, 0.5125327, 0.2062477, 0.3867039, 
    0.1057041, 0.4106168, 0.2698475, 0.1660056, 0.3462541,
  0.3695028, 0.5301396, 0.4487988, 0.449558, 0.5238662, 0.5174123, 0.4817831, 
    0.5039585, 0.5287849, 0.4890264, 0.3783997, 0.4371587, 0.435876, 
    0.457891, 0.4187365, 0.4401753, 0.4607263, 0.352772, 0.412502, 0.5223194, 
    0.5043918, 0.4133394, 0.2840298, 0.3625837, 0.2979293, 0.2657085, 
    0.1253721, 0.1129256, 0.4027112,
  0.2447793, 0.2482699, 0.2517605, 0.255251, 0.2587416, 0.2622321, 0.2657227, 
    0.3108236, 0.3259882, 0.3411528, 0.3563174, 0.371482, 0.3866466, 
    0.4018112, 0.4199027, 0.4102513, 0.4006, 0.3909486, 0.3812972, 0.3716459, 
    0.3619945, 0.2988719, 0.2898681, 0.2808644, 0.2718606, 0.2628568, 
    0.253853, 0.2448492, 0.2419869,
  0.121621, 0.2582647, 0.1880969, 0.1422658, 0.1343677, 0.2418953, 0.2660447, 
    0.2421696, 0.01639672, 0.0340244, 0.09619115, 0.1358776, 0.2206935, 
    0.0348452, 0.1787101, 0.1749964, 0.1994592, 0.1435199, 0.1427945, 
    0.1390383, 0.3092424, 0.3726681, 0.517303, 0.3417265, 0.2644976, 
    0.1982534, 0.03670898, 0.0689749, 0.1515917,
  0.2943662, 0.1586402, 0.172873, 0.05629392, 0.2728668, 0.2631553, 
    0.05378783, 0.3348631, 0.2722608, 0.2375141, 0.2403411, 0.2359125, 
    0.2522019, 0.1955614, 0.3298457, 0.4234229, 0.4148854, 0.3858494, 
    0.3734446, 0.3595178, 0.4562899, 0.443885, 0.2046124, 0.3734183, 
    0.3842672, 0.3798106, 0.6081311, 0.5375466, 0.4349023,
  0.4140736, 0.2002767, 0.1493897, 0.200436, 0.201296, 0.1786502, 0.3228639, 
    0.3014501, 0.3269188, 0.3401123, 0.3281939, 0.4065284, 0.356293, 
    0.3071327, 0.3430399, 0.3404045, 0.3893039, 0.3525213, 0.3252167, 
    0.2300918, 0.1947907, 0.1261852, 0.2266043, 0.2544447, 0.3281724, 
    0.4605314, 0.4952089, 0.5196182, 0.5571595,
  0.1739427, 0.1932555, 0.2099951, 0.1552147, 0.1442873, 0.1352336, 
    0.1101222, 0.1544093, 0.2129343, 0.2464431, 0.174704, 0.1943212, 
    0.1447227, 0.2220801, 0.2847019, 0.173403, 0.3242657, 0.4027659, 
    0.4052896, 0.2603344, 0.2146076, 0.182316, 0.1449556, 0.2173228, 
    0.09831082, 0.2092742, 0.342172, 0.3107924, 0.20266,
  0.1405092, 0.06899615, 0.01797726, 0.05191821, 0.118384, 0.1416838, 
    0.1725672, 0.2106386, 0.2175996, 0.1381013, 0.0932977, 0.04377778, 
    0.01380321, 0.09805748, 0.4129958, 0.07721203, 0.146925, 0.1965502, 
    0.1837569, 0.1349472, 0.149252, 0.09787979, 0.1157189, 0.3156742, 
    0.1073636, 0.07828802, 0.1205954, 0.131029, 0.07168567,
  0.04162803, 0.08334084, 0.01142808, 0.06204396, 0.07726143, 0.04154645, 
    0.01823625, 0.06039537, 0.05476564, 0.008878381, 0.0004795374, 
    8.62555e-05, 0.01350996, 0.01592937, 0.03989072, 0.0408275, 0.06493229, 
    0.08761652, 0.09831743, 0.07312728, 0.03895975, 0.0235202, 0.07040855, 
    0.03474358, 0.04362208, 0.05018549, 0.01826081, 0.04261937, 0.05236559,
  0.04010389, 0.02790338, 0.0001468488, 0.05145481, 0.001070264, 0.000949482, 
    0.001230901, 0.05272092, 0.01089932, 0.0001073205, 2.133989e-12, 
    -6.631827e-09, 0.01420879, 0.06835912, 0.05502977, 0.03409293, 
    0.06325978, 0.08418692, 0.01246196, 0.005011041, 0.01677249, 0.02318885, 
    0.1026965, -0.0006196392, 0.07505833, 0.03558435, 0.008937929, 
    0.005172907, 0.01137749,
  0.1699197, 0.03081857, -4.982511e-07, 0.1068625, 0.01738944, 0.006062451, 
    0.005158794, 0.01058947, 0.001000519, -0.002909607, 0.01877727, 
    0.00378845, 0.07409523, 0.01402503, 0.01244282, 0.003125791, 0.001875569, 
    0.00551632, 0.003317205, 0.003367827, 0.009667888, 0.04804116, 0.3076996, 
    0.002057002, 1.865999e-05, -7.887083e-07, -0.001885971, 0.00107718, 
    0.03398369,
  0.1696176, 0.0389967, 0.003721171, 0.0272284, 0.03202206, 0.001741678, 
    0.005817463, 0.0115563, 0.04440622, 0.02702735, 0.005077139, 0.006245915, 
    0.02311204, 0.006497436, 0.01860988, 0.004197385, 0.02395326, 0.01009817, 
    0.005734256, 0.01656391, 0.06172385, 0.1688468, 0.4087479, 0.08582112, 
    0.03265269, 0.01035503, 0.03174874, 0.01301427, 0.0318362,
  0.0003986238, 0.0002639044, 5.531082e-06, -3.60497e-06, -1.104054e-05, 
    0.0005254071, 0.05271947, 0.0005482103, -0.0006482542, 0.004428707, 
    0.009748545, 0.03893442, 0.009192527, 0.006294705, 0.01801679, 
    0.01371007, 0.01951711, 0.04618277, 0.0606226, 0.05957581, 0.05093119, 
    0.06593598, 0.09037175, 0.01342076, 0.01043379, 0.04174015, 0.06971175, 
    0.1299727, 0.0128177,
  1.055674e-06, 1.099483e-06, 4.318881e-08, 1.787786e-09, 6.761733e-09, 
    0.1611757, 0.00787676, 0.01482213, 0.08238336, 0.05618102, 0.04502672, 
    0.02660274, 0.0007332601, 0.0009265449, 0.00378964, 0.0161062, 
    0.01553489, 0.03601272, 0.1450756, 0.281813, 0.08502994, 0.02014829, 
    0.004151059, 0.0001355695, 0.001033721, 0.001432601, 0.01679306, 
    0.1053085, 3.196642e-07,
  5.374155e-07, 1.825265e-06, 9.066436e-09, 8.398816e-07, 3.578092e-07, 
    2.968172e-08, -5.774359e-06, 0.08152011, 0.3456468, 0.02370389, 
    0.2008238, 0.4109362, 0.2797685, 0.1933677, 0.2228525, 0.1282318, 
    0.1456671, 0.03097546, 0.08713336, 0.2184799, 1.308601e-07, 0.02574499, 
    0.0469728, 0.04107932, 0.0430735, 0.04168709, 0.02640113, 0.09043343, 
    0.008669874,
  -0.001325101, 0.00160208, -6.888611e-05, 0.1091326, 0.000277256, 
    -8.141425e-07, 0.02301337, 4.456933e-06, -3.576552e-05, 0.0005793346, 
    0.2803236, 0.2744903, 0.447831, 0.5342473, 0.358115, 0.261739, 0.4228236, 
    0.5666887, 0.3697389, 0.05109392, 0.006866797, 0.03103008, 0.02078974, 
    0.0424457, 0.227206, 0.2771429, 0.175192, 0.2605012, 0.1212149,
  0.1405747, 0.1329549, 0.09374265, -0.0004013341, 0.002681647, 0.003210029, 
    0.01510085, 0.1372877, 0.08171985, 0.03130833, 0.1630103, 0.1880929, 
    0.5098757, 0.3357847, 0.4866768, 0.6264524, 0.4810601, 0.4909265, 
    0.3163403, 0.1474155, 0.01660346, 0.008602389, 0.02032228, 0.1623287, 
    0.1263803, 0.2432874, 0.3733867, 0.4180714, 0.1310354,
  0.1531726, 0.04232083, 0.05290117, 0.05105821, 0.07488336, 0.0580815, 
    0.0648073, 0.05158351, 0.06038567, 0.02676941, 0.03780901, 0.1360927, 
    0.1043438, 0.1290183, 0.4049602, 0.3937535, 0.2603864, 0.3217634, 
    0.1075636, 0.007243702, 0.01057749, 0.08618414, 0.1171381, 0.1880731, 
    0.3428605, 0.2251423, 0.4860694, 0.3308874, 0.1793054,
  0.4451056, 0.4009208, 0.317891, 0.4263926, 0.2877322, 0.3247889, 0.19157, 
    0.1515767, 0.0972537, 0.1537142, 0.1295242, 0.07126479, 0.05924264, 
    0.1495684, 0.2381429, 0.162942, 0.122308, 0.2191956, 0.2690954, 
    0.3252612, 0.393275, 0.5075556, 0.1553418, 0.3796945, 0.1549329, 
    0.3564304, 0.2276816, 0.1714129, 0.4109754,
  0.60755, 0.5640274, 0.4045913, 0.3902225, 0.4226193, 0.4872241, 0.4834418, 
    0.4329187, 0.469138, 0.46328, 0.4141717, 0.4586623, 0.4713977, 0.4970443, 
    0.5463384, 0.5647354, 0.5469514, 0.4887829, 0.529652, 0.5695119, 
    0.5319236, 0.4255882, 0.3333752, 0.4015858, 0.2715828, 0.2188092, 
    0.09978164, 0.257124, 0.4920674,
  0.1370479, 0.1357534, 0.134459, 0.1331645, 0.13187, 0.1305755, 0.1292811, 
    0.1626512, 0.183018, 0.2033849, 0.2237518, 0.2441187, 0.2644855, 
    0.2848524, 0.322751, 0.3163008, 0.3098506, 0.3034003, 0.2969501, 
    0.2904999, 0.2840496, 0.2542166, 0.2415945, 0.2289723, 0.2163501, 
    0.203728, 0.1911058, 0.1784837, 0.1380835,
  0.1399632, 0.2589181, 0.1360819, 0.1266608, 0.1012153, 0.1979637, 
    0.2672009, 0.2094958, 0.009980102, 0.001687909, 0.03916633, 0.13091, 
    0.2147904, 0.01305254, 0.1958013, 0.2061466, 0.294057, 0.1897097, 
    0.1467793, 0.1436002, 0.2785613, 0.4045767, 0.4433841, 0.2852738, 
    0.2222589, 0.1858993, 0.05505071, 0.08631222, 0.1171733,
  0.2684484, 0.1300165, 0.1464578, 0.03421434, 0.1870546, 0.2276786, 
    0.03030896, 0.309542, 0.2554939, 0.2230902, 0.2277998, 0.2488437, 
    0.2296541, 0.1714018, 0.3308643, 0.4332, 0.398697, 0.3690868, 0.4002984, 
    0.3254899, 0.4507453, 0.4347454, 0.2145906, 0.3566473, 0.3715338, 
    0.4511947, 0.6962283, 0.5611659, 0.4168398,
  0.3531699, 0.1569221, 0.104126, 0.1539237, 0.1645901, 0.1310143, 0.2635827, 
    0.2411665, 0.2713726, 0.2911586, 0.2631795, 0.3356515, 0.313287, 
    0.2850365, 0.2847653, 0.33419, 0.4030688, 0.3180592, 0.3020744, 
    0.2003625, 0.1722302, 0.1018619, 0.1977675, 0.2119337, 0.288444, 
    0.4434088, 0.441216, 0.4520451, 0.5053925,
  0.1272106, 0.1541928, 0.1784922, 0.1240229, 0.1237578, 0.1162158, 
    0.08863502, 0.1347524, 0.1895716, 0.2163276, 0.1484154, 0.1720033, 
    0.106973, 0.2048784, 0.2594096, 0.1452829, 0.2696119, 0.3915859, 
    0.3854195, 0.2501795, 0.1837229, 0.1490961, 0.09542645, 0.1822287, 
    0.06401195, 0.1476057, 0.2874932, 0.2841639, 0.1681432,
  0.09821247, 0.04783489, 0.00862865, 0.03269419, 0.08087229, 0.1038362, 
    0.1249722, 0.1618785, 0.1672866, 0.08965103, 0.06202177, 0.02135432, 
    0.006205711, 0.06290402, 0.3599136, 0.06521687, 0.1299313, 0.1646533, 
    0.1428595, 0.1274601, 0.1111474, 0.05871711, 0.0805136, 0.3030625, 
    0.08158807, 0.04978366, 0.08241755, 0.08360896, 0.04266804,
  0.0210038, 0.04611214, 0.01165168, 0.03731214, 0.03953586, 0.01858334, 
    0.008317823, 0.04877558, 0.04508511, 0.004911726, 0.0002411095, 
    0.0001168342, 0.01619596, 0.01074365, 0.02965786, 0.03229839, 0.05507055, 
    0.07327063, 0.06279028, 0.0480005, 0.01955899, 0.01308816, 0.03599467, 
    0.04069915, 0.03962515, 0.02284811, 0.007606902, 0.01996899, 0.03037105,
  0.01719108, 0.02891062, 0.0003497406, 0.01863614, -0.002915844, 
    0.0004201646, 0.0003570718, 0.04597571, 0.004086859, 6.663513e-05, 
    1.612612e-12, -7.629883e-09, 0.01124957, 0.04182892, 0.02682896, 
    0.008430072, 0.01760284, 0.03337615, 0.005769922, 0.001638182, 
    0.006500053, 0.007426364, 0.03907233, 0.02908684, 0.051799, 0.05880341, 
    0.002868262, 0.001685656, 0.004129331,
  0.07552917, 0.01215622, -6.902979e-06, 0.1158718, 0.00636988, 0.001365021, 
    0.001234449, 0.003227873, 0.0003458932, -0.00221744, 0.01084583, 
    0.0006178669, 0.03878721, 0.002858898, 0.003864225, 0.0009567026, 
    0.0005285412, 0.001441595, 0.001231815, 0.001506161, 0.004329749, 
    0.01737924, 0.1321442, 0.0003856417, 1.290015e-06, -1.591403e-07, 
    -0.0006672816, 0.0004263377, 0.01474959,
  0.04687367, 0.0268383, 0.004226398, 0.01728532, 0.004637954, 0.0003592727, 
    0.001379407, 0.005412942, 0.04782136, 0.0186414, 0.0008771938, 
    0.0006157622, 0.01099443, 0.001122111, 0.008300124, 0.0003573479, 
    0.009429052, 0.0002437936, 0.0002261668, 0.001244222, 0.01101771, 
    0.03944387, 0.1922387, 0.08003605, 0.0303949, 0.004424209, 0.02518557, 
    0.002115439, 0.005773333,
  0.0001860988, 0.000109148, -1.559156e-06, -1.096505e-05, 1.010055e-05, 
    2.232434e-05, 0.0410049, 2.248909e-05, -0.0005813913, 0.0005555074, 
    0.004178981, 0.02317341, 0.00145301, 0.0008769264, 0.006188718, 
    0.002625359, 0.01012202, 0.01755157, 0.03097319, 0.0166822, 0.01228049, 
    0.0255438, 0.09987152, 0.008020001, 0.00143421, 0.01350477, 0.01901217, 
    0.05817, 0.01077589,
  9.953114e-07, 1.035044e-06, 4.244311e-08, 1.277544e-09, 5.642681e-09, 
    0.05401125, 0.00360204, 0.01233893, 0.07245561, 0.02447542, 0.01585214, 
    0.01865249, 2.839813e-05, 7.420161e-05, 0.0006711169, 0.003908505, 
    0.008589394, 0.01392649, 0.06901827, 0.1233724, 0.114823, 0.01177775, 
    0.001119539, -0.0005461635, 0.0001289391, 0.0003459814, 0.006542297, 
    0.04117791, 6.216263e-08,
  5.083438e-07, 2.639384e-07, -8.82122e-09, 8.036744e-07, 3.355283e-07, 
    2.956371e-08, -3.322749e-06, 0.07345273, 0.334464, 0.02038358, 0.1916634, 
    0.3556229, 0.3077469, 0.1065947, 0.1230809, 0.0604732, 0.09703771, 
    0.01246679, 0.04066518, 0.1815244, 1.207087e-07, 0.02229588, 0.05021536, 
    0.01438709, 0.02068838, 0.03444579, 0.0123758, 0.02887673, 0.01783552,
  -0.001175215, 0.0009431613, -9.513443e-05, 0.1121985, -5.136722e-05, 
    7.283189e-08, 0.01746144, 1.483841e-06, -3.052026e-05, -0.0004455119, 
    0.2646742, 0.2222334, 0.3610229, 0.4354296, 0.2566848, 0.2135263, 
    0.4314519, 0.3708586, 0.2743686, 0.04639498, 0.006274497, 0.02223693, 
    0.01399424, 0.03217563, 0.1851534, 0.2302359, 0.1437514, 0.1872814, 
    0.1329855,
  0.1130248, 0.1227707, 0.06731708, -0.0005332725, 0.0007488942, 0.001281229, 
    0.01176728, 0.1294278, 0.07474933, 0.02995639, 0.1596868, 0.1910574, 
    0.5360528, 0.3369311, 0.4751083, 0.5444832, 0.4877767, 0.5642455, 
    0.2754082, 0.1401846, 0.0103559, 0.005188175, 0.01767806, 0.1516076, 
    0.1285085, 0.2536377, 0.3801851, 0.3850487, 0.1583519,
  0.1725965, 0.0293889, 0.04150444, 0.04366207, 0.05850589, 0.04603998, 
    0.04626481, 0.0393174, 0.04740816, 0.02233308, 0.03602352, 0.124871, 
    0.08531689, 0.1482751, 0.4329954, 0.4162995, 0.2314211, 0.2823019, 
    0.08729225, 0.003632656, 0.007483691, 0.09079058, 0.1127682, 0.1552516, 
    0.3643004, 0.2004587, 0.4054481, 0.2649366, 0.1282373,
  0.5288747, 0.3801596, 0.2597238, 0.3925734, 0.2898463, 0.3265413, 
    0.1518694, 0.1383838, 0.07701817, 0.1301285, 0.1085505, 0.05137905, 
    0.0451984, 0.1727263, 0.2034859, 0.1614498, 0.09457308, 0.1976485, 
    0.2847002, 0.2733449, 0.2921724, 0.4240774, 0.1177813, 0.3192645, 
    0.1669164, 0.3063715, 0.1851789, 0.1780706, 0.5000083,
  0.6305339, 0.4813277, 0.2702223, 0.334919, 0.3686137, 0.4127651, 0.4573088, 
    0.4624566, 0.3936927, 0.4680094, 0.4087959, 0.3999018, 0.4521515, 
    0.4672485, 0.530253, 0.550751, 0.5157396, 0.5364575, 0.5287276, 
    0.4971167, 0.5240062, 0.394228, 0.2804624, 0.3888633, 0.2291532, 
    0.1542811, 0.1021191, 0.3683391, 0.4614212,
  0.06687903, 0.06453998, 0.06220093, 0.05986188, 0.05752283, 0.05518378, 
    0.05284473, 0.05236546, 0.06822726, 0.08408907, 0.09995087, 0.1158127, 
    0.1316745, 0.1475363, 0.1807851, 0.1780778, 0.1753706, 0.1726633, 
    0.1699561, 0.1672488, 0.1645415, 0.1318028, 0.1209873, 0.1101718, 
    0.09935634, 0.08854084, 0.07772536, 0.06690986, 0.06875028,
  0.150223, 0.233447, 0.08625349, 0.1038498, 0.06746922, 0.1578824, 
    0.2133923, 0.1674335, 0.008544817, 0.002663225, 0.002235947, 0.07342818, 
    0.2283267, 0.006563863, 0.2534513, 0.2459519, 0.3971389, 0.2215515, 
    0.1232691, 0.1661931, 0.2667904, 0.4249825, 0.3063406, 0.2320919, 
    0.159083, 0.1998864, 0.07233704, 0.0956633, 0.1152701,
  0.239791, 0.1161822, 0.1303371, 0.0207456, 0.1220955, 0.2002393, 
    0.01309073, 0.2631292, 0.2344933, 0.1965969, 0.2105916, 0.2603021, 
    0.2027335, 0.1516591, 0.3408729, 0.406676, 0.3685144, 0.3608825, 
    0.3923987, 0.3073823, 0.4610066, 0.3849004, 0.2475578, 0.3337949, 
    0.3583888, 0.5008827, 0.7031288, 0.5647407, 0.3859947,
  0.296211, 0.1126106, 0.07076733, 0.1060232, 0.1184453, 0.09371948, 
    0.2028381, 0.1841221, 0.209433, 0.2253361, 0.1953853, 0.2706467, 
    0.2564198, 0.2457967, 0.2680978, 0.2957537, 0.3769206, 0.2883371, 
    0.2533961, 0.1628878, 0.1396233, 0.07883367, 0.1708439, 0.1669228, 
    0.2431189, 0.4000273, 0.3898295, 0.3809532, 0.4281781,
  0.09905187, 0.1153873, 0.1377108, 0.09563427, 0.1037406, 0.1007403, 
    0.07434781, 0.1083169, 0.157927, 0.1821164, 0.1139594, 0.1321827, 
    0.07545243, 0.1516371, 0.2133021, 0.101912, 0.2164516, 0.3677009, 
    0.3448452, 0.2114574, 0.1524106, 0.1164313, 0.061269, 0.1453855, 
    0.04765813, 0.0964878, 0.2367029, 0.2418425, 0.1259801,
  0.06554495, 0.02883306, 0.00399426, 0.01931546, 0.04898374, 0.06254721, 
    0.07988326, 0.1162631, 0.1101496, 0.05392195, 0.03622668, 0.01011468, 
    0.003087883, 0.03684026, 0.2937941, 0.05330767, 0.09790926, 0.1240909, 
    0.1053182, 0.1035551, 0.07641993, 0.03178937, 0.0611286, 0.287636, 
    0.0550688, 0.03474091, 0.05671056, 0.05044379, 0.02600233,
  0.008477109, 0.02507726, 0.01151907, 0.01954184, 0.01641234, 0.00664791, 
    0.004181082, 0.03846848, 0.03377537, 0.003351694, 0.0001102792, 
    -7.578405e-06, 0.01607867, 0.007540764, 0.02188255, 0.0241578, 
    0.04556064, 0.05117792, 0.04362917, 0.02695292, 0.007132353, 0.004290661, 
    0.01636473, 0.02043928, 0.03211689, 0.01015354, 0.003220036, 0.008841795, 
    0.01605954,
  0.009814578, 0.03060822, 0.000164915, 0.01025482, -0.00230861, 
    0.0002604372, 0.0001787008, 0.02652708, 0.002070867, 4.6622e-05, 
    1.789292e-12, -7.597684e-09, 0.007671639, 0.01763922, 0.01102123, 
    0.00237178, 0.007864407, 0.01479638, 0.002352291, 0.0005997755, 
    0.002131064, 0.003842466, 0.02006966, 0.01726349, 0.04456296, 0.07844348, 
    0.001463833, 0.0008634939, 0.002077618,
  0.04312776, 0.004608193, -5.60584e-06, 0.09786598, 0.001476165, 
    0.0005275861, 0.0003980161, 0.001808972, 0.0001890813, -0.001172636, 
    0.006486418, 0.0002422892, 0.0152531, 0.00061097, 0.001986807, 
    0.0005119239, 0.0003108559, 0.0007585295, 0.0006470429, 0.0008675752, 
    0.002498174, 0.008861222, 0.07596237, 0.0002316123, 2.141294e-07, 
    -4.462835e-07, -0.0005160084, 0.0002315963, 0.008206352,
  0.02067177, 0.02651661, 0.003753389, 0.009069555, 0.000763436, 
    0.0001809463, 0.0006750962, 0.002740963, 0.04384656, 0.01462419, 
    0.0003435133, 0.000190006, 0.006295281, 0.0002508356, 0.002443023, 
    4.00119e-05, 0.003228145, -1.66606e-05, 6.288985e-05, 0.0002296742, 
    0.003976768, 0.01307195, 0.0888498, 0.07806593, 0.03616286, 0.001781633, 
    0.01646471, 0.0009276274, 0.002515593,
  2.864268e-05, 5.100984e-05, -6.58436e-07, -5.436673e-06, 1.205489e-07, 
    4.515451e-06, 0.02034866, 9.349724e-06, -0.0002775806, 0.0001459514, 
    0.001697371, 0.01184358, 0.0003574664, 0.0001429854, 0.001946799, 
    0.0004065347, 0.003941184, 0.00555509, 0.01145714, 0.006461321, 
    0.003877209, 0.01299495, 0.08879539, 0.008463517, 0.0004792196, 
    0.004823669, 0.007806156, 0.03191146, 0.01532818,
  9.482941e-07, 9.893394e-07, 4.254025e-08, 1.004736e-09, 5.492901e-09, 
    0.02413384, -0.0004374949, 0.001962087, 0.06202707, 0.009321654, 
    0.004803828, 0.01198724, 1.030806e-05, 2.417108e-05, 0.0003270968, 
    0.00190551, 0.004714449, 0.006361001, 0.03504134, 0.06776182, 0.08471283, 
    0.009082764, 0.0005210484, -0.0008584831, 5.384901e-05, 0.0001837478, 
    0.003432145, 0.0197862, 4.69736e-08,
  4.975157e-07, 1.599866e-06, -2.821337e-05, 7.804776e-07, 3.121804e-07, 
    2.949494e-08, -2.427721e-06, 0.06171302, 0.3124183, 0.01626298, 
    0.1633579, 0.2385498, 0.2145149, 0.02819065, 0.07163766, 0.02965339, 
    0.04723891, 0.005046643, 0.02495461, 0.1208268, 1.161744e-07, 0.01745722, 
    0.04230256, 0.005267312, 0.01026777, 0.01375054, 0.004109131, 0.01428383, 
    0.01589624,
  -0.001187833, 0.0003291701, -8.957888e-05, 0.1009187, -0.0001332192, 
    4.400293e-07, 0.01214387, 1.134695e-06, -2.426112e-05, 4.884766e-05, 
    0.2388175, 0.1693585, 0.3056759, 0.337611, 0.2053231, 0.1723962, 
    0.3929892, 0.2155127, 0.2014079, 0.03836771, 0.005679139, 0.01510092, 
    0.008150483, 0.02346623, 0.1569328, 0.1711149, 0.09425043, 0.1328939, 
    0.08660936,
  0.08957904, 0.1162154, 0.04391199, -0.0004077766, 0.00030356, 0.0002143781, 
    0.008172238, 0.119818, 0.06275676, 0.02591833, 0.1646634, 0.1734118, 
    0.5542969, 0.366338, 0.4387082, 0.4539145, 0.4206451, 0.5103244, 
    0.2176237, 0.1295266, 0.006928423, 0.002682937, 0.01466471, 0.1378353, 
    0.1290573, 0.2957572, 0.3654244, 0.3099891, 0.1613425,
  0.2216759, 0.02244406, 0.02987946, 0.03088486, 0.04291029, 0.037137, 
    0.03134855, 0.02483897, 0.04266278, 0.0194316, 0.03449929, 0.1061545, 
    0.0725093, 0.1412457, 0.4185684, 0.4298052, 0.1995083, 0.2431034, 
    0.06495615, 0.002132579, 0.006437558, 0.07670348, 0.1131907, 0.1251381, 
    0.3374245, 0.1875222, 0.3227399, 0.1883547, 0.1499448,
  0.545023, 0.3723749, 0.2120673, 0.349504, 0.2237163, 0.3430574, 0.1945017, 
    0.1169209, 0.06390455, 0.1063724, 0.09352215, 0.04166272, 0.03265224, 
    0.1609352, 0.1929848, 0.2122424, 0.0617138, 0.160019, 0.2382115, 
    0.1890274, 0.2202739, 0.3477152, 0.08925643, 0.2608138, 0.1478179, 
    0.2600305, 0.1393023, 0.1776705, 0.5214714,
  0.5452734, 0.3879451, 0.1793205, 0.3234832, 0.3542299, 0.4142577, 
    0.4609136, 0.4450128, 0.3266995, 0.4135352, 0.3815283, 0.3594055, 
    0.3941211, 0.4468693, 0.4967868, 0.4894159, 0.4802227, 0.4921913, 
    0.476295, 0.3442197, 0.4719681, 0.3267681, 0.2081494, 0.3371387, 
    0.1925529, 0.1131292, 0.08841208, 0.3602917, 0.3887067,
  0.01312607, 0.01031134, 0.007496613, 0.004681883, 0.001867154, 
    -0.0009475756, -0.003762305, -0.02450204, -0.01326158, -0.002021121, 
    0.009219341, 0.0204598, 0.03170026, 0.04294073, 0.0865261, 0.08558026, 
    0.08463442, 0.08368858, 0.08274274, 0.0817969, 0.08085106, 0.05527757, 
    0.04779768, 0.04031779, 0.0328379, 0.025358, 0.01787811, 0.01039822, 
    0.01537785,
  0.1709878, 0.138003, 0.04666971, 0.03127191, 0.01714034, 0.06984116, 
    0.0961485, 0.07282211, 0.02889867, 0.01146461, 0.01228895, 0.02177054, 
    0.1554652, 0.005366279, 0.2992078, 0.3320437, 0.4330211, 0.2271218, 
    0.09427339, 0.1827251, 0.2754481, 0.3993279, 0.2194001, 0.178379, 
    0.1428364, 0.2570027, 0.07948329, 0.0883642, 0.1470973,
  0.2290378, 0.09643407, 0.1071636, 0.01469061, 0.08063713, 0.1716352, 
    0.008248067, 0.2065335, 0.208826, 0.1658771, 0.2039787, 0.2534359, 
    0.1823862, 0.1390127, 0.3505324, 0.3915877, 0.3334623, 0.3398488, 
    0.3581639, 0.2644446, 0.3967816, 0.3442486, 0.2439599, 0.317848, 
    0.3522639, 0.5101858, 0.630806, 0.5124421, 0.3480835,
  0.233025, 0.0756368, 0.05045962, 0.07366487, 0.08353083, 0.06688915, 
    0.1503874, 0.1371438, 0.1596882, 0.1610999, 0.1292173, 0.2184371, 
    0.1922432, 0.1949126, 0.2217414, 0.2374181, 0.3123338, 0.2261992, 
    0.2082008, 0.1233957, 0.1107397, 0.06018182, 0.1384588, 0.1240345, 
    0.2011965, 0.3252361, 0.3012277, 0.3013557, 0.3283455,
  0.07527215, 0.08605608, 0.1007927, 0.0705579, 0.08550398, 0.08467328, 
    0.05960939, 0.08229531, 0.1203206, 0.1350262, 0.07370482, 0.08802474, 
    0.04763874, 0.08918432, 0.1538687, 0.05445203, 0.16635, 0.2973068, 
    0.2593368, 0.151865, 0.1159452, 0.0785421, 0.03948353, 0.1197519, 
    0.03593681, 0.05702578, 0.1815426, 0.2008043, 0.09105334,
  0.04205864, 0.01699126, 0.002269244, 0.0122023, 0.02834985, 0.0333398, 
    0.05420944, 0.07434652, 0.0682699, 0.02795352, 0.01972503, 0.005335679, 
    0.001660026, 0.01692051, 0.2333538, 0.03581658, 0.05678883, 0.0825148, 
    0.06410997, 0.06970942, 0.05150443, 0.01837128, 0.04356984, 0.266552, 
    0.03986099, 0.02214413, 0.03315408, 0.02959909, 0.0157414,
  0.003890091, 0.01579184, 0.01229637, 0.01010935, 0.00584536, 0.003036866, 
    0.002478383, 0.02463256, 0.02429504, 0.002558735, 6.200389e-05, 
    -3.787523e-05, 0.01348224, 0.004996774, 0.01328558, 0.0148113, 
    0.03183869, 0.02750394, 0.02675601, 0.0143326, 0.003279775, 0.001616138, 
    0.007238057, 0.01056278, 0.02701522, 0.004864146, 0.001678551, 
    0.003250062, 0.006438765,
  0.006633538, 0.02798114, 0.0001596453, 0.006860198, -0.001532018, 
    0.0001844261, 0.0001094749, 0.0102397, 0.001274886, 3.561588e-05, 
    1.840988e-12, -7.649242e-09, 0.003976866, 0.007519453, 0.004104218, 
    0.001095573, 0.004527162, 0.006638032, 0.0008441862, 0.0002815423, 
    0.001050019, 0.002475276, 0.0128711, 0.01144515, 0.03755703, 0.08714142, 
    0.0009953901, 0.0005472586, 0.001281925,
  0.02915776, 0.002439849, -1.057744e-05, 0.07477728, 0.000393685, 
    0.0002898061, 0.0001634586, 0.001213702, 0.0001322344, -0.0005391133, 
    0.004343932, 0.0001101172, 0.005515356, 0.0002670152, 0.00118546, 
    0.0003371136, 0.0002113283, 0.0005009471, 0.000410335, 0.0005923435, 
    0.001682192, 0.00556526, 0.04956454, 0.0004347042, 2.619903e-07, 
    -1.633589e-08, -0.0002075298, 0.0001500551, 0.005413961,
  0.01212369, 0.03009618, 0.002447255, 0.004577825, 0.0004086768, 
    0.0001159407, 0.0004267476, 0.001407638, 0.03201291, 0.01578085, 
    0.000203677, 0.0001044514, 0.002607486, 7.829035e-05, 0.0007318587, 
    1.865743e-05, 0.0009951941, 1.304952e-06, 3.46294e-05, 0.0001253291, 
    0.002174689, 0.006546376, 0.05319223, 0.05964539, 0.03712902, 
    0.0006149537, 0.008023313, 0.0005427096, 0.001561699,
  -1.2784e-05, 2.468497e-05, -5.349453e-07, -2.477959e-06, 1.104326e-06, 
    1.825619e-06, 0.007268725, 5.26253e-06, -9.627367e-05, 6.497523e-05, 
    0.0007688871, 0.005183473, 0.0001392952, 2.903027e-05, 0.000664106, 
    0.0001780909, 0.001154338, 0.002003855, 0.003782374, 0.003990437, 
    0.001867664, 0.006541948, 0.0703719, 0.01238342, 0.0003210524, 
    0.001972447, 0.003740083, 0.01523585, 0.01203822,
  9.14128e-07, 9.653257e-07, 4.296798e-08, 8.613829e-10, 5.427605e-09, 
    0.0135919, -0.001276504, 0.0003130008, 0.05296442, 0.003090089, 
    0.001554257, 0.006181011, 5.546102e-06, 1.41976e-05, 0.0002083739, 
    0.001212981, 0.002599265, 0.003570359, 0.02086501, 0.04387286, 0.0518467, 
    0.006244298, 0.0003011802, -0.0009058407, 3.084157e-05, 0.0001201779, 
    0.002182626, 0.01215596, 4.606036e-08,
  4.909242e-07, 1.788587e-06, 3.764584e-06, 7.189809e-07, 2.960749e-07, 
    2.945716e-08, -2.013805e-06, 0.0516039, 0.2853262, 0.009140283, 
    0.1088443, 0.1408698, 0.08933557, 0.009968463, 0.04578515, 0.01082028, 
    0.02030207, 0.00280988, 0.01517433, 0.07626408, 1.133142e-07, 0.013456, 
    0.03189813, 0.001807723, 0.002661276, 0.005781706, 0.002045353, 
    0.00918393, 0.01354468,
  -0.001087299, 9.394089e-05, -7.054725e-05, 0.09246992, -0.0001251452, 
    3.606557e-07, 0.009258362, 5.849558e-07, -1.951547e-05, 0.000283669, 
    0.2014153, 0.1358603, 0.250044, 0.2503338, 0.1696546, 0.1341641, 
    0.3216764, 0.1400275, 0.1300526, 0.03169211, 0.004082329, 0.008522875, 
    0.004672619, 0.04940285, 0.121786, 0.1111291, 0.0565246, 0.08089509, 
    0.06002224,
  0.0595682, 0.1013906, 0.0298971, -0.0001233593, 0.0001609358, 7.065787e-05, 
    0.006616945, 0.1076316, 0.05231669, 0.02109101, 0.1514425, 0.1446603, 
    0.4607567, 0.3359244, 0.3427094, 0.353434, 0.3148599, 0.3725698, 
    0.1565678, 0.1124219, 0.004337448, 0.001502512, 0.01351325, 0.1180609, 
    0.1242669, 0.2823227, 0.3095672, 0.2187032, 0.1348661,
  0.3110629, 0.01780094, 0.01854734, 0.02416349, 0.03265114, 0.02870324, 
    0.02447777, 0.01560482, 0.04072339, 0.01734167, 0.03066991, 0.08999851, 
    0.05900775, 0.1242728, 0.3712041, 0.3637269, 0.1631447, 0.2154182, 
    0.04764961, 0.001983368, 0.004779796, 0.05445998, 0.0984484, 0.09750435, 
    0.2830839, 0.1631721, 0.2259047, 0.1161425, 0.132152,
  0.4909719, 0.3171276, 0.1770455, 0.2797296, 0.1718966, 0.3445497, 
    0.2024923, 0.1035265, 0.05700564, 0.08684621, 0.06699596, 0.0282251, 
    0.02051595, 0.1314357, 0.1732742, 0.3090648, 0.03796107, 0.1177309, 
    0.1959593, 0.1401614, 0.1709502, 0.2951956, 0.06459152, 0.2202791, 
    0.1202366, 0.2159941, 0.1172972, 0.1491333, 0.4823712,
  0.4534509, 0.3357246, 0.1275081, 0.3013856, 0.308801, 0.3609986, 0.4225812, 
    0.375795, 0.2843617, 0.3548441, 0.3248078, 0.305717, 0.3107148, 
    0.3853801, 0.4248838, 0.415007, 0.4127392, 0.4154127, 0.4026498, 
    0.2308573, 0.3614318, 0.2442872, 0.1558582, 0.2731231, 0.1623152, 
    0.08562385, 0.07521395, 0.3453979, 0.3118494,
  0.004821852, 0.004244498, 0.003667143, 0.003089789, 0.002512434, 
    0.001935079, 0.001357725, -0.00457966, -0.001710595, 0.001158469, 
    0.004027533, 0.006896597, 0.009765661, 0.01263473, 0.01761499, 
    0.01757837, 0.01754176, 0.01750514, 0.01746853, 0.01743191, 0.01739529, 
    0.0113094, 0.009054309, 0.006799216, 0.004544123, 0.002289029, 
    3.393623e-05, -0.002221157, 0.005283736,
  0.1662404, 0.07912147, 0.03723666, 0.02472381, 0.004292083, 0.01473855, 
    0.004025264, -0.0002501011, 0.01249702, 0.007396626, 0.003884891, 
    0.004761416, 0.06418762, 0.004653354, 0.3491358, 0.3979336, 0.4103546, 
    0.2734196, 0.08482037, 0.275032, 0.2992077, 0.3867881, 0.1712199, 
    0.1399169, 0.1765267, 0.280641, 0.08487973, 0.07504754, 0.1488773,
  0.2267075, 0.08199195, 0.08787143, 0.01084224, 0.06821984, 0.1520299, 
    0.00603419, 0.1762011, 0.1895038, 0.1459503, 0.1989118, 0.2624206, 
    0.1640057, 0.1216365, 0.3307678, 0.3561999, 0.2875736, 0.316602, 
    0.3173803, 0.2382467, 0.3629751, 0.3299336, 0.2690751, 0.3051579, 
    0.3333923, 0.4671897, 0.5610815, 0.4580947, 0.3057768,
  0.1978872, 0.05734479, 0.03875284, 0.05741705, 0.06203141, 0.05239245, 
    0.1218876, 0.109527, 0.1288254, 0.1250758, 0.09661086, 0.1757844, 
    0.1470192, 0.1614894, 0.1844117, 0.1899893, 0.262339, 0.1861834, 
    0.1730863, 0.09779319, 0.08838876, 0.04780502, 0.1152221, 0.09527826, 
    0.1648248, 0.2678127, 0.2479449, 0.2472751, 0.2723844,
  0.05978972, 0.06773738, 0.07779457, 0.05678185, 0.07631456, 0.0757053, 
    0.05161058, 0.06445162, 0.0945475, 0.09979328, 0.05145172, 0.05825735, 
    0.03324904, 0.05268167, 0.10815, 0.03398632, 0.1208627, 0.222379, 
    0.190549, 0.1047571, 0.09078865, 0.05569087, 0.02820075, 0.1083174, 
    0.02651382, 0.03817787, 0.1401727, 0.164421, 0.06939813,
  0.02822194, 0.01107253, 0.001573453, 0.008392622, 0.01684725, 0.02117351, 
    0.03823482, 0.04451483, 0.04122673, 0.01633207, 0.011694, 0.003307933, 
    0.001247875, 0.007165234, 0.191872, 0.02388285, 0.03495309, 0.05125653, 
    0.03740346, 0.04355836, 0.03479163, 0.01015133, 0.0311937, 0.2551354, 
    0.03144279, 0.01214883, 0.01898391, 0.02006038, 0.01035291,
  0.002421634, 0.01152633, 0.01203402, 0.006152337, 0.003152945, 0.002098526, 
    0.001852735, 0.01394781, 0.01927161, 0.002098127, 5.509452e-05, 
    -6.530012e-05, 0.0117884, 0.003451963, 0.007702426, 0.006882862, 
    0.01773851, 0.01421743, 0.01494901, 0.01034881, 0.002114607, 0.000925565, 
    0.003717505, 0.007303815, 0.02234879, 0.003100941, 0.001129659, 
    0.001694817, 0.003274626,
  0.005048098, 0.0245423, -7.096454e-05, 0.005169513, -0.0009715512, 
    0.0001445728, 7.818858e-05, 0.004300317, 0.0009053271, 2.913108e-05, 
    1.882837e-12, -2.031926e-08, 0.002146879, 0.004027354, 0.002123173, 
    0.0006827269, 0.003182353, 0.004082454, 0.0004429811, 0.0001653645, 
    0.0006850066, 0.00182107, 0.009433139, 0.00894603, 0.03800176, 0.0842462, 
    0.0007621889, 0.0003978174, 0.0009145848,
  0.0220347, 0.001700094, -4.597732e-06, 0.05612167, 0.000185811, 
    0.0002051972, 0.0001031168, 0.0009119617, 0.0001005834, -0.0002029814, 
    0.003208844, 8.871537e-05, 0.002054247, 0.0001524479, 0.0006079094, 
    0.0002528765, 0.0001613524, 0.00037414, 0.0002988448, 0.0004377912, 
    0.001273665, 0.004035751, 0.03669678, 0.0007045873, 2.170499e-07, 
    4.138359e-08, -0.0001409159, 0.0001111724, 0.004044206,
  0.008467038, 0.02623698, 0.00257555, 0.002375926, 0.0002817804, 
    8.516837e-05, 0.0003120551, 0.0007137932, 0.02840158, 0.02749272, 
    0.0001430287, 7.296915e-05, 0.001299016, 4.817073e-05, 0.0003257729, 
    1.40061e-05, 0.0003378339, 4.33798e-06, 2.396048e-05, 8.568196e-05, 
    0.001471294, 0.004253014, 0.03730442, 0.03604165, 0.02977586, 
    0.0002634624, 0.003667502, 0.000378364, 0.001134729,
  0.0001472635, 5.890844e-06, -1.134363e-06, -4.709879e-05, 3.196698e-07, 
    1.214736e-06, 0.002977012, 3.81808e-06, -7.729507e-05, 3.788996e-05, 
    0.0004922911, 0.002397248, 8.488943e-05, 2.027463e-05, 0.0003206319, 
    0.0001128222, 0.0004751986, 0.00100617, 0.001471024, 0.002992544, 
    0.001139777, 0.003217252, 0.06787726, 0.01530296, 0.0002338025, 
    0.0008021354, 0.00214742, 0.008073134, 0.00911618,
  8.848637e-07, 9.499694e-07, 4.361305e-08, 6.624392e-10, 5.415902e-09, 
    0.009126814, -0.0007451468, 0.0001988539, 0.04941708, 0.0002373068, 
    0.0008953615, 0.002800246, 3.971607e-06, 1.021176e-05, 0.0001532234, 
    0.0008855287, 0.001788675, 0.0024198, 0.0147287, 0.03251821, 0.03582113, 
    0.004590197, 0.0002081148, -0.001007374, 2.136676e-05, 8.970563e-05, 
    0.001587526, 0.008717384, 4.536555e-08,
  4.850423e-07, 1.69634e-06, 0.0004496074, 7.28983e-07, 2.888339e-07, 
    2.941519e-08, -1.802433e-06, 0.04706916, 0.2588615, 0.005190894, 
    0.06556414, 0.08482513, 0.04739414, 0.004583234, 0.02948764, 0.00679847, 
    0.01008031, 0.001970108, 0.009077347, 0.05188895, 1.102939e-07, 
    0.01045637, 0.02556509, 0.001130742, 0.00145375, 0.003506088, 0.00141422, 
    0.006761974, 0.01180573,
  -0.0009191409, 2.970155e-05, -5.109078e-05, 0.09156384, -0.0001134218, 
    3.989144e-07, 0.007998796, 1.545653e-07, -1.597785e-05, 0.0001994361, 
    0.1688724, 0.1095832, 0.2079912, 0.187282, 0.1352247, 0.09820063, 
    0.2550473, 0.09700944, 0.08887362, 0.02563873, 0.003323867, 0.004721736, 
    0.0022534, 0.0370202, 0.08316647, 0.06558249, 0.03446733, 0.04331589, 
    0.04682869,
  0.03966174, 0.08594826, 0.02002753, 2.855661e-05, 9.857874e-05, 
    3.993939e-05, 0.006236521, 0.1000723, 0.04602255, 0.01879681, 0.1309007, 
    0.121217, 0.3820892, 0.2656112, 0.2513844, 0.2609824, 0.2283285, 
    0.2627645, 0.1220689, 0.1028256, 0.003400626, 0.001009013, 0.01458828, 
    0.1007394, 0.1190863, 0.2661823, 0.2173901, 0.1377425, 0.09281383,
  0.301486, 0.01368098, 0.01302111, 0.01807741, 0.0268177, 0.02310697, 
    0.02393831, 0.01161827, 0.04296475, 0.01949732, 0.02777528, 0.07551862, 
    0.04544854, 0.1079509, 0.2914695, 0.2664847, 0.1348968, 0.1909619, 
    0.0387283, 0.002007857, 0.003201985, 0.03992473, 0.09019451, 0.07606933, 
    0.227468, 0.142873, 0.1562327, 0.07203569, 0.1002755,
  0.4139046, 0.2903087, 0.1543667, 0.222281, 0.1384032, 0.317339, 0.2010919, 
    0.1076128, 0.05741071, 0.07023415, 0.05161146, 0.02014524, 0.01334951, 
    0.1089631, 0.1541761, 0.3540257, 0.02518076, 0.09810451, 0.1632659, 
    0.1067482, 0.1409157, 0.2591049, 0.04716182, 0.190451, 0.0957708, 
    0.1848599, 0.1087592, 0.1321736, 0.4084273,
  0.3744468, 0.2903448, 0.09694233, 0.2420348, 0.2348708, 0.2974199, 
    0.3442414, 0.3157582, 0.239132, 0.3004722, 0.2657618, 0.2404088, 
    0.2501464, 0.301408, 0.3591503, 0.3651477, 0.3570538, 0.3427451, 
    0.3502753, 0.1832211, 0.3033555, 0.1946401, 0.125468, 0.2343265, 
    0.1452479, 0.06999604, 0.06103561, 0.322912, 0.2419153,
  0.003101829, 0.003021918, 0.002942007, 0.002862095, 0.002782184, 
    0.002702273, 0.002622361, -0.002654138, -0.001223312, 0.0002075136, 
    0.001638339, 0.003069165, 0.004499991, 0.005930817, 0.006071579, 
    0.005788084, 0.005504589, 0.005221094, 0.004937598, 0.004654103, 
    0.004370608, 0.005591964, 0.004524544, 0.003457125, 0.002389706, 
    0.001322286, 0.0002548669, -0.0008125525, 0.003165758,
  0.1139426, 0.06065706, 0.02608033, 0.01800037, 0.00226133, 0.009067209, 
    0.003730393, 0.004076627, 0.01167819, 0.001752928, 0.0004934887, 
    0.003274766, 0.05330605, 0.005528295, 0.4514134, 0.3101855, 0.3517537, 
    0.3145308, 0.09126353, 0.3695453, 0.3574361, 0.4156448, 0.1549391, 
    0.1246343, 0.1483443, 0.2921789, 0.1017774, 0.07607947, 0.124138,
  0.2266357, 0.08379359, 0.08203021, 0.008664012, 0.05809554, 0.1424995, 
    0.004764386, 0.1600276, 0.1815369, 0.1381171, 0.2132749, 0.2582998, 
    0.1576981, 0.1129877, 0.3094626, 0.335844, 0.2726706, 0.2904983, 
    0.2977206, 0.2165921, 0.3475657, 0.3133765, 0.2698301, 0.2782935, 
    0.3091095, 0.4269277, 0.492166, 0.4212394, 0.2791926,
  0.1764769, 0.04892945, 0.03324956, 0.04963687, 0.05220741, 0.04530503, 
    0.1060851, 0.09682041, 0.111129, 0.1051409, 0.07978206, 0.1495496, 
    0.1214891, 0.1342483, 0.1545475, 0.1645828, 0.2306461, 0.1626978, 
    0.1503648, 0.08521318, 0.0746778, 0.04123511, 0.1008463, 0.08068553, 
    0.1398121, 0.2387093, 0.2255305, 0.2193235, 0.2459071,
  0.05176079, 0.05820234, 0.06523571, 0.04952841, 0.0678772, 0.06638562, 
    0.04670164, 0.05606445, 0.07807735, 0.08318667, 0.04031178, 0.04348994, 
    0.02681958, 0.0399126, 0.07742097, 0.02569414, 0.09430323, 0.1756736, 
    0.1458812, 0.07615202, 0.07017437, 0.04413902, 0.02261118, 0.139383, 
    0.02051791, 0.03058494, 0.1177801, 0.1386998, 0.05758491,
  0.02052585, 0.008362202, 0.001275334, 0.006516748, 0.01203067, 0.01587848, 
    0.02828122, 0.03029612, 0.03051828, 0.01162902, 0.008343868, 0.002558574, 
    0.001053172, 0.004125926, 0.1740034, 0.01788875, 0.02429065, 0.03467795, 
    0.02672753, 0.03189638, 0.02545396, 0.007187481, 0.0224278, 0.2617121, 
    0.0222778, 0.008204751, 0.01305687, 0.01504913, 0.00799269,
  0.001828763, 0.009425484, 0.01478113, 0.003918653, 0.002319777, 
    0.001734299, 0.001576124, 0.00713783, 0.01342212, 0.001843006, 
    1.951608e-05, -7.186066e-05, 0.01580936, 0.002616844, 0.005467587, 
    0.004537822, 0.009010388, 0.008240452, 0.009971046, 0.00569056, 
    0.001789946, 0.0006954657, 0.002447506, 0.005729835, 0.03137, 
    0.002405778, 0.000923522, 0.001251215, 0.002278901,
  0.004258203, 0.02113734, -0.0002283554, 0.004303757, -0.0008136022, 
    0.0001253265, 6.551999e-05, 0.00255654, 0.0007353714, 2.590227e-05, 
    1.756996e-12, -1.847218e-08, 0.00123606, 0.002858893, 0.001492146, 
    0.0005134483, 0.002500346, 0.003112839, 0.0003215973, 0.0001221255, 
    0.0005354031, 0.001501797, 0.00777347, 0.007717735, 0.04649362, 
    0.09154331, 0.0006401189, 0.0003286903, 0.0007454079,
  0.01847047, 0.00135086, -2.968293e-06, 0.04645842, 0.0001297272, 
    0.0001692541, 8.623351e-05, 0.0007644776, 8.719815e-05, -0.0001563408, 
    0.002663253, 7.915871e-05, 0.001378101, 0.000110272, 0.0004029695, 
    0.000212229, 0.0001364312, 0.00032859, 0.000247306, 0.0003797404, 
    0.0010784, 0.003335758, 0.03021387, 0.002654247, -4.210221e-07, 
    2.369362e-08, -0.0001339515, 9.414924e-05, 0.00340075,
  0.006757699, 0.03891043, 0.003979358, 0.002406392, 0.000238953, 
    7.099806e-05, 0.0002500856, 0.0005205091, 0.04680521, 0.06871002, 
    0.0001158743, 5.79384e-05, 0.0008908649, 3.669813e-05, 0.0002187265, 
    1.326547e-05, 0.0002113166, 4.423695e-06, 1.972962e-05, 7.27145e-05, 
    0.001149835, 0.003257747, 0.02977743, 0.05247298, 0.03901488, 
    0.0001826577, 0.001911754, 0.0003050457, 0.0009307992,
  0.01465327, -6.037871e-07, -0.0001079729, -8.82099e-05, 3.12057e-07, 
    1.008255e-06, 0.01871198, 3.111304e-06, -0.002306401, 2.910378e-05, 
    0.0003899459, 0.0014593, 6.490617e-05, 1.65432e-05, 0.0002185663, 
    8.992497e-05, 0.0002980459, 0.000699393, 0.0009005973, 0.002425765, 
    0.000866873, 0.001922405, 0.1193626, 0.02549918, 0.000178867, 
    0.0004762434, 0.001532245, 0.005665075, 0.02579089,
  8.693813e-07, 9.428806e-07, 4.41533e-08, 6.829673e-10, 5.461555e-09, 
    0.007154076, -0.0005581517, 0.0001585386, 0.1098948, -0.0002488044, 
    0.0006683022, 0.001522608, 3.338973e-06, 8.540887e-06, 0.0001273794, 
    0.0007229635, 0.001418189, 0.0018994, 0.01179335, 0.02682675, 0.02823167, 
    0.004799603, 0.0001646532, -0.001825556, 1.748594e-05, 7.591245e-05, 
    0.001321196, 0.007107859, 4.486099e-08,
  4.813256e-07, 1.719834e-06, 4.346689e-06, 7.366094e-07, 2.908706e-07, 
    2.926676e-08, -1.681835e-06, 0.04956224, 0.2565667, 0.005346994, 
    0.04230832, 0.05297459, 0.02860038, 0.00252896, 0.01620572, 0.00387339, 
    0.0063284, 0.001617512, 0.00632219, 0.03927647, 1.103555e-07, 0.016793, 
    0.05486586, 0.0008869563, 0.001044728, 0.002721711, 0.001146592, 
    0.00559053, 0.01019658,
  -0.0007548711, -5.84857e-05, -4.941957e-05, 0.09898495, -0.000111495, 
    4.574203e-07, 0.008412395, 4.228278e-07, -1.342908e-05, 0.0004698283, 
    0.1739841, 0.08611467, 0.1681137, 0.1463211, 0.1031319, 0.06845154, 
    0.2010871, 0.0703662, 0.06676417, 0.02265024, 0.003073066, 0.003633665, 
    0.002220723, 0.02688838, 0.05281664, 0.03910423, 0.02298985, 0.02402077, 
    0.04082531,
  0.0300843, 0.09109193, 0.01609222, 0.0006301084, 6.719002e-05, 
    2.587476e-05, 0.007585032, 0.1002485, 0.05155092, 0.0285674, 0.1383029, 
    0.1235195, 0.3329932, 0.2226735, 0.198713, 0.2036291, 0.1701877, 
    0.2057322, 0.09241719, 0.1177361, 0.004349855, 0.0006940773, 0.0199948, 
    0.115285, 0.1294764, 0.2375127, 0.1694481, 0.09578189, 0.06418771,
  0.2635828, 0.01362056, 0.01100034, 0.02546432, 0.03134891, 0.03619752, 
    0.04537862, 0.02979602, 0.07983128, 0.0476287, 0.03977362, 0.07426008, 
    0.03346899, 0.1090686, 0.220997, 0.2054532, 0.154143, 0.1867561, 
    0.04217591, 0.006036929, 0.007458689, 0.03115033, 0.08099094, 0.06261717, 
    0.1885105, 0.1238969, 0.1199812, 0.04970997, 0.08037597,
  0.3623294, 0.2557249, 0.1465703, 0.1765603, 0.1154619, 0.321972, 0.2008918, 
    0.1276606, 0.07452619, 0.08053355, 0.04444643, 0.01774721, 0.01229031, 
    0.09199896, 0.1466549, 0.3284869, 0.01976082, 0.09013387, 0.1550411, 
    0.08781437, 0.1216161, 0.2354953, 0.0342505, 0.1717933, 0.08062723, 
    0.1642389, 0.1154028, 0.1195241, 0.3261597,
  0.3322743, 0.2421519, 0.08196965, 0.1953124, 0.1989774, 0.2571159, 
    0.2939459, 0.2762956, 0.2175041, 0.2505496, 0.2273219, 0.1960485, 
    0.1978529, 0.2506857, 0.2954805, 0.3067698, 0.3148738, 0.2987885, 
    0.3190962, 0.1616397, 0.2608035, 0.1691426, 0.1077325, 0.2128884, 
    0.1329461, 0.0621626, 0.05556951, 0.3071523, 0.2019845,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, -6.28338e-05, -8.629723e-06, 0, 0, 0.0001934205, 
    -1.707569e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0001458001, 0, -1.743515e-06, 0, 0, 0, 
    0, 0, 0, 0, 0, -1.608895e-05, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, -5.27651e-05, -0.0001208161, 0, 0, 0.007828182, 
    0.0003190515, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001130097, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0004424294, 0.0003436588, -4.934978e-05, 
    -2.821005e-06, 0, 0, 0, -3.426819e-06, 0, -2.462264e-05, -1.461686e-05, 
    -5.642043e-05, 0, -2.893673e-06, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0.001146988, 0.0004760596, -2.320508e-05, -2.459766e-05, 
    0.01787085, 0.001463385, -4.877928e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -6.467927e-06, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0.0009526605, -1.651027e-05, 0, 0, 1.198454e-05, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0.0001409429, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -7.429572e-05, -5.412493e-05, 
    0.002992075, 0, 0, 0, 0, 0, 0, 0, 0, -4.084597e-06, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.002681999, 0.00137432, 0.002825239, 
    -1.948753e-05, -1.492971e-05, 0, -1.451148e-05, 3.43776e-05, 
    0.0005897764, 0.002527683, 4.89005e-05, 0.0002536713, 0, -1.49598e-05, 0, 
    0, -4.852951e-05, 0,
  0, 0, 0, 0, 0, 0, 0.00562779, 0.001094137, -0.0001021127, 0.0005365978, 
    0.02457816, 0.00548337, 0.0007564643, 0.0001285487, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.0001292268, -4.982855e-05, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0.001347379, -8.711516e-05, 0, -4.596034e-06, 
    5.22651e-05, 2.341247e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, -5.71078e-05, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0.0001257202, 2.23359e-05, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -6.753331e-06, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, -4.726824e-08, 0, 0, 0, 0.0007324474, -1.48585e-05, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, -6.218539e-06, 0, -1.244392e-05, -0.0001317939, 
    0.0002166405, 0.008075136, 0, 0, 0, 0, 0, 0, 0, 0, 3.904219e-05, 0, 0, 0, 
    0, 0,
  0, 0, 0, -6.947599e-06, 0.0002030726, 0, 0, 0, 0, 0, -1.667745e-05, 
    0.00846437, 0.003115781, 0.004019106, 0.0009368486, 0.0002129918, 
    0.0003704293, 0.0009309053, 0.001363005, 0.00250411, 0.005496522, 
    0.002865284, 0.0004920645, 0, -2.06906e-05, -3.787769e-07, 0.000470624, 
    0.0007487769, 0,
  0, 0, 0, 0, 0, 0, 0.009280074, 0.001362807, 0.006339668, 0.0008706662, 
    0.03547078, 0.02610384, 0.002929782, 0.003476928, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.0005991394, -0.0001088128, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0.0006754693, 0.001608004, -0.0001956011, 0, 
    -1.838414e-05, 0.001761366, -1.396076e-05, -2.754645e-05, 0, 0, 0, 0, 0, 
    0, 0, 0, -0.0002828915, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6.143925e-05, 0, -8.413726e-05, 0.002118088, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    7.062357e-05, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2.29401e-05, 0, 0, 0, 
    -1.185415e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, -3.789182e-05, 0, 0, 0, 0.002535175, -9.631352e-05, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, -1.856363e-05, 0.0001972788, -2.188268e-05, 
    0.000670007, 0.003062993, 0.0118305, -4.431267e-07, -2.4266e-05, 0, 0, 0, 
    0, 0, 0, -4.555637e-05, 0, 0, 0, 0, 0,
  0, 0.0001376049, 0, 4.489469e-05, 0.001844709, 0, 0, 0, 0, -7.236312e-06, 
    -5.28009e-05, 0.01189264, 0.009340597, 0.01088191, 0.001918999, 
    0.001409692, 0.001638925, 0.002913821, 0.005950653, 0.008065159, 
    0.008738504, 0.008176462, 0.004430135, 0, -2.28261e-05, 0.0001570634, 
    0.0008131437, 0.003821552, 0.0004226483,
  0, 0, 0, 0, 0, 0, 0.02426068, 0.0039194, 0.01421744, 0.001179463, 
    0.06395964, 0.04687455, 0.007084331, 0.007223499, -2.969004e-06, 0, 0, 0, 
    0, 0, 0, -1.388265e-05, -7.841987e-06, 0.001007903, -0.0001452343, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0.001576479, 0.00311996, 0.001104591, 0.0002262865, 
    0.0005733153, 0.002986177, 0.0002048386, -5.703494e-05, 4.727015e-05, 0, 
    0, 0, 0, 0, -6.596902e-06, 0, 0.0003082208, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0008845687, -9.724401e-06, 0.004879666, 
    0.005071064, 0.0003955568, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0001520907, 
    -1.642998e-05, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.868039e-06, 0.0002530304, -1.755382e-05, 
    0, 0, 0, 0, 0, 0, 0, 0, 1.347897e-05, -5.459624e-05, -4.108468e-06, 
    0.001989478, -6.050042e-08, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001223503, 0, 
    -4.563156e-06, 0.0002712327, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.005164639, 0.001880931, 0, 0, 
    0.0006156432, 0.001280135, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9.946139e-05, -1.462195e-05, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, -3.434668e-05, 0.0004633008, 0, 0, 0, 0.005437088, 
    0.001084134, 0, 0, 0, 0, 0, 0, 0, -3.452107e-07, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, -8.124457e-06, -4.243408e-06, -5.576159e-05, 
    0.0006654775, 0.001386545, 0.006438669, 0.01026451, 0.01797092, 
    -4.377747e-06, 0.0002429864, 0, 0, 0, 0, 0, 0, -0.0001601965, 0, 0, 0, 0, 0,
  -2.922517e-06, 0.0003205948, -1.263975e-05, 0.0007877595, 0.005754255, 0, 
    -1.891255e-05, -8.477698e-05, -2.210494e-05, -6.682849e-05, 0.004860885, 
    0.01903849, 0.01690854, 0.01917987, 0.003498205, 0.004013139, 
    0.002354892, 0.005879439, 0.01499141, 0.01512846, 0.01382349, 0.01564124, 
    0.009477846, 0, -0.0001030755, 0.003513292, 0.003668943, 0.01200788, 
    0.001223441,
  0, 0, 0, 0, 0, 0.005516998, 0.06695677, 0.01305154, 0.02662143, 
    0.005749776, 0.09777068, 0.06514635, 0.01729619, 0.01141995, 
    -4.737719e-06, 0, 0, 0, 0, 0, -5.468321e-06, -5.441241e-05, 
    -4.710928e-05, 0.0008594771, -0.000212111, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0.003747493, 0.005035531, 0.007809978, 0.001019526, 
    0.0005897277, 0.009255996, 0.009511703, 0.003123751, 0.001805496, 0, 0, 
    0, 0, 0, 0.0001580757, 0, 0.002703699, 0, -4.181559e-07, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 4.387855e-06, 0.0003111984, 0.006367152, 
    -8.584918e-06, 0.01419747, 0.007501562, 0.002291491, -1.030895e-05, 0, 0, 
    0, 0, -3.280895e-06, 0.0001993859, 0, 4.847069e-05, 0.0008980603, 
    0.003959763, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0.0001033828, 0.003790178, 0.0007580266, 
    -2.087398e-05, 0, 0, 0, 0, 0, 0, 0, 0.001274536, 0.002159558, 
    0.002701509, 0.005646841, 0.001391481, 5.167232e-05, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, -4.700647e-06, 0, 0.0001407927, 0, 
    -2.783961e-05, -1.52406e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, -2.003004e-05, 0,
  0, 0, -2.394434e-07, -4.019539e-07, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -3.429497e-05, 0.004611813, -5.881321e-05, -6.670784e-05, 0.0007409515, 
    -2.792044e-05, 0, 0, 0, 0, -8.337207e-08, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01294249, 0.01192356, 
    0.002338709, 0.0011167, 0.002060574, 0.002079786, 0, 0, 0, 0, 0, 
    0.00103843, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.000852009, -6.285207e-05, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, -8.172032e-05, 3.444403e-05, 0.001123708, -3.717363e-07, 
    -2.099676e-05, -2.453797e-05, 0.02132214, 0.004019374, -8.047056e-05, 0, 
    0, 0, 0, 0, 0, -1.860258e-07, 0, 0, 0, 0, -4.892072e-10, 0, 0,
  0, -8.560212e-06, -3.694723e-06, 0, 0, 7.311113e-06, 1.476455e-05, 
    6.356668e-05, -1.784521e-05, 0.0001014465, 0.0009641726, 0.002525612, 
    0.01737639, 0.02334521, 0.02635051, -3.234981e-05, 0.002661986, 0, 0, 0, 
    0, 7.176009e-05, 0, -0.0002344546, -1.878941e-09, -1.676127e-05, 0, 0, 0,
  0.0004524451, 0.002333335, 0.0009836829, 0.007959343, 0.009779528, 0, 
    0.001178256, 0.001563307, 0.001276962, 0.001871678, 0.01001753, 
    0.03591429, 0.03572326, 0.02796761, 0.01268886, 0.01089575, 0.006851308, 
    0.01157747, 0.02418694, 0.02271047, 0.02620289, 0.03662795, 0.02718753, 
    7.810823e-06, -2.800646e-05, 0.01498921, 0.01058683, 0.04475218, 
    0.004582541,
  0, 0, 0, 2.773822e-06, -3.76775e-06, 0.01576406, 0.1016146, 0.03369742, 
    0.06112952, 0.01113806, 0.1337394, 0.1027842, 0.03662008, 0.03170984, 
    -1.495201e-05, 0, -3.869046e-05, 0, 0, 0, -3.405531e-05, 0.002046571, 
    -0.0001271344, 0.002462605, -2.763913e-05, 0, 0, 0, 0,
  0, 0, 0, 0, 0, -6.765873e-06, 0.02346103, 0.009297996, 0.02401189, 
    0.002320722, 0.006442212, 0.02540692, 0.0301429, 0.01420689, 0.003734327, 
    0, 0, 0, 0, 0, 0.0003484835, -2.146713e-05, 0.01208285, 0.000429508, 
    -1.813241e-06, -4.545216e-06, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0.005778482, 0.002721773, 0.01832076, 0.001655139, 
    0.03566513, 0.01330792, 0.008597168, 0.004496753, -1.08646e-05, 0, 0, 0, 
    -1.849614e-05, 0.002268869, 0, 0.0001109004, 0.005566, 0.006708546, 0, 0, 0,
  0, -2.029994e-05, 0, 0, 0, 0, 0, -5.580542e-06, 0, 0.0002317591, 
    -0.0001678206, 0.009001845, 0.006571886, 0.009038785, 0, -1.295184e-05, 
    0, 0, 0, 0, 5.838199e-05, 0.002063119, 0.005390918, 0.006558724, 
    0.01970495, 0.005804842, 0.004941931, -4.141194e-05, 0,
  0, 0, 0, 0, 0, -0.0001295162, -9.099916e-06, -4.120385e-05, 0, 
    0.0002474748, 0.0008376695, 0.007877238, 0.004566151, 0.001704187, 
    -2.737396e-05, 2.552625e-08, -7.437325e-09, 0, 0, 0, 0, 0, -3.497059e-06, 
    -1.163554e-06, 0, -0.0001059993, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8.992914e-09, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0.0001762788, -4.229623e-05, 0, -9.965818e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.002682467, 0, 0, 0, 0, 0, 0, 0, 0, 2.575733e-05, 0, 0, -1.807419e-06, 
    0, 0.0003727373, 0,
  0, 0, -2.605591e-05, 0.001665838, -8.100762e-05, -2.420327e-05, 0, 
    0.0001230266, 0, 0, 0, 0, 0, 0.0004760941, 0.0001294327, 0, 0.0002795268, 
    0.0136219, -0.0002698824, 0.004702603, 0.00764016, 6.635425e-05, 
    0.001278745, 0, 0, 0, -5.848669e-06, -9.834055e-06, -3.38871e-05,
  0, 0, 0, 0, 0, 0, 0, 0, -4.864349e-12, 0, 0, 0, 0, 0, 0.01623799, 
    0.0296455, 0.01168417, 0.00238724, 0.004297304, 0.004747861, 
    -2.607084e-05, 0, 0, 0, -3.653833e-05, 0.00245214, 0, 1.592137e-05, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0004293644, 0.01319632, 
    -0.0001213074, 0.00107071, 0.0001012296, -1.437408e-06, 0, 0, 0, 0, 
    -4.442752e-10, 0.0004694382, 0, 0, 0, 2.06238e-07, 0,
  1.782186e-07, 0, 0, 0, 0, 0, -4.536528e-05, 0.003981834, 0.001459856, 
    9.535122e-06, 0.0003718219, 0.006107567, 0.03999959, 0.01941706, 
    -0.0001041519, 0, 0, 0, 0, 0, -2.084042e-08, -1.947771e-07, 0, 
    0.0004193676, -1.345481e-07, 3.752604e-07, 1.584049e-08, 0, 0,
  -1.079602e-05, -1.97062e-05, -2.986569e-05, 1.987748e-07, -3.04234e-07, 
    0.001161354, 0.001944231, 0.003523564, 0.000261255, 0.004653475, 
    0.007012425, 0.008581677, 0.03803472, 0.05638516, 0.03281837, 
    0.0001002889, 0.003930574, 0, 0, -8.102423e-08, 0, 0.001654451, 
    3.822326e-08, 0.002511052, -1.60079e-05, -0.0001413762, -2.303923e-06, 
    -1.376821e-09, 0,
  0.003552187, 0.004743248, 0.003494937, 0.02054979, 0.01146712, 5.79844e-06, 
    0.01266109, 0.009626685, 0.008517086, 0.0132176, 0.02558063, 0.07341082, 
    0.09385099, 0.04810854, 0.03494493, 0.02453109, 0.01465241, 0.02097778, 
    0.03738094, 0.03262697, 0.04487862, 0.0562309, 0.05724802, 0.0008891657, 
    0.005467962, 0.03829711, 0.02370473, 0.08983359, 0.00932215,
  0, 0, 0.0002839758, 0.0008788122, 0.0005658746, 0.1079858, 0.156628, 
    0.1403124, 0.1212239, 0.04465181, 0.2076851, 0.1608419, 0.08986003, 
    0.05028285, -6.829656e-05, -1.666436e-06, 0.0005576788, 0.006567571, 0, 
    -2.623197e-08, -0.0002067861, 0.005944473, -0.0001373638, 0.01285619, 
    -0.0001206509, 0, 0, 0, 0,
  0, -6.174647e-07, 0, 1.20743e-06, -1.172033e-06, -0.0001619029, 0.1640414, 
    0.02061147, 0.03501025, 0.06698795, 0.02447334, 0.0420013, 0.08032356, 
    0.03122638, 0.01572666, 0.0003176497, 0, 0, 0, 0, 0.0002960222, 
    0.001219714, 0.05640476, 0.0005185692, 0.0001258706, -4.661581e-05, 0, 0, 
    -8.609346e-05,
  0, 6.872423e-06, -7.4021e-05, 0, -4.905631e-09, 2.968995e-06, 
    -8.509742e-10, 3.511265e-10, 0.0151889, 0.00610084, 0.04918268, 
    0.01180731, 0.0688106, 0.04082193, 0.01578525, 0.01152615, -6.062925e-05, 
    0, 0, 0, 0.001184455, 0.005325648, 0.002543789, -9.835403e-05, 0.0106415, 
    0.01256683, 0.0003286779, 0, 0,
  0, -4.678657e-05, 0, 0.001080067, -7.158734e-07, -1.107811e-05, 
    -6.298503e-07, 0.0007070848, 0.00152249, 0.004072124, 0.007639678, 
    0.03722601, 0.02792483, 0.02528142, -1.083921e-05, -4.709251e-05, 
    0.0005735728, 0, 0, 0, 0.005030392, 0.005414588, 0.009939325, 0.02012805, 
    0.03944101, 0.02040493, 0.01240453, 0.006222283, 0,
  0, 0, 0, 0, -9.050358e-05, -0.000151535, 1.486193e-05, 0.002128899, 
    -0.0006078418, 0.007104998, 0.005802928, 0.02504925, 0.01565741, 
    0.005330005, -4.550687e-05, 1.697304e-07, 0.0004797651, 0, 0, 0, 
    -2.017386e-05, -5.048061e-06, -0.0001162154, -6.10377e-06, -4.617824e-05, 
    0.00214931, 2.939659e-05, 0, -7.090023e-05,
  0, 0, 0, 0, -7.926265e-05, 0, 0, -2.620212e-06, 0.002657401, 0.000723612, 
    0, -2.427672e-05, 0, -4.388082e-06, -2.357685e-05, 0, 0, 0, 0, 0, 0, 0, 
    -2.134458e-05, 0, 0, 0, 0, 0, -4.499013e-05,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, -1.661794e-05, 0, 0, 0, -1.252192e-05, 0, 0, 0, 
    0, 0, 0, 0, 0, -3.367939e-05, 0, 0, 0, 0, 0, 0,
  0.003311124, 0.003706268, -6.28613e-07, -7.916218e-05, 1.283343e-05, 
    -5.034168e-05, -1.017747e-06, 0, 0, 3.311539e-05, 0, 0, -3.303785e-06, 
    0.004764292, 0, 0, 0, 0, 0, 0, -3.008775e-05, 0, 0.002198206, 
    -9.258125e-06, 0, 0.0010733, 0, 0.002540175, 0,
  -0.0001454081, 0, 4.798028e-06, 0.006483726, 0.004169419, -6.262999e-05, 
    -8.291546e-05, 0.00869623, 2.683007e-05, -2.134151e-10, 0, -3.977579e-12, 
    0, 0.006692448, 0.0024512, 0.0003199274, 0.004695989, 0.03114854, 
    0.008360047, 0.01929272, 0.02841163, 0.003047283, 0.001985769, 
    -6.544934e-07, -6.163474e-06, 0, 1.850244e-05, 3.146288e-05, 0.002809272,
  0.002535769, 0, 0, -7.259366e-09, -0.0001704931, 0, 0.001066188, 
    -2.099334e-09, -4.023896e-06, 1.526007e-07, 2.694769e-09, -3.688057e-09, 
    0, -1.056586e-06, 0.02223909, 0.06520909, 0.04037989, 0.01567744, 
    0.01748785, 0.01611078, 0.001691632, 0, 0, 0, 0.0008298552, 0.002777549, 
    1.472479e-05, 0.007980067, -3.181688e-06,
  -7.248552e-07, -3.789936e-11, 0, 5.09947e-09, 0, 1.752028e-08, 6.07801e-07, 
    7.844241e-06, 1.198745e-06, 2.181236e-07, 7.7872e-07, 3.033683e-07, 
    0.002471176, 0.03117898, 0.00325353, 0.00834275, 0.005104079, 
    0.0005493409, 4.177554e-06, 0, 0, -5.816984e-06, -5.33344e-06, 
    0.0007671958, 0, 0, 3.897958e-05, 3.368932e-06, -3.089379e-07,
  0.0001141715, 7.925149e-09, 0, 0, 0, 6.403773e-07, 0.0002700512, 
    0.02935988, 0.002350533, 0.00389712, 0.007349081, 0.02919992, 0.08162378, 
    0.1075807, 0.01502933, 8.067733e-07, -3.207303e-05, 9.145056e-09, 0, 0, 
    -1.146691e-05, 0.001034456, 1.36421e-05, 0.0001016586, 0.000273961, 
    0.001001735, -2.673537e-06, 4.207835e-06, 8.179735e-10,
  8.678203e-05, 0.000103032, 0.0001012028, 0.0001772854, 3.909007e-06, 
    0.004998447, 0.01590715, 0.05824615, 0.00120054, 0.02030612, 0.1724261, 
    0.2801974, 0.1827772, 0.1916786, 0.1289465, 0.0004315297, 0.008900394, 
    1.136349e-05, 2.052441e-06, -1.134513e-06, 2.824832e-06, 0.004342062, 
    -8.332656e-07, 0.01303612, 0.001895845, -0.0002316925, -1.234699e-05, 
    5.634897e-05, -3.692982e-06,
  0.01461315, 0.02034537, 0.01852738, 0.02724013, 0.01943077, 0.01343044, 
    0.2115763, 0.5048127, 0.4200841, 0.3551604, 0.3461486, 0.3674308, 
    0.322501, 0.2367308, 0.1624757, 0.09083331, 0.04423827, 0.08815744, 
    0.1188724, 0.09806691, 0.131298, 0.1321331, 0.1265633, 0.02524571, 
    0.01706997, 0.06032063, 0.03759809, 0.1364621, 0.0315036,
  1.413427e-05, 0.0001393962, 0.0045976, 0.01681546, 0.1557019, 0.1989823, 
    0.3246053, 0.1497194, 0.3872986, 0.1345125, 0.3476554, 0.2735767, 
    0.2616019, 0.09468197, 0.002500925, 0.0009387957, 0.001602737, 
    0.01255274, -4.556838e-06, -2.092267e-05, 0.01285984, 0.07084312, 
    0.003696087, 0.04071485, 0.003604172, -1.431902e-07, 0, 5.80309e-07, 
    7.68278e-05,
  -2.804598e-11, -6.904737e-05, -2.393078e-09, 3.273866e-06, 0.0007824103, 
    0.00305851, 0.1272031, 0.03080701, 0.05454367, 0.125347, 0.06493344, 
    0.1556427, 0.2772499, 0.1286449, 0.04923804, 0.01314277, -5.917155e-07, 
    0.00037722, -3.386767e-11, 0.000131474, 0.005108346, 0.0224381, 
    0.2019198, 0.03387262, 0.002738313, 0.0001352231, -2.389785e-07, 0, 
    0.002401103,
  1.218747e-08, 0.003173276, 0.0003162043, -1.252587e-10, 1.294028e-07, 
    3.180052e-05, -3.501493e-07, -4.532394e-05, 0.03584703, 0.05548437, 
    0.1619724, 0.1022207, 0.1573303, 0.09442831, 0.05768564, 0.03389199, 
    0.001223648, 0.000912696, -2.752181e-06, 0, 0.001243041, 0.009576556, 
    0.01100448, 0.004510919, 0.02088426, 0.01776913, 5.724666e-05, 
    -3.062439e-05, 0,
  -4.562987e-05, -8.198916e-06, 2.449489e-06, 0.005330303, 0.0001423614, 
    0.002199926, 0.0002216308, 0.004488032, 0.009346136, 0.006229437, 
    0.01564057, 0.07543732, 0.08582463, 0.07729958, 0.0324804, 0.003157102, 
    0.002868925, 0.001453483, 0.002143434, 0, 0.007646037, 0.01141385, 
    0.01722163, 0.03410749, 0.05200616, 0.04881223, 0.0256404, 0.01095676, 
    0.002145847,
  -3.081081e-09, 0, 0.0001061039, -1.023765e-05, 0.01015409, 0.01077153, 
    2.978741e-05, 0.01866242, -0.001514381, 0.01826051, 0.0115761, 
    0.03679036, 0.03610884, 0.02232292, 0.000373237, -0.0001198468, 
    0.001161789, 0, -3.110301e-08, 0, -0.0002237537, -3.216742e-05, 
    0.001251815, 0.00129264, -0.0003931711, 0.004788273, 0.005913823, 
    -9.623852e-05, 0.001609454,
  0, 0, 0, 0, 0.0005822234, -5.982965e-05, 0.0001610334, 3.050467e-05, 
    0.005149806, 0.001721388, 7.276926e-06, -4.24394e-05, -0.000326774, 
    2.910765e-05, 0.002230137, 0, 0, 0, 0, 0, 0, 0.0005068814, 0.0004908458, 
    -2.982372e-05, 0, 0, 0, -2.861259e-07, 0.001916011,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, -3.765411e-05, 0, 0, 0, -2.504384e-05, 0, 
    1.234681e-05, 0, 0, 0, 0, 0, -3.590361e-06, 0.007405255, -3.533451e-05, 
    0, 0.0009830742, -3.47601e-05, 0, -2.415013e-05,
  0.004997895, 0.01008977, 0.002748933, 0.00300405, 0.0003446835, 
    0.001545624, 0.00126449, 0.0004656149, 0.001492765, 0.0004265535, 
    7.227373e-05, 0, -1.669641e-05, 0.005017828, 0.0004787359, 0, 0, 0, 0, 
    -1.078186e-05, 0.001677731, 4.070203e-06, 0.008746437, 0.002375735, 0, 
    0.003093804, -9.597838e-06, 0.007876838, 8.470886e-06,
  0.005769238, 0, 0.004304593, 0.02305552, 0.02010026, 0.004796817, 
    0.003387797, 0.01257673, 0.0006699455, 4.209747e-06, -4.282081e-05, 
    -1.252798e-05, -1.128763e-05, 0.009846429, 0.01029501, 0.004794996, 
    0.01336559, 0.05310992, 0.02864052, 0.041162, 0.06460004, 0.01574712, 
    0.007341051, -2.545688e-05, 0.002702848, -1.978809e-07, -0.0001455867, 
    0.003931769, 0.0118987,
  0.01733702, -2.816758e-06, 0.000751406, -1.738564e-07, -7.52826e-05, 
    7.137354e-05, 0.009541092, 6.405926e-09, 3.763298e-05, 2.367401e-06, 
    4.879563e-06, -1.803142e-06, -1.857448e-08, -6.834754e-05, 0.04138709, 
    0.1310723, 0.09727878, 0.0419454, 0.05367801, 0.0369624, 0.00717484, 
    0.0002043677, 2.636033e-05, -4.647474e-07, 0.003437898, 0.003317301, 
    5.031152e-05, 0.02469626, 0.002424895,
  0.0002230556, 0.001533086, 0, 5.05499e-07, -2.442127e-11, 0, -7.016756e-07, 
    6.710159e-06, 2.500818e-07, 4.552101e-08, 3.21575e-07, 1.151981e-06, 
    0.001473365, 0.05426798, 0.03498132, 0.06132545, 0.03709366, 0.01229562, 
    0.009151012, -6.520027e-06, -2.991651e-09, 2.045224e-05, 0.00555556, 
    0.0004642414, 0.01511135, -5.701571e-07, 0.003953077, 0.0006166633, 
    1.186801e-05,
  0.007291486, -2.839141e-05, 3.231284e-05, -7.763354e-09, 4.360633e-08, 
    8.732673e-05, 0.07115214, 0.07124776, 0.003698175, 0.01069466, 
    0.01711163, 0.03160019, 0.09183551, 0.1151853, 0.01808211, 6.065735e-05, 
    -5.272174e-05, 1.316483e-07, 3.800566e-08, -2.37531e-09, 8.065868e-05, 
    0.005218796, 1.742378e-05, 0.03299342, 0.02036639, 0.01415872, 
    0.0003747215, 0.02836001, 0.0161887,
  0.01109751, 0.06973586, 0.1945474, 0.01733859, 0.01166599, 0.03873343, 
    0.2079234, 0.3812582, 0.1379707, 0.4092163, 0.2149495, 0.270796, 
    0.1433786, 0.1519724, 0.1099954, 0.0001619911, 0.009857835, 1.201556e-05, 
    3.373728e-05, -8.400017e-05, 0.002615265, 0.02433028, 0.0006218035, 
    0.04598448, 0.02910015, 0.009392165, 0.01263338, 0.07708835, 0.02508802,
  0.1896576, 0.3164671, 0.3563547, 0.03961189, 0.05167792, 0.02819913, 
    0.2433646, 0.5020753, 0.368412, 0.2329828, 0.261601, 0.3009609, 0.279681, 
    0.1817862, 0.2193549, 0.1521563, 0.06071734, 0.1005297, 0.1426969, 
    0.1303347, 0.2199166, 0.2290065, 0.3996212, 0.1619765, 0.09360505, 
    0.1603789, 0.08293732, 0.2762375, 0.3100674,
  0.002304302, 0.0006912366, 0.002110851, 0.02473275, 0.1421606, 0.2187144, 
    0.3212684, 0.1221859, 0.3967678, 0.1190754, 0.3271185, 0.2246025, 
    0.2352231, 0.1344383, 0.1139528, 0.06211125, 0.05681775, 0.09941343, 
    0.003140542, 0.005145196, 0.0210638, 0.09919591, 0.07107449, 0.1015683, 
    0.1002941, 0.006383257, 0.001051555, 0.01016515, 0.002603062,
  0.00160397, 0.001234713, 0, 2.136047e-06, 0.01514537, 0.003871831, 
    0.08959877, 0.05398087, 0.09081387, 0.09384304, 0.05309939, 0.1141245, 
    0.3363467, 0.2808177, 0.2261212, 0.05043139, 0.02342801, 0.01796843, 
    0.003511715, 0.003341652, 0.05034491, 0.1398124, 0.2733876, 0.2101427, 
    0.1186211, 0.09304833, 0.0001655857, 1.711062e-05, 0.01244291,
  0.004424498, 0.009137676, 0.002544341, -1.283486e-07, 5.180592e-07, 
    -5.255835e-07, 5.540767e-07, 0.006923228, 0.06370121, 0.1740445, 
    0.2287424, 0.1600429, 0.2749702, 0.1829689, 0.07466482, 0.1033669, 
    0.0428558, 0.05810714, 0.005795237, 8.108807e-06, 0.002471575, 0.1096826, 
    0.1024169, 0.1183482, 0.103639, 0.09663263, 0.04482479, 0.01055795, 
    0.001587903,
  0.003700919, 0.0001908688, 0.0003490002, 0.01550862, 0.01925142, 
    0.02118443, 0.005235905, 0.007950686, 0.01307026, 0.01155539, 0.033556, 
    0.1887297, 0.1537543, 0.1864566, 0.1608708, 0.1012157, 0.07462866, 
    0.04571921, 0.02070213, 0, 0.01026839, 0.02288297, 0.0282483, 0.07062474, 
    0.1246073, 0.1246566, 0.08052147, 0.02450869, 0.01641002,
  5.737486e-05, 1.069532e-05, 0.0005452425, 0.0005528031, 0.01711321, 
    0.01677512, 0.01492253, 0.08873424, 0.01119624, 0.02864683, 0.0182466, 
    0.05198845, 0.09652048, 0.1055108, 0.07959504, 0.04170112, 0.006900629, 
    -8.874741e-05, -1.462594e-05, 0.003031576, 0.002472029, 0.0003813927, 
    0.004632617, 0.002750454, -0.0008005302, 0.02386038, 0.0499048, 
    0.02592661, 0.00549137,
  -3.626713e-05, 0.0002523622, -4.325601e-05, 0.002737256, 0.003868374, 
    0.001102975, 0.003331579, 0.001049918, 0.01124643, 0.008999045, 
    0.000263949, 0.001631824, 0.007198213, 0.02541541, 0.02943451, 
    0.003782746, -3.540638e-06, -9.919708e-09, -1.942714e-05, -1.107037e-06, 
    0.001007225, 0.002277442, 0.01159213, 0.003289116, 1.502316e-05, 0, 
    -8.459752e-07, 0.001020218, 0.007548573,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2.377861e-09, -4.198415e-06, 
    -2.892306e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -6.797101e-05, 0.002177022, 
    0.0001542102, 0, 0, 0, 0, 0, 0, 0, -3.155488e-05, 0, 0, 0, 0, 0,
  -7.782054e-05, -5.224259e-07, -3.611115e-06, -2.145057e-06, 0, 0, 0, 0, 0, 
    -3.772381e-05, 3.843028e-05, -8.409232e-05, 0, 0.000528163, 1.489162e-05, 
    0.0003837064, 0, 0, 0, 0, 0, -1.419945e-05, 0.01078923, 0.006060364, 
    -5.666232e-05, 0.001667921, -4.23221e-05, 0, -5.461966e-05,
  0.009929203, 0.01690405, 0.006280002, 0.01121526, 0.003264417, 0.007417372, 
    0.004720997, 0.00299369, 0.00899701, 0.007367638, 0.007346666, 
    -6.833619e-05, -2.741248e-05, 0.005774882, 0.01526907, 0, -2.1283e-06, 0, 
    0.00197347, -4.342036e-05, 0.005163949, 0.01018195, 0.0238316, 
    0.01074513, 0.0003926987, 0.005067551, -6.424593e-05, 0.01565997, 
    0.007721891,
  0.01679822, -0.0001108111, 0.01198136, 0.03334731, 0.03507973, 0.02165777, 
    0.01194671, 0.01916042, 0.01051467, 0.01169839, 0.0004585949, 
    9.396679e-05, -0.0002291494, 0.01163683, 0.03589231, 0.02803731, 
    0.03872331, 0.07107214, 0.05590286, 0.07104263, 0.1061558, 0.04543018, 
    0.02496803, -0.0001373598, 0.005480977, 0.002883012, 0.001005316, 
    0.01154654, 0.02660427,
  0.005116649, 0.00133357, 0.00192171, 6.940064e-05, 0.001340296, 
    0.003053527, 0.01697125, 1.477949e-07, 0.005966074, 0.0003432972, 
    0.0008913651, 0.001466195, -1.787057e-05, 0.001718122, 0.07553124, 
    0.1799271, 0.1835369, 0.2097973, 0.179245, 0.1940784, 0.1115935, 
    0.04729268, 0.01544623, -2.884958e-05, 0.005825225, 0.01272464, 
    0.007817396, 0.04865678, 0.0006625202,
  1.805171e-06, 0.0001505827, 2.202669e-06, 5.786396e-07, -3.675062e-10, 0, 
    -1.324543e-05, 1.350538e-06, 9.525143e-08, 3.106902e-07, 3.195169e-07, 
    9.415752e-07, 1.198621e-05, 0.05792637, 0.05009044, 0.07521088, 
    0.04532911, 0.0274657, 0.01199191, 0.003161692, 0.0001092307, 
    -4.099534e-06, 0.0006448762, -1.113577e-06, 0.0020819, 0.007815426, 
    0.0004164683, 7.772706e-05, -0.0001074373,
  0.000615061, -3.16819e-07, 2.575003e-05, 1.128997e-09, 1.08429e-08, 
    4.72342e-05, 0.03746836, 0.04879901, 0.004422716, 0.003671527, 
    0.00966026, 0.02195081, 0.1010995, 0.1099743, 0.008301176, 0.000204938, 
    5.793918e-06, 1.191865e-08, 1.649182e-08, 0, 1.01944e-05, 0.0007984589, 
    3.507739e-05, 0.04417666, 0.003662826, 0.003015669, 0.004764284, 
    0.02004841, 0.000467992,
  0.004387743, 0.03254641, 0.1067114, 0.01084873, 0.003479085, 0.01706746, 
    0.1356611, 0.2523268, 0.08116747, 0.3457611, 0.1592309, 0.2160627, 
    0.123992, 0.1317806, 0.08244979, 0.0002605421, 0.01005976, 4.812769e-07, 
    1.755281e-05, 1.945291e-05, 6.52144e-05, 0.02388756, 0.003611645, 
    0.03908293, 0.01301865, 0.004883323, 0.01088334, 0.04917068, 0.02463305,
  0.1303897, 0.275056, 0.3114762, 0.1690706, 0.04155293, 0.00631445, 
    0.1568402, 0.4161921, 0.322546, 0.126767, 0.1957363, 0.2553411, 
    0.2839445, 0.1468977, 0.1377279, 0.1208202, 0.03802374, 0.06885883, 
    0.09388506, 0.09176905, 0.1592578, 0.1852002, 0.3313145, 0.09640259, 
    0.0585541, 0.1250979, 0.07105335, 0.2462837, 0.2325677,
  0.0002948885, 1.290909e-05, 0.001540515, 0.03280275, 0.1477968, 0.2279613, 
    0.3335218, 0.09610019, 0.4043781, 0.118884, 0.3040932, 0.2023912, 
    0.1998093, 0.1147053, 0.07528671, 0.05636414, 0.02336753, 0.05808853, 
    0.01068153, 0.004947087, 0.01502612, 0.05556765, 0.047831, 0.06859775, 
    0.06212114, 0.002629478, 0.0001557054, 0.007175948, 0.001836066,
  0.01878209, 0.008339281, -3.478771e-08, 1.973965e-06, 0.006788534, 
    0.001312109, 0.07614331, 0.1415153, 0.1327406, 0.08456755, 0.04701028, 
    0.09373911, 0.2900227, 0.2649984, 0.2102402, 0.173705, 0.1498033, 
    0.01537336, 0.02070716, 0.002283651, 0.1123398, 0.1458628, 0.179044, 
    0.1480662, 0.09500748, 0.09100778, 0.008207573, -0.00010503, 0.03649233,
  0.07668594, 0.04943966, 0.00708817, 6.351954e-05, 1.077629e-05, 
    5.421459e-07, 6.10606e-06, 0.01934836, 0.09742226, 0.1830325, 0.1802155, 
    0.1195868, 0.2674761, 0.2189578, 0.089986, 0.2131165, 0.1135501, 
    0.1401112, 0.008083697, 0.009681066, 0.04934508, 0.09983067, 0.08316147, 
    0.1107161, 0.1110854, 0.1110776, 0.1626669, 0.1039397, 0.04196738,
  0.04531786, 0.008239051, 0.00295159, 0.03744152, 0.05892623, 0.06719326, 
    0.0215132, 0.02174511, 0.02993888, 0.05979269, 0.1177901, 0.2443594, 
    0.2074196, 0.2027213, 0.2072903, 0.1781254, 0.1099966, 0.07224984, 
    0.08036268, 0.005099773, 0.04280003, 0.1057478, 0.09437398, 0.1290809, 
    0.1621765, 0.1678345, 0.1392203, 0.1109954, 0.07779676,
  0.06908289, 0.0169632, 0.01126723, 0.009860572, 0.01961753, 0.03513796, 
    0.07969813, 0.17751, 0.08744002, 0.08929168, 0.07070779, 0.1459441, 
    0.2137088, 0.1484524, 0.1043251, 0.0924072, 0.04600183, 0.0420618, 
    0.002100948, 0.01883325, 0.0115859, 0.01032716, 0.02581957, 0.01580576, 
    0.0257408, 0.05500497, 0.07867012, 0.0830196, 0.07310948,
  0.02033776, 0.00170011, 0.002024278, 0.005395428, 0.01110559, 0.01002553, 
    0.02925233, 0.05393535, 0.05759883, 0.05105656, 0.03298813, 0.03251905, 
    0.02059732, 0.09035941, 0.05815836, 0.03104685, 0.01326017, 0.003418212, 
    0.005154031, 0.005028402, 0.007291919, 0.005995872, 0.023324, 0.0113341, 
    0.002525733, 0, 4.691778e-06, 0.01788063, 0.02753977,
  0.0003722826, -0.0001213788, 1.912137e-05, 0, -0.0001514097, 0.002470593, 
    0.0006898592, 0.006157306, 0.001358047, -0.0001413086, 0, -1.868563e-06, 
    -8.980042e-06, -9.736249e-13, 5.926786e-07, 7.159558e-05, -0.0001020808, 
    -5.743989e-05, -2.594481e-10, -3.380612e-09, 0, 0, -3.910572e-06, 
    8.317669e-06, -5.26471e-07, 0, 0, -1.266017e-07, -3.278077e-05,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0.0004570957, -1.224161e-05, -6.571705e-07, 0, 0, 0, 0, 0, 0, 
    -1.153697e-05, -2.188027e-05, 0, 0, -0.0001214064, 0.004429416, 
    0.002173402, 0, 0, 0, 0, 0, 0, 0, 0.0002198435, 0.00259037, 0.0001587242, 
    -3.229779e-06, 0, 0,
  0.000209943, 0.002734302, 0.0006366629, 0.0008903795, 0, 0, 0, 
    6.023765e-06, 0, 0.0008692254, 0.0007530207, 0.004205023, 0.00330498, 
    0.006251751, 0.001613427, 0.002256141, 0.0002031148, 0, 0, 0.0005945398, 
    0, -2.83989e-05, 0.01993833, 0.02022206, 0.0008344341, 0.006012806, 
    0.009559529, 0.0004700672, -0.0001201145,
  0.025465, 0.03916915, 0.01357786, 0.02521553, 0.01277239, 0.01641542, 
    0.005631629, 0.006087118, 0.01981656, 0.03120768, 0.02706319, 
    0.008213017, 0.002501206, 0.006163338, 0.02193064, 0.0003063721, 
    0.0003779769, 0.0003492042, 0.005295906, 0.01146194, 0.0220263, 
    0.04281238, 0.0765807, 0.04567027, 0.007189944, 0.01626136, 0.0007987912, 
    0.02301689, 0.03150997,
  0.05505132, 0.02445546, 0.02200607, 0.05348443, 0.05032658, 0.03335393, 
    0.02696526, 0.03165041, 0.04557042, 0.02702647, 0.008253162, 0.02070731, 
    0.008907436, 0.01983079, 0.0503437, 0.06490634, 0.05859921, 0.09573849, 
    0.0914444, 0.1293635, 0.163363, 0.1302308, 0.1524805, 0.002906353, 
    0.02775278, 0.03418186, 0.02741421, 0.03816424, 0.08398675,
  0.0007294529, 1.979913e-05, 0.002525837, 0.003513594, 0.007070043, 
    0.01039337, 0.0177327, -4.590772e-05, 0.006446204, 0.003704931, 
    0.02208453, 0.01232525, 0.002755862, 0.01225351, 0.08999176, 0.2027574, 
    0.2012301, 0.1887074, 0.2300429, 0.2366566, 0.1553838, 0.06839827, 
    0.02340217, 0.0001951762, 0.009902279, 0.03957289, 0.03869067, 
    0.08323538, 0.0005049198,
  6.939222e-07, 5.485914e-05, 1.312778e-07, 5.048732e-07, -2.576899e-11, 
    -8.675887e-11, 0.000177693, 3.703095e-06, 1.038251e-07, 8.532759e-09, 
    3.53598e-07, 9.05367e-07, 0.001551969, 0.0548136, 0.06523357, 0.07105223, 
    0.04921236, 0.02833553, 0.01178335, 0.001738762, 1.06459e-05, 
    -5.497093e-07, 8.521138e-05, 2.396365e-06, 0.0002171932, 0.0001409441, 
    3.335242e-05, 1.04936e-07, -3.798808e-07,
  4.202571e-05, 3.35832e-07, 1.979103e-06, -7.914632e-10, -2.982359e-10, 
    1.947356e-05, 0.01580483, 0.03893176, 0.005655798, 0.01001588, 
    0.008764671, 0.004210231, 0.1107971, 0.09997758, 0.01027292, 
    0.0004392668, 0.0003792788, -3.48066e-11, -1.480643e-09, -1.065616e-09, 
    5.076e-07, 0.0006932988, 1.079206e-06, 0.03814777, 5.812934e-05, 
    0.0001511594, 0.0001969702, 0.00883447, 9.320822e-05,
  0.002736944, 0.01010622, 0.05751846, 0.00350885, 0.0003168762, 0.01412775, 
    0.05879282, 0.1207967, 0.05965385, 0.2658007, 0.1245452, 0.1887507, 
    0.1193348, 0.1237422, 0.0665746, 0.0007152508, 0.008697631, 1.093672e-06, 
    1.283445e-05, 0.002209034, 8.864853e-06, 0.01180495, 0.0007476903, 
    0.03945484, 0.01368938, 0.006735562, 0.02064543, 0.03425501, 0.008260514,
  0.1126864, 0.2696992, 0.2923191, 0.1395025, 0.04686907, 0.005492663, 
    0.1241649, 0.2603641, 0.3051794, 0.09634786, 0.1561524, 0.2244263, 
    0.2621857, 0.1349202, 0.09524026, 0.09075214, 0.0380925, 0.06068778, 
    0.08178178, 0.08175628, 0.1259272, 0.1700055, 0.2885486, 0.08029516, 
    0.05660223, 0.1072068, 0.06718194, 0.2249213, 0.18212,
  0.001216152, 1.311012e-05, 0.0004389511, 0.04058949, 0.1563636, 0.2450462, 
    0.3571401, 0.08427345, 0.3946447, 0.09709056, 0.2878497, 0.188261, 
    0.173704, 0.1024397, 0.05262281, 0.04867479, 0.009296229, 0.03476504, 
    0.0123854, 0.003805554, 0.008753616, 0.04554932, 0.03888701, 0.05853637, 
    0.04421468, 0.001819236, 0.0001087651, 0.004914534, 0.002240512,
  0.01253012, 0.01472797, -2.500713e-08, 9.232189e-07, 0.0003534002, 
    0.0002468908, 0.05410605, 0.1407889, 0.1385254, 0.06501216, 0.04108923, 
    0.07849351, 0.2763989, 0.2551247, 0.2107809, 0.1618611, 0.1213581, 
    0.008490068, 0.001454079, 2.265006e-05, 0.1150013, 0.1649494, 0.1340583, 
    0.1352479, 0.08324671, 0.05667194, 0.02170937, -3.062786e-05, 0.03348753,
  0.108873, 0.07061797, 0.01513991, 0.001055713, 0.000287917, 3.608186e-07, 
    9.320053e-06, 0.06044916, 0.1675286, 0.1780262, 0.1331813, 0.08728632, 
    0.2353541, 0.22561, 0.08167277, 0.2042367, 0.1447606, 0.1270605, 
    0.006537124, 0.01081587, 0.1039134, 0.07726569, 0.06889457, 0.1087165, 
    0.1209133, 0.09215028, 0.1376008, 0.07682995, 0.06048714,
  0.1082496, 0.09528967, 0.05537981, 0.204083, 0.1208987, 0.1705034, 
    0.108602, 0.07473686, 0.1162911, 0.1450002, 0.09733376, 0.2189495, 
    0.2037071, 0.1591535, 0.1938559, 0.230402, 0.1487483, 0.09982128, 
    0.1173034, 0.05490564, 0.07335141, 0.1270853, 0.1233698, 0.1525232, 
    0.1588756, 0.1685549, 0.1368276, 0.1444533, 0.09062897,
  0.126065, 0.1224129, 0.08108628, 0.09152155, 0.1075111, 0.1241013, 
    0.1802656, 0.2979858, 0.1769934, 0.1682747, 0.1201014, 0.2557065, 
    0.2733824, 0.1795253, 0.115862, 0.1133242, 0.1056919, 0.1400469, 
    0.07941505, 0.1131449, 0.07234583, 0.08737481, 0.09211881, 0.06566107, 
    0.1059818, 0.09777865, 0.105268, 0.1666397, 0.2040845,
  0.0999102, 0.09283518, 0.09423015, 0.06104857, 0.05533126, 0.04148327, 
    0.05305089, 0.07535153, 0.1244296, 0.1566454, 0.08058819, 0.03437912, 
    0.1081209, 0.1845883, 0.1436657, 0.1487943, 0.1265061, 0.07954372, 
    0.03776034, 0.02241971, 0.01096232, 0.02186535, 0.03186971, 0.03259239, 
    0.02732349, -0.0001463751, 0.001239303, 0.1334361, 0.1286188,
  0.01037244, 0.01800403, 0.02342978, 0.01323268, 0.001942684, 0.02871606, 
    0.009491215, 0.0140173, 0.01014964, 0.001756925, 0.03563028, 0.07055202, 
    0.06102526, 0.06554796, 0.02754235, 0.0334697, 0.03759678, 0.04319886, 
    0.03799191, 0.03237258, 0.008869038, 0.002928424, 0.0001197175, 
    -0.0009473164, 0.00121198, 0.0003077658, -0.0003805066, -0.002351096, 
    0.0277497,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0001893045, 0, 0, 0, 0, 0,
  0.002783546, 0.006327305, 0.005528532, 0.0005743282, -0.0001217364, 0, 0, 
    0, 0, -2.307395e-05, -4.376053e-05, 0, 0.001357814, -0.0001908352, 
    0.01555108, 0.007888172, 0, -2.936371e-05, 0, -2.469644e-06, 0, 
    0.002192683, -1.034569e-05, 0.003511951, 0.01431796, 0.00789043, 
    0.003553004, 0, 0,
  0.02856104, 0.03565698, 0.03564135, 0.03141202, -1.512165e-05, 
    -4.852383e-06, 0, 9.908135e-05, 2.935406e-05, 0.004393737, 0.008263066, 
    0.009002537, 0.008979709, 0.01467026, 0.01506855, 0.01310856, 
    0.004038169, 0.005017293, 0, 0.002256945, -1.541276e-05, -0.0002643421, 
    0.02277894, 0.03601475, 0.02160856, 0.02266213, 0.01805369, 0.01025683, 
    0.01547056,
  0.1005492, 0.0901259, 0.07852981, 0.0861755, 0.04642895, 0.04270079, 
    0.0101794, 0.02229617, 0.03626435, 0.0629207, 0.04601372, 0.02325682, 
    0.02339514, 0.006761429, 0.043833, -0.0002512302, 0.01029628, 0.03127948, 
    0.02733967, 0.045183, 0.06424923, 0.1053949, 0.1639623, 0.1217366, 
    0.09579777, 0.1234919, 0.06495385, 0.04663298, 0.07529835,
  0.09375394, 0.09178737, 0.08405849, 0.09226181, 0.1092114, 0.09616726, 
    0.08707014, 0.0646947, 0.06871719, 0.05765259, 0.046727, 0.04189295, 
    0.02882685, 0.03244415, 0.07138133, 0.10115, 0.0850397, 0.1205471, 
    0.09862323, 0.1323511, 0.2124779, 0.1775382, 0.1829584, 0.07159851, 
    0.111875, 0.1071291, 0.05569885, 0.1126255, 0.1488799,
  -0.0001106212, 0.002543527, 0.003394897, 0.01512164, 0.006284994, 
    0.01093393, 0.01937415, 0.001792924, 0.002585602, 0.003098866, 
    0.04838292, 0.02285134, 0.003512602, 0.01631785, 0.08926596, 0.205378, 
    0.1980165, 0.1584248, 0.2025135, 0.1838346, 0.1210401, 0.04265872, 
    0.00535169, 0.0003230863, 0.0144755, 0.04859594, 0.05155434, 0.09003446, 
    0.001699353,
  1.187272e-07, 1.007498e-05, 3.879242e-07, 8.402322e-08, 0, -1.335918e-10, 
    6.488971e-07, 4.203118e-06, 6.783969e-08, -3.271917e-09, 1.407105e-07, 
    -4.694602e-05, 0.01515401, 0.07670143, 0.0831136, 0.08194999, 0.02551843, 
    0.0183407, 0.004714693, 0.001310168, 3.810656e-07, -7.033744e-08, 
    8.432266e-06, 1.359207e-06, 3.28666e-05, 2.786766e-05, -7.110831e-06, 
    -1.169281e-08, 4.016479e-07,
  5.959518e-06, 5.904179e-08, 2.018675e-06, -1.032362e-10, -4.55507e-10, 
    1.098172e-05, 0.005743038, 0.05130031, 0.01282614, 0.0154179, 
    0.008997231, 0.001187099, 0.1231102, 0.1118632, 0.009960076, 
    0.0006821376, 0.0001003255, -1.074128e-09, 0, -2.661364e-10, 
    9.905573e-09, 4.895555e-06, 2.700976e-08, 0.02194529, -3.494142e-05, 
    2.063211e-05, -4.740011e-06, 0.0001356302, 1.603513e-05,
  0.0004360388, 0.005196803, 0.02543126, 0.0007595759, 7.145487e-05, 
    0.009195089, 0.02457168, 0.04487025, 0.03996445, 0.1754881, 0.09086487, 
    0.1571899, 0.1270814, 0.1094636, 0.05504552, 0.0007539514, 0.00681671, 
    8.282595e-06, 1.544398e-05, 0.002693211, 1.549562e-06, 0.004911566, 
    0.0003856921, 0.03495805, 0.006243599, 0.009263845, 0.01190944, 
    0.02378497, 0.0005758219,
  0.09268485, 0.2491986, 0.2411998, 0.1477866, 0.05296393, 0.005957639, 
    0.1146392, 0.1077033, 0.2810161, 0.0753296, 0.1125895, 0.2029306, 
    0.2426331, 0.1220025, 0.07780211, 0.07849924, 0.05397704, 0.05850437, 
    0.06923296, 0.06497524, 0.1157234, 0.1388791, 0.2062554, 0.05778025, 
    0.04618943, 0.08857215, 0.06641093, 0.2078719, 0.1327742,
  0.002405241, 0.0003663572, 4.079935e-05, 0.04205085, 0.155905, 0.257337, 
    0.358478, 0.07753585, 0.377557, 0.07684701, 0.2733507, 0.1783379, 
    0.1229568, 0.09179818, 0.03893887, 0.04803754, 0.002792674, 0.02921325, 
    0.009621147, 0.001955387, 0.006135502, 0.03314791, 0.02420065, 
    0.04612814, 0.02638124, 0.00470341, -0.0001786272, 0.003535943, 
    0.002344953,
  0.009710118, 0.01377099, 0, 3.05458e-07, 0.000115887, 0.0005018357, 
    0.03806377, 0.1332091, 0.1394291, 0.04388193, 0.03807366, 0.08045415, 
    0.2576101, 0.2384821, 0.1976925, 0.1639116, 0.1093295, 0.006931101, 
    -4.401494e-05, 1.143692e-05, 0.143373, 0.1704732, 0.08929477, 0.1028399, 
    0.06896047, 0.04373147, 0.03259615, 0.000150842, 0.02655274,
  0.083624, 0.06743941, 0.00745663, 0.002123705, 0.003893762, -1.539266e-05, 
    -5.466815e-05, 0.07732686, 0.1520641, 0.1864766, 0.1153864, 0.07903044, 
    0.2091012, 0.2417323, 0.09372322, 0.1867146, 0.1377186, 0.1036356, 
    0.001545009, 0.005208418, 0.09508915, 0.06733563, 0.06130461, 0.1070539, 
    0.1117236, 0.09253784, 0.1208385, 0.0568676, 0.05088931,
  0.06663998, 0.09553896, 0.06607381, 0.1984435, 0.113979, 0.1731365, 
    0.06878959, 0.1441478, 0.1651668, 0.1092283, 0.06258462, 0.1963173, 
    0.194647, 0.1364348, 0.1678274, 0.2088075, 0.1704361, 0.1511734, 
    0.116424, 0.05919199, 0.05839756, 0.1193211, 0.12357, 0.1633113, 
    0.1588585, 0.1587775, 0.1299628, 0.1159549, 0.07835115,
  0.1013242, 0.100801, 0.09589151, 0.12919, 0.1620906, 0.1174604, 0.2652901, 
    0.2591974, 0.1450583, 0.1376442, 0.1111334, 0.2282532, 0.2478954, 
    0.1705776, 0.116607, 0.194781, 0.1561869, 0.2349349, 0.2588457, 0.170516, 
    0.158692, 0.1348821, 0.1378339, 0.09416159, 0.1033755, 0.1222116, 
    0.1568125, 0.1766543, 0.1715981,
  0.1607534, 0.1570926, 0.1791068, 0.1195737, 0.102281, 0.1466744, 
    0.08221591, 0.09593071, 0.13695, 0.1721779, 0.09719133, 0.1205709, 
    0.1722852, 0.1730567, 0.1413271, 0.1720868, 0.17223, 0.1003058, 0.13619, 
    0.1938956, 0.1409428, 0.1061249, 0.05508498, 0.05141355, 0.1764701, 
    0.005864965, 0.003633973, 0.2136976, 0.1904179,
  0.09163361, 0.09056525, 0.11484, 0.07727187, 0.07879312, 0.1115304, 
    0.134455, 0.1552227, 0.1169786, 0.1223858, 0.1367351, 0.178634, 
    0.2139661, 0.1420912, 0.09775732, 0.1544473, 0.160881, 0.1901452, 
    0.1556778, 0.1522766, 0.08156843, 0.1053179, 0.04883818, 0.01914199, 
    0.09180223, 0.008196322, -0.003934813, 0.0813252, 0.1029584,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0005797151, 0.005047776, 2.900135e-07, 0, 0, 0, 0,
  0.01302656, 0.02237858, 0.02785476, 0.0149491, -0.0003061512, 0, 0, 0, 0, 
    0.0004232075, -0.000174086, -5.894474e-05, 0.004438455, 0.01161216, 
    0.05082813, 0.02393362, 0.002301523, -7.296447e-05, 0.0008718786, 
    0.0003772554, 0.004767455, 0.01031946, -3.399582e-05, 0.01495383, 
    0.02434579, 0.02461928, 0.01215466, -0.000524591, -0.0001495348,
  0.03769139, 0.06664235, 0.1061471, 0.1051962, 0.04424767, 0.01652736, 
    0.006832727, 0.003620227, 0.004418473, 0.007523188, 0.02187308, 
    0.02789192, 0.04235687, 0.04457284, 0.04935874, 0.0388595, 0.03409573, 
    0.01437114, -9.7809e-05, 0.01595975, 0.03954254, 0.04556724, 0.06932309, 
    0.08563897, 0.06674853, 0.08013219, 0.08489671, 0.06713355, 0.02535435,
  0.160562, 0.2031242, 0.1841008, 0.1800178, 0.1595106, 0.1079956, 
    0.05562292, 0.09779439, 0.08547811, 0.1051738, 0.1130497, 0.09549785, 
    0.1005702, 0.05684493, 0.1116529, 0.1142319, 0.06952623, 0.1005306, 
    0.07502152, 0.09220389, 0.1541501, 0.1614125, 0.2521779, 0.2205608, 
    0.1463986, 0.164615, 0.1682791, 0.1173017, 0.1548779,
  0.09572803, 0.08936848, 0.08401915, 0.1009865, 0.1032647, 0.1440382, 
    0.1151745, 0.1033564, 0.06277421, 0.06803874, 0.08865263, 0.08888828, 
    0.1012562, 0.1636331, 0.1312054, 0.191989, 0.1708018, 0.1812114, 
    0.1166836, 0.1530054, 0.2295205, 0.173316, 0.1857868, 0.1229625, 
    0.1166702, 0.09464408, 0.07579593, 0.1713066, 0.1674551,
  0.0009321115, 0.01254178, 0.004020844, 0.01532585, 0.006304388, 0.01753172, 
    0.01787329, 0.01374742, 1.12908e-05, 0.006031007, 0.02556863, 0.01725922, 
    0.01012866, 0.01531817, 0.07467029, 0.2000448, 0.1844518, 0.1274041, 
    0.1469614, 0.1263053, 0.08468156, 0.03028752, 0.001881968, 0.005353016, 
    0.01916858, 0.05310196, 0.05849459, 0.09025833, 0.009324415,
  1.629542e-07, 2.688857e-06, 1.451341e-07, 4.915632e-08, -6.525318e-12, 
    -4.343179e-09, -1.267467e-08, 1.782651e-05, 2.397732e-08, 4.298767e-10, 
    3.358704e-09, -0.0001823486, 0.04380215, 0.09434027, 0.09133475, 
    0.08053798, 0.008476278, 0.004657646, 6.056617e-05, 0.0002979427, 
    4.589357e-09, -3.481126e-06, 1.327409e-06, 3.79979e-07, 0.0002806529, 
    1.167472e-05, -9.588077e-05, -1.465193e-10, 7.275006e-08,
  6.796655e-07, 6.703006e-08, 2.09947e-06, 0, 1.124371e-08, 1.145525e-05, 
    0.002080074, 0.03499844, 0.01447365, 0.02265125, 0.01314072, 0.001332929, 
    0.1358762, 0.1066949, 0.009743664, 0.0004191964, 0.0001046182, 
    3.532503e-10, 0, 0, -2.132972e-12, 3.320006e-08, -1.643327e-10, 
    0.0006833655, -5.342874e-06, 4.631848e-06, 9.581436e-08, 1.690539e-06, 
    5.832442e-07,
  0.0006284056, 0.001204704, 0.008497918, 0.001862869, 0.0001857095, 
    0.006673412, 0.01457968, 0.01605439, 0.02014706, 0.1035013, 0.06683248, 
    0.1201072, 0.1332565, 0.08876682, 0.04713361, 0.0008295941, 0.004638187, 
    1.175915e-05, -4.706464e-05, 0.00140786, 6.594217e-07, 0.0003634437, 
    4.668548e-07, 0.02795129, 0.01640387, 0.01564731, 0.006075722, 
    0.00645813, 0.0001132026,
  0.07113375, 0.2033178, 0.1872999, 0.1760364, 0.06408617, 0.004553258, 
    0.09322744, 0.04346485, 0.2420627, 0.06341198, 0.06452511, 0.1628126, 
    0.2314414, 0.1095771, 0.06172048, 0.07212232, 0.07250248, 0.06876481, 
    0.07314745, 0.06630526, 0.1094343, 0.1252808, 0.1600817, 0.04373236, 
    0.03675003, 0.07948788, 0.07065223, 0.1881575, 0.1007296,
  0.001513584, 0.0009613274, 0.000155174, 0.04021969, 0.1627816, 0.2275752, 
    0.3931607, 0.07360701, 0.3563294, 0.05864768, 0.2783085, 0.1791577, 
    0.08331633, 0.08627035, 0.02961539, 0.04378777, 0.003444419, 0.02115092, 
    0.008117342, 0.0004300015, 0.006266909, 0.02330201, 0.0166004, 
    0.03571233, 0.01758915, 0.0007757916, 0.0007644391, 0.002391406, 
    0.0005877407,
  0.01370112, 0.01864209, -1.980462e-11, 6.577693e-08, 0.0003617499, 
    0.001105538, 0.02797294, 0.120623, 0.1376977, 0.03092592, 0.03548947, 
    0.08343213, 0.2324737, 0.204518, 0.1944764, 0.1792033, 0.1103235, 
    0.005375037, 0.001944435, 0.001056537, 0.1415259, 0.1484888, 0.0646553, 
    0.06522263, 0.05495575, 0.03222836, 0.02597782, 2.104322e-06, 0.01853553,
  0.06463838, 0.057782, 0.00494475, 0.00373318, 0.01191364, 0.001487637, 
    0.001071451, 0.06677337, 0.1382694, 0.1936602, 0.1163706, 0.0807182, 
    0.2012674, 0.2303519, 0.135605, 0.1611355, 0.1241713, 0.09885487, 
    0.0006975108, 0.001532797, 0.06836848, 0.05824775, 0.04837314, 
    0.09274152, 0.09650445, 0.09750675, 0.1000635, 0.03994517, 0.03152821,
  0.04488623, 0.05809236, 0.05237738, 0.176312, 0.1063215, 0.1634963, 
    0.05622107, 0.2037948, 0.1372014, 0.08498145, 0.04622037, 0.1778204, 
    0.1807727, 0.1292431, 0.1417546, 0.1916007, 0.1671368, 0.1431816, 
    0.1257474, 0.06276165, 0.04809356, 0.1184306, 0.112458, 0.1515172, 
    0.154089, 0.1518486, 0.1182365, 0.1188882, 0.05937989,
  0.09453364, 0.08161122, 0.09244902, 0.1118181, 0.1699016, 0.1019538, 
    0.2092943, 0.2210482, 0.1236128, 0.1223513, 0.09188264, 0.1929098, 
    0.2346636, 0.1596232, 0.1199474, 0.2025057, 0.1852817, 0.2606792, 
    0.3171627, 0.1356918, 0.1365401, 0.1243516, 0.1205317, 0.108756, 
    0.1085248, 0.1496995, 0.1619991, 0.1848687, 0.142327,
  0.1617819, 0.1465133, 0.1726224, 0.1238245, 0.1435553, 0.1575149, 
    0.1164231, 0.108504, 0.1202616, 0.1465719, 0.1351581, 0.1180833, 
    0.1565763, 0.1908163, 0.182895, 0.2092998, 0.170778, 0.1147689, 
    0.1311944, 0.1769236, 0.1550434, 0.1606504, 0.1874254, 0.1432887, 
    0.2097283, 0.08415665, 0.01619929, 0.216641, 0.1965463,
  0.1136844, 0.1068844, 0.2084064, 0.119759, 0.09259786, 0.1689287, 
    0.2488101, 0.2652025, 0.2248475, 0.195075, 0.2070775, 0.2266542, 
    0.2398589, 0.1534151, 0.1112072, 0.1742506, 0.1764297, 0.2050355, 
    0.2070829, 0.2045664, 0.1406348, 0.1432584, 0.1872177, 0.0808959, 
    0.2781037, 0.05258118, 0.07549562, 0.0876694, 0.1038769,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -8.795099e-05, -1.952153e-05, 0, 
    0, 0, 0, -4.011335e-05, -8.196748e-05, 0.002769854, 0.02111701, 
    0.01326348, 0.002978988, 0.009273157, -7.090277e-05, 0,
  0.07632558, 0.09373024, 0.1296002, 0.07794879, 1.867044e-05, -5.205857e-05, 
    0.0006614882, 0, 0, 0.0008987535, -0.000128198, -2.427491e-05, 
    0.005523335, 0.1119176, 0.1184832, 0.06427522, 0.03461882, 0.01254438, 
    0.009998848, 0.003297875, 0.0312478, 0.05298066, 0.0790533, 0.08234383, 
    0.08750699, 0.0524373, 0.0323539, 0.02991978, 0.05864473,
  0.1358258, 0.1038281, 0.2152012, 0.2359548, 0.1640995, 0.06279811, 
    0.03961529, 0.01982567, 0.02994264, 0.06810221, 0.09744716, 0.1832322, 
    0.1936079, 0.1122867, 0.2072251, 0.1380866, 0.11183, 0.09583615, 
    0.04156885, 0.0965462, 0.1095975, 0.1230111, 0.1372801, 0.1452823, 
    0.1548368, 0.142633, 0.1324743, 0.1326973, 0.1345539,
  0.19802, 0.2440645, 0.1944422, 0.192827, 0.1588948, 0.1529142, 0.09902544, 
    0.1318413, 0.1443648, 0.1558116, 0.1472118, 0.189243, 0.2687609, 
    0.1889465, 0.160393, 0.1441741, 0.1363662, 0.1186821, 0.1141443, 
    0.1479715, 0.1870585, 0.2022386, 0.2596201, 0.2616989, 0.1507192, 
    0.1638955, 0.1903585, 0.16016, 0.209668,
  0.09519793, 0.0559449, 0.05978814, 0.088509, 0.0974775, 0.1363082, 
    0.1046987, 0.1016258, 0.0818285, 0.06857742, 0.09157545, 0.1153211, 
    0.1152944, 0.2110422, 0.1946698, 0.2080432, 0.1728224, 0.1788476, 
    0.1309341, 0.1579776, 0.2295489, 0.1833514, 0.2003099, 0.1175605, 
    0.08787248, 0.06712504, 0.06712721, 0.1522049, 0.1658043,
  0.003592436, 0.009310861, 0.005073902, 0.01898805, 0.007020629, 0.02776561, 
    0.01690936, 0.01787562, 0.000333523, 0.0003486192, 0.004205473, 
    0.009998378, 0.0115991, 0.01082167, 0.05968481, 0.1760395, 0.1866126, 
    0.1252358, 0.1436639, 0.1102408, 0.06681582, 0.015683, 0.001552914, 
    0.002761421, 0.01912642, 0.05235373, 0.0591726, 0.07766334, 0.01349775,
  4.034316e-08, 1.771818e-07, 1.842882e-08, 2.546242e-08, 4.339927e-09, 
    -4.77702e-07, 1.171135e-06, -0.0002629207, 2.096193e-08, 2.510177e-09, 
    -3.320119e-10, -0.0001758142, 0.02951435, 0.09824754, 0.09651758, 
    0.05998993, 0.002076364, 0.004183434, -0.0001072086, 1.44231e-06, 
    8.776539e-11, -3.219222e-05, 6.201636e-07, 6.403106e-08, 0.002414546, 
    3.100742e-06, -0.0001914177, 1.666707e-08, 7.819813e-08,
  1.541493e-07, 3.70373e-08, 3.830438e-06, -3.367196e-11, 1.443285e-07, 
    1.236693e-05, 0.001618295, 0.03528565, 0.01027861, 0.02277293, 
    0.01117766, 0.01603438, 0.1431177, 0.1056913, 0.009706721, 0.001020026, 
    9.975747e-05, -1.013428e-08, 0, 0, -1.491948e-14, -1.02832e-09, 
    -3.556926e-11, 0.0001234806, -1.87501e-06, 1.192833e-06, 1.319262e-08, 
    1.715081e-06, 1.263835e-07,
  3.2855e-05, 0.0009230119, 0.007349466, 0.002831757, 0.0007194778, 
    0.005403069, 0.01058393, 0.008397758, 0.02191547, 0.06373107, 0.05167194, 
    0.09314629, 0.1332779, 0.07956535, 0.04312865, 0.0009865653, 0.0029407, 
    0.002364665, -6.582235e-05, 0.0005200187, 3.992139e-07, 2.976902e-05, 
    -1.142734e-06, 0.01516113, 0.02983012, 0.0247178, 0.006588136, 
    0.003015063, 6.71416e-06,
  0.05906409, 0.1599925, 0.1482778, 0.2072443, 0.0702305, 0.01120994, 
    0.06383244, 0.01795187, 0.2203047, 0.05394259, 0.0432329, 0.1402763, 
    0.215158, 0.1108627, 0.05391086, 0.08838045, 0.0888915, 0.08415446, 
    0.07548653, 0.06390091, 0.1104175, 0.1127006, 0.1335299, 0.03556848, 
    0.03558847, 0.07721069, 0.08024622, 0.1725807, 0.0895331,
  0.0006866236, 5.822786e-05, 0.0003461208, 0.03959025, 0.1726479, 0.1905751, 
    0.4214438, 0.07727851, 0.3612051, 0.05444334, 0.2859395, 0.1753598, 
    0.0710153, 0.07665186, 0.01988757, 0.03407465, 0.000305704, 0.009163367, 
    0.003236738, 0.0001219928, 0.01207296, 0.01497053, 0.01203943, 
    0.02943858, 0.01213636, 0.0005824927, -0.0002875885, 0.002593693, 
    0.001818109,
  0.04505276, 0.02348698, -4.221841e-11, 4.186445e-10, 0.001213599, 
    0.00281707, 0.02165263, 0.1130674, 0.143116, 0.02165741, 0.03177254, 
    0.08539247, 0.2021567, 0.1717487, 0.1915654, 0.1435767, 0.06896211, 
    0.003748022, 0.007409859, 0.003002742, 0.1172385, 0.1005042, 0.05274748, 
    0.0411224, 0.03862952, 0.01590534, 0.02613097, -3.420539e-05, 0.01348807,
  0.06244715, 0.06270484, 0.004136729, 0.003670339, 0.01858404, 0.004418822, 
    0.002384323, 0.06222624, 0.1198238, 0.1782615, 0.1000851, 0.08355924, 
    0.2037181, 0.188674, 0.1000868, 0.1490422, 0.1477674, 0.08945873, 
    0.001072821, 0.0002663063, 0.06491989, 0.04536779, 0.03473537, 0.0895721, 
    0.07757773, 0.08409976, 0.07384095, 0.0277723, 0.01450201,
  0.04091546, 0.05310359, 0.04369451, 0.1646906, 0.1053937, 0.1440142, 
    0.05752327, 0.2101013, 0.122281, 0.07994586, 0.03862081, 0.1589617, 
    0.1789118, 0.1210006, 0.1299341, 0.1768904, 0.154643, 0.1376216, 
    0.122956, 0.06930892, 0.04316162, 0.1088808, 0.1086224, 0.1365276, 
    0.1522631, 0.1473738, 0.113438, 0.1336774, 0.05103942,
  0.09173655, 0.06872262, 0.08912586, 0.09711742, 0.1424503, 0.07605505, 
    0.1712822, 0.1945181, 0.1101565, 0.1115725, 0.07481044, 0.1800601, 
    0.2112172, 0.1530834, 0.1292628, 0.2219931, 0.1702757, 0.2764211, 
    0.3030842, 0.1165662, 0.1159655, 0.1019913, 0.1083225, 0.1331306, 
    0.1102616, 0.1521177, 0.1541865, 0.1782876, 0.1191915,
  0.1711867, 0.1414307, 0.1721453, 0.1389726, 0.1343392, 0.141879, 0.1281724, 
    0.0972279, 0.09935334, 0.1181652, 0.1197127, 0.103616, 0.1484008, 
    0.1866279, 0.1942739, 0.1968741, 0.1515853, 0.10431, 0.1282884, 
    0.1717566, 0.1537526, 0.1762476, 0.2230684, 0.2048889, 0.2272173, 
    0.1931489, 0.06888556, 0.2079592, 0.197512,
  0.109565, 0.1057205, 0.215217, 0.1262406, 0.08155844, 0.1849255, 0.2466902, 
    0.2550972, 0.202786, 0.1921147, 0.203675, 0.2011542, 0.2070815, 0.124545, 
    0.09100681, 0.1588682, 0.1764967, 0.1753159, 0.2137766, 0.2059631, 
    0.1378685, 0.1374436, 0.1954603, 0.1030079, 0.2842447, 0.1926461, 
    0.1253368, 0.08190265, 0.09285085,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.181253e-05, 0.006338023, 
    0.01441222, 0.001062291, 0.0007494933, 1.539195e-05, -3.681653e-05, 
    -0.0004357036, 0.001465617, 0.009630959, 0.03117377, 0.04119095, 
    0.03426726, 0.03836599, 0.000638695, 0,
  0.1596545, 0.2609697, 0.2206123, 0.1443285, 0.001149208, -0.001992023, 
    0.007950237, 0, -4.944576e-05, 0.0007305306, 0.001617035, 0.001479325, 
    0.05880309, 0.2176391, 0.2248282, 0.1591946, 0.1242567, 0.08101693, 
    0.06077673, 0.1051381, 0.110721, 0.1373257, 0.1313713, 0.163172, 
    0.139066, 0.06848828, 0.05333175, 0.07602634, 0.1283427,
  0.1878568, 0.1708546, 0.3005297, 0.2619541, 0.1794994, 0.1057048, 
    0.1213985, 0.04874421, 0.06953546, 0.1344259, 0.14715, 0.2734385, 
    0.2865607, 0.1970628, 0.2913685, 0.1570769, 0.1507341, 0.09025124, 
    0.06196135, 0.1283615, 0.1699971, 0.167089, 0.1624576, 0.1827669, 
    0.2004257, 0.2233078, 0.2284716, 0.1508329, 0.1934348,
  0.200432, 0.2532054, 0.1830178, 0.1875174, 0.1615589, 0.1592675, 
    0.09891643, 0.1522127, 0.1722319, 0.184583, 0.1848281, 0.2542018, 
    0.2910738, 0.1697125, 0.1481466, 0.1536361, 0.1445267, 0.1121651, 
    0.1257112, 0.154016, 0.1939822, 0.2096167, 0.2730907, 0.2373472, 
    0.1329967, 0.1603083, 0.1987184, 0.1766616, 0.2098019,
  0.0942588, 0.04371687, 0.05737522, 0.09166212, 0.09927239, 0.1413812, 
    0.1088545, 0.1040662, 0.08728475, 0.07015481, 0.098235, 0.1208533, 
    0.1119674, 0.195524, 0.1888981, 0.1993313, 0.1656254, 0.1697736, 
    0.1345937, 0.1542715, 0.2244311, 0.1827763, 0.2063149, 0.08695659, 
    0.05917302, 0.05306182, 0.06462275, 0.1382953, 0.1573859,
  0.00183778, 0.00542563, 0.006927919, 0.02524361, 0.009460703, 0.02678306, 
    0.01726355, 0.01824321, 3.190802e-06, 3.025026e-05, 8.152393e-06, 
    0.002654971, 0.009176365, 0.01460469, 0.05137999, 0.1522158, 0.176788, 
    0.1145815, 0.1427207, 0.1181243, 0.07618687, 0.01134843, 0.002507911, 
    0.0008782007, 0.01907676, 0.04423803, 0.04913102, 0.06651624, 0.0211262,
  -7.872725e-11, -6.418117e-09, -3.160754e-08, 2.131547e-09, -2.126909e-07, 
    -6.791951e-07, 0.0001888248, 0.000600185, -2.012158e-05, 0, 3.601084e-09, 
    0.004540802, 0.02665911, 0.09176781, 0.08794444, 0.05499938, 
    0.0006687865, 0.007321968, -2.085412e-05, 1.401648e-08, 1.976654e-08, 
    -0.0002586395, 1.090922e-07, 1.204275e-07, 0.001244026, 3.277214e-06, 
    -0.0001565672, 1.851476e-08, -3.187814e-10,
  1.394308e-08, -3.139908e-09, 8.222055e-06, -1.660571e-10, 3.980513e-07, 
    0.0005166347, 0.002612952, 0.0315081, 0.02127505, 0.007550607, 
    0.02813076, 0.02969547, 0.16361, 0.09188038, 0.01670907, 0.002519151, 
    0.000294154, -3.83222e-08, -8.590516e-11, 0, 0, 3.968676e-14, 
    3.227234e-09, 6.445703e-05, -7.321173e-07, 3.422269e-07, 2.782955e-07, 
    1.901218e-06, 2.170521e-08,
  0.0001774863, 0.001559422, 0.00917198, 0.002340453, 0.001050847, 
    0.005542514, 0.009574297, 0.007840479, 0.01448229, 0.03948498, 0.042869, 
    0.07592208, 0.1302517, 0.07723559, 0.04599093, 0.00291452, 0.002920062, 
    0.005204886, -5.312826e-08, 0.0002271796, -1.278644e-07, 0.0005153414, 
    -4.961379e-05, 0.007490606, 0.03445868, 0.04049765, 0.006800561, 
    0.005700409, 2.974677e-07,
  0.05782802, 0.146483, 0.1275919, 0.2622249, 0.08016578, 0.01390377, 
    0.05799511, 0.01190836, 0.1893139, 0.06212695, 0.03310052, 0.13121, 
    0.1958866, 0.101901, 0.06443229, 0.09798791, 0.09196091, 0.09495327, 
    0.08037371, 0.06492344, 0.1125675, 0.1026653, 0.1231143, 0.03050868, 
    0.03721014, 0.07707185, 0.09675641, 0.1712744, 0.07705319,
  0.01032181, 6.642304e-06, 0.00203157, 0.0214028, 0.1675746, 0.1374085, 
    0.4651225, 0.08548947, 0.3573627, 0.04600407, 0.2629194, 0.1804946, 
    0.06294139, 0.06487788, 0.01286199, 0.0154419, 0.0005790778, 0.01620845, 
    0.0002675957, -1.49556e-05, 0.01833596, 0.01200979, 0.008887595, 
    0.02438718, 0.00986993, 0.01088119, 0.01183324, 0.004716009, 0.02046628,
  0.1063712, 0.04668168, 0, -3.257917e-11, 0.005448626, 0.001896144, 
    0.02490395, 0.1105372, 0.1631976, 0.01346202, 0.02756761, 0.07863564, 
    0.1917923, 0.1732616, 0.1734364, 0.09840293, 0.03737281, 0.004254647, 
    0.0004122895, 0.004742058, 0.1097057, 0.05187857, 0.04790368, 0.0317998, 
    0.02835313, 0.01418689, 0.02305331, -1.711549e-05, 0.01289413,
  0.05717225, 0.06585562, 0.005373692, 0.003748564, 0.00786676, 0.004621924, 
    0.002936627, 0.05219829, 0.1108241, 0.1585965, 0.08001548, 0.07347933, 
    0.2047729, 0.1808147, 0.09986952, 0.1050903, 0.09593633, 0.1018428, 
    0.0001352766, 0.0004088765, 0.06127168, 0.03945331, 0.0258533, 
    0.07735761, 0.05990004, 0.07374666, 0.06021338, 0.01927812, 0.005420213,
  0.04280349, 0.06315466, 0.03118614, 0.1521421, 0.09510062, 0.1281644, 
    0.05588437, 0.2004794, 0.1157774, 0.07374483, 0.03844382, 0.1488888, 
    0.1521375, 0.1269839, 0.1248759, 0.1702414, 0.1371893, 0.1360845, 
    0.1361683, 0.05794974, 0.04143995, 0.09208177, 0.1047931, 0.1223696, 
    0.1330113, 0.1427476, 0.1237829, 0.1212258, 0.04753818,
  0.07793747, 0.06895482, 0.08903091, 0.07224328, 0.1295109, 0.06500608, 
    0.1564832, 0.1738524, 0.1000201, 0.1048782, 0.06375276, 0.181202, 
    0.1992629, 0.1704365, 0.1412875, 0.1844325, 0.1484466, 0.2788464, 
    0.2934394, 0.1032875, 0.1029777, 0.09160105, 0.08784918, 0.1508919, 
    0.1145665, 0.1411279, 0.1425126, 0.1458615, 0.1055522,
  0.1703516, 0.1463557, 0.1709195, 0.153419, 0.1342445, 0.1425871, 0.1266251, 
    0.08364676, 0.09024917, 0.1075311, 0.1098357, 0.08876399, 0.1364011, 
    0.1885005, 0.2140947, 0.1823081, 0.1410842, 0.08115812, 0.1305274, 
    0.1592175, 0.1576674, 0.1712585, 0.2161908, 0.2125638, 0.2341424, 
    0.323635, 0.1819648, 0.1923282, 0.2105923,
  0.0947618, 0.1001106, 0.2076809, 0.1260542, 0.07994983, 0.1818654, 
    0.247601, 0.2619915, 0.1988027, 0.178343, 0.190976, 0.1766737, 0.1743295, 
    0.1186477, 0.07174139, 0.1469041, 0.1494051, 0.1649664, 0.234878, 
    0.2117942, 0.1339039, 0.1369295, 0.1991137, 0.1065544, 0.2579204, 
    0.1824559, 0.1161866, 0.08135056, 0.09053622,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.007538422, 0.03765026, 0.05281661, 
    0.02890601, 0.03396554, 0.004730321, -0.0003002975, 0.0008142233, 
    0.004647113, 0.02517042, 0.1048981, 0.08557108, 0.06323671, 0.07893871, 
    0.02393248, 0,
  0.2631797, 0.3402656, 0.3052508, 0.1787934, 0.01017334, 0.01032661, 
    0.01749001, -0.000183558, -0.0003325595, 0.0001019984, 0.005928797, 
    0.01127607, 0.1785893, 0.2346301, 0.2359778, 0.1555877, 0.1344087, 
    0.08166666, 0.07091612, 0.1339002, 0.1822963, 0.1904702, 0.1876337, 
    0.2475181, 0.2091946, 0.1169123, 0.1186869, 0.1374286, 0.1932519,
  0.2343567, 0.2007391, 0.3423262, 0.2601999, 0.2093282, 0.166631, 0.162479, 
    0.1221898, 0.116273, 0.2030167, 0.260058, 0.3122831, 0.3276757, 
    0.2083412, 0.2849487, 0.1480423, 0.1614063, 0.09224798, 0.08542369, 
    0.1422397, 0.2230058, 0.2106692, 0.2028899, 0.2272209, 0.2276008, 
    0.2738764, 0.2968212, 0.207097, 0.2544895,
  0.1910654, 0.2389772, 0.1640327, 0.1789604, 0.1439255, 0.157347, 0.1111404, 
    0.1522285, 0.1774574, 0.214485, 0.2190268, 0.2747956, 0.2947184, 
    0.1620343, 0.1342182, 0.1537808, 0.1471083, 0.1241322, 0.1313209, 
    0.1685428, 0.1870921, 0.1896911, 0.240033, 0.2184246, 0.1263408, 
    0.1320938, 0.196698, 0.2319572, 0.2205397,
  0.1067588, 0.04461997, 0.06107322, 0.08988738, 0.1042137, 0.1480705, 
    0.1094224, 0.1084028, 0.08560167, 0.06426512, 0.1030302, 0.1267, 
    0.09905846, 0.1739489, 0.1816295, 0.200125, 0.1553074, 0.1452177, 
    0.1311313, 0.1444359, 0.2065356, 0.182903, 0.1777842, 0.0696918, 
    0.04229632, 0.04940609, 0.06526095, 0.1317416, 0.1366201,
  0.002013327, 0.009013304, 0.009780935, 0.03298802, 0.01622503, 0.02858243, 
    0.0159832, 0.01562695, -3.948771e-05, 0.0003041686, -2.436341e-05, 
    0.0001402905, 0.00721211, 0.01795808, 0.0497391, 0.1436834, 0.1480219, 
    0.1036783, 0.1438648, 0.07730562, 0.06086993, 0.01185179, 0.001944115, 
    0.002377458, 0.02255455, 0.04763792, 0.04293248, 0.06603028, 0.02753596,
  -7.033093e-13, -1.661238e-09, -9.456487e-05, 4.312455e-10, -2.600007e-07, 
    -5.47629e-06, 0.000510947, 2.466239e-05, -0.0001875892, 1.081753e-10, 
    1.458662e-08, 0.0002974789, 0.03267083, 0.08086471, 0.0751885, 
    0.03609886, 0.0007043501, 0.01549209, -1.941103e-06, -8.761648e-09, 
    2.586033e-10, 0.001609077, 1.434262e-09, 2.253284e-07, 0.0003135742, 
    2.472903e-05, 0.0005253503, -1.296339e-10, 0,
  3.644611e-08, 2.17385e-08, 6.617646e-06, -1.258027e-11, 4.022319e-07, 
    0.00720477, 0.001093011, 0.02619378, 0.0296212, 0.003688121, 0.0332555, 
    0.04471543, 0.1539686, 0.08463163, 0.02134001, 0.0054456, 0.0010265, 
    -1.412117e-07, 0, 4.30863e-13, -2.360261e-12, 1.134291e-10, 6.440633e-09, 
    9.367153e-05, 5.941537e-06, 1.785715e-06, 8.628808e-08, 9.198973e-08, 
    1.35071e-10,
  0.0004668768, 0.002135692, 0.0290547, 0.001845868, 0.001505474, 
    0.007903181, 0.008409785, 0.00636518, 0.01028231, 0.01869669, 0.02748782, 
    0.05871478, 0.1192376, 0.07993005, 0.04320469, 0.00826771, 0.003500061, 
    0.01314275, 0.01814402, 0.003585316, -8.723414e-06, 0.0002178161, 
    1.798205e-05, 0.008987864, 0.04299719, 0.07002521, 0.007050985, 
    0.01030636, -3.424271e-06,
  0.05033524, 0.1338428, 0.1186777, 0.2958798, 0.1558209, 0.02023017, 
    0.05141725, 0.01209443, 0.148729, 0.08764651, 0.03294862, 0.1229653, 
    0.1984284, 0.1070378, 0.06331438, 0.09115045, 0.08571596, 0.1093709, 
    0.08445057, 0.07648886, 0.1350288, 0.1027805, 0.1215145, 0.02990312, 
    0.02727253, 0.07037188, 0.09887596, 0.1563264, 0.077783,
  0.05762905, 0.001280884, 0.0003180692, 0.005228029, 0.1214958, 0.1031482, 
    0.5017723, 0.09338322, 0.3918933, 0.04173926, 0.2784975, 0.1842875, 
    0.05805294, 0.04794, 0.01166132, 0.004118938, 0.0001361175, 0.001588773, 
    0.0002145568, 0.002488898, 0.0213145, 0.01151684, 0.007038485, 
    0.02048508, 0.008457617, 0.01729129, 0.005527017, 0.02027491, 0.0283798,
  0.08141846, 0.03508931, -1.966941e-10, 1.660177e-10, 0.0009050465, 
    0.0005721511, 0.03132406, 0.1237195, 0.1882635, 0.01652347, 0.03416107, 
    0.07584549, 0.1830308, 0.1744167, 0.156565, 0.06089897, 0.01886745, 
    0.000184819, 4.431758e-06, 0.01287255, 0.0827715, 0.03389223, 0.05093726, 
    0.0252483, 0.02840716, 0.01309515, 0.01731761, -4.827996e-06, 0.01149512,
  0.04989621, 0.06365258, 0.004221104, 0.004191344, 0.00453966, 0.004030039, 
    0.006937591, 0.03633433, 0.0875411, 0.1603645, 0.07046016, 0.06803546, 
    0.2022848, 0.1823648, 0.07226618, 0.08545075, 0.08435318, 0.08251077, 
    -3.060787e-06, 0.000135844, 0.07557832, 0.04277251, 0.02398504, 
    0.07045876, 0.05482115, 0.07081521, 0.0662726, 0.009606082, 0.001167273,
  0.0332531, 0.06155834, 0.01876632, 0.143821, 0.09238713, 0.1091705, 
    0.0546457, 0.1802957, 0.1088678, 0.06705272, 0.04686748, 0.1439655, 
    0.138401, 0.1175249, 0.1039349, 0.1574841, 0.1349697, 0.1185795, 
    0.1472339, 0.04324874, 0.04097622, 0.08903711, 0.09507071, 0.1001801, 
    0.1189935, 0.1503099, 0.1339417, 0.1261999, 0.05178076,
  0.07842536, 0.07204339, 0.09285075, 0.0588006, 0.1057002, 0.05579596, 
    0.1664093, 0.1548612, 0.1004284, 0.1128086, 0.05735035, 0.1684308, 
    0.1972463, 0.1554322, 0.1322097, 0.1773406, 0.1522714, 0.2709951, 
    0.276142, 0.1096501, 0.09736111, 0.09738571, 0.0911369, 0.1570976, 
    0.1218013, 0.1529246, 0.2026948, 0.1750431, 0.1282053,
  0.1868008, 0.2047367, 0.1838266, 0.1676174, 0.1260945, 0.1412315, 
    0.1235891, 0.07868841, 0.0845961, 0.09853665, 0.08847867, 0.08127089, 
    0.1414735, 0.2059089, 0.2188963, 0.1924302, 0.143338, 0.06923326, 
    0.1225954, 0.1245176, 0.1763239, 0.1807604, 0.2233746, 0.2279373, 
    0.2517796, 0.2926745, 0.2011828, 0.1686553, 0.1855432,
  0.1247683, 0.1334431, 0.2089003, 0.1271378, 0.08955732, 0.1688604, 
    0.257804, 0.2738855, 0.2149034, 0.1816481, 0.1744962, 0.1533593, 
    0.1696727, 0.1111235, 0.06749683, 0.1574481, 0.166593, 0.1767232, 
    0.2391096, 0.1931245, 0.1145126, 0.1452461, 0.2182743, 0.1159234, 
    0.2452084, 0.1840317, 0.1283929, 0.1098864, 0.1232698,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  -4.819941e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.500025e-06, 0.03211579, 
    0.06479277, 0.07442254, 0.04979835, 0.06037658, 0.03063703, 0.01549769, 
    0.01191671, 0.01274871, 0.04307376, 0.2726077, 0.1434346, 0.07828052, 
    0.1323161, 0.06085199, 0.00496636,
  0.3138412, 0.4246641, 0.3479908, 0.23885, 0.03849317, 0.04064019, 
    0.02168219, -0.001080759, 0.0009088151, 0.02867486, 0.03297396, 
    0.05539041, 0.2744912, 0.2678492, 0.2303818, 0.1517041, 0.116193, 
    0.08017636, 0.07813921, 0.1538415, 0.1999697, 0.2310994, 0.2506982, 
    0.3597952, 0.2897564, 0.1441354, 0.153185, 0.1527208, 0.2561479,
  0.2408442, 0.2088721, 0.3431506, 0.2706255, 0.2137941, 0.1794857, 
    0.1991121, 0.1768703, 0.1252308, 0.2491749, 0.2734303, 0.3448447, 
    0.3187724, 0.2130475, 0.2646535, 0.1525639, 0.1692458, 0.08151925, 
    0.08361271, 0.1536073, 0.2370036, 0.2276553, 0.2300608, 0.2208759, 
    0.2188875, 0.2721499, 0.2707715, 0.2288673, 0.2584653,
  0.2159545, 0.2426263, 0.1475949, 0.1800412, 0.1363823, 0.1589638, 
    0.1198337, 0.1555219, 0.2133278, 0.2419295, 0.2290633, 0.2824814, 
    0.271652, 0.1564368, 0.1224566, 0.127892, 0.1451088, 0.1236253, 
    0.1176649, 0.1727826, 0.1911033, 0.2007301, 0.2202828, 0.2008774, 
    0.1216233, 0.1198058, 0.2180621, 0.238264, 0.2128771,
  0.1073934, 0.04548934, 0.06506584, 0.08928761, 0.1003684, 0.1307684, 
    0.10452, 0.1207397, 0.08535232, 0.06900106, 0.1076293, 0.1177662, 
    0.1044215, 0.1660742, 0.1787555, 0.1950561, 0.1453492, 0.135797, 
    0.1376079, 0.1436139, 0.1859733, 0.1733937, 0.1787049, 0.05978447, 
    0.03649537, 0.04801547, 0.06004015, 0.1284026, 0.127177,
  0.009385579, 0.01019599, 0.01597754, 0.04335926, 0.01955852, 0.03156033, 
    0.01532931, 0.01217074, -0.0001185374, 0.0007744576, -3.631438e-05, 
    0.0001410852, 0.009845247, 0.01630642, 0.05103691, 0.1250912, 0.1233715, 
    0.09153163, 0.1470813, 0.07779518, 0.05246265, 0.01324691, 0.005205084, 
    0.003641679, 0.03208897, 0.04287639, 0.0452997, 0.06409912, 0.02843559,
  9.482514e-10, 4.238971e-10, -0.0001274504, -3.798093e-08, -8.87336e-07, 
    -4.635163e-05, 0.0009364653, 0.001831192, -0.000566171, 1.093766e-08, 
    6.065342e-08, 0.001976169, 0.0370537, 0.08265497, 0.0774366, 0.02022682, 
    0.001387696, 0.02306101, -2.274158e-06, 4.072607e-08, 1.550989e-09, 
    0.003952771, 8.432708e-10, 3.024032e-06, 0.0005971267, 0.0006016409, 
    0.001342277, 2.11776e-08, 1.598986e-08,
  7.951409e-08, 2.344218e-07, 5.573036e-06, 3.443526e-11, -8.583351e-06, 
    0.01212408, 0.002269255, 0.02559935, 0.04529158, 0.002133216, 0.05524505, 
    0.03595201, 0.1467449, 0.08201255, 0.02031906, 0.004819986, 0.001196277, 
    2.611198e-07, -1.263856e-11, -3.678966e-12, 3.681538e-11, 4.32635e-10, 
    5.154293e-09, 0.001306218, 5.414916e-05, 7.009959e-07, 2.56608e-06, 
    -6.958543e-07, 3.320225e-09,
  0.00661554, 0.00296011, 0.0508207, 0.01533702, 0.0005057947, 0.007234311, 
    0.006956982, 0.007081044, 0.008572118, 0.01009526, 0.0258174, 0.0677579, 
    0.1264983, 0.0843723, 0.04857633, 0.01901173, 0.003000603, 0.0127595, 
    0.02520433, 0.009737287, 3.941335e-05, 4.720675e-05, 0.0001740308, 
    0.02700335, 0.06231272, 0.085867, 0.01824839, 0.007602519, -3.828096e-06,
  0.04518059, 0.1089322, 0.1196496, 0.3615955, 0.1927694, 0.01838393, 
    0.06424384, 0.01454523, 0.1165164, 0.1302429, 0.05183981, 0.1354527, 
    0.2073793, 0.1280408, 0.06169931, 0.1094439, 0.09351954, 0.1300261, 
    0.1016657, 0.07625877, 0.1868882, 0.101155, 0.1304661, 0.03073391, 
    0.02579085, 0.06771299, 0.1051897, 0.1493637, 0.09175823,
  0.02118338, 1.656652e-05, -1.814719e-05, 0.0001207718, 0.08857059, 
    0.1083186, 0.5658917, 0.1319288, 0.4401376, 0.05102551, 0.2922335, 
    0.1992758, 0.07405262, 0.03455146, 0.0112851, 0.003393904, 0.0002733319, 
    0.0004721617, 0.01286694, 0.006351158, 0.01940189, 0.01475985, 
    0.006350588, 0.01994317, 0.009144773, 0.002681893, 0.004447875, 
    0.01419542, 0.03533715,
  0.02904928, 0.0132854, 1.271844e-07, 1.49603e-08, 4.747261e-05, 
    0.0001795375, 0.04142593, 0.124968, 0.2003244, 0.02360601, 0.0340252, 
    0.09069623, 0.2045839, 0.1726332, 0.1424406, 0.05570224, 0.02741469, 
    0.0009745395, -2.302344e-06, 0.006306706, 0.06558605, 0.0307204, 
    0.06007609, 0.01952899, 0.02453927, 0.00950386, 0.01191865, 
    -6.829694e-08, 0.01166052,
  0.0517815, 0.06516465, 0.00685959, 0.005601169, 0.005341465, 0.001643507, 
    0.02647459, 0.02378334, 0.06951064, 0.1618105, 0.06822579, 0.07544338, 
    0.2043507, 0.240246, 0.07736735, 0.06532335, 0.07690684, 0.07982779, 
    -1.003061e-05, 0.0005961761, 0.08992756, 0.05805025, 0.01991139, 
    0.06972477, 0.05738233, 0.063042, 0.06990796, 0.009121968, 0.0006792609,
  0.02362832, 0.05663585, 0.02053033, 0.1296237, 0.08993808, 0.1110172, 
    0.05672506, 0.1742455, 0.1100314, 0.05889195, 0.05486791, 0.1457209, 
    0.1208121, 0.1161819, 0.08842362, 0.1438056, 0.1216573, 0.1172117, 
    0.1340653, 0.03423051, 0.0401082, 0.08298485, 0.10181, 0.09439892, 
    0.1104398, 0.1264092, 0.1479113, 0.1339473, 0.05736785,
  0.05065053, 0.06830654, 0.09247793, 0.05207308, 0.1067519, 0.05278843, 
    0.1584069, 0.1415903, 0.09309028, 0.1211424, 0.05835029, 0.1585769, 
    0.2019233, 0.1712728, 0.1007822, 0.1668048, 0.1406532, 0.297646, 
    0.2553439, 0.1091587, 0.07855482, 0.09143183, 0.1032826, 0.166573, 
    0.1474039, 0.1480341, 0.1810676, 0.1554868, 0.1248288,
  0.2151963, 0.1444605, 0.1777119, 0.1948862, 0.122158, 0.1461009, 0.1185991, 
    0.07920538, 0.07346569, 0.0904687, 0.08961193, 0.1002675, 0.1670867, 
    0.2336379, 0.2572785, 0.1784322, 0.1558984, 0.06500024, 0.103324, 
    0.09788896, 0.1904799, 0.2007003, 0.2267514, 0.2555195, 0.2687652, 
    0.2738178, 0.2306818, 0.1817145, 0.240623,
  0.1097577, 0.1341966, 0.1855187, 0.1625345, 0.1168639, 0.204916, 0.2877861, 
    0.3514002, 0.2370026, 0.2266854, 0.1750429, 0.130855, 0.1660717, 
    0.1104676, 0.1051164, 0.1940707, 0.2035201, 0.2154418, 0.2675326, 
    0.2146333, 0.1335774, 0.174128, 0.2303474, 0.1237978, 0.2416342, 
    0.1644435, 0.1658015, 0.1116142, 0.1069454,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0.0002964842, -0.0002347901, 
    -0.000173096, -0.0001114019, -4.970775e-05, 1.198637e-05, 7.368049e-05, 
    0.0002066753, 0.0001449812, 8.328706e-05, 2.159294e-05, -4.010117e-05, 
    -0.0001017953, -0.0001634894, 0,
  0.007347177, -0.0001837689, -2.305369e-06, 0, -9.871556e-06, 0.0002249186, 
    0, 0, 0, 0, 0, 0, 5.578863e-06, 0.04694335, 0.06512734, 0.09476645, 
    0.06337351, 0.07550213, 0.07679788, 0.02959025, 0.03316778, 0.03459539, 
    0.0952637, 0.3076118, 0.1648062, 0.09736492, 0.1590398, 0.1263372, 
    0.04435923,
  0.3471883, 0.4349149, 0.3385206, 0.2400831, 0.06996578, 0.081123, 
    0.02169081, 0.01080264, 0.04132573, 0.09397265, 0.1040537, 0.1529929, 
    0.3146679, 0.268217, 0.2303373, 0.1476759, 0.106167, 0.0902239, 
    0.1118365, 0.1914218, 0.2905188, 0.3003486, 0.2715821, 0.3990395, 
    0.2797021, 0.1424071, 0.1537993, 0.1287784, 0.2751257,
  0.2683767, 0.1934931, 0.3387697, 0.2616794, 0.2219367, 0.1831958, 
    0.2111987, 0.1905899, 0.1465416, 0.2396286, 0.2717786, 0.319885, 
    0.286066, 0.2210855, 0.2607028, 0.161146, 0.1873158, 0.07251552, 
    0.1018258, 0.1778474, 0.2174602, 0.2400132, 0.2021577, 0.2245805, 
    0.2025034, 0.2450065, 0.2665608, 0.2296409, 0.3066576,
  0.2038051, 0.2245985, 0.1460534, 0.1687328, 0.1321218, 0.153955, 0.1312771, 
    0.1843878, 0.2108034, 0.250967, 0.2356074, 0.2773087, 0.2598586, 
    0.1607381, 0.1092269, 0.1214171, 0.1286495, 0.1163606, 0.1087695, 
    0.1840099, 0.189915, 0.1991435, 0.2084807, 0.1797629, 0.1078896, 
    0.09724391, 0.2146738, 0.246138, 0.2110335,
  0.1160804, 0.07503965, 0.07291046, 0.09875759, 0.08620115, 0.1324844, 
    0.106274, 0.117796, 0.09312189, 0.07970777, 0.1177629, 0.1140643, 
    0.1140234, 0.1737988, 0.1673995, 0.1833108, 0.1355433, 0.1362427, 
    0.1497677, 0.1427092, 0.189172, 0.1663664, 0.1479813, 0.05261964, 
    0.04122676, 0.04581978, 0.06367023, 0.1432735, 0.142991,
  0.01177548, 0.0130788, 0.02954789, 0.04671416, 0.02364998, 0.02807847, 
    0.0140407, 0.01642244, -2.945743e-06, 0.00209727, 0.0002493944, 
    0.004996358, 0.01799044, 0.01763155, 0.0533312, 0.1189117, 0.1155581, 
    0.09131649, 0.1399206, 0.06904449, 0.04939297, 0.01682901, 0.009604386, 
    0.003160588, 0.04658645, 0.03988596, 0.04502557, 0.07349931, 0.02850068,
  1.225959e-07, 1.410866e-08, -1.5661e-05, 1.029296e-07, 2.378072e-05, 
    -0.0001478767, 0.006840086, 0.002059474, -0.0004766519, 6.19796e-08, 
    2.078993e-07, 0.0005067266, 0.02803493, 0.08482723, 0.08792682, 
    0.02394709, 0.002416355, 0.02799896, -1.926602e-06, 7.521918e-08, 
    2.543747e-07, 0.007573408, 1.622829e-09, 7.460707e-06, 0.0009929114, 
    0.0007694178, 0.0005391301, -1.076829e-06, 2.01126e-07,
  3.590923e-07, 1.000713e-06, 2.06509e-06, 8.608642e-08, 7.273375e-05, 
    0.01962779, 0.00740434, 0.03288529, 0.04863484, 0.000981806, 0.0461337, 
    0.02941197, 0.1474275, 0.09432893, 0.02360534, 0.004881487, 0.001023221, 
    3.539692e-05, -1.495349e-10, 2.811357e-11, 1.225887e-10, 7.023831e-10, 
    4.719292e-07, 0.001350337, 5.065493e-05, 2.529376e-07, 1.546567e-06, 
    2.931262e-07, -1.036895e-07,
  0.03247477, 0.02926744, 0.06044719, 0.02301012, 0.00174661, 0.008592196, 
    0.009794304, 0.0140043, 0.01054603, 0.01064258, 0.03655829, 0.09160059, 
    0.1318084, 0.08332898, 0.05538488, 0.02990612, 0.007116681, 0.009645111, 
    0.02424278, 0.003377479, 2.491529e-05, 3.277503e-05, 0.001729723, 
    0.0628864, 0.06015233, 0.07480794, 0.01743474, 0.002692871, 0.00582862,
  0.05245778, 0.1036648, 0.1498735, 0.4296079, 0.179365, 0.01768977, 
    0.1026553, 0.02835638, 0.1070288, 0.1869796, 0.09452904, 0.1728175, 
    0.2390953, 0.1443563, 0.07466529, 0.1193915, 0.1172406, 0.1458252, 
    0.1272914, 0.09217615, 0.2196377, 0.1375923, 0.1514839, 0.03826916, 
    0.03795008, 0.07479688, 0.1188207, 0.1784479, 0.1365956,
  0.005957138, 2.294927e-06, -9.813041e-06, -2.064682e-05, 0.05786302, 
    0.1126329, 0.6536289, 0.1699485, 0.4844373, 0.06858824, 0.3052654, 
    0.2258227, 0.09305833, 0.02735661, 0.01274041, 0.00383775, 0.0006097132, 
    0.0001427718, 0.003187893, 0.008338768, 0.03617631, 0.02735479, 
    0.0102475, 0.02528972, 0.01333247, 0.001271426, 0.005877757, 0.01270171, 
    0.008256259,
  0.001669037, 0.003867964, 7.942022e-08, 2.761526e-08, 1.371212e-05, 
    0.000308579, 0.05510987, 0.1395017, 0.2393298, 0.03662794, 0.03661907, 
    0.1314564, 0.2454524, 0.1738019, 0.1407703, 0.06433474, 0.02331362, 
    0.02580356, -8.574892e-06, 0.003235124, 0.07333609, 0.03359663, 
    0.0864312, 0.02281115, 0.02481459, 0.004049613, 0.02342508, 1.519928e-06, 
    0.005418483,
  0.05585465, 0.06652552, 0.01012316, 0.007419268, 0.003547357, 0.0002804457, 
    0.05746217, 0.01751591, 0.04961105, 0.1786624, 0.07982445, 0.08397903, 
    0.2055169, 0.2161115, 0.08972644, 0.08524654, 0.07880554, 0.07857493, 
    0.0008729649, 0.0004913062, 0.05807914, 0.05130587, 0.01833366, 
    0.08401975, 0.06274409, 0.0659238, 0.05898778, 0.01860618, 0.003151855,
  0.01897911, 0.06034923, 0.02761378, 0.1256406, 0.08825695, 0.09637222, 
    0.05072728, 0.1763618, 0.1111606, 0.05463919, 0.05398879, 0.1518612, 
    0.1153269, 0.1247738, 0.1078162, 0.1581868, 0.1363834, 0.1277454, 
    0.1254093, 0.02986686, 0.04087697, 0.09336622, 0.1121403, 0.08609926, 
    0.1003274, 0.1196821, 0.1307795, 0.1211499, 0.06842935,
  0.08045439, 0.06505831, 0.08505021, 0.06822369, 0.1155149, 0.05072459, 
    0.1733803, 0.1275369, 0.09380974, 0.1544466, 0.06137339, 0.1578562, 
    0.2091965, 0.1644261, 0.1108387, 0.1665065, 0.1501951, 0.3386031, 
    0.255956, 0.1040404, 0.06804026, 0.0757083, 0.08573313, 0.1514588, 
    0.1374904, 0.1647506, 0.1226062, 0.1751834, 0.1115396,
  0.2236087, 0.1673449, 0.2313782, 0.1778717, 0.1251868, 0.1381264, 
    0.1365298, 0.05469934, 0.07547282, 0.07846823, 0.06567498, 0.0854255, 
    0.1507286, 0.2516888, 0.2592065, 0.2300808, 0.1833179, 0.07771919, 
    0.1350043, 0.09277646, 0.2002484, 0.2618696, 0.2577322, 0.2797472, 
    0.2617896, 0.2980791, 0.2451439, 0.1616642, 0.1979757,
  0.07587407, 0.1149499, 0.1465332, 0.1236747, 0.08415253, 0.1973625, 
    0.2972801, 0.3021668, 0.2330795, 0.187849, 0.1605066, 0.1743165, 
    0.1699791, 0.140844, 0.1080878, 0.220928, 0.2223451, 0.2367836, 
    0.3123575, 0.226823, 0.1568005, 0.1862392, 0.2617811, 0.1416467, 
    0.2333396, 0.1531953, 0.1794835, 0.1321824, 0.1124198,
  0.001665664, 0.0009907245, 0.0003157849, -0.0003591548, -0.001034094, 
    -0.001709034, -0.002383974, -2.928824e-06, -1.847284e-06, -7.657441e-07, 
    3.157957e-07, 1.397335e-06, 2.478875e-06, 3.560415e-06, -0.00243741, 
    -0.001784925, -0.001132439, -0.0004799544, 0.0001725308, 0.0008250159, 
    0.001477501, -0.002445885, -0.002424512, -0.002403139, -0.002381766, 
    -0.002360394, -0.00233902, -0.002317647, 0.002205616,
  0.04188894, -0.001239319, 7.270479e-05, 0, -2.577557e-05, 0.003863742, 
    0.000210953, -4.634671e-06, 0, 0, -2.36745e-08, -4.91409e-06, 
    0.0006181891, 0.04457829, 0.0585419, 0.09928618, 0.07602967, 0.1122077, 
    0.140772, 0.06700775, 0.04012215, 0.0658159, 0.1560393, 0.2990254, 
    0.1510129, 0.09276594, 0.1611152, 0.188651, 0.08422847,
  0.3504385, 0.4432698, 0.329939, 0.2397791, 0.1103997, 0.09690622, 
    0.02761214, 0.0323054, 0.09144775, 0.2062189, 0.2150687, 0.2875343, 
    0.3252932, 0.2598791, 0.2357133, 0.1462331, 0.1117933, 0.1068593, 
    0.1537281, 0.2381292, 0.3162705, 0.3450754, 0.2890674, 0.4179721, 
    0.2779084, 0.1397329, 0.159841, 0.1198971, 0.2808702,
  0.2590558, 0.1830236, 0.3160676, 0.2428457, 0.2252085, 0.2018976, 
    0.2093275, 0.1998781, 0.1440479, 0.2047015, 0.2643238, 0.2966772, 
    0.268944, 0.2177976, 0.2152491, 0.1526306, 0.1900053, 0.08568822, 
    0.1181756, 0.2012052, 0.2242788, 0.2453017, 0.2001218, 0.2144777, 
    0.2023031, 0.2341867, 0.2632382, 0.2059408, 0.2933687,
  0.2154844, 0.2022146, 0.147139, 0.1566299, 0.1281092, 0.1651174, 0.1274761, 
    0.1459117, 0.2185939, 0.2446447, 0.2405826, 0.2773394, 0.2568274, 
    0.1579453, 0.1086794, 0.1138346, 0.1383286, 0.1134109, 0.1341742, 
    0.1943911, 0.1863231, 0.2012378, 0.2087139, 0.1575399, 0.08897203, 
    0.1071135, 0.201602, 0.2562636, 0.2313154,
  0.1285353, 0.1018482, 0.07982233, 0.1024802, 0.08424401, 0.1233628, 
    0.1145642, 0.117328, 0.09147621, 0.09600074, 0.1411162, 0.1219919, 
    0.1240434, 0.155265, 0.1600582, 0.1661163, 0.1251905, 0.1418708, 
    0.1448291, 0.148725, 0.1897088, 0.1698688, 0.1182319, 0.05207954, 
    0.05969479, 0.04580729, 0.0718344, 0.1404154, 0.1467959,
  0.01388812, 0.014129, 0.0317965, 0.04605232, 0.02724267, 0.02791668, 
    0.01582032, 0.02716338, 0.001222101, 0.004011369, 0.01174592, 0.01042356, 
    0.01898354, 0.01954531, 0.05264231, 0.1093514, 0.09726884, 0.1020165, 
    0.1348414, 0.0769363, 0.05798326, 0.02429356, 0.01285707, 0.003403788, 
    0.04437985, 0.03910075, 0.04617366, 0.09462355, 0.03403863,
  1.220783e-07, 5.812673e-08, 3.044709e-05, 2.560447e-05, -1.060299e-05, 
    -0.0002496027, 0.01196639, 0.003253269, -3.967109e-05, 2.450119e-07, 
    2.409554e-07, 0.002064894, 0.008811773, 0.06630251, 0.1150366, 
    0.03387685, 0.002527342, 0.0332412, -1.005091e-05, 2.411926e-07, 
    -3.342764e-06, 0.01292272, 3.919749e-09, 3.729932e-06, 0.001886243, 
    0.0008576731, 0.008163912, -3.018989e-06, 2.031479e-07,
  3.211871e-07, 3.110648e-07, 2.749123e-06, 6.867833e-07, 0.004137722, 
    0.025258, 0.006494103, 0.04239355, 0.04754603, 0.001057604, 0.03314145, 
    0.04243687, 0.171922, 0.09466571, 0.02570283, 0.003930014, 0.002411823, 
    0.0001185338, 3.251929e-09, 4.32138e-10, 1.288652e-11, 2.923392e-09, 
    2.685663e-06, 0.001933417, 3.055108e-05, 7.654844e-07, 1.426139e-06, 
    7.570637e-07, -3.327066e-06,
  0.02605362, 0.02816611, 0.1000968, 0.01899544, 0.0006471734, 0.01139483, 
    0.01097233, 0.01381331, 0.01599668, 0.01982987, 0.04550301, 0.1135294, 
    0.1393845, 0.08288789, 0.05402698, 0.0343046, 0.006604592, 0.006994789, 
    0.02770399, 0.002923213, -5.614714e-05, 5.026153e-05, 0.001947709, 
    0.08241448, 0.07598473, 0.04761796, 0.01222839, 0.002209766, 0.007278648,
  0.04935496, 0.1262029, 0.1903358, 0.4585755, 0.1364124, 0.03881847, 
    0.1399968, 0.0481091, 0.1024737, 0.2056693, 0.1240689, 0.1885739, 
    0.2580377, 0.1580821, 0.08296657, 0.1210848, 0.1381527, 0.1625571, 
    0.1453401, 0.1193141, 0.2585413, 0.1628335, 0.1771564, 0.05908441, 
    0.05049854, 0.08783594, 0.1293996, 0.2166388, 0.1681922,
  0.001431822, 3.702005e-07, 2.554482e-05, -7.92507e-07, 0.02199227, 
    0.1083139, 0.6886118, 0.1769583, 0.5323683, 0.07246237, 0.3001554, 
    0.2338102, 0.09779271, 0.02877649, 0.0130768, 0.006036224, 0.0008243439, 
    7.959472e-05, 0.01525102, 0.004071725, 0.0421332, 0.03528018, 0.0125245, 
    0.02989456, 0.01493406, 0.003289445, 0.002281999, 0.01201321, 0.0008006368,
  7.511292e-05, 0.0004125593, 7.089889e-08, 2.09179e-08, 7.272994e-06, 
    0.0005752338, 0.06281052, 0.1654301, 0.2563238, 0.04839418, 0.03759573, 
    0.1272564, 0.2659085, 0.2156322, 0.1417916, 0.0725291, 0.02372973, 
    0.007952549, 0.0004063417, -4.624621e-05, 0.07479481, 0.04577286, 
    0.1054548, 0.0351548, 0.02921898, 0.002627475, 0.006035063, 4.609058e-06, 
    0.0009219155,
  0.05492174, 0.0834462, 0.01156504, 0.01160121, 8.105944e-05, 2.785799e-06, 
    0.05887427, 0.007970532, 0.03270773, 0.1883093, 0.08986204, 0.07131943, 
    0.2505755, 0.2347627, 0.1128855, 0.0691442, 0.08270491, 0.07646032, 
    0.0003087173, 0.0005281101, 0.02710525, 0.05793451, 0.02814151, 0.104887, 
    0.06977279, 0.06002209, 0.06487001, 0.008500527, 0.02269787,
  0.04104097, 0.0739282, 0.04213218, 0.1413265, 0.07893009, 0.08514448, 
    0.06466996, 0.1829359, 0.1165735, 0.06064795, 0.06558412, 0.1780591, 
    0.1062108, 0.1444265, 0.1166939, 0.1851919, 0.1674033, 0.1463364, 
    0.185607, 0.02254945, 0.04240748, 0.08183349, 0.1238873, 0.09324956, 
    0.1066635, 0.1280559, 0.1411767, 0.1242456, 0.05331618,
  0.05921194, 0.06697308, 0.09184527, 0.04898812, 0.1021652, 0.05349367, 
    0.1770735, 0.1348073, 0.10036, 0.1508532, 0.06716213, 0.1667511, 
    0.2189378, 0.1854035, 0.1256497, 0.1782264, 0.1503444, 0.341277, 
    0.307083, 0.09518027, 0.06067485, 0.09282281, 0.09993681, 0.1730799, 
    0.1417831, 0.1604574, 0.1419147, 0.1755165, 0.1511399,
  0.2230674, 0.1901469, 0.2317823, 0.1529663, 0.1041709, 0.1586324, 
    0.1746111, 0.0840346, 0.06819595, 0.07726602, 0.08432478, 0.09231793, 
    0.1835574, 0.227284, 0.2805041, 0.2215057, 0.1885576, 0.08905378, 
    0.1232079, 0.09492989, 0.1881327, 0.2510801, 0.2761202, 0.3364899, 
    0.2531437, 0.2940874, 0.2646833, 0.1253785, 0.1827769,
  0.08286488, 0.1140838, 0.1865501, 0.1828789, 0.1925725, 0.2872108, 
    0.2876683, 0.3190179, 0.26777, 0.1870317, 0.1634646, 0.2221814, 
    0.2234639, 0.1362755, 0.09184634, 0.1427946, 0.1879443, 0.2121973, 
    0.1913035, 0.1194019, 0.08851761, 0.1562245, 0.2585797, 0.1266254, 
    0.2193535, 0.1613896, 0.2161442, 0.1542201, 0.1059252,
  0.02388384, 0.02115944, 0.01843505, 0.01571065, 0.01298626, 0.01026186, 
    0.007537468, 0.01402848, 0.01423109, 0.01443369, 0.0146363, 0.0148389, 
    0.01504151, 0.01524411, 0.009035141, 0.01134411, 0.01365307, 0.01596204, 
    0.018271, 0.02057997, 0.02288894, 0.02601385, 0.02622668, 0.0264395, 
    0.02665233, 0.02686515, 0.02707797, 0.0272908, 0.02606335,
  0.04975493, 0.00279889, 0.005217889, -0.0001508479, 0.0007124855, 
    0.01095153, 0.003865619, 0.001301014, -4.677615e-08, 3.948568e-06, 
    0.000551165, -2.722231e-05, 0.01241486, 0.03798392, 0.05322285, 
    0.09803265, 0.08392055, 0.1238957, 0.1586632, 0.1163837, 0.08935896, 
    0.1118092, 0.2401415, 0.2798717, 0.171707, 0.1074539, 0.1789361, 
    0.2004602, 0.1305017,
  0.3831985, 0.4529211, 0.3202178, 0.2413524, 0.1348893, 0.09070169, 
    0.03448511, 0.07805908, 0.1631929, 0.2730699, 0.2747796, 0.3885804, 
    0.3389992, 0.2781536, 0.2381759, 0.1487325, 0.1189058, 0.125573, 
    0.1820767, 0.2779817, 0.3043161, 0.3061667, 0.2844365, 0.4249909, 
    0.2814994, 0.1286007, 0.1494865, 0.1091327, 0.2623738,
  0.2725483, 0.1908851, 0.3069762, 0.2432182, 0.2237453, 0.2049552, 
    0.2196988, 0.2008457, 0.1567765, 0.213948, 0.2524197, 0.2880411, 
    0.2606326, 0.2280248, 0.1910975, 0.1763944, 0.1666612, 0.06592732, 
    0.128877, 0.2064209, 0.2122336, 0.2408828, 0.2005443, 0.2078713, 
    0.1910466, 0.2657989, 0.2429056, 0.2077812, 0.2992581,
  0.2119436, 0.1984306, 0.16512, 0.1755579, 0.1651785, 0.142075, 0.1422345, 
    0.1696419, 0.236659, 0.2651919, 0.2534495, 0.2861601, 0.2506217, 
    0.1668934, 0.1084446, 0.1102519, 0.1154794, 0.1174082, 0.1479935, 
    0.2009352, 0.1885147, 0.2070016, 0.2097641, 0.155977, 0.0885089, 
    0.09682454, 0.2127162, 0.2351463, 0.2089781,
  0.1393223, 0.07993613, 0.08757235, 0.1004085, 0.08781181, 0.1210074, 
    0.1225534, 0.1237356, 0.09450285, 0.09750762, 0.1289955, 0.1270847, 
    0.1305491, 0.1725222, 0.1639874, 0.1638959, 0.1233525, 0.1397181, 
    0.1421496, 0.1618998, 0.1772969, 0.1635638, 0.09568661, 0.05342326, 
    0.07408899, 0.04641563, 0.07111005, 0.1433684, 0.1596368,
  0.01728451, 0.01663961, 0.03576639, 0.04782587, 0.03033476, 0.02866448, 
    0.02653521, 0.03487283, 0.005783312, 0.006159049, 0.04050106, 0.01400166, 
    0.02207596, 0.0296151, 0.06081617, 0.1014855, 0.08760879, 0.09902055, 
    0.1315817, 0.08473323, 0.05911799, 0.03362754, 0.01651177, 0.002766516, 
    0.04035374, 0.04123749, 0.05605789, 0.09914932, 0.03300229,
  1.451473e-07, 1.083378e-07, 0.0003132776, 0.0009678106, 0.000241275, 
    0.0006602454, 0.01219595, 0.005388756, 0.0002837504, -3.740568e-06, 
    0.0001138826, 0.001194609, 0.001654216, 0.04047475, 0.1381874, 
    0.04378769, 0.003770876, 0.03651197, 6.34146e-06, 8.664595e-06, 
    -1.651873e-05, 0.01661645, 3.498428e-09, 1.646055e-06, 0.001217392, 
    0.001196442, 0.01977061, 9.480969e-05, 1.401359e-07,
  3.387877e-07, -3.100408e-06, 1.987019e-06, 0.0004107646, 0.01332089, 
    0.04124265, 0.005590334, 0.04628469, 0.04819421, 0.002083703, 0.0157074, 
    0.05013639, 0.1643467, 0.08703467, 0.02771898, 0.004516368, 0.002351296, 
    7.927306e-05, -3.622113e-07, 8.184753e-10, 8.751412e-11, 1.131259e-08, 
    1.998514e-06, 0.002374453, 3.220001e-05, -6.415054e-07, 6.653044e-06, 
    6.663585e-07, -2.5604e-08,
  0.01116255, 0.02099566, 0.1414078, 0.01207484, 0.0006217007, 0.006216553, 
    0.01007885, 0.01279948, 0.01578227, 0.02349419, 0.03464385, 0.06780993, 
    0.1086801, 0.07397529, 0.05419526, 0.02896512, 0.004756584, 0.007831793, 
    0.02794864, 0.005879691, -4.409703e-05, 0.0008106442, 0.008415899, 
    0.1072212, 0.09580354, 0.03621987, 0.01918779, 0.003421713, 0.003941212,
  0.03978504, 0.1389776, 0.2140076, 0.4669966, 0.05712774, 0.03048308, 
    0.1486379, 0.03271131, 0.04560024, 0.1464063, 0.05653692, 0.1220395, 
    0.1835213, 0.1263039, 0.081474, 0.1223118, 0.1382607, 0.1591349, 
    0.1557527, 0.1414004, 0.27043, 0.142419, 0.1832988, 0.06911379, 
    0.03779421, 0.1075564, 0.1239527, 0.1967684, 0.1842534,
  0.0001456563, 5.384439e-08, 1.394617e-06, 4.879751e-07, 0.0003365885, 
    0.0956675, 0.5758546, 0.186161, 0.5571743, 0.07408863, 0.2483656, 
    0.1830532, 0.08013915, 0.02609133, 0.01339534, 0.006633537, 0.001443819, 
    -1.901389e-05, 0.006859304, 0.0006390305, 0.02722512, 0.02842309, 
    0.01097056, 0.02180312, 0.01551505, 0.001578806, 0.00011869, 0.009272358, 
    6.557778e-05,
  2.994852e-05, 5.264928e-05, 2.661906e-08, 6.266488e-09, 3.412732e-06, 
    0.0005920657, 0.06614338, 0.2116618, 0.3002819, 0.05300214, 0.03274223, 
    0.09419294, 0.2191333, 0.2072747, 0.1396087, 0.06901028, 0.01560605, 
    0.001243888, 0.001104316, -5.367691e-07, 0.05273913, 0.04003564, 
    0.08435488, 0.03424243, 0.02591718, 0.00192777, 0.000748676, 
    7.423798e-06, 0.0004399137,
  0.05495218, 0.05163659, 0.01945241, 0.01388321, -7.956092e-05, 
    7.297644e-07, 0.03014648, 0.006399103, 0.01466049, 0.1913172, 0.08223162, 
    0.06911595, 0.2670984, 0.23631, 0.1274747, 0.06615572, 0.08655836, 
    0.07587331, 0.0004480835, 0.0006926758, 0.01411794, 0.0383793, 
    0.03244177, 0.1110431, 0.07377411, 0.06747935, 0.08572032, 0.01827118, 
    0.02911767,
  0.02068992, 0.08506694, 0.04677493, 0.1525512, 0.1100336, 0.07607669, 
    0.07767823, 0.1951521, 0.1030336, 0.05967527, 0.07364868, 0.206484, 
    0.1228802, 0.1572355, 0.1497238, 0.1926207, 0.1950169, 0.1622613, 
    0.1724511, 0.02179932, 0.05580641, 0.04708986, 0.1326981, 0.1099077, 
    0.110038, 0.148995, 0.1474065, 0.1406139, 0.04169415,
  0.06528109, 0.08031911, 0.1028673, 0.06368498, 0.1161043, 0.0675102, 
    0.1816673, 0.132811, 0.1168528, 0.1748528, 0.0711806, 0.1703001, 
    0.2332146, 0.2053835, 0.1354945, 0.245054, 0.1374323, 0.3592083, 
    0.314479, 0.09280296, 0.06945881, 0.09029051, 0.1134091, 0.1728758, 
    0.1325363, 0.1554086, 0.1024863, 0.173987, 0.1402559,
  0.2258493, 0.1424607, 0.2402551, 0.1767059, 0.1199637, 0.1518547, 0.140715, 
    0.07215207, 0.08163187, 0.06898723, 0.06906283, 0.1006932, 0.1779081, 
    0.2574375, 0.3152182, 0.2373689, 0.1857379, 0.09224482, 0.09316504, 
    0.1017228, 0.1650525, 0.2857159, 0.2360926, 0.3415288, 0.2352709, 
    0.3345815, 0.2703446, 0.1400621, 0.1942311,
  0.08831993, 0.08807055, 0.1747143, 0.1599746, 0.1521947, 0.2239272, 
    0.2641135, 0.274539, 0.2654886, 0.2074221, 0.2404442, 0.3189353, 
    0.2317604, 0.13116, 0.1124465, 0.2005378, 0.1538693, 0.2482584, 
    0.2398777, 0.09910046, 0.0875755, 0.1685797, 0.2378191, 0.1170747, 
    0.196963, 0.2106339, 0.2399231, 0.1794095, 0.09408903,
  0.0499032, 0.04821989, 0.04653659, 0.04485329, 0.04316999, 0.04148668, 
    0.03980338, 0.0388468, 0.03841291, 0.03797903, 0.03754515, 0.03711127, 
    0.03667739, 0.03624351, 0.04334953, 0.04600516, 0.04866078, 0.0513164, 
    0.05397203, 0.05662765, 0.05928327, 0.05031749, 0.04977905, 0.04924061, 
    0.04870217, 0.04816373, 0.04762529, 0.04708685, 0.05124984,
  0.07182139, 0.03350017, 0.02272072, 0.005075698, 0.009918905, 0.03821428, 
    0.03037602, 0.02712945, 0.01341297, 0.006483639, 0.009704929, 
    0.001366593, 0.01112551, 0.02411522, 0.02448378, 0.08336163, 0.07635378, 
    0.1265818, 0.1710798, 0.1295678, 0.1570093, 0.3050327, 0.297882, 
    0.272889, 0.1741299, 0.1183823, 0.1984785, 0.2093006, 0.1859515,
  0.4151387, 0.4517686, 0.3202672, 0.2472208, 0.1339902, 0.0804897, 
    0.03829278, 0.1315934, 0.2459091, 0.3142164, 0.3135507, 0.399426, 
    0.3388601, 0.2786869, 0.25404, 0.1676876, 0.124687, 0.1395357, 0.194788, 
    0.2960759, 0.3169557, 0.3740648, 0.3014144, 0.4573137, 0.317717, 
    0.167078, 0.1955783, 0.1471065, 0.3299303,
  0.3276822, 0.1982021, 0.3160209, 0.2422759, 0.2285194, 0.233525, 0.1979779, 
    0.226128, 0.1930865, 0.2529712, 0.2985134, 0.2822614, 0.2482683, 
    0.2268485, 0.1977277, 0.1643455, 0.1723408, 0.08450759, 0.1425972, 
    0.2266598, 0.2501574, 0.2487328, 0.2038363, 0.2206215, 0.1904534, 
    0.2676295, 0.2359766, 0.2171761, 0.2900924,
  0.2223317, 0.1855816, 0.1682134, 0.1859962, 0.1480579, 0.1443593, 
    0.1670724, 0.2033518, 0.2797536, 0.2786035, 0.2838553, 0.2671245, 
    0.2402858, 0.1904912, 0.1217558, 0.09413223, 0.119225, 0.1070272, 
    0.1898366, 0.192859, 0.1930267, 0.2013834, 0.2032617, 0.1584543, 
    0.0840183, 0.1003359, 0.1991768, 0.2354161, 0.2312821,
  0.1667376, 0.1015276, 0.09911969, 0.1005445, 0.09398723, 0.1438286, 
    0.1280769, 0.1254248, 0.1117276, 0.1194475, 0.1236922, 0.1302787, 
    0.1355888, 0.1610534, 0.1702395, 0.1719722, 0.1541175, 0.1549426, 
    0.1497507, 0.1556928, 0.1906144, 0.1665106, 0.07658911, 0.05467453, 
    0.09125043, 0.05101439, 0.08048663, 0.1579197, 0.1601632,
  0.02263561, 0.02064892, 0.0500689, 0.04584202, 0.04113375, 0.03073978, 
    0.04411577, 0.04984574, 0.005908308, 0.008543095, 0.0300791, 0.01171072, 
    0.01772643, 0.04341875, 0.0731812, 0.09500435, 0.08084025, 0.0923908, 
    0.1358354, 0.09671998, 0.07141496, 0.03690216, 0.01701566, 0.002415167, 
    0.04756305, 0.04696227, 0.06153525, 0.09788699, 0.03785125,
  6.729441e-08, 7.666919e-08, 0.0005047769, 0.00435554, 0.004100084, 
    0.002465101, 0.01759518, 0.01018886, 0.02785559, -2.282639e-05, 
    0.00242715, -0.0008255339, -0.0003716486, 0.02429716, 0.1291003, 
    0.05795036, 0.004630613, 0.03206233, 0.001079654, 0.0006236525, 
    0.000274114, 0.01711361, 6.844356e-10, 5.341493e-07, 0.001091345, 
    0.00241563, 0.05150571, 0.0009855729, 8.978414e-08,
  1.568957e-07, -7.579457e-05, 6.651381e-07, 0.006126864, 0.01651789, 
    0.04778777, 0.005271778, 0.04442504, 0.04743611, 0.0009783886, 
    0.003557373, 0.05380064, 0.1799216, 0.08928415, 0.03123726, 0.006046916, 
    0.0036026, 0.0007531003, 0.0001293573, 9.726207e-08, 3.172794e-09, 
    2.468498e-08, 3.435176e-07, 0.004000662, 0.001504142, 0.0006209126, 
    0.001403319, 3.471547e-07, 7.867168e-08,
  0.003952362, 0.01422776, 0.1351838, 0.02188906, 0.0006959777, 0.002944442, 
    0.009002135, 0.014763, 0.0177849, 0.01838744, 0.02488937, 0.03727375, 
    0.08992934, 0.0689119, 0.05125483, 0.02857199, 0.01204887, 0.004915903, 
    0.02093035, 0.003586312, 0.0006308525, 0.0005302511, 0.01904827, 
    0.1322106, 0.1139223, 0.0231326, 0.0261098, 0.007343098, 0.0004027689,
  0.02570806, 0.07564961, 0.1340178, 0.4911284, 0.02252175, 0.01661518, 
    0.1496366, 0.02826894, 0.01739234, 0.09593804, 0.02487067, 0.08857137, 
    0.145296, 0.104222, 0.0771306, 0.1119578, 0.1354616, 0.1653831, 
    0.1647545, 0.1589913, 0.2564474, 0.1382865, 0.1637804, 0.06266294, 
    0.0299575, 0.09208096, 0.1211816, 0.1514273, 0.1440704,
  9.111729e-06, 9.803547e-09, 1.430127e-07, 7.200329e-07, 3.574532e-05, 
    0.06668142, 0.4845566, 0.2036702, 0.4650767, 0.0850822, 0.2158158, 
    0.1390456, 0.0672477, 0.02020508, 0.01325574, 0.008990526, 0.0008035164, 
    4.628346e-06, 0.009922696, 5.541254e-05, 0.01997682, 0.02685837, 
    0.01024841, 0.01762487, 0.01758965, 0.0007518449, 3.972333e-05, 
    0.001962037, -3.413526e-07,
  1.253889e-05, 2.255298e-05, 1.218578e-08, 1.929967e-09, 1.533526e-06, 
    0.0002747609, 0.06284138, 0.2035471, 0.3604055, 0.06772871, 0.03790655, 
    0.07087503, 0.1616133, 0.1341983, 0.123504, 0.06343336, 0.007749423, 
    2.264017e-05, 0.001183525, 7.605105e-07, 0.02418003, 0.01911923, 
    0.07942751, 0.02861777, 0.01081717, 0.002196043, 0.0003855481, 
    5.141887e-06, 1.141596e-05,
  0.06391197, 0.03459374, 0.02845835, 0.01751934, -6.189797e-05, 
    1.833571e-07, 0.0129133, 0.001646846, 0.004273904, 0.1487506, 0.07357961, 
    0.06984696, 0.2378952, 0.230802, 0.1438724, 0.103909, 0.1001772, 
    0.07862818, 0.001139054, 0.0003676541, 0.006308501, 0.01060465, 
    0.02239602, 0.07161637, 0.06182911, 0.064652, 0.06457137, 0.01983922, 
    0.01726463,
  0.03511606, 0.0911384, 0.05858267, 0.1842182, 0.1037318, 0.08058676, 
    0.07261369, 0.2344209, 0.1021123, 0.05596146, 0.07787431, 0.221999, 
    0.09995287, 0.1629609, 0.1411707, 0.2585323, 0.2240226, 0.2162122, 
    0.1980635, 0.02817411, 0.05838388, 0.03794419, 0.1316843, 0.1180874, 
    0.1153094, 0.1366396, 0.1549153, 0.155819, 0.04721359,
  0.06607038, 0.08516088, 0.1007525, 0.1028308, 0.174337, 0.0832319, 
    0.1918604, 0.1368823, 0.1347934, 0.2062518, 0.09388244, 0.1920111, 
    0.2410169, 0.2215254, 0.1386008, 0.2719499, 0.1504285, 0.3856755, 
    0.3133677, 0.1009461, 0.08671597, 0.1144164, 0.1257146, 0.1641111, 
    0.1373635, 0.1703703, 0.1316999, 0.1752989, 0.1717671,
  0.2256483, 0.2132217, 0.2792103, 0.1633764, 0.1290816, 0.1432075, 0.137336, 
    0.05503481, 0.1054682, 0.09067692, 0.1026657, 0.1605077, 0.1704254, 
    0.2555698, 0.3021362, 0.1666482, 0.1845595, 0.1281028, 0.1019968, 
    0.09939408, 0.2030073, 0.2722383, 0.3027902, 0.3461272, 0.2303425, 
    0.3731565, 0.3503708, 0.1604468, 0.2093402,
  0.1663582, 0.1178791, 0.258922, 0.1904377, 0.2255507, 0.2427646, 0.3057017, 
    0.3173164, 0.2497141, 0.1506484, 0.219848, 0.2346669, 0.2642115, 
    0.1928591, 0.1459526, 0.1576548, 0.1766684, 0.2482059, 0.2327468, 
    0.1316479, 0.1354203, 0.1594655, 0.2387925, 0.1024268, 0.2064734, 
    0.1888339, 0.2085714, 0.1850755, 0.119932,
  0.08085403, 0.07733684, 0.07381966, 0.07030248, 0.06678529, 0.06326811, 
    0.05975093, 0.06507412, 0.06479787, 0.06452163, 0.06424538, 0.06396914, 
    0.0636929, 0.06341665, 0.05894035, 0.06400046, 0.06906057, 0.07412069, 
    0.0791808, 0.08424091, 0.08930103, 0.07180566, 0.07053898, 0.06927229, 
    0.06800561, 0.06673892, 0.06547223, 0.06420555, 0.08366777,
  0.1194001, 0.07778943, 0.06537564, 0.02206232, 0.01743705, 0.06352977, 
    0.0480464, 0.04941972, 0.02305329, 0.0383653, 0.009639305, 0.01575303, 
    0.02126198, 0.01455517, 0.009038932, 0.06838615, 0.0727092, 0.1126934, 
    0.169838, 0.1228978, 0.1850453, 0.4395719, 0.3499011, 0.2693197, 
    0.186513, 0.1175132, 0.2413989, 0.2236508, 0.2047852,
  0.4872804, 0.4950539, 0.3241335, 0.2535706, 0.1374974, 0.07134117, 
    0.0547134, 0.1408719, 0.2851982, 0.3403605, 0.3590285, 0.4492536, 
    0.3255285, 0.2802909, 0.2641619, 0.1517635, 0.1102859, 0.134848, 
    0.1949186, 0.3342776, 0.3375933, 0.3642102, 0.2773851, 0.4654158, 
    0.3261651, 0.1558893, 0.1764086, 0.1593657, 0.3632447,
  0.3372477, 0.2120526, 0.3379532, 0.2331759, 0.2460686, 0.270198, 0.2180182, 
    0.2546099, 0.248704, 0.2819125, 0.3284942, 0.2922247, 0.300413, 
    0.2461433, 0.2656065, 0.1809649, 0.185769, 0.1077795, 0.1817352, 
    0.2246944, 0.3062701, 0.2623, 0.2094095, 0.2276035, 0.2049622, 0.2811204, 
    0.2667723, 0.2680234, 0.2845125,
  0.2540118, 0.1998403, 0.1873121, 0.1983927, 0.1732928, 0.1509478, 
    0.1805092, 0.2221477, 0.2736505, 0.2703308, 0.2935791, 0.2585135, 
    0.2522378, 0.2062792, 0.1240398, 0.1185028, 0.1466113, 0.1427869, 
    0.1958983, 0.1770429, 0.1885718, 0.2098248, 0.2123201, 0.1737704, 
    0.08593606, 0.1089124, 0.2106041, 0.2508627, 0.2399668,
  0.1907303, 0.1184955, 0.1155588, 0.1013774, 0.1071965, 0.1578298, 0.147424, 
    0.1400443, 0.1217209, 0.1351366, 0.1293634, 0.1460837, 0.1383378, 
    0.1595215, 0.176473, 0.1839661, 0.1778613, 0.1608171, 0.1635307, 
    0.1521732, 0.1999289, 0.1858694, 0.0778674, 0.05943211, 0.09333132, 
    0.06736178, 0.1095741, 0.1762733, 0.1849353,
  0.04020014, 0.03375218, 0.05579365, 0.04261701, 0.06182458, 0.0362026, 
    0.0497461, 0.06506847, 0.01407399, 0.01131054, 0.01305726, 0.00292976, 
    0.01631319, 0.05954371, 0.08885364, 0.09486046, 0.08558501, 0.0932796, 
    0.1380913, 0.1031304, 0.09507236, 0.05609325, 0.01700719, 0.001620205, 
    0.06344522, 0.05947479, 0.07793265, 0.1082594, 0.04796222,
  -2.608377e-07, 2.711052e-08, 6.351082e-05, 0.01452984, 0.02357305, 
    0.008778517, 0.0234806, 0.01596106, 0.05094697, 0.05762776, 0.0002966821, 
    -0.0001029963, 0.003815544, 0.01652525, 0.1097961, 0.1131508, 0.02478507, 
    0.02718528, 0.007763691, 0.002388119, 0.003271157, 0.01439375, 
    9.09123e-08, 2.290391e-07, 0.009979444, 0.00370258, 0.06245562, 
    0.002045717, 9.558094e-06,
  1.095281e-07, -4.032418e-06, 1.901755e-07, 0.04292428, 0.03232195, 
    0.0543486, 0.002879109, 0.0401696, 0.04486328, 0.001901989, 0.01683525, 
    0.05919546, 0.2014183, 0.09105173, 0.03663085, 0.01385382, 0.008429754, 
    0.00709302, 0.002792013, 6.332321e-05, 6.071086e-07, 3.040785e-08, 
    1.289366e-07, 0.005790813, 0.05906192, 0.008985235, 0.01896685, 
    3.91951e-05, 3.108154e-08,
  0.000494846, 0.01078837, 0.1438312, 0.03727178, 0.001472424, 0.003269629, 
    0.01012511, 0.01606649, 0.02309202, 0.01744835, 0.02206223, 0.0246032, 
    0.08080009, 0.06399532, 0.0516329, 0.04246769, 0.02525551, 0.005625714, 
    0.01977205, 0.001715654, 0.0009792703, 0.001392293, 0.02838073, 
    0.1531084, 0.1474317, 0.0202215, 0.01517901, 0.003145061, 0.001051446,
  0.02402831, 0.04595203, 0.08309077, 0.4715319, 0.01269907, 0.009583371, 
    0.1479142, 0.02639512, 0.01161542, 0.06119429, 0.01113496, 0.06899563, 
    0.1166679, 0.08723599, 0.08085339, 0.1089422, 0.1324943, 0.1767968, 
    0.1783534, 0.1668106, 0.2421809, 0.1372217, 0.1631297, 0.05764098, 
    0.02441516, 0.08441902, 0.1280562, 0.1404149, 0.1425351,
  2.284834e-06, 3.076275e-09, 1.591646e-08, 5.979118e-07, 1.875962e-06, 
    0.04878817, 0.4149407, 0.2460088, 0.4365859, 0.09679168, 0.1963017, 
    0.1181641, 0.06047346, 0.02584697, 0.01818675, 0.01283918, 0.0004414817, 
    7.011909e-06, 0.0126789, 2.173313e-05, 0.01636089, 0.03123934, 
    0.01021181, 0.01682987, 0.02152238, 0.002937647, 2.476528e-05, 
    0.0003518218, -2.297078e-06,
  5.913839e-06, 1.118169e-05, 8.134543e-09, 1.128716e-09, 9.655508e-07, 
    8.706714e-05, 0.05660001, 0.2026461, 0.3745982, 0.08088862, 0.03895599, 
    0.05828641, 0.1257911, 0.09452105, 0.09483174, 0.04347359, 0.01003746, 
    9.08731e-06, 0.0003911119, 2.886755e-07, 0.00767839, 0.02133005, 
    0.09026991, 0.02547086, 0.007912739, 0.003584442, 0.0007723966, 
    1.095083e-05, 1.771865e-06,
  0.04910366, 0.02976318, 0.02503226, 0.0222782, -2.556034e-05, 4.313328e-08, 
    0.003753262, 2.03e-05, 0.001526399, 0.1123208, 0.07404581, 0.07660472, 
    0.2282968, 0.1732767, 0.09521052, 0.1222359, 0.1184305, 0.08272429, 
    0.01852026, 0.0002367162, 0.002968239, 0.003827349, 0.02303769, 
    0.06257134, 0.05134759, 0.06442229, 0.05283284, 0.01103893, 0.00465558,
  0.03826183, 0.1075713, 0.07171481, 0.1932655, 0.07824391, 0.07949557, 
    0.08422114, 0.2417793, 0.1210023, 0.03912299, 0.07135858, 0.2326651, 
    0.07605286, 0.1577056, 0.1566076, 0.2911361, 0.2480629, 0.1856697, 
    0.2012919, 0.04077043, 0.05219514, 0.02884492, 0.1251318, 0.1359303, 
    0.1224805, 0.1302301, 0.1469479, 0.1587122, 0.0466213,
  0.06801858, 0.106198, 0.1346343, 0.1784511, 0.175547, 0.09241056, 
    0.1853369, 0.1852082, 0.1569103, 0.2216298, 0.1159848, 0.2300741, 
    0.2703424, 0.2408703, 0.1590011, 0.2765438, 0.1660171, 0.4001263, 
    0.349066, 0.1127801, 0.132071, 0.1754774, 0.1550251, 0.1925344, 
    0.1628308, 0.1770111, 0.1383689, 0.1743174, 0.1779754,
  0.2776181, 0.216122, 0.3394124, 0.2346317, 0.1723274, 0.1410119, 0.1510419, 
    0.07073457, 0.1575494, 0.0957863, 0.118744, 0.1633354, 0.1843824, 
    0.2923654, 0.3291096, 0.2004247, 0.2113698, 0.1194892, 0.1105412, 
    0.1249231, 0.2012173, 0.2652593, 0.2594052, 0.3670338, 0.2226206, 
    0.3992048, 0.3451746, 0.1748089, 0.2428194,
  0.1644105, 0.1967767, 0.3272951, 0.2192471, 0.1852945, 0.1988638, 
    0.2643213, 0.2933468, 0.2527376, 0.1441348, 0.1939871, 0.2291018, 
    0.2005535, 0.2157597, 0.1874844, 0.1565273, 0.2044907, 0.23659, 
    0.2188737, 0.07852653, 0.1022925, 0.1585774, 0.2051911, 0.09536128, 
    0.1642791, 0.179083, 0.2261657, 0.2057568, 0.1749441,
  0.1517885, 0.1415054, 0.1312223, 0.1209391, 0.110656, 0.1003729, 
    0.09008975, 0.1107574, 0.1120048, 0.1132521, 0.1144994, 0.1157468, 
    0.1169941, 0.1182414, 0.1437705, 0.155001, 0.1662314, 0.1774618, 
    0.1886922, 0.1999226, 0.211153, 0.2151315, 0.2129369, 0.2107423, 
    0.2085477, 0.206353, 0.2041584, 0.2019638, 0.160015,
  0.1371081, 0.1055079, 0.1076041, 0.02945217, 0.0391835, 0.08818945, 
    0.05582544, 0.06072592, 0.04535293, 0.05347211, 0.02822234, 0.02402824, 
    0.02227536, 0.01152533, 0.007044737, 0.06062346, 0.06862225, 0.100134, 
    0.1492109, 0.1078398, 0.2109481, 0.4806925, 0.3603082, 0.24951, 
    0.1798909, 0.1233137, 0.294752, 0.2316951, 0.2258357,
  0.5072373, 0.5120538, 0.3556292, 0.2481799, 0.1331668, 0.07393526, 
    0.0552828, 0.162048, 0.3079028, 0.3632942, 0.3979449, 0.4544295, 
    0.3143775, 0.2545081, 0.2446725, 0.1339669, 0.1171861, 0.1602294, 
    0.2084059, 0.3070534, 0.3492515, 0.3176575, 0.2593345, 0.4404603, 
    0.2947781, 0.1251087, 0.1523839, 0.1769551, 0.3966967,
  0.3223525, 0.2221972, 0.3195148, 0.2128775, 0.2724209, 0.2607007, 
    0.1847659, 0.2739003, 0.2494965, 0.2879849, 0.2756606, 0.2979283, 
    0.2954006, 0.2318444, 0.2834642, 0.2927344, 0.2480325, 0.1682803, 
    0.2221904, 0.2636018, 0.3215813, 0.2743544, 0.20987, 0.2554646, 
    0.1856228, 0.2672874, 0.2793418, 0.2949437, 0.2850246,
  0.2436845, 0.2115854, 0.2057654, 0.211362, 0.1976955, 0.1877537, 0.1853923, 
    0.2558917, 0.2666329, 0.2779318, 0.2771163, 0.241174, 0.2483897, 
    0.2058056, 0.1528841, 0.1434679, 0.1651513, 0.1509078, 0.21839, 
    0.1856637, 0.1883561, 0.2199931, 0.1997442, 0.2040244, 0.09011932, 
    0.1216317, 0.2328006, 0.2696456, 0.2625994,
  0.1975486, 0.1528696, 0.129954, 0.1166322, 0.1227143, 0.1734599, 0.1677279, 
    0.1697035, 0.1517444, 0.1401049, 0.1467643, 0.1696311, 0.1397428, 
    0.168924, 0.1950206, 0.1932471, 0.1978341, 0.1873049, 0.1919799, 
    0.1650487, 0.2053778, 0.1901487, 0.102331, 0.07018371, 0.08317079, 
    0.1003839, 0.1461956, 0.1920862, 0.2204416,
  0.05336695, 0.03150215, 0.04531569, 0.04539063, 0.0529073, 0.04495775, 
    0.05477669, 0.06253074, 0.04151062, 0.02357508, 0.01514394, 0.001417213, 
    0.01082908, 0.07089927, 0.09692748, 0.0969954, 0.1031185, 0.07728354, 
    0.1289099, 0.1123685, 0.09911697, 0.07807749, 0.01860516, 0.002037834, 
    0.06946743, 0.07171498, 0.08835147, 0.1198481, 0.06300282,
  1.219813e-05, 2.236307e-08, 0.0001011991, 0.03051867, 0.06646946, 
    0.02356681, 0.02936594, 0.01056082, 0.06815293, 0.04716923, 3.095647e-06, 
    1.863574e-05, 0.006424204, 0.009338493, 0.09493703, 0.1207088, 
    0.02780998, 0.02768607, 0.01969676, 0.007660451, 0.01430037, 0.01154599, 
    3.27377e-07, 1.537368e-07, 0.01568576, 0.005057419, 0.08759142, 
    0.01428331, 0.002283605,
  5.5701e-08, -1.120189e-06, -1.725128e-05, 0.159635, 0.0399251, 0.05408945, 
    0.005128162, 0.04053682, 0.04698127, 0.005430223, 0.03891258, 0.05462567, 
    0.2198016, 0.08923477, 0.0391045, 0.02245838, 0.01941395, 0.01757208, 
    0.01394375, 0.003580932, 0.0001843968, 2.70952e-08, 2.884289e-08, 
    0.007767473, 0.0437627, 0.01700182, 0.03648629, 0.001839805, 3.300508e-07,
  3.601955e-05, 0.009207645, 0.1135959, 0.05276747, 0.005847665, 0.004457247, 
    0.01252199, 0.01668078, 0.02473373, 0.02118934, 0.02400924, 0.01942267, 
    0.0748497, 0.05664105, 0.05439494, 0.05382721, 0.02539074, 0.007393965, 
    0.01735652, 0.0004775804, 0.0002251639, 0.002185662, 0.02252265, 
    0.1801262, 0.1368441, 0.01918494, 0.01679997, 0.005984039, 4.554696e-05,
  0.0259526, 0.03138559, 0.05826298, 0.4022018, 0.01015853, 0.01031464, 
    0.1349514, 0.02592722, 0.009381882, 0.04097822, 0.009155819, 0.05595847, 
    0.09675525, 0.07385184, 0.0894409, 0.1139486, 0.1336695, 0.1888191, 
    0.1889038, 0.1539372, 0.2359513, 0.1341775, 0.1598346, 0.05921327, 
    0.02237649, 0.0842132, 0.1427661, 0.1385549, 0.1392766,
  9.689063e-07, 1.148017e-09, 2.024693e-09, 1.816921e-07, 5.142043e-07, 
    0.02058404, 0.3797132, 0.2911924, 0.4283025, 0.1093409, 0.1936894, 
    0.1068228, 0.05380206, 0.02429082, 0.02073197, 0.02289198, 0.001621826, 
    0.0002422228, 0.01641249, 4.190199e-06, 0.0151885, 0.03918774, 
    0.01119413, 0.01772073, 0.03020085, 0.01060468, 0.0005128465, 
    4.166191e-05, -9.056466e-07,
  2.684619e-06, 6.296511e-06, -8.006622e-07, 2.406501e-10, 6.242943e-07, 
    3.824049e-05, 0.04740914, 0.2133285, 0.373971, 0.09273235, 0.04466455, 
    0.0521018, 0.1041892, 0.06429645, 0.0842416, 0.03701308, 0.0153197, 
    0.0009562852, 2.622318e-06, 1.147163e-07, 0.002997538, 0.01178819, 
    0.08690886, 0.0241066, 0.01054128, 0.01399428, 0.0008444107, 
    0.0001354942, 2.059294e-06,
  0.02850099, 0.02258964, 0.01694537, 0.03125361, 2.186236e-05, 8.884016e-09, 
    0.000783055, 4.554994e-07, 0.001098949, 0.07199424, 0.08738802, 
    0.09391328, 0.2414897, 0.1617928, 0.08314632, 0.1352712, 0.1146448, 
    0.06759843, 0.0342441, 0.0001554238, 0.0006536928, 0.002797424, 
    0.02438303, 0.05707765, 0.0482498, 0.07574423, 0.03932297, 0.004247006, 
    0.01458587,
  0.03692898, 0.1234359, 0.07481999, 0.1744595, 0.03877192, 0.0505437, 
    0.1049188, 0.2482434, 0.1346115, 0.02518303, 0.06815899, 0.2259334, 
    0.07748104, 0.1711325, 0.1473718, 0.2637492, 0.2821152, 0.2177744, 
    0.2060543, 0.04201138, 0.03901743, 0.02415727, 0.1076188, 0.1669452, 
    0.1298655, 0.1375694, 0.1356873, 0.1419198, 0.04069633,
  0.0553914, 0.1061374, 0.1474324, 0.1488395, 0.1885744, 0.08763348, 
    0.192625, 0.1957694, 0.1541678, 0.2120643, 0.1137096, 0.2615603, 
    0.3022088, 0.2629929, 0.1425897, 0.293037, 0.1821026, 0.4205216, 
    0.3810499, 0.1215762, 0.1530398, 0.1601478, 0.1395856, 0.2244942, 
    0.167167, 0.1881035, 0.1962266, 0.2042673, 0.1697064,
  0.2580709, 0.2620392, 0.3998565, 0.247747, 0.1803322, 0.2162493, 0.1794962, 
    0.09361441, 0.2520105, 0.1291362, 0.1167637, 0.2203433, 0.2368895, 
    0.3419348, 0.3738095, 0.1937269, 0.2293011, 0.1295916, 0.1344318, 
    0.1294517, 0.1944035, 0.2898684, 0.2344287, 0.4092049, 0.2308524, 
    0.3935305, 0.2957329, 0.2087649, 0.2777725,
  0.1693327, 0.2497879, 0.3019583, 0.2538325, 0.1839653, 0.2241965, 0.329751, 
    0.3891225, 0.336751, 0.229061, 0.1960091, 0.2128696, 0.217904, 0.1938745, 
    0.1875967, 0.1469403, 0.2338427, 0.2964484, 0.2164117, 0.07539257, 
    0.08236737, 0.1583646, 0.1970246, 0.1007972, 0.1589682, 0.1246083, 
    0.1568981, 0.1958714, 0.2207163,
  0.3133529, 0.3057201, 0.2980872, 0.2904544, 0.2828216, 0.2751888, 0.267556, 
    0.2644531, 0.2642198, 0.2639865, 0.2637531, 0.2635198, 0.2632865, 
    0.2630532, 0.2762856, 0.284901, 0.2935164, 0.3021317, 0.3107471, 
    0.3193625, 0.3279779, 0.2999263, 0.299177, 0.2984278, 0.2976785, 
    0.2969292, 0.29618, 0.2954307, 0.3194591,
  0.1468954, 0.1349598, 0.1261354, 0.04744729, 0.06065214, 0.0934947, 
    0.1158564, 0.1095218, 0.06999896, 0.06044986, 0.03829031, 0.02444267, 
    0.01774875, 0.01879283, 0.03243168, 0.06192395, 0.07201827, 0.09222794, 
    0.1341496, 0.1257155, 0.2477844, 0.5409208, 0.3943177, 0.258714, 
    0.1769766, 0.1521766, 0.2685771, 0.26076, 0.2356339,
  0.5212163, 0.5035238, 0.3593956, 0.2415617, 0.1394327, 0.07778603, 
    0.08077269, 0.1712121, 0.324949, 0.3744895, 0.4121276, 0.4525426, 
    0.301756, 0.2533889, 0.2328566, 0.1225504, 0.117899, 0.1312325, 0.219566, 
    0.2657067, 0.3407953, 0.3021755, 0.2564465, 0.423649, 0.2681382, 
    0.1307671, 0.1364713, 0.1759282, 0.446309,
  0.3045209, 0.2316549, 0.349901, 0.2501311, 0.2794529, 0.282957, 0.2317178, 
    0.2568131, 0.2567574, 0.2864034, 0.2678388, 0.294014, 0.2677117, 
    0.2560256, 0.2157963, 0.2512748, 0.3009492, 0.250338, 0.2272656, 
    0.2926757, 0.3270234, 0.2699597, 0.2255544, 0.2369868, 0.1613214, 
    0.2411608, 0.2405629, 0.2930369, 0.3258691,
  0.2514958, 0.233913, 0.2569652, 0.2273885, 0.2206826, 0.2018813, 0.1891525, 
    0.2778521, 0.2723487, 0.2866369, 0.2756749, 0.2709584, 0.269811, 
    0.2091077, 0.15827, 0.1929576, 0.2216004, 0.1976827, 0.2370601, 
    0.1914773, 0.2246531, 0.2483747, 0.2253181, 0.2171089, 0.1002497, 
    0.1333962, 0.2371035, 0.2932445, 0.2781147,
  0.2371562, 0.1651672, 0.1451832, 0.1518161, 0.1304159, 0.1722635, 
    0.1758248, 0.1968407, 0.1792805, 0.167654, 0.1514708, 0.1731531, 
    0.1408325, 0.1806371, 0.2046765, 0.1967021, 0.2353017, 0.2125869, 
    0.2217402, 0.1834588, 0.2173578, 0.1864673, 0.1258215, 0.08278993, 
    0.07684651, 0.1277854, 0.1847097, 0.2179585, 0.2401729,
  0.05373195, 0.02986632, 0.04137202, 0.05316193, 0.0586531, 0.05290724, 
    0.06852604, 0.06483153, 0.1017145, 0.05158572, 0.01557344, 0.009387049, 
    0.00248773, 0.07936369, 0.08815102, 0.1187279, 0.1233454, 0.07130224, 
    0.1285168, 0.1319715, 0.09505384, 0.09144413, 0.03466509, 0.002280553, 
    0.0437722, 0.09010236, 0.1103215, 0.1245676, 0.08597891,
  0.001657141, -8.314601e-08, 0.0293898, 0.03761641, 0.05965536, 0.03566553, 
    0.04008355, 0.01589134, 0.08003534, 0.02908677, 1.001288e-07, 
    -2.397135e-05, 0.01315969, 0.01186335, 0.09325226, 0.1072145, 0.02398029, 
    0.03487443, 0.03868166, 0.02722135, 0.03635297, 0.01364345, 
    -3.119767e-05, 8.529612e-08, 0.006086224, 0.02732597, 0.1070949, 
    0.04953681, 0.02071233,
  5.538102e-08, -2.003549e-08, -3.879249e-06, 0.2328577, 0.03404751, 
    0.04578409, 0.01465029, 0.04574164, 0.04899948, 0.01461405, 0.04893259, 
    0.06562459, 0.2409544, 0.07567281, 0.03663534, 0.02237075, 0.02257527, 
    0.02781106, 0.01528642, 0.008428785, 0.001669117, -2.671141e-07, 
    7.479406e-09, 0.01137275, 0.01717682, 0.0007394752, 0.05438546, 
    0.009845537, 3.810336e-06,
  0.0001029285, 0.01235045, 0.074317, 0.02272065, 0.01571777, 0.006539719, 
    0.01227959, 0.01635787, 0.02603886, 0.03497402, 0.0232665, 0.01539061, 
    0.06352235, 0.04883973, 0.04932121, 0.0489543, 0.02604696, 0.01333492, 
    0.007297355, 0.0005814339, 0.0009587735, 0.0006825824, 0.009069324, 
    0.180427, 0.1259188, 0.01429156, 0.01905773, 0.001253714, 2.552992e-05,
  0.03597644, 0.02957065, 0.04607359, 0.301006, 0.006017389, 0.01091614, 
    0.1146896, 0.0261278, 0.008337151, 0.02589923, 0.008507113, 0.04534638, 
    0.0750792, 0.06185851, 0.08174057, 0.1234282, 0.1296445, 0.1962319, 
    0.1724267, 0.1354147, 0.2152976, 0.1217295, 0.1503603, 0.07234347, 
    0.02027309, 0.0771571, 0.1528523, 0.1277474, 0.1244848,
  5.985353e-07, 5.719504e-10, 7.843643e-10, 3.251434e-08, 4.64168e-07, 
    0.002235201, 0.3690267, 0.3117213, 0.4085166, 0.1156673, 0.1631596, 
    0.09993932, 0.04556739, 0.02149309, 0.02035565, 0.02879049, 0.01318343, 
    0.00632512, 0.01930677, -5.243107e-06, 0.01808808, 0.04104895, 
    0.01129889, 0.01798686, 0.0341468, 0.03393012, 0.0009355597, 
    4.915796e-06, 2.376209e-08,
  7.541169e-07, 4.044463e-06, -1.289763e-06, 1.220956e-10, 4.270413e-07, 
    6.539518e-06, 0.04010815, 0.1752363, 0.3296965, 0.1058762, 0.05271721, 
    0.05242449, 0.1009114, 0.04472899, 0.07618421, 0.0343519, 0.03237598, 
    0.01210602, 0.0002196693, 6.54661e-08, 0.001500868, 0.006162699, 
    0.0816433, 0.0229811, 0.016607, 0.03527187, 0.003520614, 0.001863951, 
    1.675933e-06,
  0.01715211, 0.0173664, 0.01527965, 0.04013744, -6.968416e-05, 2.883879e-09, 
    0.0002000429, 3.50298e-06, 0.0001418592, 0.05440011, 0.1146195, 
    0.08659291, 0.243922, 0.159914, 0.06708512, 0.0944506, 0.1276003, 
    0.07715891, 0.02851675, 7.513824e-05, 0.0003676275, 0.002234417, 
    0.0243954, 0.05927737, 0.04890293, 0.07159115, 0.04569035, 0.004299174, 
    0.003464758,
  0.05048059, 0.1511988, 0.07250857, 0.156954, 0.0244477, 0.03223224, 
    0.1064404, 0.2256859, 0.1306524, 0.01452119, 0.06080357, 0.2295691, 
    0.08521065, 0.1670518, 0.1900579, 0.2521881, 0.2669797, 0.2353576, 
    0.2155372, 0.05352264, 0.01732422, 0.02088647, 0.07894623, 0.1819081, 
    0.1642663, 0.1571102, 0.1381832, 0.1338705, 0.04502675,
  0.05802276, 0.1232813, 0.1319626, 0.1166805, 0.206805, 0.09588575, 
    0.1813671, 0.1328926, 0.1314285, 0.2002461, 0.1076204, 0.2648632, 
    0.301993, 0.271618, 0.1608862, 0.2941616, 0.219123, 0.4207198, 0.3830958, 
    0.1290609, 0.1656824, 0.158069, 0.1751141, 0.2753312, 0.1718748, 
    0.2014515, 0.213318, 0.2174421, 0.1714594,
  0.2642754, 0.2531, 0.4168542, 0.2305018, 0.1830679, 0.2192239, 0.1759485, 
    0.09737396, 0.2326396, 0.1666901, 0.1421006, 0.2234303, 0.2197411, 
    0.3656517, 0.4006101, 0.1675477, 0.2652988, 0.1474114, 0.134939, 
    0.1480255, 0.1782556, 0.3134344, 0.2734519, 0.3838579, 0.2327161, 
    0.3780854, 0.2571353, 0.2322968, 0.3155882,
  0.1654459, 0.1932764, 0.2683648, 0.1926354, 0.165735, 0.2539687, 0.4066486, 
    0.4426842, 0.3489651, 0.201898, 0.1805777, 0.2172844, 0.2708086, 
    0.1977925, 0.1897122, 0.191842, 0.2128689, 0.3341396, 0.221699, 
    0.1167556, 0.09246305, 0.1669998, 0.1887849, 0.1118564, 0.1501374, 
    0.1302651, 0.1538237, 0.2264196, 0.2200213,
  0.3800527, 0.377435, 0.3748172, 0.3721994, 0.3695817, 0.366964, 0.3643462, 
    0.390067, 0.3864025, 0.3827381, 0.3790736, 0.3754091, 0.3717446, 
    0.3680802, 0.3495966, 0.3583671, 0.3671375, 0.375908, 0.3846784, 
    0.3934488, 0.4022192, 0.3781036, 0.3756153, 0.3731271, 0.3706389, 
    0.3681507, 0.3656625, 0.3631743, 0.3821469,
  0.1548824, 0.1613692, 0.1496453, 0.08457264, 0.08760451, 0.1143617, 
    0.177661, 0.15209, 0.06059615, 0.06522011, 0.04840487, 0.02290847, 
    0.03548265, 0.02848264, 0.0370223, 0.0524875, 0.06698272, 0.09769896, 
    0.1379959, 0.1220616, 0.2955105, 0.5607806, 0.4280182, 0.2912837, 
    0.1795377, 0.157326, 0.2699974, 0.2417366, 0.2346026,
  0.566232, 0.5148947, 0.4004277, 0.2443478, 0.1462655, 0.08751066, 
    0.08120905, 0.1901682, 0.3389916, 0.4106745, 0.422149, 0.457308, 
    0.2905559, 0.2756881, 0.2264886, 0.1396924, 0.1131011, 0.1547805, 
    0.2166589, 0.2837351, 0.3791154, 0.3251709, 0.2331039, 0.4160253, 
    0.2424114, 0.1435723, 0.1156604, 0.215433, 0.4260848,
  0.3308083, 0.2741126, 0.4044685, 0.3073878, 0.2883156, 0.3086101, 
    0.3043357, 0.2041605, 0.2601303, 0.3141633, 0.3166028, 0.2840038, 
    0.2819599, 0.3119029, 0.2659388, 0.327882, 0.3037472, 0.2742982, 
    0.2786508, 0.2960972, 0.3047737, 0.2846234, 0.2253734, 0.2685409, 
    0.1913928, 0.2795688, 0.2576736, 0.2775273, 0.3254278,
  0.2633538, 0.2924571, 0.3284214, 0.2606772, 0.2356047, 0.2465239, 
    0.2506739, 0.287063, 0.2959754, 0.3013392, 0.2848379, 0.2820098, 
    0.2842794, 0.2405843, 0.1643919, 0.1823236, 0.2841488, 0.2382964, 
    0.3200125, 0.3032432, 0.2578369, 0.2829214, 0.2933109, 0.2457252, 
    0.1134912, 0.1703347, 0.325922, 0.3174732, 0.298159,
  0.2618821, 0.203736, 0.1590871, 0.1598958, 0.1436867, 0.1875702, 0.2001619, 
    0.2342384, 0.1948756, 0.1811384, 0.1583526, 0.1726958, 0.1398141, 
    0.1898038, 0.2321923, 0.1894461, 0.2505385, 0.2394785, 0.2361911, 
    0.2114473, 0.2465552, 0.2186902, 0.1445638, 0.1040511, 0.0887541, 
    0.1654251, 0.1959744, 0.2717044, 0.2502875,
  0.09509423, 0.03950943, 0.05419122, 0.1211538, 0.08524776, 0.07013451, 
    0.08733846, 0.08568615, 0.1165614, 0.09423848, 0.007152982, 0.004643521, 
    0.0009772702, 0.09769681, 0.1198484, 0.1254603, 0.128132, 0.1246823, 
    0.1369421, 0.1645758, 0.1203897, 0.1128603, 0.0685015, 0.001914971, 
    0.02946489, 0.12807, 0.1364429, 0.1379783, 0.1218932,
  0.02086104, -3.911035e-07, 0.009854835, 0.07312171, 0.05884545, 0.06555159, 
    0.09275528, 0.08187705, 0.1480149, 0.0228708, 5.143674e-09, 
    -2.416555e-06, 0.02616978, 0.03931568, 0.1061725, 0.1009205, 0.02252296, 
    0.03766081, 0.03598624, 0.0642594, 0.1242278, 0.1101535, 0.007234973, 
    9.073633e-08, 0.004547757, 0.06023469, 0.1217951, 0.2043684, 0.07276952,
  6.094203e-07, 3.674544e-07, -1.728978e-05, 0.1582179, 0.02107788, 
    0.03910922, 0.04196094, 0.05310474, 0.047989, 0.02234463, 0.06586961, 
    0.07964924, 0.2881429, 0.06440537, 0.03346634, 0.02167654, 0.01901301, 
    0.01914385, 0.02000862, 0.01032301, 0.002555107, 6.949993e-06, 
    3.348066e-09, 0.0128214, 0.001421856, 9.742144e-06, 0.05269827, 
    0.02854596, 0.002108179,
  3.887586e-05, 0.02604479, 0.04578539, 0.007929928, 0.02101141, 0.01036536, 
    0.01376093, 0.01736913, 0.02801052, 0.04892399, 0.02777249, 0.0136652, 
    0.05009101, 0.04301485, 0.04391031, 0.03458083, 0.02340175, 0.02056163, 
    0.009871156, 0.004170533, 0.002908037, 0.001284278, 0.005839472, 
    0.1682843, 0.1382358, 0.01102998, 0.02044473, 0.008033514, 0.001206426,
  0.03660142, 0.03115927, 0.04165577, 0.2449216, 0.001006233, 0.01244278, 
    0.08965637, 0.0248504, 0.008266172, 0.01889718, 0.007927658, 0.03767263, 
    0.05656533, 0.05021727, 0.07526056, 0.1158708, 0.1275494, 0.19547, 
    0.1377715, 0.1134244, 0.206154, 0.11177, 0.1474991, 0.08134274, 
    0.01889978, 0.06950489, 0.148505, 0.1293212, 0.1201323,
  3.906244e-07, 3.939612e-10, 4.672713e-10, 1.043511e-08, 3.459306e-07, 
    0.005723031, 0.364729, 0.2907824, 0.3826881, 0.1015562, 0.1278197, 
    0.08522904, 0.03777052, 0.02126983, 0.02443235, 0.0414086, 0.02481967, 
    0.02192271, 0.02073158, -1.315005e-05, 0.02097191, 0.04704963, 
    0.01096697, 0.01816668, 0.0372317, 0.04369661, 0.0101451, 2.671351e-06, 
    2.500401e-07,
  3.866521e-07, 3.055446e-06, 4.722009e-10, 5.282953e-10, 3.092954e-07, 
    -1.713134e-06, 0.03040327, 0.1534699, 0.2926041, 0.1106967, 0.05432497, 
    0.05626314, 0.09070084, 0.03377874, 0.05936771, 0.03259614, 0.04150837, 
    0.05192717, 0.003078383, 7.332293e-08, 0.000679596, 0.006554276, 
    0.07128345, 0.02206284, 0.02119217, 0.04598108, 0.03152468, 0.006722864, 
    1.301835e-06,
  0.0100622, 0.01764127, 0.00514084, 0.05535626, -6.449646e-05, 2.446394e-10, 
    1.003895e-05, 2.427596e-06, -3.924327e-05, 0.05761281, 0.1793483, 
    0.08517993, 0.2573541, 0.1756629, 0.06175797, 0.122862, 0.1582387, 
    0.1314868, 0.04435207, -1.217266e-05, 0.0001410797, 0.001676, 0.02351799, 
    0.06301126, 0.04821366, 0.08395623, 0.06655719, 0.01211735, 0.0007490873,
  0.1092759, 0.1971658, 0.07515636, 0.143464, 0.007026942, 0.02202729, 
    0.06431308, 0.2490516, 0.1143015, 0.009063011, 0.05973035, 0.2392514, 
    0.1055109, 0.175878, 0.2032818, 0.269193, 0.2730905, 0.243713, 0.2637341, 
    0.04748729, 0.01279713, 0.01724531, 0.06935512, 0.1735208, 0.1487879, 
    0.1438646, 0.1781362, 0.1501259, 0.08938888,
  0.07720102, 0.1409673, 0.1560348, 0.1783637, 0.222227, 0.1042973, 0.193735, 
    0.1463588, 0.1433177, 0.1902687, 0.1052755, 0.2686219, 0.3371267, 
    0.2811952, 0.1583065, 0.3197022, 0.2502712, 0.4115867, 0.395194, 
    0.1343194, 0.1110707, 0.1693712, 0.157787, 0.3099042, 0.1669535, 
    0.2194148, 0.2457535, 0.2339983, 0.1859852,
  0.2808079, 0.2721575, 0.4243201, 0.2569589, 0.2607942, 0.3181231, 
    0.2207681, 0.1116846, 0.1835937, 0.1577799, 0.1601163, 0.2372455, 
    0.2985204, 0.3846693, 0.4155904, 0.1581686, 0.2578287, 0.1748387, 
    0.1524564, 0.1427738, 0.2166066, 0.3704014, 0.3760447, 0.3983443, 
    0.220439, 0.3921001, 0.2729436, 0.2411948, 0.3275988,
  0.1970226, 0.2842891, 0.32264, 0.1696122, 0.1661003, 0.2557706, 0.4062746, 
    0.4137938, 0.4050953, 0.2256212, 0.2640317, 0.2876951, 0.2898021, 
    0.2147173, 0.176178, 0.2234202, 0.2623319, 0.3892703, 0.2515785, 
    0.1608506, 0.1628832, 0.1841321, 0.209064, 0.1282585, 0.1350714, 
    0.1840595, 0.1370948, 0.2700732, 0.2869329,
  0.4115606, 0.4109752, 0.4103899, 0.4098045, 0.4092192, 0.4086339, 
    0.4080485, 0.4346605, 0.4290607, 0.423461, 0.4178612, 0.4122614, 
    0.4066617, 0.4010619, 0.4080335, 0.4173872, 0.4267409, 0.4360946, 
    0.4454483, 0.454802, 0.4641557, 0.4297926, 0.4266241, 0.4234554, 
    0.4202869, 0.4171183, 0.4139497, 0.4107811, 0.4120288,
  0.1654784, 0.1634051, 0.1692608, 0.1154973, 0.1096254, 0.164056, 0.2140146, 
    0.1790332, 0.06191596, 0.07317775, 0.06399082, 0.02653444, 0.04275079, 
    0.02760895, 0.03852824, 0.04120924, 0.06849363, 0.08700077, 0.1284237, 
    0.1344077, 0.3563176, 0.5668674, 0.4744848, 0.2945427, 0.2091114, 
    0.2007136, 0.2425236, 0.2276258, 0.2450833,
  0.5947822, 0.4854546, 0.4166095, 0.216889, 0.154872, 0.08482692, 
    0.08344254, 0.2150855, 0.3619866, 0.4309402, 0.4434986, 0.4552067, 
    0.2662404, 0.2891268, 0.235515, 0.1474943, 0.1266844, 0.1929945, 
    0.2952568, 0.2859932, 0.3493247, 0.284804, 0.2391577, 0.4540417, 
    0.227969, 0.1423124, 0.1133326, 0.2680214, 0.4367922,
  0.4003985, 0.3480289, 0.4674751, 0.3407776, 0.3693264, 0.4420871, 
    0.3255621, 0.2358695, 0.2813828, 0.349048, 0.3824039, 0.279791, 0.309084, 
    0.3319177, 0.3588105, 0.3506111, 0.3519554, 0.4108124, 0.4010079, 
    0.3399578, 0.2941897, 0.2375828, 0.2258706, 0.315755, 0.301372, 
    0.3662771, 0.2872024, 0.3176405, 0.3316086,
  0.3461192, 0.3610771, 0.3599479, 0.3076137, 0.2631666, 0.2507662, 
    0.2934355, 0.3274331, 0.2792782, 0.2621795, 0.2546788, 0.2618477, 
    0.2843186, 0.2628838, 0.2306244, 0.2094124, 0.3098339, 0.278973, 
    0.3055871, 0.3516207, 0.2772895, 0.3647128, 0.341633, 0.2479884, 
    0.1189222, 0.2617149, 0.4112729, 0.3587809, 0.3167843,
  0.3076019, 0.2049766, 0.1825352, 0.1794283, 0.2244134, 0.2076994, 
    0.1933376, 0.2225038, 0.1833586, 0.1684071, 0.1555178, 0.1514341, 
    0.1251903, 0.1786223, 0.2847391, 0.1836891, 0.2423442, 0.2737859, 
    0.2488525, 0.2412399, 0.2472438, 0.2724135, 0.1703747, 0.130795, 
    0.1138597, 0.1914571, 0.2427086, 0.2694894, 0.2514273,
  0.150207, 0.07640245, 0.04981263, 0.1465148, 0.1496208, 0.1633123, 
    0.1478768, 0.2293316, 0.1958617, 0.136046, 0.0007544381, 0.0002934271, 
    0.0006036076, 0.1023538, 0.09610333, 0.1201078, 0.1006996, 0.09725092, 
    0.1367272, 0.1531035, 0.1689643, 0.1785547, 0.1139221, 0.001497333, 
    0.04718078, 0.1002777, 0.1098193, 0.1930108, 0.2115428,
  0.1656363, -2.7623e-06, 0.001485541, 0.1346037, 0.07685819, 0.08111931, 
    0.1154288, 0.1686515, 0.2865485, 0.05027104, 2.558035e-09, -1.033827e-07, 
    0.1159294, 0.1638423, 0.1256646, 0.1085579, 0.03275977, 0.0432764, 
    0.03920467, 0.07317695, 0.1620897, 0.2278921, 0.1349016, 1.34593e-07, 
    0.006885813, 0.04808723, 0.1011483, 0.3252634, 0.4519317,
  0.0001700947, 5.804145e-06, -0.0001700073, 0.0377951, 0.0239363, 
    0.03629715, 0.05955491, 0.0610376, 0.0524688, 0.02783359, 0.08727518, 
    0.08389249, 0.3123775, 0.05718749, 0.03218196, 0.02495561, 0.02017511, 
    0.018265, 0.02200495, 0.02695038, 0.01675214, 0.004059118, 3.638501e-07, 
    0.01562976, 0.0001713698, -1.854016e-06, 0.07039291, 0.03403917, 0.0329051,
  0.003838011, 0.08302879, 0.02828957, 0.006394078, 0.0253431, 0.01990623, 
    0.02457964, 0.0207138, 0.03051353, 0.0612733, 0.0285191, 0.01516053, 
    0.04343272, 0.03988555, 0.03777048, 0.02608059, 0.01787577, 0.02006348, 
    0.01787917, 0.009501779, 0.01137601, 0.000239469, 0.00242713, 0.179801, 
    0.1503441, 0.01038679, 0.02575574, 0.0175666, 0.01116608,
  0.04382998, 0.03795469, 0.03219978, 0.2206696, -0.0004430183, 0.0129283, 
    0.07354469, 0.0252548, 0.00791625, 0.01772269, 0.007292614, 0.03190652, 
    0.0449679, 0.04547553, 0.0659282, 0.1037911, 0.1191519, 0.1813743, 
    0.115434, 0.1007935, 0.1784105, 0.09410384, 0.1340883, 0.0768297, 
    0.01971281, 0.06674521, 0.1318644, 0.1342667, 0.1186834,
  2.803612e-07, 1.834091e-10, 3.050274e-10, 5.685973e-09, 2.128223e-07, 
    0.0249347, 0.3478626, 0.2527398, 0.352503, 0.08096375, 0.09985001, 
    0.06737965, 0.04089415, 0.02606298, 0.03074628, 0.0494226, 0.06104566, 
    0.03959696, 0.02271389, 5.942755e-05, 0.01949638, 0.05255375, 0.01376402, 
    0.02060952, 0.04689411, 0.068331, 0.05190685, 2.528783e-06, 2.355479e-07,
  2.411787e-07, 2.482095e-06, 7.529223e-09, 4.187853e-10, 2.401572e-07, 
    -1.71545e-06, 0.02045849, 0.1482661, 0.3065953, 0.09737671, 0.05320406, 
    0.06947501, 0.07626475, 0.03145571, 0.05537131, 0.03840333, 0.05066568, 
    0.07702126, 0.00663532, 1.436499e-07, 0.0002135902, 0.007530245, 
    0.06012698, 0.02247235, 0.03188643, 0.05518319, 0.09208895, 0.01543456, 
    1.201263e-06,
  0.003061653, 0.01388687, 0.003064215, 0.0729993, 9.985684e-05, 
    1.609225e-10, 4.878771e-07, 2.393412e-06, -4.80105e-05, 0.043888, 
    0.2218095, 0.07713784, 0.2497305, 0.1840008, 0.06619015, 0.1363292, 
    0.2277933, 0.185223, 0.1203395, -9.948391e-06, -5.639188e-05, 
    0.001186331, 0.02541547, 0.05694189, 0.06008833, 0.1091795, 0.1079597, 
    0.02688778, 0.004966705,
  0.1390122, 0.2040391, 0.07052691, 0.1273691, 0.001961637, 0.0111272, 
    0.04232142, 0.2426779, 0.09308802, 0.008072671, 0.04849982, 0.2549992, 
    0.1182628, 0.2389549, 0.209296, 0.2876523, 0.2974178, 0.2344441, 
    0.2741777, 0.03777593, 0.00506928, 0.01583329, 0.06714214, 0.1895544, 
    0.1708323, 0.141383, 0.250475, 0.1719289, 0.1061453,
  0.1155743, 0.133988, 0.08769143, 0.1511798, 0.1761769, 0.1354045, 
    0.2318487, 0.1583007, 0.1658474, 0.1772679, 0.1801707, 0.2965789, 
    0.3759921, 0.2905644, 0.2027922, 0.3125341, 0.3001029, 0.3982199, 
    0.3935731, 0.1197357, 0.07260977, 0.1473556, 0.1594885, 0.3049614, 
    0.1596884, 0.2310795, 0.3037051, 0.2767126, 0.1813295,
  0.3216685, 0.3496852, 0.441123, 0.2776057, 0.3049515, 0.3636532, 0.2316251, 
    0.1668235, 0.2404881, 0.1858142, 0.2269264, 0.2833925, 0.3235425, 
    0.3801129, 0.3770826, 0.1641772, 0.2856793, 0.1638755, 0.1483321, 
    0.1603193, 0.4287504, 0.4211519, 0.4620505, 0.4760342, 0.2130688, 
    0.3914858, 0.3087103, 0.2497787, 0.3405862,
  0.3886762, 0.4379748, 0.4041964, 0.2421265, 0.2034399, 0.355791, 0.5342992, 
    0.4798355, 0.4279902, 0.2950676, 0.3219521, 0.3285092, 0.2956803, 
    0.2184703, 0.1965994, 0.2190775, 0.3444676, 0.4122322, 0.2695881, 
    0.2313265, 0.2189631, 0.2449138, 0.2777937, 0.1518654, 0.1454845, 
    0.2168199, 0.1534622, 0.2823373, 0.3815597,
  0.4590726, 0.4590345, 0.4589964, 0.4589583, 0.4589202, 0.4588821, 
    0.4588439, 0.4722054, 0.4665974, 0.4609895, 0.4553815, 0.4497736, 
    0.4441657, 0.4385577, 0.4613092, 0.4703952, 0.4794812, 0.4885672, 
    0.4976532, 0.5067392, 0.5158252, 0.4655696, 0.4621297, 0.4586897, 
    0.4552497, 0.4518098, 0.4483698, 0.4449298, 0.4591031,
  0.1793326, 0.1650474, 0.1715545, 0.1392134, 0.1074049, 0.1834987, 
    0.2266273, 0.1902586, 0.06706682, 0.0702081, 0.06874046, 0.03063908, 
    0.05126024, 0.02212904, 0.03978762, 0.03563727, 0.06668389, 0.07616467, 
    0.125525, 0.1517708, 0.3902988, 0.542482, 0.4891895, 0.3025157, 
    0.2462326, 0.2356068, 0.235899, 0.2048863, 0.2414315,
  0.5804593, 0.4493321, 0.4320178, 0.178799, 0.1463487, 0.08980293, 
    0.05719498, 0.247412, 0.3890055, 0.4539008, 0.4516488, 0.4497268, 
    0.2314386, 0.2968342, 0.2624217, 0.1700487, 0.138411, 0.2403911, 
    0.3162031, 0.3098326, 0.3582908, 0.2695005, 0.2408517, 0.4702717, 
    0.230627, 0.1489418, 0.1795886, 0.244248, 0.4366402,
  0.4251462, 0.4518175, 0.4422669, 0.3209437, 0.4153073, 0.5147516, 
    0.3216658, 0.283728, 0.3317266, 0.364278, 0.4286606, 0.3100985, 
    0.3393435, 0.3460513, 0.3504995, 0.328878, 0.4293961, 0.374168, 
    0.3460635, 0.2693655, 0.2345019, 0.1968907, 0.2267378, 0.2779665, 
    0.3446717, 0.3655447, 0.2861519, 0.3477829, 0.378311,
  0.3378104, 0.3650085, 0.3710038, 0.3567841, 0.2912815, 0.2693534, 
    0.2931706, 0.2439621, 0.2254392, 0.2316657, 0.2390559, 0.2503985, 
    0.2889176, 0.2493361, 0.2756007, 0.2329821, 0.2627479, 0.285511, 
    0.3142873, 0.3383441, 0.2557177, 0.2898194, 0.3062687, 0.2559471, 
    0.1404802, 0.2942767, 0.4040808, 0.3548495, 0.3264052,
  0.3004868, 0.2155129, 0.1598275, 0.1967006, 0.2572449, 0.1949598, 
    0.2141478, 0.211395, 0.1650434, 0.1904259, 0.1418643, 0.1087309, 
    0.09420812, 0.1313938, 0.3553113, 0.1925251, 0.2353602, 0.2259232, 
    0.2272782, 0.1909979, 0.2148337, 0.2430524, 0.2140033, 0.1564246, 
    0.1110744, 0.1774871, 0.1611279, 0.2060262, 0.2207279,
  0.1818115, 0.07349476, 0.04867544, 0.1136163, 0.1383207, 0.1640332, 
    0.2052623, 0.2440908, 0.2535735, 0.09038907, 5.381481e-05, -1.594535e-06, 
    0.0001823818, 0.03678822, 0.06256515, 0.116248, 0.09227678, 0.09839493, 
    0.1135525, 0.1279448, 0.1448864, 0.182848, 0.2010859, 0.003381463, 
    0.02998627, 0.06759685, 0.07439347, 0.1194744, 0.1876414,
  0.346688, -0.0004502993, 0.0001314466, 0.164815, 0.06438896, 0.06045974, 
    0.120658, 0.1329305, 0.2897331, 0.01936293, 1.750656e-09, 9.657069e-09, 
    0.1042074, 0.1439673, 0.1346108, 0.1403488, 0.06051934, 0.05468409, 
    0.07027277, 0.1113838, 0.1693819, 0.3699039, 0.3032727, -1.368368e-07, 
    0.004301465, 0.0425052, 0.0702019, 0.1939926, 0.4506766,
  0.02094815, 8.372337e-05, -0.0001357999, 0.02264612, 0.04552276, 
    0.05327195, 0.05252624, 0.05475255, 0.07230959, 0.04669321, 0.1284477, 
    0.1382508, 0.2795999, 0.05452678, 0.04755805, 0.0414852, 0.03553194, 
    0.04455435, 0.06462863, 0.09445346, 0.127447, 0.05923451, 3.471988e-06, 
    0.01841467, 3.13656e-05, -3.379634e-07, 0.09200203, 0.064184, 0.1618613,
  0.04367311, 0.1657441, 0.02167086, 0.004148404, 0.0403873, 0.1074497, 
    0.08708499, 0.03388428, 0.02266829, 0.05850593, 0.03476461, 0.01867761, 
    0.03984167, 0.04868081, 0.03548, 0.02309416, 0.01539729, 0.01444086, 
    0.01594299, 0.01295068, 0.0216231, 0.002406091, 0.0006727564, 0.217598, 
    0.115477, 0.01410967, 0.05612638, 0.04189987, 0.05724899,
  0.05521909, 0.04333945, 0.02402891, 0.2190976, -0.0004650034, 0.0105408, 
    0.06342651, 0.02967058, 0.006571879, 0.01857962, 0.005354041, 0.03363502, 
    0.04003794, 0.03778505, 0.06053923, 0.09273479, 0.1020995, 0.1663654, 
    0.1032939, 0.09619743, 0.1492921, 0.08150006, 0.1278189, 0.06238338, 
    0.02539231, 0.06670506, 0.116724, 0.1291893, 0.1064734,
  2.109563e-07, 1.663353e-10, 2.200486e-10, 2.775432e-09, 1.343758e-07, 
    0.04005906, 0.2718025, 0.213593, 0.3245111, 0.06178814, 0.09441812, 
    0.05855858, 0.0485796, 0.0371513, 0.03763299, 0.06095111, 0.1151495, 
    0.1112472, 0.03970629, 0.0006869527, 0.008266519, 0.05534329, 0.02337705, 
    0.02270021, 0.05332794, 0.0851974, 0.1061834, 1.724634e-05, 1.778412e-07,
  1.830537e-07, 2.108737e-06, -1.675788e-07, 3.473468e-11, 1.982231e-07, 
    -9.185405e-07, 0.01046412, 0.1661586, 0.3154364, 0.08240382, 0.05296834, 
    0.08633979, 0.06821129, 0.03336216, 0.06555285, 0.04630392, 0.08819612, 
    0.1398833, 0.07348157, 1.267256e-07, 6.881056e-05, 0.006612807, 
    0.04914207, 0.02748386, 0.03748351, 0.07833225, 0.1603737, 0.05662455, 
    -6.761288e-06,
  0.0008538844, 0.008160323, 0.0009725721, 0.1168947, -6.954226e-05, 
    2.809003e-11, 6.92025e-06, 2.233673e-06, -3.862287e-05, 0.03678623, 
    0.236947, 0.07654949, 0.2675047, 0.2032091, 0.1556171, 0.2155878, 
    0.3416018, 0.2811219, 0.1775092, -1.999183e-06, -0.0003102481, 
    0.0006392756, 0.01751821, 0.05241658, 0.0594984, 0.1945843, 0.2065963, 
    0.07822527, 0.009538637,
  0.1144776, 0.1792744, 0.05720705, 0.1080113, 0.0001305997, 0.006955252, 
    0.03025695, 0.2222313, 0.07118251, 0.004518882, 0.03356254, 0.2446255, 
    0.1551308, 0.2870285, 0.2574916, 0.3683084, 0.3456712, 0.3837442, 
    0.3286495, 0.02955441, 0.001035781, 0.01085337, 0.07300584, 0.1943218, 
    0.1512167, 0.1380673, 0.3737141, 0.2769575, 0.1214559,
  0.1591004, 0.08878966, 0.07526362, 0.1293415, 0.1533961, 0.1002902, 
    0.2055725, 0.1544004, 0.1763279, 0.1511752, 0.1172121, 0.2925345, 
    0.3859378, 0.300225, 0.2048921, 0.3174272, 0.3236472, 0.3838176, 
    0.3560849, 0.06105333, 0.04522407, 0.1263859, 0.1383492, 0.3203634, 
    0.1470593, 0.2443287, 0.3176273, 0.3390265, 0.2406202,
  0.4381697, 0.449619, 0.4470052, 0.3337723, 0.3085316, 0.3219521, 0.2184283, 
    0.2453927, 0.2735847, 0.2625848, 0.2404322, 0.4198308, 0.3477145, 
    0.3968909, 0.3611198, 0.1756594, 0.319681, 0.1443399, 0.1419342, 
    0.1924764, 0.489639, 0.4246067, 0.5436376, 0.5039298, 0.2076222, 
    0.4066684, 0.3075362, 0.2393621, 0.3797896,
  0.4524936, 0.4898471, 0.4292863, 0.3665286, 0.3425702, 0.4908524, 
    0.6022769, 0.5536057, 0.4399625, 0.3657796, 0.3630459, 0.4244512, 
    0.3328923, 0.278955, 0.2531728, 0.2832864, 0.3927805, 0.3852558, 
    0.2616633, 0.2433599, 0.2795731, 0.2489794, 0.3350773, 0.236825, 
    0.1607946, 0.3213769, 0.181072, 0.3646951, 0.4489101,
  0.4964442, 0.497359, 0.4982738, 0.4991887, 0.5001035, 0.5010183, 0.5019331, 
    0.5019032, 0.4954969, 0.4890907, 0.4826843, 0.476278, 0.4698717, 
    0.4634654, 0.5085719, 0.5174382, 0.5263045, 0.5351709, 0.5440372, 
    0.5529035, 0.5617698, 0.5069106, 0.5035357, 0.5001609, 0.496786, 
    0.4934112, 0.4900363, 0.4866615, 0.4957123,
  0.1812605, 0.1707458, 0.1701986, 0.1564195, 0.1180832, 0.1972276, 
    0.2402415, 0.2056525, 0.07318781, 0.06525917, 0.08566636, 0.03513468, 
    0.0540992, 0.01315624, 0.02013427, 0.04668522, 0.0621812, 0.05632624, 
    0.127562, 0.1409688, 0.3951787, 0.5236706, 0.5069607, 0.2957096, 
    0.237708, 0.2409528, 0.2064052, 0.1898482, 0.2358328,
  0.541477, 0.4186948, 0.449297, 0.1246723, 0.1306385, 0.105202, 0.0242558, 
    0.3032918, 0.4330108, 0.4586753, 0.4637522, 0.4151065, 0.2087002, 
    0.2887414, 0.2794101, 0.2100466, 0.1486948, 0.2871469, 0.3212054, 
    0.3176594, 0.3791421, 0.257608, 0.2390647, 0.4632376, 0.255449, 
    0.2535251, 0.2195359, 0.269301, 0.4388863,
  0.4496145, 0.4496028, 0.3920155, 0.3530392, 0.3569428, 0.4370988, 0.341343, 
    0.3504968, 0.4456198, 0.3014865, 0.3519961, 0.3129676, 0.3408004, 
    0.3463918, 0.4264548, 0.327059, 0.3888134, 0.3213799, 0.2982729, 
    0.1978602, 0.1873277, 0.2181418, 0.2201281, 0.2485342, 0.3168382, 
    0.4131854, 0.3362022, 0.4025007, 0.4646249,
  0.3302567, 0.3370016, 0.3541585, 0.3809029, 0.3298355, 0.3291374, 
    0.2809227, 0.1807553, 0.1700472, 0.2129692, 0.2244597, 0.2409247, 
    0.2680364, 0.240409, 0.2423509, 0.1713304, 0.1848845, 0.2746876, 
    0.270465, 0.2863064, 0.2510188, 0.2603821, 0.29868, 0.2737257, 0.2246393, 
    0.2239414, 0.3512754, 0.3426326, 0.3323243,
  0.2762094, 0.2081813, 0.1207672, 0.1893865, 0.1997974, 0.1482098, 
    0.1502477, 0.1926158, 0.1831457, 0.1647149, 0.1103063, 0.07721581, 
    0.05815059, 0.07909504, 0.3891111, 0.1790328, 0.1956211, 0.2133522, 
    0.1795252, 0.183741, 0.181204, 0.2577789, 0.2419143, 0.1747269, 
    0.0666288, 0.1652382, 0.1156803, 0.1734301, 0.1870605,
  0.1967304, 0.04173893, 0.04122229, 0.05467142, 0.09792659, 0.1008062, 
    0.1704493, 0.2015504, 0.1537471, 0.04022841, -3.376207e-05, 1.366443e-06, 
    4.795414e-05, 0.01231489, 0.03997758, 0.06113169, 0.09333251, 0.09496825, 
    0.07337288, 0.1060642, 0.09950306, 0.1451387, 0.2374994, 0.0112142, 
    0.02417408, 0.03858512, 0.06073093, 0.06917088, 0.1174745,
  0.2757769, 0.001301232, -5.510289e-05, 0.04673217, 0.04205962, 0.0488814, 
    0.1171725, 0.101936, 0.1727896, 0.01388456, 1.026224e-09, 5.88957e-09, 
    0.02796717, 0.1354483, 0.1301146, 0.1584243, 0.08816896, 0.1046632, 
    0.1337692, 0.08609468, 0.180033, 0.3279709, 0.4604791, -1.555082e-05, 
    0.001563461, 0.08075212, 0.05613675, 0.1366877, 0.2472933,
  0.5388756, 0.002893795, -2.059144e-05, 0.01404135, 0.03471287, 0.04529741, 
    0.08800948, 0.1194052, 0.08417676, 0.08092234, 0.07522999, 0.08139087, 
    0.2091386, 0.07606427, 0.05114783, 0.04047873, 0.02532083, 0.03326632, 
    0.02601763, 0.08780453, 0.2086444, 0.4428118, 0.001032614, 0.01394656, 
    7.403914e-06, -7.156327e-07, 0.04699115, 0.04641208, 0.2646886,
  0.2027737, 0.2127843, 0.007159233, 0.007314834, 0.04398428, 0.05429692, 
    0.1439315, 0.09797178, 0.02167646, 0.04738506, 0.06148674, 0.02424468, 
    0.08594595, 0.04692484, 0.03742317, 0.02828303, 0.01784208, 0.01513077, 
    0.01594238, 0.01100129, 0.03740992, 0.02113993, 0.007312594, 0.1667415, 
    0.06953157, 0.04767467, 0.06508479, 0.09211777, 0.1068462,
  0.07536155, 0.0440866, 0.01129295, 0.2200456, -0.0002299915, 0.01114243, 
    0.05920791, 0.03434256, 0.004881299, 0.01735036, 0.004379713, 0.03460005, 
    0.04352336, 0.04243383, 0.05908405, 0.08972271, 0.1043764, 0.1514697, 
    0.1151111, 0.09675222, 0.1233471, 0.08177599, 0.122917, 0.05068207, 
    0.04758409, 0.08610237, 0.09966794, 0.1321112, 0.08875695,
  1.71539e-07, 1.494863e-10, 1.881009e-10, 1.420236e-09, 8.942257e-08, 
    0.05898186, 0.2705248, 0.1631064, 0.3097333, 0.05079378, 0.08330116, 
    0.05675095, 0.0422507, 0.03969675, 0.04588524, 0.05990126, 0.1123951, 
    0.2151443, 0.1580697, 0.02493651, 0.009397528, 0.07512365, 0.06243068, 
    0.02434443, 0.05111324, 0.08894651, 0.2140775, 0.001573741, 1.466376e-07,
  1.512967e-07, 1.350931e-06, -6.924317e-06, -2.073039e-09, 1.731781e-07, 
    -4.64575e-07, 0.005355488, 0.1783659, 0.3160849, 0.05770702, 0.06257054, 
    0.06943141, 0.06719081, 0.07501285, 0.1058173, 0.06196658, 0.1067103, 
    0.1390738, 0.1953502, 5.875067e-06, 4.317965e-05, 0.006147364, 
    0.03885119, 0.03432183, 0.04541116, 0.103726, 0.2032345, 0.334484, 
    -0.0002204577,
  -5.186467e-05, 0.007027728, 0.0002397783, 0.1687675, -9.385931e-05, 
    1.972392e-11, 7.906915e-06, 1.947402e-06, -2.961118e-05, 0.03667311, 
    0.2383284, 0.07407617, 0.3304066, 0.2598167, 0.2591489, 0.3592387, 
    0.4345167, 0.3524537, 0.2796168, 8.74239e-05, -0.000245391, 0.001535664, 
    0.01593076, 0.07420538, 0.07396302, 0.2448637, 0.2363927, 0.2510948, 
    0.02741557,
  0.1349581, 0.1806558, 0.03207161, 0.09869922, 5.623367e-05, 0.005342302, 
    0.02613413, 0.2230057, 0.06010359, 0.003556254, 0.02876039, 0.2318842, 
    0.2360136, 0.369964, 0.388978, 0.4938194, 0.4482587, 0.4720454, 
    0.4263903, 0.03262212, 0.0003894611, 0.007629022, 0.06173418, 0.1568996, 
    0.1462952, 0.1578279, 0.4057072, 0.4336522, 0.1933775,
  0.1746063, 0.07831182, 0.05261356, 0.1083868, 0.1173566, 0.06021286, 
    0.1543495, 0.13976, 0.1727692, 0.1335496, 0.08179292, 0.269133, 
    0.3837505, 0.302217, 0.2296089, 0.3808943, 0.2997707, 0.3705537, 
    0.3291765, 0.04226621, 0.0299671, 0.09394323, 0.1295936, 0.3009101, 
    0.1607427, 0.2585769, 0.3414882, 0.4117139, 0.2889209,
  0.4688095, 0.5244871, 0.4278736, 0.3583362, 0.343864, 0.3638406, 0.2397454, 
    0.2028819, 0.2446963, 0.2254598, 0.2845547, 0.4439852, 0.4051208, 
    0.3952662, 0.3939224, 0.2553476, 0.3817885, 0.1667166, 0.1721017, 
    0.2604239, 0.4596839, 0.5638077, 0.4656525, 0.527551, 0.2452145, 
    0.4149444, 0.3280486, 0.2377481, 0.3977704,
  0.4135458, 0.4218167, 0.5152508, 0.4347166, 0.5671725, 0.6922894, 
    0.6276155, 0.5905841, 0.5507405, 0.4478893, 0.4585131, 0.569976, 
    0.4501019, 0.4584276, 0.381108, 0.3445961, 0.3250748, 0.387912, 
    0.3371882, 0.3829121, 0.4497441, 0.2573511, 0.3435049, 0.3273624, 
    0.2109745, 0.2346913, 0.2591669, 0.4508516, 0.4391621,
  0.5531421, 0.5556651, 0.5581881, 0.560711, 0.563234, 0.565757, 0.56828, 
    0.5721695, 0.5655715, 0.5589734, 0.5523753, 0.5457773, 0.5391791, 
    0.5325811, 0.552763, 0.5599717, 0.5671805, 0.5743892, 0.581598, 
    0.5888067, 0.5960155, 0.5334653, 0.5303317, 0.5271981, 0.5240644, 
    0.5209308, 0.5177972, 0.5146635, 0.5511238,
  0.1793602, 0.1831701, 0.1883988, 0.1891377, 0.1619752, 0.2122969, 
    0.2509711, 0.2033872, 0.06895217, 0.07755145, 0.1047394, 0.06579016, 
    0.0606335, 0.00791894, 0.01632708, 0.07048429, 0.05993231, 0.05349089, 
    0.1203648, 0.109966, 0.3679912, 0.5289307, 0.5117778, 0.2969895, 
    0.1988276, 0.2598341, 0.1664843, 0.1640416, 0.2263988,
  0.5248144, 0.3820548, 0.4453025, 0.08683501, 0.1056618, 0.1054785, 
    0.008796287, 0.3217965, 0.4455738, 0.4554766, 0.4646307, 0.4049024, 
    0.179655, 0.2629269, 0.2868885, 0.254577, 0.1897437, 0.3520409, 
    0.3629252, 0.3616977, 0.4146, 0.2735611, 0.2434752, 0.4590874, 0.2637381, 
    0.2770714, 0.2788191, 0.29219, 0.4780154,
  0.5466233, 0.4770662, 0.3710031, 0.3190448, 0.2975199, 0.3589932, 
    0.3304653, 0.4118247, 0.3730453, 0.2267731, 0.3007612, 0.2983167, 
    0.3288504, 0.3759556, 0.4475572, 0.3594014, 0.3399193, 0.3585887, 
    0.2518193, 0.1415743, 0.1743058, 0.1914119, 0.189744, 0.2690542, 
    0.2616935, 0.446657, 0.4081293, 0.4795683, 0.503671,
  0.3363329, 0.3746754, 0.3310013, 0.3868814, 0.3848042, 0.3640358, 
    0.2456978, 0.137581, 0.1460649, 0.1934162, 0.2188362, 0.236008, 
    0.2138309, 0.1840625, 0.2234214, 0.1372467, 0.132339, 0.1625128, 
    0.1922453, 0.2248808, 0.2198077, 0.2500281, 0.3495895, 0.2837046, 
    0.186387, 0.2129331, 0.343015, 0.3093356, 0.3287745,
  0.2432628, 0.1135165, 0.06679933, 0.1529131, 0.1236433, 0.1141826, 
    0.1266436, 0.1700453, 0.1743373, 0.1288051, 0.07769725, 0.0547046, 
    0.02754319, 0.05144857, 0.4161397, 0.1166257, 0.1718655, 0.1823325, 
    0.1462917, 0.1555502, 0.1833414, 0.2322884, 0.2419482, 0.204711, 
    0.0411435, 0.1331105, 0.1040808, 0.1661858, 0.1861978,
  0.09192054, 0.01467551, 0.03502577, 0.03427841, 0.05217427, 0.04179683, 
    0.07864869, 0.114485, 0.1002276, 0.01024178, -3.295835e-06, 5.094819e-07, 
    -0.0001698525, 0.004949218, 0.02598429, 0.06063714, 0.08448356, 
    0.08755975, 0.07030219, 0.07894047, 0.05540191, 0.1186395, 0.1546819, 
    0.0189558, 0.02184991, 0.04016078, 0.02159799, 0.05070477, 0.04412323,
  0.1184005, 0.009573177, -7.760255e-05, 0.01344938, 0.001076726, 0.01840165, 
    0.04257405, 0.04658487, 0.05691196, 0.004698239, 5.40662e-10, 
    4.897082e-09, 0.009867216, 0.05491135, 0.080328, 0.1437834, 0.1089172, 
    0.1485685, 0.04832289, 0.03764783, 0.04889127, 0.1411173, 0.3365573, 
    0.002521246, 0.001128877, 0.06993857, 0.0224234, 0.07318999, 0.1030296,
  0.3299836, 0.04892978, -2.145872e-05, 0.00710182, 0.01187214, 0.02051206, 
    0.02627013, 0.07045699, 0.03162587, 0.04783706, 0.03517522, 0.03019948, 
    0.1491265, 0.04586744, 0.01769806, 0.01027245, 0.007524677, 0.008621074, 
    0.006588238, 0.02374279, 0.07236096, 0.254613, 0.1285563, 0.006770845, 
    1.330117e-06, -2.55785e-07, 0.005366822, 0.007033807, 0.09117571,
  0.4346142, 0.1144292, 0.002778855, 0.007805247, 0.03079742, 0.01347181, 
    0.02884562, 0.05013349, 0.02143792, 0.03081155, 0.05719792, 0.04887456, 
    0.03002269, 0.02575737, 0.02556882, 0.01842471, 0.01741009, 0.0129919, 
    0.01317218, 0.01283905, 0.07428867, 0.1862711, 0.0252635, 0.06375448, 
    0.04328369, 0.02459975, 0.01981196, 0.04803019, 0.1222294,
  0.04186317, 0.0487211, 0.006111868, 0.2227083, -0.000141068, 0.007970573, 
    0.06313614, 0.009693396, 0.0008346002, 0.007414706, 0.001911621, 
    0.02884176, 0.046884, 0.04967564, 0.04382049, 0.06153341, 0.08350525, 
    0.1270826, 0.1203469, 0.1024772, 0.1380419, 0.1062522, 0.1462616, 
    0.03555026, 0.05803317, 0.073744, 0.1558127, 0.1716061, 0.0588575,
  1.462559e-07, 1.252541e-10, 1.819752e-10, 6.016984e-10, 5.254603e-08, 
    0.03634045, 0.2990795, 0.1093039, 0.3083421, 0.04061846, 0.1039057, 
    0.04558576, 0.01552134, 0.005567019, 0.01026552, 0.01433614, 0.02850876, 
    0.1052659, 0.4060569, 0.2326923, 0.08818062, 0.08005232, 0.009825617, 
    0.005547582, 0.02197438, 0.02701012, 0.1534928, 0.08535275, 1.328644e-07,
  1.387422e-07, -3.263041e-05, -3.256937e-05, -4.993774e-08, 1.57804e-07, 
    -2.230844e-07, 0.001445346, 0.1728397, 0.3192399, 0.04318134, 0.1211354, 
    0.07694876, 0.07028682, 0.07101425, 0.1190517, 0.06899358, 0.07247901, 
    0.2084582, 0.3091416, 0.002281259, 1.40891e-05, 0.008112092, 0.01829713, 
    0.06653934, 0.06652103, 0.06440878, 0.09126636, 0.352562, -0.0009140769,
  -0.0007425143, 0.006096787, -4.788326e-06, 0.2235943, -8.624391e-05, 
    2.251463e-11, 7.610734e-06, 1.64878e-06, -2.179805e-05, 0.03723561, 
    0.2794448, 0.07015032, 0.4276898, 0.3843224, 0.4042735, 0.449815, 
    0.4808276, 0.3783599, 0.3704862, 0.00641515, -0.0002128258, 0.008507892, 
    0.009081734, 0.06429335, 0.137541, 0.2658738, 0.1974082, 0.3852276, 
    0.09610933,
  0.1124843, 0.1384506, 0.02696737, 0.08504412, 4.761e-05, 0.00461174, 
    0.02423124, 0.2333306, 0.0509393, 0.002646292, 0.02012573, 0.2153567, 
    0.3185032, 0.4336892, 0.5222884, 0.5918713, 0.5415158, 0.515622, 
    0.5096251, 0.03023867, 0.001167364, 0.005295634, 0.06022328, 0.1318203, 
    0.1436111, 0.2588147, 0.3712548, 0.4633608, 0.2856788,
  0.2505697, 0.05675537, 0.03355753, 0.1098321, 0.09175931, 0.03555196, 
    0.1453027, 0.1261515, 0.1301238, 0.1190704, 0.05382064, 0.2317975, 
    0.4179361, 0.2904561, 0.2790176, 0.4962313, 0.2795355, 0.3414662, 
    0.3095241, 0.0390104, 0.02160153, 0.07026291, 0.1210373, 0.2684505, 
    0.1726348, 0.2628489, 0.3758926, 0.408117, 0.3967778,
  0.5002823, 0.552771, 0.3953169, 0.3645308, 0.419224, 0.3965726, 0.2263891, 
    0.1108091, 0.1605701, 0.1420912, 0.2483271, 0.4031413, 0.4695687, 
    0.4216475, 0.4553332, 0.4076489, 0.3505268, 0.1735364, 0.1977035, 
    0.3515784, 0.3934077, 0.5625222, 0.3868725, 0.5244135, 0.3317097, 
    0.4147133, 0.3187971, 0.2489921, 0.514493,
  0.4095618, 0.4724112, 0.5603195, 0.568583, 0.6741715, 0.7336739, 0.6857122, 
    0.625369, 0.6727837, 0.5522594, 0.6876796, 0.6857191, 0.6825291, 
    0.6217757, 0.6380476, 0.6252319, 0.5674562, 0.5668328, 0.5748953, 
    0.6511965, 0.5927877, 0.368174, 0.3011892, 0.5043235, 0.2972056, 
    0.1930058, 0.261583, 0.4790885, 0.4684502,
  0.5002319, 0.4986661, 0.4971004, 0.4955347, 0.493969, 0.4924032, 0.4908375, 
    0.4989586, 0.4968937, 0.4948288, 0.4927639, 0.4906991, 0.4886342, 
    0.4865693, 0.5055794, 0.5138975, 0.5222156, 0.5305337, 0.5388518, 
    0.5471699, 0.555488, 0.5706394, 0.565952, 0.5612645, 0.556577, 0.5518895, 
    0.5472021, 0.5425146, 0.5014845,
  0.1927524, 0.2122944, 0.2075101, 0.2179234, 0.2240735, 0.2109681, 
    0.2429603, 0.2020059, 0.05384609, 0.1004908, 0.09033147, 0.0497913, 
    0.1003541, 0.00363986, 0.01575578, 0.07084827, 0.07709739, 0.06114937, 
    0.1233144, 0.09976692, 0.3573178, 0.5532531, 0.4949792, 0.3016467, 
    0.1989567, 0.2315162, 0.1370185, 0.155284, 0.2127501,
  0.5264474, 0.3289409, 0.3867749, 0.05449733, 0.08313394, 0.09410242, 
    0.003252823, 0.307166, 0.4478724, 0.4304871, 0.44719, 0.3834164, 
    0.1292136, 0.2205371, 0.2807502, 0.2792989, 0.2191321, 0.4277253, 
    0.4174523, 0.4043307, 0.4524351, 0.3231147, 0.2460029, 0.433344, 
    0.2687748, 0.3506168, 0.3534892, 0.3192764, 0.5200554,
  0.608493, 0.4879602, 0.318509, 0.2804173, 0.2484224, 0.300582, 0.3289091, 
    0.3652618, 0.2857262, 0.1592944, 0.2673296, 0.3180561, 0.3343211, 
    0.392841, 0.4633597, 0.3296074, 0.3425752, 0.3438819, 0.2046729, 
    0.1012838, 0.153165, 0.1512676, 0.1598049, 0.2541828, 0.2418551, 0.44255, 
    0.4632923, 0.5038628, 0.574963,
  0.3138264, 0.4011015, 0.3341872, 0.4173392, 0.3524778, 0.2873342, 
    0.1973422, 0.1118319, 0.1329254, 0.1800862, 0.2032566, 0.2233457, 
    0.1980845, 0.1532401, 0.1761051, 0.1021136, 0.09108549, 0.08959147, 
    0.1500433, 0.1748138, 0.2105976, 0.2788748, 0.3473732, 0.2768176, 
    0.1603948, 0.2204132, 0.3189965, 0.2793538, 0.3152593,
  0.2398426, 0.06479137, 0.02982443, 0.1070795, 0.08373081, 0.09467581, 
    0.1047658, 0.1410467, 0.1242365, 0.08066761, 0.04614415, 0.03212208, 
    0.01068775, 0.03464554, 0.3705768, 0.08478341, 0.1353317, 0.1482778, 
    0.1188528, 0.1302621, 0.1779041, 0.2178559, 0.2257528, 0.2231196, 
    0.02644799, 0.06343905, 0.08847817, 0.128672, 0.1844835,
  0.04198858, 0.00589289, 0.03262972, 0.01783754, 0.02520998, 0.02164763, 
    0.05630274, 0.04914175, 0.07294477, 0.004195368, -4.866793e-07, 
    -4.753543e-07, 0.000104372, 0.001897508, 0.0190591, 0.03428936, 
    0.06258452, 0.08457961, 0.06097427, 0.06557339, 0.03615805, 0.07019125, 
    0.08589572, 0.02929798, 0.030058, 0.01789436, 0.01332255, 0.03174654, 
    0.01975612,
  0.05828966, 0.01224533, -5.977921e-05, 0.005634002, -0.001817795, 
    0.003092513, 0.01183503, 0.01203201, 0.0231873, 0.002523029, 
    3.968861e-10, 4.26438e-09, 0.002924037, 0.02668726, 0.04350137, 
    0.07867336, 0.04744865, 0.05894928, 0.009521834, 0.007011716, 0.01424531, 
    0.04767621, 0.1270659, 0.02625767, 0.0003659258, 0.07766867, 0.01430541, 
    0.02235084, 0.0362358,
  0.1421079, 0.2226499, -3.525451e-05, 0.00576409, 0.002739683, 0.003325184, 
    0.003487421, 0.01837141, 0.009341418, 0.005979428, 0.01804981, 0.0073128, 
    0.1135867, 0.02389267, 0.003162079, 0.0005681132, 0.0004796286, 
    0.0006022378, 0.0008429325, 0.00704248, 0.02033147, 0.08498064, 
    0.2398048, 0.001443319, 2.146826e-07, -6.791995e-08, -0.002747558, 
    0.0006455141, 0.03423383,
  0.1515986, 0.06641266, 0.002018101, 0.003029417, 0.01559811, 0.00291108, 
    0.005436233, 0.01126113, 0.04916859, 0.02184621, 0.01431, 0.01073392, 
    0.02098293, 0.01186195, 0.01752872, 0.003430148, 0.006719552, 
    0.004524442, 0.003839199, 0.009484251, 0.0398524, 0.3947894, 0.2795689, 
    0.02207055, 0.03112626, 0.002758882, 0.002565854, 0.01086347, 0.06028322,
  0.03067053, 0.04373294, 0.003567181, 0.2308923, -6.360174e-05, 0.001458152, 
    0.0732564, 0.0007976187, -0.0005579251, 0.001139841, 0.0005820753, 
    0.01493283, 0.03094363, 0.0217338, 0.01858055, 0.03894835, 0.06674682, 
    0.08505917, 0.07277611, 0.06905349, 0.1040946, 0.1087624, 0.1956334, 
    0.02328235, 0.008667259, 0.03100104, 0.09866264, 0.100807, 0.05258339,
  1.302469e-07, 1.180817e-10, 1.794345e-10, 1.680937e-10, 2.817847e-08, 
    0.01342056, 0.2683751, 0.0528865, 0.3240095, 0.03586905, 0.04800847, 
    0.03291954, 0.003645337, 0.0005778844, 0.001161105, 0.001816119, 
    0.005861019, 0.03143943, 0.213448, 0.4501146, 0.2283119, 0.06832261, 
    0.002153048, 0.00166177, 0.006832281, 0.005063207, 0.05686431, 
    0.08718795, 1.271989e-07,
  1.327835e-07, -0.0001508606, -7.188729e-06, -1.070398e-06, 1.477375e-07, 
    -7.113568e-08, -0.001679976, 0.1809506, 0.3224863, 0.03867283, 0.1064989, 
    0.06110116, 0.07671358, 0.03920198, 0.09749652, 0.06096813, 0.03572865, 
    0.08471384, 0.2023928, 0.1927831, 4.156905e-06, 0.004528729, 0.00948757, 
    0.007982449, 0.01760472, 0.0111597, 0.01909516, 0.1484403, -0.00131712,
  -0.001578362, 0.002865556, -3.880183e-05, 0.2464095, -6.687072e-05, 
    2.670584e-11, 6.922999e-06, 1.530176e-06, -1.708473e-05, 0.03556927, 
    0.3273299, 0.08624556, 0.5000964, 0.5551542, 0.456201, 0.5261889, 
    0.5152928, 0.2611146, 0.3772746, 0.002484932, -0.0002026781, 0.009719701, 
    0.006529036, 0.0654323, 0.1819403, 0.2350529, 0.1297356, 0.2774076, 
    0.1382828,
  0.133085, 0.1123563, 0.02362335, 0.05846898, 1.189658e-05, 0.002187516, 
    0.01883761, 0.2307762, 0.04048296, 0.002218123, 0.02039645, 0.2027457, 
    0.4234655, 0.6117585, 0.7331904, 0.6404013, 0.7139853, 0.5394904, 
    0.3918267, 0.03321411, 0.000326203, 0.002310885, 0.06443318, 0.1092874, 
    0.1611518, 0.4164126, 0.3705923, 0.4594984, 0.2197368,
  0.2902099, 0.03962373, 0.01692711, 0.08063615, 0.07941973, 0.01912458, 
    0.1434534, 0.1161722, 0.105998, 0.1046984, 0.04466688, 0.2211276, 
    0.440446, 0.305416, 0.3320787, 0.6572358, 0.2628381, 0.3124007, 
    0.2742646, 0.03097856, 0.0180894, 0.06692115, 0.1276851, 0.2265688, 
    0.1945623, 0.2461072, 0.3437325, 0.4107052, 0.4394945,
  0.5289808, 0.4680775, 0.3951489, 0.3607263, 0.4131682, 0.3646356, 
    0.1879611, 0.06638651, 0.1146959, 0.07668001, 0.1995042, 0.3306161, 
    0.4314563, 0.3799428, 0.4650504, 0.4463432, 0.298979, 0.1828079, 
    0.2645406, 0.3082838, 0.3401373, 0.4821396, 0.3230598, 0.515191, 
    0.3159426, 0.4070437, 0.2892678, 0.2958018, 0.618288,
  0.5078288, 0.4872628, 0.5460719, 0.6555972, 0.7016723, 0.7367828, 
    0.7079265, 0.667078, 0.7439076, 0.7237198, 0.8244943, 0.7294193, 
    0.7250437, 0.6322338, 0.6848707, 0.7181044, 0.7009531, 0.6883082, 
    0.7751109, 0.8044645, 0.6425376, 0.4520831, 0.2983404, 0.5950755, 
    0.3540643, 0.1917995, 0.2764509, 0.5146587, 0.5918204,
  0.3106402, 0.3028205, 0.2950008, 0.2871811, 0.2793614, 0.2715417, 
    0.2637219, 0.2682148, 0.278383, 0.2885512, 0.2987194, 0.3088876, 
    0.3190558, 0.329224, 0.3858169, 0.3936033, 0.4013898, 0.4091763, 
    0.4169627, 0.4247492, 0.4325356, 0.4633153, 0.4531803, 0.4430454, 
    0.4329104, 0.4227755, 0.4126405, 0.4025055, 0.316896,
  0.215673, 0.1980826, 0.1950289, 0.2064826, 0.2924828, 0.1742962, 0.2166511, 
    0.2097372, 0.04917222, 0.04251159, 0.08899663, 0.05176216, 0.1223163, 
    0.001325506, 0.03877483, 0.08430272, 0.130111, 0.09385211, 0.1223993, 
    0.1022459, 0.3484782, 0.573041, 0.4672077, 0.292242, 0.215272, 0.2527889, 
    0.1982738, 0.1477693, 0.1985183,
  0.4672927, 0.2674193, 0.2834018, 0.02540819, 0.06865007, 0.08709653, 
    -0.0004661477, 0.2666146, 0.4470713, 0.3747864, 0.4065438, 0.3714087, 
    0.09055406, 0.1839138, 0.2865348, 0.2911864, 0.2776225, 0.4600759, 
    0.4186199, 0.4533705, 0.4886808, 0.3379676, 0.2507014, 0.4288642, 
    0.2843599, 0.4023176, 0.4300411, 0.4169224, 0.5260981,
  0.6064748, 0.4607402, 0.2635027, 0.2572047, 0.2095816, 0.2274825, 
    0.3092926, 0.3847156, 0.231404, 0.124947, 0.2207382, 0.3097802, 
    0.3308662, 0.3669846, 0.4435141, 0.3127653, 0.3089937, 0.2960203, 
    0.1678139, 0.06922188, 0.1203195, 0.1268572, 0.1375617, 0.2242883, 
    0.2231447, 0.3996634, 0.475694, 0.4716238, 0.5833434,
  0.2640284, 0.3599767, 0.3201314, 0.3982563, 0.3070936, 0.2225946, 
    0.1611669, 0.09161111, 0.1140778, 0.1575995, 0.1722637, 0.1820223, 
    0.1764868, 0.1262408, 0.1449999, 0.08644568, 0.06518205, 0.05829279, 
    0.1215321, 0.1423733, 0.2035292, 0.2829798, 0.3195498, 0.2479439, 
    0.122006, 0.1718277, 0.2811806, 0.2556462, 0.289271,
  0.2019581, 0.03674224, 0.01529625, 0.07340018, 0.05100587, 0.06850295, 
    0.07525899, 0.09385329, 0.08176287, 0.05145173, 0.02302849, 0.0195392, 
    0.004273907, 0.02324913, 0.3080374, 0.05429394, 0.09770456, 0.1146847, 
    0.08540077, 0.1091486, 0.1533662, 0.1993524, 0.1808303, 0.2306011, 
    0.01850311, 0.0315017, 0.05986353, 0.09543393, 0.134785,
  0.01978324, 0.001616309, 0.02868346, 0.01163464, 0.01398473, 0.01366047, 
    0.04126747, 0.02665158, 0.05091251, 0.002517833, -4.056402e-07, 
    -4.840974e-07, 0.0001820695, 0.0007455628, 0.01350931, 0.02206101, 
    0.04424382, 0.06550112, 0.04392613, 0.049025, 0.02363762, 0.03391535, 
    0.04677612, 0.02202167, 0.02999166, 0.007055159, 0.009010725, 0.01494183, 
    0.009050519,
  0.02351608, 0.01277605, -3.724978e-05, 0.003000733, -0.001802212, 
    0.0006190055, 0.002660871, 0.00443069, 0.0096879, 0.0006827483, 
    4.140582e-10, 3.762765e-09, 0.001522114, 0.01233061, 0.01961708, 
    0.0345206, 0.01223736, 0.01163253, 0.00349652, 0.002700532, 0.005787798, 
    0.01765646, 0.05317046, 0.034564, 9.155666e-05, 0.09110621, 0.005033458, 
    0.008000071, 0.01390432,
  0.06509008, 0.1509921, -4.034514e-05, 0.005271009, 9.384006e-05, 
    0.000441683, 0.0008280374, 0.005754505, 0.002811071, 0.001393283, 
    0.007427079, 0.001821628, 0.07426403, 0.01238135, 0.0004854675, 
    0.0001386594, 4.825948e-05, 0.0001903813, 0.0003504575, 0.002957402, 
    0.00738973, 0.03291276, 0.1124905, 0.0005288917, 3.922555e-08, 
    3.138948e-09, -0.001662107, 0.0002117337, 0.01523105,
  0.05780242, 0.04437316, 0.002337859, 0.001203341, 0.002283473, 
    0.0007744441, 0.002298765, 0.002347444, 0.05397449, 0.01499543, 
    0.002703479, 0.0009870613, 0.01572351, 0.01270547, 0.01337639, 
    0.000458741, 0.0003307356, 0.0003921596, 8.21353e-05, 0.0003392582, 
    0.00703237, 0.182563, 0.1410702, 0.009675381, 0.02663376, 0.0004077554, 
    0.0001428568, 0.001945313, 0.009515715,
  0.01414479, 0.03677743, 0.002412527, 0.2537289, -1.951503e-05, 
    4.710038e-05, 0.06952158, 1.854594e-05, -0.0004843723, 4.467845e-05, 
    6.37565e-05, 0.004653439, 0.01077679, 0.007799756, 0.008132715, 
    0.0255922, 0.04351654, 0.05707223, 0.04036889, 0.02968797, 0.06889509, 
    0.03562888, 0.2702688, 0.01905573, 0.001464466, 0.01403177, 0.04289085, 
    0.04044614, 0.05618877,
  1.195135e-07, 1.190726e-10, 1.818009e-10, -6.368889e-11, 2.261169e-08, 
    0.0008574034, 0.1998791, 0.01848852, 0.3352317, 0.0169067, 0.02322102, 
    0.01788696, 0.0005945081, -1.437662e-05, 0.0001528191, 0.0004079202, 
    0.001938595, 0.01079572, 0.1089742, 0.2429907, 0.06248381, 0.05375376, 
    0.0008184951, 0.0007307805, 0.001718421, 0.0007125633, 0.01895251, 
    0.03501749, 1.236164e-07,
  1.301802e-07, -0.0001231974, -8.624714e-07, -1.73561e-06, 1.410105e-07, 
    -1.154229e-09, -0.002736607, 0.1713365, 0.3144962, 0.03190707, 
    0.03833226, 0.01470578, 0.04811549, 0.01759311, 0.02302883, 0.01240416, 
    0.01304446, 0.02958084, 0.08796245, 0.239523, 2.103915e-06, 0.0009895198, 
    0.003215123, 0.001536346, 0.002553923, 0.00257108, 0.00666668, 
    0.06499813, 0.0007121539,
  -0.00151132, 0.0009280588, -0.0001700192, 0.2558618, -7.053163e-05, 
    2.983313e-11, 6.209465e-06, 1.445052e-06, -1.35946e-05, 0.03168101, 
    0.3556481, 0.1553731, 0.5704978, 0.6202014, 0.4614365, 0.5056608, 
    0.4236867, 0.1645765, 0.2246156, 0.001618152, -0.0002297916, 0.009158247, 
    0.004890086, 0.07265659, 0.09160106, 0.175569, 0.09145928, 0.1536541, 
    0.1462167,
  0.1309177, 0.09662378, 0.01560598, 0.03639026, -1.724355e-06, 0.0009844964, 
    0.01269311, 0.2082967, 0.03126473, 0.002603873, 0.01899791, 0.1947187, 
    0.5030614, 0.7023736, 0.7807146, 0.6464053, 0.7117001, 0.4797027, 
    0.2897075, 0.03817422, 0.002092004, 0.0009800004, 0.06169726, 0.09302918, 
    0.1676037, 0.4297295, 0.3664915, 0.427079, 0.1653762,
  0.2747344, 0.0294489, 0.008769901, 0.05321686, 0.06894307, 0.01201317, 
    0.1305767, 0.1053995, 0.09128579, 0.09966373, 0.04502556, 0.2148423, 
    0.4384635, 0.297655, 0.3923284, 0.7525395, 0.2508893, 0.2881032, 
    0.2486608, 0.02471987, 0.01393172, 0.06656688, 0.1573223, 0.1923965, 
    0.2343869, 0.2493682, 0.3095589, 0.3978907, 0.4626899,
  0.5922025, 0.3986933, 0.3593754, 0.2881512, 0.3563576, 0.3354994, 
    0.1344283, 0.04644588, 0.09232702, 0.04728046, 0.1534369, 0.2759735, 
    0.3585422, 0.3663007, 0.412349, 0.3938221, 0.2487022, 0.1988035, 
    0.2698119, 0.2312467, 0.2646882, 0.4589528, 0.26347, 0.5045041, 
    0.3688784, 0.3687263, 0.254503, 0.3302431, 0.6448188,
  0.5899056, 0.4061948, 0.554144, 0.6736379, 0.6518468, 0.7274455, 0.745528, 
    0.7552239, 0.7638382, 0.7375149, 0.7599838, 0.6875851, 0.6773783, 
    0.6062374, 0.6932244, 0.6913312, 0.7299448, 0.7246093, 0.738542, 
    0.7295401, 0.626053, 0.3978318, 0.2188589, 0.5445231, 0.3151225, 
    0.1998744, 0.2897486, 0.5616896, 0.6940376,
  0.1824317, 0.1766734, 0.1709152, 0.165157, 0.1593987, 0.1536405, 0.1478823, 
    0.1262592, 0.1352835, 0.1443078, 0.1533321, 0.1623564, 0.1713806, 
    0.1804049, 0.1864895, 0.1934193, 0.200349, 0.2072788, 0.2142085, 
    0.2211383, 0.2280681, 0.25168, 0.2414842, 0.2312884, 0.2210926, 
    0.2108968, 0.200701, 0.1905051, 0.1870382,
  0.21429, 0.1708363, 0.1177971, 0.1881295, 0.2323073, 0.145801, 0.1754809, 
    0.1904949, 0.03309298, 0.03338964, 0.06982041, 0.09250019, 0.1135427, 
    0.004358326, 0.09383953, 0.09850153, 0.2044274, 0.1471221, 0.1316578, 
    0.1050728, 0.3407155, 0.5792033, 0.4321436, 0.2755395, 0.1993959, 
    0.3093791, 0.2107833, 0.1356543, 0.1868677,
  0.4058149, 0.2040445, 0.2055663, 0.01444073, 0.04834439, 0.08273284, 
    -0.0009077392, 0.2169347, 0.4435938, 0.337678, 0.362843, 0.3750267, 
    0.06905518, 0.1490589, 0.2938959, 0.2791459, 0.321476, 0.4922826, 
    0.4116831, 0.5018615, 0.4491194, 0.3787672, 0.2804622, 0.4155576, 
    0.2728834, 0.4239068, 0.4597276, 0.4904873, 0.4822504,
  0.510604, 0.4168741, 0.2165105, 0.2049248, 0.166852, 0.1605993, 0.2942797, 
    0.3345908, 0.1877068, 0.09992747, 0.1718908, 0.2682475, 0.2800055, 
    0.3331154, 0.3927857, 0.2826478, 0.2509769, 0.2332906, 0.1366633, 
    0.04576589, 0.1010824, 0.0870818, 0.1158941, 0.1821466, 0.1875806, 
    0.349397, 0.4248672, 0.450087, 0.5197064,
  0.2247003, 0.301527, 0.2910612, 0.3576985, 0.2520632, 0.1648042, 0.1321468, 
    0.07178736, 0.09344572, 0.1242992, 0.1274973, 0.1307841, 0.1238135, 
    0.09161378, 0.1156385, 0.07363066, 0.04499536, 0.03473642, 0.09599572, 
    0.1130303, 0.1801201, 0.2686703, 0.2682707, 0.218197, 0.06850883, 
    0.1078449, 0.2263718, 0.211701, 0.2690964,
  0.1463173, 0.01872747, 0.0080803, 0.04416978, 0.02931768, 0.043663, 
    0.04263892, 0.05423148, 0.04735772, 0.03463645, 0.01327465, 0.01060312, 
    0.001781453, 0.01439502, 0.247457, 0.03627406, 0.06920762, 0.0855496, 
    0.06073318, 0.07928175, 0.120183, 0.154637, 0.113627, 0.222535, 
    0.01469467, 0.02039793, 0.03408242, 0.06380015, 0.09522015,
  0.01108166, 0.0009188852, 0.02539571, 0.007195329, 0.004864176, 
    0.009678279, 0.02522582, 0.01480249, 0.03671163, 0.001772184, 
    -2.954066e-07, -1.961288e-07, 0.0002144028, 0.00037212, 0.009403645, 
    0.01583627, 0.03188608, 0.05171996, 0.02886695, 0.02995155, 0.01540516, 
    0.01340176, 0.02424872, 0.01583844, 0.02269411, 0.004013652, 0.005775738, 
    0.006480937, 0.004694513,
  0.01401748, 0.01290655, -4.608682e-05, 0.001750632, -0.001612163, 
    0.0002642119, 0.001019083, 0.002208356, 0.004140846, 0.0002426405, 
    4.165426e-10, 1.510181e-09, 0.0009712242, 0.004850458, 0.008546079, 
    0.01419143, 0.003199779, 0.004321225, 0.002032228, 0.001525959, 
    0.002600957, 0.008329006, 0.02950679, 0.03298808, 5.262472e-05, 
    0.08884269, 0.001882892, 0.003846426, 0.007157161,
  0.03664028, 0.07702064, -2.80079e-05, 0.00465733, 3.189917e-05, 
    0.0001117345, 0.000451827, 0.001891896, 0.00112202, 0.0006667975, 
    0.003236458, 0.0007331115, 0.03876973, 0.005251249, 0.0002100338, 
    7.721569e-05, 2.136333e-05, 0.0001106302, 0.0001931469, 0.00157125, 
    0.003672895, 0.01707764, 0.06131114, 0.0003556974, 4.643837e-08, 
    7.344683e-09, -0.001093508, 0.0001018603, 0.008501216,
  0.02893026, 0.04434452, 0.002018272, 9.728134e-05, 0.0001677869, 
    0.0004214507, 0.001322866, 0.0009744808, 0.03928697, 0.01267492, 
    0.0006022408, 0.000249623, 0.009738751, 0.00864688, 0.007620716, 
    9.771841e-05, 2.279002e-05, 2.773009e-05, 1.714998e-05, 3.706129e-05, 
    0.002567596, 0.07294498, 0.06914728, 0.005835742, 0.02946903, 
    0.000202238, 6.644911e-05, 0.0009538047, 0.003518024,
  0.006014039, 0.02745075, 0.0009564455, 0.2504074, -5.836826e-06, 
    2.904238e-06, 0.05599853, 7.191529e-06, -0.0001897148, 9.542608e-06, 
    4.924865e-06, 0.001470633, 0.004449532, 0.002447973, 0.00305395, 
    0.01745137, 0.01998518, 0.03506994, 0.02294008, 0.01118704, 0.03742946, 
    0.01385, 0.2475225, 0.01694043, 0.0005618529, 0.007025633, 0.0192924, 
    0.01853436, 0.04092629,
  1.10271e-07, 1.145066e-10, 1.817571e-10, -1.926451e-10, 2.242221e-08, 
    0.0003798977, 0.104546, 0.00384361, 0.3140387, 0.002692347, 0.01148081, 
    0.007816714, 0.0001758761, -1.144319e-05, 7.573803e-05, 0.0001940264, 
    0.001003688, 0.00541774, 0.06047364, 0.1180178, 0.03119867, 0.04543811, 
    0.0004696527, -3.618982e-05, 0.0005857681, 0.0002862313, 0.008009935, 
    0.01232369, 1.209158e-07,
  1.282576e-07, -5.588038e-06, 4.531151e-05, -3.067732e-06, 1.364648e-07, 
    5.366209e-09, -0.003410204, 0.1519774, 0.2969581, 0.01737085, 0.01520915, 
    0.004737876, 0.02068684, 0.005002494, 0.006851531, 0.002527412, 
    0.006510044, 0.01452054, 0.04556566, 0.1689532, 1.06689e-06, 
    0.0002797751, 0.00106039, 0.0006823611, 0.0009418033, 0.001175566, 
    0.003557747, 0.03015965, 0.002015861,
  -0.00104171, 0.0001891178, -0.0001713924, 0.2301247, -6.515768e-05, 
    3.232073e-11, 5.707247e-06, 1.400897e-06, -1.011499e-05, 0.02532843, 
    0.3405862, 0.2545649, 0.6476256, 0.5241212, 0.3761846, 0.4610384, 
    0.3268666, 0.1351356, 0.1453903, 0.001419214, -0.0002084693, 0.006210175, 
    0.004430361, 0.073501, 0.04817265, 0.1002279, 0.0437876, 0.07523052, 
    0.1253016,
  0.1140388, 0.07602142, 0.01056379, 0.01971275, -8.480118e-06, 0.0002102684, 
    0.006753494, 0.1833114, 0.02648687, 0.003998617, 0.02268297, 0.1780305, 
    0.6010256, 0.690618, 0.6989489, 0.6164558, 0.6345968, 0.4013511, 
    0.2285884, 0.03732563, 0.002788963, 0.0002796363, 0.05466696, 0.07849605, 
    0.1727236, 0.4379918, 0.3639056, 0.3759989, 0.1300867,
  0.1925354, 0.02378184, 0.004638867, 0.03307385, 0.05958468, 0.008181606, 
    0.1174272, 0.09790164, 0.08421218, 0.09635998, 0.0443076, 0.1982761, 
    0.4280686, 0.2777027, 0.446205, 0.7627456, 0.2284264, 0.2606622, 
    0.1985902, 0.02789385, 0.00971341, 0.07168625, 0.2068882, 0.1553217, 
    0.2241884, 0.2458758, 0.2647678, 0.364332, 0.4253062,
  0.5694719, 0.3604665, 0.3088867, 0.2340965, 0.3403727, 0.3409763, 
    0.1004945, 0.03177177, 0.07535886, 0.03138348, 0.1207533, 0.2292056, 
    0.3033331, 0.3246668, 0.3689264, 0.3724851, 0.2156759, 0.2380453, 
    0.2372099, 0.1646458, 0.1933365, 0.4204463, 0.2196623, 0.4727894, 
    0.3902463, 0.3227303, 0.2069456, 0.3316634, 0.5839799,
  0.6702647, 0.3762229, 0.5158728, 0.6659769, 0.5609642, 0.7312171, 
    0.8159826, 0.7848464, 0.7927262, 0.7694405, 0.6992024, 0.6791965, 
    0.6567651, 0.6221851, 0.6508035, 0.6608775, 0.7060143, 0.7509662, 
    0.6867545, 0.6517804, 0.5639144, 0.3236109, 0.1745465, 0.4704233, 
    0.2801257, 0.1812162, 0.2928094, 0.5773346, 0.7253532,
  0.1078733, 0.1031233, 0.09837333, 0.09362333, 0.08887332, 0.08412331, 
    0.07937331, 0.06800117, 0.07074249, 0.0734838, 0.07622512, 0.07896643, 
    0.08170775, 0.08444905, 0.08735736, 0.09391793, 0.1004785, 0.107039, 
    0.1135996, 0.1201602, 0.1267207, 0.125754, 0.1212021, 0.1166503, 
    0.1120984, 0.1075465, 0.1029947, 0.09844279, 0.1116733,
  0.1589639, 0.122722, 0.09375569, 0.1323944, 0.09869929, 0.1099753, 
    0.131665, 0.1275226, 0.05068134, 0.02670457, 0.02360626, 0.09717391, 
    0.1067703, 0.004344345, 0.1367391, 0.1972742, 0.2932443, 0.1827246, 
    0.1256073, 0.1098801, 0.3923734, 0.5531359, 0.3792595, 0.2163536, 
    0.2380323, 0.3757893, 0.2265854, 0.117572, 0.1855955,
  0.3156371, 0.1693328, 0.1539192, 0.009533782, 0.03955067, 0.07669723, 
    -0.0009398494, 0.1856846, 0.4346073, 0.3069507, 0.3457949, 0.3927671, 
    0.05419525, 0.1104232, 0.2896887, 0.2550217, 0.2864547, 0.3951788, 
    0.3714889, 0.5400417, 0.3754801, 0.3792551, 0.3047951, 0.4036642, 
    0.268612, 0.4053724, 0.4316685, 0.4780741, 0.4064429,
  0.4131348, 0.3486371, 0.1660752, 0.1466951, 0.1109548, 0.1188841, 
    0.2672419, 0.2863131, 0.1548095, 0.07398655, 0.1218485, 0.2241047, 
    0.2107007, 0.271547, 0.3124642, 0.2325209, 0.1874311, 0.1731612, 
    0.1057924, 0.03216368, 0.07858916, 0.05986374, 0.08765954, 0.1337747, 
    0.1453485, 0.2816211, 0.3642636, 0.3886179, 0.4385986,
  0.196624, 0.2430479, 0.2623111, 0.3002172, 0.199583, 0.122615, 0.1030259, 
    0.05308598, 0.0706079, 0.09098754, 0.08938827, 0.07860361, 0.06688374, 
    0.05598003, 0.07322452, 0.05587987, 0.02981335, 0.02113255, 0.07053852, 
    0.07925709, 0.1464913, 0.1988272, 0.2003716, 0.1875042, 0.03589467, 
    0.06530885, 0.1623499, 0.1624651, 0.2525839,
  0.1016608, 0.009852494, 0.004690345, 0.02444266, 0.01683575, 0.02474944, 
    0.02517497, 0.03318088, 0.02470516, 0.02018519, 0.006941046, 0.005913537, 
    0.001045112, 0.008372768, 0.2007321, 0.02136314, 0.04565666, 0.05738539, 
    0.0413653, 0.04903542, 0.08305568, 0.1056428, 0.06648814, 0.2133046, 
    0.009527651, 0.01045453, 0.01801819, 0.03584156, 0.06005892,
  0.007134829, 0.0006454772, 0.02006934, 0.004663681, 0.002011576, 
    0.005801275, 0.0154868, 0.009212196, 0.01820449, 0.001361924, 
    -2.302478e-07, -7.154267e-08, 5.535613e-05, 0.00025888, 0.005016967, 
    0.008139598, 0.01826655, 0.03402961, 0.0142703, 0.01415476, 0.005097442, 
    0.006272135, 0.01518776, 0.01147827, 0.0175307, 0.002605553, 0.002066377, 
    0.00261666, 0.002784352,
  0.009577096, 0.009328283, -3.524243e-05, 0.00126268, -0.001330154, 
    0.0002091427, 0.0006267217, 0.001393, 0.0022828, 0.0001395581, 
    4.178905e-10, 1.480607e-09, 0.0006994452, 0.002512558, 0.003387752, 
    0.005761201, 0.001707918, 0.002520319, 0.001397663, 0.00102125, 
    0.00160335, 0.005021572, 0.01986704, 0.02929701, 3.585554e-05, 0.0779161, 
    0.0008994961, 0.002326023, 0.00451166,
  0.02446408, 0.04099413, -1.879172e-05, 0.003150879, 1.741762e-05, 
    4.357268e-05, 0.0002961851, 0.0009947758, 0.0005674089, 0.0004880323, 
    0.001681481, 0.0003981956, 0.01652456, 0.001723411, 0.0001277367, 
    5.359739e-05, 1.254238e-05, 7.545351e-05, 0.0001255292, 0.001006089, 
    0.00227296, 0.0109207, 0.03948141, 0.0001946804, 3.944956e-08, 
    8.909136e-09, -0.0006037909, 6.095533e-05, 0.005598574,
  0.01827615, 0.03703563, 0.001341838, -0.0002916098, 5.586159e-05, 
    0.0002797629, 0.0008929686, 0.0006125347, 0.02145564, 0.01344176, 
    0.0002977086, 0.0001224082, 0.004589871, 0.004462597, 0.003503215, 
    2.447863e-05, 1.041651e-05, 1.447736e-05, 9.212639e-06, 1.62513e-05, 
    0.001410101, 0.03771378, 0.04377099, 0.005279738, 0.03378166, 
    0.0001383498, 4.19328e-05, 0.0005906582, 0.002025684,
  0.004040186, 0.01864851, 0.0002875862, 0.2188768, -2.526719e-06, 
    1.445071e-06, 0.03607065, 3.628912e-06, -5.925733e-05, 4.283177e-06, 
    3.825734e-06, 0.0005880972, 0.001815299, 0.0009375393, 0.0009771071, 
    0.008754878, 0.008416134, 0.01908319, 0.01072651, 0.004316276, 0.0166313, 
    0.005743366, 0.2060851, 0.02290839, 0.0003234395, 0.003512804, 
    0.008080659, 0.007807379, 0.02893484,
  1.048723e-07, 1.207626e-10, 1.826691e-10, -3.890251e-10, 2.258391e-08, 
    0.0001693317, 0.03140135, 0.001011421, 0.2416253, 0.000816563, 
    0.00497747, 0.001788939, 8.409756e-05, -5.527806e-06, 4.529718e-05, 
    0.0001153739, 0.000617013, 0.002889835, 0.03583733, 0.06625959, 
    0.01557119, 0.03797925, 0.000313072, -0.0004755513, 0.0001675426, 
    0.0001688015, 0.004586175, 0.006736741, 1.190639e-07,
  1.279438e-07, 6.862975e-06, 0.0001022486, -3.351344e-06, 1.333852e-07, 
    5.063961e-09, -0.004485493, 0.1282093, 0.2628396, 0.009169026, 
    0.005964471, 0.002136181, 0.006539888, 0.002571462, 0.003510792, 
    0.001350323, 0.003930077, 0.008912082, 0.02768429, 0.1243074, 
    9.839869e-07, 0.0003395706, 0.0003632869, 0.0004172696, 0.000532098, 
    0.0007220649, 0.002364938, 0.01824287, 0.002190139,
  -0.0006378325, -8.753657e-05, -0.0001684777, 0.207013, -5.568781e-05, 
    3.425691e-11, 5.32385e-06, 1.3713e-06, -7.926708e-06, 0.01638216, 
    0.3081199, 0.275115, 0.6042143, 0.4228815, 0.3075178, 0.4253776, 
    0.235943, 0.1068198, 0.1018572, 0.0009516253, -0.0001289198, 0.003506809, 
    0.003776671, 0.09449072, 0.02548622, 0.04850688, 0.01679912, 0.03857427, 
    0.0982926,
  0.0922286, 0.05254711, 0.01205886, 0.009006116, -4.211722e-06, 4.87153e-05, 
    0.003658778, 0.1658392, 0.02286669, 0.003232148, 0.02590622, 0.1542263, 
    0.6033717, 0.6366022, 0.6113579, 0.5237566, 0.5008883, 0.3081276, 
    0.1499038, 0.03437825, 0.004267931, 0.0001191033, 0.04275221, 0.0585972, 
    0.1849614, 0.3733016, 0.2860521, 0.2881967, 0.09766044,
  0.1409332, 0.01719048, 0.002711867, 0.02091441, 0.0490083, 0.009548294, 
    0.09572068, 0.09071866, 0.08220322, 0.0839356, 0.03958232, 0.1705545, 
    0.3906381, 0.2445096, 0.4701238, 0.6484795, 0.1932595, 0.2325344, 
    0.1379832, 0.02430959, 0.005586172, 0.06284908, 0.2124407, 0.1249164, 
    0.1861992, 0.2257463, 0.1958264, 0.2834808, 0.3258488,
  0.4539506, 0.2871065, 0.2606724, 0.1858326, 0.3341519, 0.4287219, 
    0.07624175, 0.02195622, 0.06093479, 0.01940551, 0.09705806, 0.1879222, 
    0.2656894, 0.2702869, 0.3389268, 0.3524367, 0.1752455, 0.2350605, 
    0.222358, 0.1266634, 0.1405535, 0.3687106, 0.1762493, 0.4253956, 
    0.3611464, 0.274218, 0.1770571, 0.3147669, 0.5212353,
  0.6836019, 0.3541081, 0.4360135, 0.6110986, 0.4825419, 0.6661838, 
    0.7994158, 0.8253083, 0.7920077, 0.7465153, 0.6521013, 0.6304242, 
    0.6160914, 0.607716, 0.5749515, 0.6070834, 0.6537879, 0.669006, 
    0.5676551, 0.5486228, 0.4806301, 0.2531697, 0.1462686, 0.3942811, 
    0.2560838, 0.1619289, 0.2727583, 0.5277892, 0.722822,
  0.06280475, 0.0592671, 0.05572946, 0.05219181, 0.04865415, 0.0451165, 
    0.04157886, 0.01481379, 0.01534458, 0.01587538, 0.01640617, 0.01693697, 
    0.01746776, 0.01799856, 0.03316036, 0.03641255, 0.03966474, 0.04291693, 
    0.04616912, 0.04942131, 0.0526735, 0.0594155, 0.05917016, 0.05892483, 
    0.0586795, 0.05843416, 0.05818883, 0.0579435, 0.06563488,
  0.152738, 0.1112433, 0.04055041, 0.07306843, 0.05106652, 0.08105221, 
    0.08258934, 0.0375369, 0.0347288, 0.02367296, 0.02023496, 0.08263542, 
    0.08429301, 0.002860357, 0.1968048, 0.2566608, 0.2921907, 0.2279511, 
    0.1132297, 0.2036583, 0.4536539, 0.5541665, 0.3497598, 0.1718717, 
    0.3676457, 0.4556513, 0.253722, 0.09570386, 0.1326005,
  0.2520731, 0.1334419, 0.1236507, 0.006859567, 0.02360948, 0.07130838, 
    -0.001141631, 0.1673189, 0.4154786, 0.2749804, 0.3182407, 0.3947141, 
    0.04863392, 0.09606442, 0.2831696, 0.2452364, 0.2318289, 0.3125016, 
    0.3078764, 0.4721248, 0.3249315, 0.3565952, 0.2906112, 0.3848901, 
    0.2610956, 0.3639303, 0.387121, 0.3955691, 0.3273375,
  0.349612, 0.2775654, 0.1312435, 0.1158645, 0.08233403, 0.09672957, 
    0.2391709, 0.2487746, 0.1330893, 0.05974842, 0.09487391, 0.1895344, 
    0.1628535, 0.2242837, 0.2335844, 0.1781754, 0.1421207, 0.1373786, 
    0.08752704, 0.02523579, 0.06350344, 0.04744032, 0.0698302, 0.1000107, 
    0.1161548, 0.2319354, 0.3106225, 0.3259055, 0.3717851,
  0.1763688, 0.2034115, 0.2250682, 0.249473, 0.1612402, 0.0979532, 
    0.08447228, 0.03979566, 0.05663007, 0.07047681, 0.06472105, 0.0501864, 
    0.04171041, 0.03573115, 0.05255033, 0.03693132, 0.02177201, 0.01538417, 
    0.04612952, 0.0575561, 0.110158, 0.1458053, 0.142676, 0.177156, 
    0.02590861, 0.04611417, 0.1264426, 0.1336335, 0.2267414,
  0.06644248, 0.006606597, 0.003323128, 0.01369214, 0.01087328, 0.01475595, 
    0.01468329, 0.02217202, 0.01531729, 0.0132641, 0.003911326, 0.003687061, 
    0.0007559583, 0.005568746, 0.1675527, 0.01180048, 0.02751127, 0.03609264, 
    0.02603497, 0.03251319, 0.05346001, 0.07582049, 0.04337798, 0.2006693, 
    0.006747274, 0.005673332, 0.01017985, 0.02076626, 0.03700419,
  0.005398344, 0.0005064534, 0.01802641, 0.002935792, 0.001378239, 
    0.00242552, 0.009519539, 0.006791842, 0.008921826, 0.001110857, 
    -1.818635e-07, -2.430976e-08, 0.0001154634, 0.0002074928, 0.002143338, 
    0.004431881, 0.009091981, 0.01909084, 0.005923274, 0.007058396, 
    0.002618708, 0.004039542, 0.0113266, 0.009279064, 0.01421229, 
    0.001886478, 0.001070627, 0.001794758, 0.002096166,
  0.007333498, 0.006656447, -2.684965e-05, 0.001013632, -0.0009698174, 
    0.0001786167, 0.0004590249, 0.001020932, 0.001538155, 9.934913e-05, 
    4.205257e-10, 1.471899e-09, 0.0005526416, 0.001791595, 0.001798719, 
    0.003079932, 0.00116875, 0.001782356, 0.001072551, 0.0007674272, 
    0.001178826, 0.003563246, 0.01505366, 0.02613172, 2.83318e-05, 
    0.07045618, 0.000529101, 0.001637605, 0.003269734,
  0.01847407, 0.02524411, -1.230417e-05, 0.002326172, 1.206967e-05, 
    2.560744e-05, 0.0002200093, 0.0006873937, 0.0003747036, 0.0004549189, 
    0.001201285, 0.000293158, 0.008127244, 0.0007542147, 9.411973e-05, 
    4.128947e-05, 9.344987e-06, 5.77192e-05, 9.308697e-05, 0.0007376574, 
    0.001633292, 0.007996696, 0.02919396, 0.0006729316, 3.692117e-08, 
    1.05348e-08, -0.0002890496, 4.269931e-05, 0.004188107,
  0.01328486, 0.03048387, 0.0003836858, -0.0002764567, 2.983256e-05, 
    0.0002106847, 0.0006741066, 0.0004482927, 0.01730785, 0.02737865, 
    0.0001928211, 8.4258e-05, 0.002330119, 0.002139087, 0.00147727, 
    1.972896e-05, 6.35042e-06, 9.696136e-06, 5.820447e-06, 9.465234e-06, 
    0.0009379177, 0.0249417, 0.03185019, 0.004336744, 0.03308025, 
    0.0001057006, 3.092027e-05, 0.0004260633, 0.001403923,
  0.008163763, 0.01363805, 6.115073e-05, 0.1879372, -1.389153e-06, 
    8.942868e-07, 0.02369895, 2.598947e-06, -4.671215e-05, 2.966088e-06, 
    3.16445e-06, 0.0002893312, 0.001003954, 0.0004781004, 0.0004140915, 
    0.004223715, 0.003965969, 0.009381312, 0.004968614, 0.001929815, 
    0.006677322, 0.002438778, 0.1816465, 0.02772808, 0.0002215361, 
    0.001810121, 0.003580276, 0.003858503, 0.02125167,
  1.010254e-07, 1.197135e-10, 1.856693e-10, -4.760051e-10, 2.213681e-08, 
    9.844166e-05, 0.01056618, 0.0004980977, 0.1502732, 0.0003181246, 
    0.002286894, 0.0007304913, 5.565282e-05, -3.447296e-06, 3.197107e-05, 
    8.051822e-05, 0.0004412434, 0.002037574, 0.02433763, 0.04480691, 
    0.01022893, 0.03187586, 0.000233785, -0.0007793798, 8.607082e-05, 
    0.0001150384, 0.003137063, 0.004429558, 1.177535e-07,
  1.277267e-07, -2.296544e-06, 0.0001947613, -2.286727e-06, 1.316939e-07, 
    4.871638e-09, -0.004431816, 0.1135545, 0.2331715, 0.005256595, 
    0.003196345, 0.001355211, 0.003014361, 0.001766714, 0.002458082, 
    0.0009338815, 0.002784234, 0.006317742, 0.01992823, 0.09994958, 
    9.519865e-07, 0.001605247, 0.003657347, 0.0002955391, 0.0003722196, 
    0.0005202256, 0.001695631, 0.01305896, 0.002153076,
  -0.0001933204, -0.0001864354, -0.0001486931, 0.187059, -4.785371e-05, 
    3.812192e-11, 5.019267e-06, 1.354249e-06, -6.348304e-06, 0.0111254, 
    0.2702593, 0.246916, 0.5074316, 0.3222165, 0.2522444, 0.3492777, 
    0.1618555, 0.07086328, 0.06985319, 0.0006490608, -8.906339e-05, 
    0.001780362, 0.003303477, 0.0621459, 0.01161887, 0.0234008, 0.007090523, 
    0.02308646, 0.07815745,
  0.07709971, 0.03830884, 0.01306796, 0.004929168, -1.796181e-06, 
    2.128945e-05, 0.002161256, 0.1551636, 0.02057425, 0.00320908, 0.02949208, 
    0.1346326, 0.5803137, 0.5563152, 0.5038207, 0.3676927, 0.370773, 
    0.216657, 0.09351167, 0.03088157, 0.004420883, 4.929385e-05, 0.03538533, 
    0.04727314, 0.1901824, 0.3151968, 0.210972, 0.2111616, 0.0688403,
  0.1114586, 0.01166961, 0.001977388, 0.01387343, 0.04286103, 0.01556853, 
    0.08070086, 0.08377703, 0.0886226, 0.07500897, 0.03558911, 0.1465328, 
    0.3418018, 0.2066628, 0.4293758, 0.4784106, 0.1642053, 0.2076082, 
    0.1002889, 0.02133004, 0.003277237, 0.05668948, 0.2075877, 0.1033474, 
    0.1524505, 0.1814177, 0.1508598, 0.2033734, 0.2254018,
  0.3311231, 0.2133776, 0.2294396, 0.1392494, 0.3204045, 0.4882177, 
    0.05737195, 0.01535372, 0.05042423, 0.0153511, 0.08058939, 0.1571626, 
    0.2349124, 0.2356953, 0.3073968, 0.3168153, 0.148107, 0.2487923, 
    0.2047959, 0.1352628, 0.1094818, 0.3214078, 0.1426376, 0.3816589, 
    0.2885219, 0.236397, 0.1610297, 0.2793491, 0.3980663,
  0.6479748, 0.3603064, 0.4006427, 0.5235876, 0.4006683, 0.567077, 0.6850292, 
    0.7437103, 0.7221592, 0.6525257, 0.5650055, 0.544745, 0.5247322, 
    0.5455204, 0.480097, 0.5171471, 0.5439091, 0.5271821, 0.466875, 0.455274, 
    0.4149494, 0.2129374, 0.1263499, 0.3498506, 0.2300633, 0.1478539, 
    0.2462754, 0.4880478, 0.6727296,
  0.02716677, 0.02403313, 0.0208995, 0.01776586, 0.01463223, 0.0114986, 
    0.008364962, 0.008004916, 0.009385442, 0.01076597, 0.0121465, 0.01352702, 
    0.01490755, 0.01628807, 0.02260991, 0.02462888, 0.02664785, 0.02866683, 
    0.0306858, 0.03270477, 0.03472374, 0.03191519, 0.03164933, 0.03138346, 
    0.0311176, 0.03085173, 0.03058587, 0.03032, 0.02967368,
  0.09622999, 0.06526627, 0.02328075, 0.02135875, 0.004396209, 0.05858721, 
    0.06648326, 0.02048876, 0.02338203, 0.02176799, 0.0142569, 0.06383775, 
    0.07595282, 0.003044721, 0.3749366, 0.2552382, 0.2288624, 0.2307392, 
    0.1408904, 0.2796127, 0.4643455, 0.5564777, 0.3058521, 0.1689578, 
    0.3174032, 0.5330403, 0.2776205, 0.1054292, 0.09991155,
  0.2140725, 0.1139818, 0.1042604, 0.005592216, 0.03499286, 0.07509637, 
    -0.001095829, 0.1583802, 0.3957831, 0.2670464, 0.3058015, 0.3879873, 
    0.04614004, 0.08862416, 0.2775335, 0.234274, 0.2086934, 0.2842482, 
    0.255328, 0.421641, 0.292305, 0.3468848, 0.2676034, 0.357361, 0.2466821, 
    0.3340033, 0.3490661, 0.3518332, 0.2979723,
  0.3100312, 0.2443619, 0.1112351, 0.1003488, 0.06891142, 0.08572555, 
    0.2202123, 0.2317347, 0.1210972, 0.05121883, 0.07949118, 0.1635685, 
    0.1402391, 0.1885229, 0.1853219, 0.1480757, 0.1191555, 0.1158068, 
    0.07737088, 0.02193773, 0.05485212, 0.04144246, 0.05888345, 0.0842548, 
    0.1016567, 0.2057104, 0.2836249, 0.285293, 0.3301179,
  0.1480512, 0.1768593, 0.1900882, 0.2082415, 0.1328737, 0.08470193, 
    0.07189627, 0.03371635, 0.04923601, 0.06129522, 0.05342919, 0.03835213, 
    0.03167425, 0.02579748, 0.03868593, 0.02634095, 0.01716676, 0.01280586, 
    0.03356716, 0.04613459, 0.08533067, 0.1136508, 0.1115652, 0.2058178, 
    0.02143728, 0.03797245, 0.1067223, 0.1143287, 0.195987,
  0.04694566, 0.00526628, 0.002751236, 0.0094976, 0.008614925, 0.01017296, 
    0.01034707, 0.01649744, 0.01165003, 0.01016336, 0.002821061, 0.002791305, 
    0.0006323395, 0.004409984, 0.1548177, 0.008190244, 0.0189264, 0.02517539, 
    0.01893839, 0.02488788, 0.03920891, 0.05784047, 0.03306389, 0.2006082, 
    0.00400297, 0.004228577, 0.006924296, 0.01428133, 0.02719941,
  0.00456324, 0.0004419036, 0.0219034, 0.002147681, 0.001160337, 0.001712467, 
    0.006751463, 0.005728232, 0.005771465, 0.0009301668, -1.45945e-07, 
    -3.851816e-09, 0.001641757, 0.000180765, 0.001139339, 0.002996559, 
    0.005517223, 0.01231854, 0.003265483, 0.004454619, 0.001913638, 
    0.003195786, 0.009528771, 0.007942005, 0.01367948, 0.001545583, 
    0.0007783597, 0.001516048, 0.001788388,
  0.006220866, 0.006210451, -2.29267e-05, 0.0008801724, -0.0009476612, 
    0.0001460299, 0.0003874559, 0.0008517159, 0.001242, 8.091701e-05, 
    4.272656e-10, 3.275129e-09, 0.0004786764, 0.001498549, 0.001248054, 
    0.002254083, 0.0009301184, 0.00143116, 0.0009045143, 0.0006414574, 
    0.0009736657, 0.002889568, 0.01264852, 0.0239704, 2.128617e-05, 
    0.07560944, 0.0003945378, 0.00131701, 0.002696525,
  0.01549873, 0.02131854, -8.096014e-06, 0.00266196, 1.100985e-05, 
    1.937302e-05, 0.0001923423, 0.0005578372, 0.0002972808, 0.0003454064, 
    0.0009850791, 0.0002493502, 0.005391991, 0.0004998935, 7.798668e-05, 
    3.503453e-05, 7.894827e-06, 4.954028e-05, 7.982105e-05, 0.0006134247, 
    0.001344518, 0.006620166, 0.02404363, 0.00137437, 8.711852e-08, 
    1.444327e-08, -0.0002125296, 3.481401e-05, 0.003502982,
  0.01081974, 0.04790808, 0.000439427, -0.0002300104, 2.201966e-05, 
    0.0001764307, 0.0005606035, 0.0003678101, 0.0286246, 0.06061198, 
    0.0001483884, 6.586485e-05, 0.001572995, 0.00136767, 0.000819649, 
    1.64915e-05, 5.096273e-06, 8.670251e-06, 4.758845e-06, 7.326665e-06, 
    0.0007198701, 0.01922213, 0.02583573, 0.03297696, 0.03289891, 
    8.869143e-05, 2.652063e-05, 0.000349469, 0.001122958,
  0.1180803, 0.01340267, 0.0003749004, 0.1912645, -9.016425e-07, 6.31561e-07, 
    0.03207821, 2.201899e-06, -0.002234968, 2.390266e-06, 2.427781e-06, 
    0.0001982866, 0.0007098458, 0.0003395428, 0.0002729621, 0.002501211, 
    0.002287986, 0.00540412, 0.003132241, 0.001244151, 0.003888919, 
    0.00145206, 0.2300706, 0.03454095, 0.0001708002, 0.00117796, 0.00218805, 
    0.002584993, 0.04695446,
  1.046612e-07, 1.154241e-10, 1.878693e-10, -4.775371e-10, 2.224857e-08, 
    7.789314e-05, 0.005202638, 0.00033597, 0.165887, -0.0006306556, 
    0.001432934, 0.0004496932, 4.505686e-05, -2.674971e-06, 2.649039e-05, 
    7.115563e-05, 0.0003518908, 0.001677907, 0.01798579, 0.03491428, 
    0.007850205, 0.02895676, 0.0001929252, -0.001735831, 5.947997e-05, 
    8.803757e-05, 0.002504781, 0.003487439, 1.170259e-07,
  1.281877e-07, -6.391745e-06, 1.114566e-05, -1.55139e-06, 1.310316e-07, 
    4.701651e-09, -0.002853116, 0.1107714, 0.2376961, 0.003722986, 
    0.002132744, 0.001056536, 0.001882334, 0.001409182, 0.001833631, 
    0.0007427509, 0.002238017, 0.005111984, 0.01622188, 0.08568668, 
    9.317701e-07, 0.01913831, 0.04493248, 0.0002371408, 0.0003072536, 
    0.0004230813, 0.001364097, 0.01068138, 0.002222427,
  -0.0001213426, -0.000345925, -0.0003395222, 0.1886565, -4.466375e-05, 
    3.990785e-11, -4.222233e-07, 1.339765e-06, -5.396441e-06, 0.008700059, 
    0.2564796, 0.1953751, 0.3886872, 0.2192048, 0.1722461, 0.286761, 
    0.1172651, 0.05014636, 0.04737808, 0.0002257912, -0.0001148244, 
    0.001100916, 0.009944619, 0.04004722, 0.006108129, 0.0134062, 
    0.004342732, 0.01609456, 0.07194415,
  0.0657567, 0.03348245, 0.02288717, 0.003064779, -9.688702e-07, 
    1.523582e-05, 0.001593035, 0.1695349, 0.03247335, 0.005605727, 
    0.07640129, 0.1635723, 0.500808, 0.457817, 0.4023402, 0.2682071, 
    0.2753415, 0.1616576, 0.06407866, 0.02976249, 0.005469401, -9.429608e-06, 
    0.04814642, 0.07642603, 0.1951486, 0.2677092, 0.1558073, 0.1635051, 
    0.04472065,
  0.09139559, 0.01528429, 0.001537448, 0.01219481, 0.05850838, 0.06497072, 
    0.109627, 0.1126717, 0.1424109, 0.1047922, 0.05846587, 0.1531975, 
    0.3229937, 0.1861966, 0.3492835, 0.3593968, 0.1699127, 0.1865637, 
    0.1016157, 0.02863265, 0.00464728, 0.06313977, 0.1726369, 0.1089025, 
    0.1164782, 0.152392, 0.123224, 0.1603977, 0.1755205,
  0.2659776, 0.1747615, 0.2305582, 0.1010905, 0.2969962, 0.5329599, 
    0.05707375, 0.01616574, 0.04773021, 0.02253462, 0.0745846, 0.1432364, 
    0.222383, 0.2411757, 0.3044652, 0.2677439, 0.1397602, 0.2983676, 
    0.2094107, 0.1279118, 0.09288386, 0.3005816, 0.1167327, 0.3521221, 
    0.2297025, 0.2153905, 0.1523473, 0.2448617, 0.3173593,
  0.5782069, 0.3518932, 0.3723981, 0.4644617, 0.3464134, 0.4955551, 0.596207, 
    0.659005, 0.6279385, 0.5593383, 0.4679066, 0.457278, 0.4429329, 
    0.4717559, 0.4166838, 0.4451783, 0.4546587, 0.4449654, 0.4106057, 
    0.4036275, 0.3561233, 0.1916557, 0.1145167, 0.3220415, 0.2161426, 
    0.1395693, 0.2278906, 0.4615752, 0.5741177,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0003189293, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, -0.0001276253, 0, 0, 0, 0.0002736177, 0.002610958, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, -1.989404e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0002370221, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -3.627659e-07, 0.0002432738, 0, 0, 0, 0, 
    0, -3.426955e-06, 0, 0, -3.454027e-05, -3.012281e-05, 0, 0, 0, 0, 0, 
    -2.218017e-05,
  0, 0, 0, 0, 0, 0, -5.296645e-05, 0, 0, 0, 0.0009332126, 0.004437122, 
    -8.361066e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0002854862, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, -0.0001233017, 0, 0, 0, 0, 0, 0, 0.0004877745, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, -8.46496e-06, 0, 0, 0, 0.001415581, 0, -2.337635e-05, 
    0.004096721, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0.0001818172, 0, 0, 0, 0, 0, 0, 0, 0, 0.0004967339, 0.002228575, 
    -0.0001232411, 0, 0.0007935438, 0.0002693002, -7.569623e-06, 
    -6.605864e-05, 0, 0.0003391352, -7.467179e-05, -3.899561e-05, 
    -4.2552e-06, 0, -2.191227e-05, 0, 0.003263406, 0.0002124966,
  0, 0, 0, 0, 0, -1.366042e-05, 0.001171925, 0, 0.0009017009, 0, 0.001606328, 
    0.01212407, 8.389082e-05, 0, 0, 0, 0, 0, 0, 0, 0, -1.975131e-05, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0.0004063836, -0.0001890663, 0, 0.001052102, 
    -5.438351e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, -1.204163e-05, 0.001738098, 0, 0, 0, -1.98015e-07, 0, 
    -5.947681e-06, 0.0004321328, -5.534468e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0,
  0, 0, 0, 0, 0, 5.962342e-05, 0, 0, 0, 0.004385331, 0, -5.363559e-05, 
    0.01890539, -4.370258e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0.003806117, 0, 0, 0, 0, 0, 0, 0, 0, 0.001403772, 0.005849476, 
    0.00286469, -5.119598e-05, 0.003033371, 0.001131109, -1.513925e-05, 
    -0.0001904746, 0, 0.002389373, 0.003601474, 0.0002245685, -1.421919e-05, 
    -5.615969e-05, -0.0002190236, -1.151961e-05, 0.007322912, 0.001761751,
  0, 0, 0, -1.461395e-06, 0.0002392186, -7.625474e-05, 0.007219065, 
    -1.239233e-09, 0.002761136, 0, 0.004095673, 0.02346612, 0.0004972934, 
    0.0009634614, 0, 0, 0, 0, 0, 0, 0.0001534252, -0.0001179234, 
    -2.335468e-05, 0, -1.852685e-07, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0.002339099, 0.000615367, -1.739236e-05, 0.003675967, 
    0.001858193, -2.437779e-06, -4.113736e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, -7.072874e-06, 0, 0, -1.595827e-06, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.931195e-07, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -1.521692e-07, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, -1.204163e-05, 0.004850963, 0, 0, 0, -1.98015e-07, 
    -3.092267e-05, -7.296885e-05, 0.0006152716, -1.343702e-05, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0.003933013, 0, 9.429435e-05, 0.0001895866, 0.008478956, 
    -4.282485e-05, -2.120586e-05, 0.03333626, 6.174092e-05, 0, -1.344526e-06, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0.004746581, -1.251522e-06, 0, 0, 0, 0, 0, 0, -2.439225e-05, 
    0.00320335, 0.02100506, 0.008594606, -0.0001214943, 0.007352732, 
    0.002506363, 5.457134e-05, 6.91934e-05, 0, 0.006748445, 0.006210878, 
    0.0008655984, -3.896051e-05, -8.650965e-05, -0.0002127788, -9.181879e-05, 
    0.01183879, 0.007036389,
  0, 0, 0, 0.0002305084, 0.0003449336, -0.0001029104, 0.01442938, 
    -2.17858e-05, 0.00569069, 0, 0.01240945, 0.04132438, 0.002052475, 
    0.006215124, 0, 0, 0, 0, 0, 0, 0.0004050588, 0.0008707627, -3.532159e-05, 
    0, -1.325181e-05, 0, 0, 0, 0,
  0, 0, 0, 0, -1.40921e-08, -8.816309e-06, 0.00369811, 0.004552383, 
    0.0005823159, 0.01259294, 0.01073118, -2.973354e-05, -0.000157236, 
    0.001811637, 0.000276023, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0001611703, 0.0009904961, -1.854668e-06, 
    -4.347356e-05, -1.204539e-05, 0.001342478, -3.194176e-05, 0, 0, 0, 0, 0, 
    -2.577013e-05, -0.0001175643, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -3.805062e-05, -2.196552e-05, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, -1.692852e-06, -6.093385e-05, 0.0005287575, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2.147278e-05, 0, 0, 0, 
    0, 0, 0, 0, -6.670797e-07, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0001079901, 
    -1.147765e-07, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, -4.177957e-07, 7.665619e-05, -9.980973e-05, 0.0148891, 0, 0, 0, 
    -0.0001296274, -7.550243e-05, 0.0001534913, 0.001016615, -2.096953e-05, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, -2.109051e-06, 0, 0, 0.00829991, -4.571861e-05, 9.508995e-05, 
    0.000388178, 0.01843463, -1.010774e-05, 0.0006072574, 0.04469664, 
    0.001928244, 7.303923e-06, -1.155828e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0,
  0.0008499934, 0.001316279, 0.01098291, 0.0005583882, 0, -1.619632e-06, 0, 
    0.0003167357, 8.982826e-06, -4.07947e-05, 1.208298e-05, 0.00427568, 
    0.04556783, 0.01553976, -0.0001137125, 0.01647941, 0.00803666, 
    0.0004166311, 0.002566998, 0.0005294397, 0.01111055, 0.01284125, 
    0.002517974, 8.374333e-06, -0.0002017409, -9.787347e-05, -0.0002123583, 
    0.01453895, 0.01691449,
  0, 0, 0, 0.002270184, 0.004559128, 0.0008531929, 0.03437382, 0.001403065, 
    0.009854834, 0.0005734381, 0.03540093, 0.05694156, 0.01155101, 
    0.01349788, -4.1796e-06, 0, 0, 0, 0, 0, 0.0007868175, 0.003231976, 
    -3.805099e-05, 0, -3.723175e-05, 0, 0, 0, 0,
  0, 0, 0, 0, 2.628361e-06, -3.121133e-05, 0.009166763, 0.007002217, 
    0.008297989, 0.02098192, 0.03621236, 0.0001325255, 0.00077356, 
    0.003096809, 0.0006810069, 0, 0, 0, 0, 0, 0, 0, 0, 0, -4.57215e-06, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, -3.726685e-05, 0.003794518, 0.006626804, 
    0.00603862, 0.0003788462, 0.001652649, 0.004689252, -5.893426e-05, 0, 0, 
    0, 0, 0, 8.337587e-05, 0.003932909, 0, 5.568992e-05, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, -9.014039e-06, -0.0003891536, -0.000125662, 0, 
    -2.384196e-07, 0, 0, 0, 0, 0, 0, 0, 3.935921e-05, 0.004380444, 
    0.002014096, -1.697905e-08, -1.246066e-05, -8.721036e-06, -4.544175e-05, 0,
  0, 0, -4.357877e-06, 0, 0, 0, 0, 0, 0, 0, 0, -3.190386e-06, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 8.727704e-06, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0001247091, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -6.941761e-05, 0, 
    -7.142796e-06, 2.000811e-05, 0, 0, 0, 0, -2.223432e-05, -6.796319e-05, 
    -5.594465e-05, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.006304761, 0.0002027811, 
    2.670748e-07, -6.45837e-06, 0, 0, 0, 0, 0.001120214, 0.002844317, 
    -1.093867e-08, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4.56309e-06, 0, 9.745677e-06, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, -8.247403e-06, 5.851777e-05, 0.0005020108, 0.02829837, 
    0.0001060831, 0, -2.607035e-08, 0.004374191, -0.0002419529, 0.0004346996, 
    0.004093439, -6.598144e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 1.522691e-05, 0, 0, 0.01572085, -0.0003877064, 0.0007819839, 
    0.001504335, 0.0285574, 0.0006613435, 0.003691625, 0.062995, 0.00903082, 
    -8.382065e-06, 1.353359e-05, 0, 0, 0, 0, 0, 0, 0, 1.898679e-05, 
    -2.259877e-05, 0, 0, 0, -9.15442e-06,
  0.002344498, 0.002109458, 0.01845891, 0.001389175, 0, -5.731073e-06, 
    0.0002105022, 0.0005659808, 0.0002582691, 0.0001248538, 0.001176841, 
    0.007724806, 0.07606573, 0.02637182, 0.000888286, 0.02752621, 0.02137465, 
    0.001846156, 0.008398887, 0.002390119, 0.02362964, 0.0279914, 0.01753213, 
    0.0002172708, -5.550538e-05, 0.002168583, 8.285451e-06, 0.02736784, 
    0.02736839,
  0, -2.104019e-09, -6.475401e-11, 0.01299602, 0.01071544, 0.01575566, 
    0.07676837, 0.004589782, 0.01626863, 0.00323041, 0.07517926, 0.08528116, 
    0.02580977, 0.02431865, 0.0003979543, 0, 0, 0, 0, 0.003635295, 
    0.008191403, 0.01038853, 0.0003478324, -1.913213e-05, 0.0001185278, 0, 0, 
    0, 0,
  0, 0, 0, -6.391064e-11, 0.0009055862, 0.001377223, 0.01976899, 0.009745033, 
    0.01532821, 0.04198844, 0.05229673, 0.004229643, 0.008459798, 
    0.006546457, 0.00611937, 0, 0, 0, 0, -5.873908e-05, -2.459103e-05, 0, 
    0.0002359277, 6.76722e-05, 8.318092e-05, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0.0002146319, 0.007339189, 0.01236616, 0.01057496, 
    0.008148362, 0.01241958, 0.0148144, -0.0003190635, 0, -6.088123e-06, 
    -2.129594e-08, 0, -1.032151e-05, 0.00417544, 0.007770297, -6.010026e-06, 
    0.0008116015, -3.128163e-05, 0, 0.00161421, 0,
  0.0007607659, -4.511431e-06, 0, 0, 0, 0, 0, 0, 0.0005441883, 0.000649463, 
    0.005753193, 0.0002820065, 0.0006953019, 0.004639525, -4.796678e-05, 
    -5.509391e-06, -2.014678e-08, 0, 0, 0, -2.134346e-07, -1.140446e-05, 
    0.02116923, 0.008652858, 0.005741573, -0.0002757575, -7.811313e-05, 
    -0.0001441199, -1.516495e-05,
  0, 0, 7.073847e-06, 0, -2.319807e-06, 0, 0, 0, -4.753651e-06, 0.001062658, 
    -0.0001798256, 0.006272113, 0, -2.254516e-06, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0002171151, -3.525455e-06, -2.103952e-05, -1.264642e-05, 4.641914e-05, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -4.9641e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0.0005600011, 0.000156852, -3.037241e-06, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, -3.188583e-05, 0, 0.0002664997, 0, 0, 0, 0.0002599332, 
    0, 0,
  -6.21302e-05, 0, 0, 0.0001533406, 7.084804e-06, -1.0248e-05, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.000622101, -4.911407e-05, 0.001932229, -2.039183e-05, 
    6.384838e-05, 0.001019348, 0.0006536924, 0, 0, 0, 0.005768114, 
    0.001889068, 0.0005472246, 0,
  0, 0, 0, 0, 0, 0, 0, 0, -2.363653e-10, 0, 0, 0, 0, 0, 3.645507e-07, 
    -9.034143e-05, 0.0171599, 0.005301883, 0.0008529955, 0.001513853, 0, 0, 
    0, 0, 0.005023094, 0.02008925, -1.294003e-06, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -6.404428e-06, -8.781381e-07, 
    0.004961599, -1.659171e-07, 0.002992552, 0, 0, 0, -7.74851e-06, 0, 0, 0, 
    -1.604861e-07, 0, 0, 0,
  0, 0, 0, 0, -1.309252e-05, 4.370717e-05, 0.003961864, 0.06101735, 
    -8.774857e-06, 7.280476e-05, -8.754934e-05, 0.01701731, 0.0002674592, 
    0.004577743, 0.008976619, 0.000147797, 6.108066e-09, 0, 0, 0, 
    -7.025197e-10, -5.744026e-10, -1.142317e-10, -3.91675e-06, 9.89773e-10, 
    5.683149e-07, 0, -1.355606e-09, 0,
  -3.495672e-08, 0.0002911048, 0.0003999472, 0, -6.53629e-10, 0.02636519, 
    0.004216527, 0.007699802, 0.007487059, 0.04587008, 0.005928379, 
    0.01164078, 0.09520397, 0.029553, 0.0006964777, 0.0004457255, 0, 0, 
    -1.014328e-07, 0, -2.301715e-05, -1.511134e-06, 1.029211e-06, 
    -4.113156e-05, 5.625529e-05, -2.994316e-05, -1.17674e-06, 0, 8.496058e-06,
  0.004198816, 0.00537512, 0.02665804, 0.008468867, 5.388098e-05, 
    -7.334244e-05, 0.002486887, 0.01878192, 0.004990606, 0.005878497, 
    0.003306088, 0.0179843, 0.1392708, 0.04068002, 0.01561945, 0.04103428, 
    0.04578357, 0.008650163, 0.01904074, 0.008664276, 0.05224641, 0.04245486, 
    0.06085015, 0.004681496, 0.000563067, 0.007313287, 0.002675779, 
    0.05095991, 0.04707859,
  -8.417966e-08, -1.637512e-06, -3.829207e-05, 0.03443049, 0.04307478, 
    0.09149158, 0.130917, 0.03237768, 0.05748678, 0.01518428, 0.1317284, 
    0.1266771, 0.05460073, 0.04731343, 0.004374088, -8.311301e-06, 0, 0, 0, 
    0.007078578, 0.01051527, 0.03149866, 0.002723176, -0.0001306794, 
    0.004022708, -1.165793e-09, 0, 1.153453e-06, 0,
  0, 0, 0, -2.233867e-06, 0.002604802, 0.004595739, 0.1188679, 0.01352742, 
    0.0266904, 0.09898813, 0.08989356, 0.02617853, 0.01953407, 0.009840533, 
    0.01008989, 0, 0, 0, 0, -9.678332e-05, 0.000160767, 0.0004344392, 
    0.01109362, 0.002541861, 0.0004683592, 0, 0, 0, 0,
  0, 0, 0.001008073, 1.210918e-09, 1.119857e-05, 9.727487e-05, -2.995266e-08, 
    6.998991e-08, 0.005274882, 0.01290429, 0.03570786, 0.0243111, 0.01813423, 
    0.02607736, 0.02517266, 0.00397423, 0.0003368149, 0.001076457, 
    -5.442331e-05, 0, -6.314199e-05, 0.009961295, 0.01050813, 0.002823812, 
    0.004894693, 0.0001451587, -5.037464e-05, 0.007118333, 0,
  0.004213766, 1.121661e-05, 4.145383e-05, 0, 0, 4.146969e-11, 0, 
    0.0004158066, 0.001935776, 0.009894723, 0.01498746, 0.01331263, 
    0.0125887, 0.01295408, -0.0004351791, -1.40658e-05, 0.007510545, 
    8.296892e-05, 0, 0, -4.672581e-06, 0.0009423197, 0.03506519, 0.01773079, 
    0.01669677, 0.001813931, 0.004224753, 0.001056396, 0.001984325,
  5.938891e-05, 0.001395429, 0.001448083, -1.07832e-06, 0.001451883, 
    -5.539522e-05, -8.090678e-05, 0.000494775, 0.0007551229, 0.001276087, 
    -0.0004611249, 0.01765682, 0, -4.917264e-05, -6.525954e-06, 0.0006576843, 
    0, 0, 0, 0, 0, -9.342146e-05, 0.002448687, -9.208101e-06, 0.005478222, 
    0.002991044, 0.001449526, 0, 0,
  0, 0, 0, 0, 0, 0, -7.422464e-06, 0, 0, 0, -4.849616e-05, -8.637708e-05, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0.0009111594, 0.0003754975, 0, -2.276775e-05, 0.001689147, 0.0001382344, 
    -1.611784e-05, -2.598708e-05, -1.135504e-06, 0, 0, 0, 0, 0, 0, 0, 
    -4.826169e-06, 0, 0, 0, 0.002578374, -6.058186e-07, 0.0009407158, 
    -6.40789e-06, 0, 0, 0.0004889165, 0, 0,
  0.0007713826, 0, 0, 0.001835304, 0.00667397, 0.01014438, 9.06697e-05, 0, 0, 
    3.386519e-10, 0, 0, 0, -1.967968e-05, -7.295958e-06, 0.007566699, 
    0.0002306266, 0.01002089, 0.001064996, 0.01485148, 0.00407325, 
    0.002799142, 0, 0, -6.169452e-06, 0.0113604, 0.006434601, 0.004684981, 
    -2.73663e-05,
  0, 0, 0, -2.278888e-10, 0, 3.206793e-10, 3.519596e-07, 0, -1.184751e-06, 
    3.192003e-07, -2.1165e-09, 0, -2.120102e-11, -1.450287e-08, 0.002757863, 
    0.006971669, 0.02794541, 0.01809433, 0.008304759, 0.004449298, 0, 
    -8.847807e-11, 0, -2.218473e-07, 0.01132332, 0.03524306, 0.0003519724, 
    5.027575e-07, 0,
  0, -1.022602e-08, 0, 5.07033e-09, 9.814893e-08, 5.896377e-07, 2.512446e-07, 
    7.660326e-07, -2.492215e-06, 3.015542e-07, 3.610957e-05, -5.06949e-08, 
    -5.358778e-05, 0.001888428, 0.001189057, 0.02076063, 0.005975209, 
    0.007146296, 0, 7.710391e-05, 0, -7.14773e-07, 0, 4.140085e-11, 
    8.40807e-05, -2.027534e-07, -1.298227e-11, 0, 0,
  0, -1.153948e-05, -9.183014e-06, -1.018739e-08, -1.647354e-05, 0.004905454, 
    0.01564646, 0.09694834, 0.00281448, 0.006977509, 0.005894351, 0.06931332, 
    0.01013282, 0.02863512, 0.02747639, 0.003859324, 2.453668e-06, 
    -1.529634e-08, 0, 0, 0.0003482456, -1.475439e-06, 2.271418e-06, 
    0.000144173, 5.17715e-05, -8.175904e-07, -1.470584e-07, 4.3185e-05, 
    -2.711994e-11,
  0.0001702798, 0.004813298, 0.005512323, -4.154549e-07, 4.635055e-07, 
    0.04125156, 0.01976764, 0.0262307, 0.04009651, 0.0803814, 0.09516272, 
    0.1354764, 0.1673237, 0.08093547, 0.03452142, 0.006709215, 0.0007677069, 
    -1.954436e-09, 2.324456e-05, -7.381882e-08, 7.583594e-05, 0.001350749, 
    0.0007102431, -0.0002440223, 0.0008769963, -1.213083e-05, 4.152066e-05, 
    0.0002433108, 0.004516276,
  0.02345029, 0.02764297, 0.06685419, 0.02758677, 0.001250559, 0.01728244, 
    0.2339084, 0.4859846, 0.3807731, 0.2343725, 0.2905758, 0.273027, 
    0.3560461, 0.1206771, 0.1408585, 0.1159343, 0.1074817, 0.04520806, 
    0.03832778, 0.04457454, 0.1304652, 0.1064821, 0.143983, 0.01886011, 
    0.003720151, 0.01923322, 0.007457065, 0.08695862, 0.08429052,
  9.902808e-07, 0.0002013689, 0.01806935, 0.1379665, 0.2022899, 0.2360538, 
    0.3761455, 0.1459673, 0.3208122, 0.1793617, 0.3294455, 0.3280225, 
    0.2534883, 0.1187948, 0.00740466, 0.0008779865, -1.129227e-09, 0, 
    1.992299e-07, 0.01543179, 0.1134949, 0.1256687, 0.03629926, 0.006463256, 
    0.01457937, -3.072669e-05, 7.030484e-05, 0.0008246647, -2.995107e-07,
  5.546873e-06, 0, -1.011358e-07, 0.001358277, 0.01896768, 0.02792969, 
    0.1241078, 0.02585003, 0.03893094, 0.2089216, 0.1638243, 0.1368536, 
    0.1096554, 0.06852244, 0.02141323, 3.846705e-05, 0, -5.497584e-06, 0, 
    -0.0001619036, 0.004142228, 0.0009270856, 0.07863943, 0.006813938, 
    0.005336625, 7.314009e-05, 3.742177e-08, 0, -1.542678e-08,
  2.171105e-05, -1.32524e-09, 0.003983915, 2.750205e-07, 0.001042495, 
    0.002844155, 3.548332e-06, 0.002187091, 0.03108039, 0.03263478, 
    0.1270811, 0.131508, 0.1001967, 0.09050431, 0.06992226, 0.02007046, 
    0.004709819, 0.004199055, -0.0001094159, 0, -5.974459e-06, 0.01945982, 
    0.02197528, 0.01351352, 0.02698968, 0.0001854769, 5.7535e-05, 0.01154581, 0,
  0.007606061, -9.862365e-05, 0.0001587546, -6.415397e-05, 0.0004070538, 
    -3.550291e-05, -2.982332e-05, 0.001503959, 0.01155607, 0.02798313, 
    0.03895089, 0.04285548, 0.04518441, 0.03009227, 0.007430896, 0.0060837, 
    0.02570985, 0.01213171, -7.341492e-06, 0, -9.08457e-05, 0.009710341, 
    0.05687824, 0.03898435, 0.02751432, 0.01661156, 0.01178983, 0.01249344, 
    0.01162642,
  0.005861313, 0.002802942, 0.005025994, 0.001801316, 0.003447606, 
    -0.0001179079, 0.003080937, 0.0006320348, 0.003696541, 0.005431448, 
    0.006579003, 0.02585087, -9.667448e-05, -0.0002978756, 0.0002248935, 
    0.003789292, -8.31559e-06, 0.0002019329, 0, 0, 0, 0.001586511, 
    0.02293502, 1.916501e-05, 0.01325214, 0.006930677, 0.01376251, 
    0.001249752, 0.0003878329,
  0, 0, 0, 0, 0, -2.189201e-05, 0.0007558673, 0.005828068, 0, 0, 
    -0.0001816507, -0.0001799444, 0, 0, 0, 0, -1.297471e-06, 0, 0, 
    0.0001790373, -7.460253e-05, 0.0005308425, 0, 0, 0, 0, 0, 0, 0.0008325417,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, -1.684141e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5.579184e-05, -6.330743e-05, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0.005424412, 0.00225989, -1.058075e-05, -6.320509e-05, 0.00526439, 
    0.002870471, 0.002149517, -2.920057e-05, 0.001991594, 4.829329e-06, 
    -5.415915e-06, 0.00155436, -6.400538e-05, 1.859685e-05, 0.002674947, 
    2.178519e-05, 0.003209432, 0.001999433, -1.713267e-05, -0.0001220369, 
    0.00856681, 0.0006753154, 0.006365424, -0.0001683013, 1.120567e-05, 0, 
    0.002271062, 0, -1.632948e-05,
  0.001111667, 0, -1.812731e-09, 0.006835407, 0.01691677, 0.0171377, 
    0.005381915, -5.661642e-06, 9.809936e-08, 4.504176e-08, 6.356658e-10, 
    -1.912791e-06, 0, 0.0005728411, 0.003355953, 0.01403823, 0.004466335, 
    0.0257882, 0.01308489, 0.05376492, 0.04102608, 0.01498252, 0.00154498, 
    0.002602894, -4.17665e-05, 0.02050998, 0.01625982, 0.01291025, 0.005577252,
  6.713325e-07, 3.57682e-05, 0, -5.274433e-08, -6.192853e-10, 1.337186e-08, 
    3.66005e-05, -2.156873e-10, -3.366989e-05, 0.000126333, 2.534563e-05, 
    -1.549824e-06, 5.010254e-07, 3.200453e-06, 0.00887078, 0.01856988, 
    0.04343116, 0.06243442, 0.04460525, 0.00775417, -0.000141614, 
    -5.412472e-07, 9.357189e-10, 0.0002770908, 0.02010283, 0.05023308, 
    0.007857842, 4.053969e-05, 0.0001036359,
  6.963004e-06, 2.390791e-06, 3.775659e-07, 7.092771e-10, 1.033451e-08, 
    -1.152337e-08, 1.380966e-05, 2.991456e-06, 1.992977e-05, 7.914684e-07, 
    2.86279e-05, 3.23101e-07, -0.0002782761, 0.004477701, 0.007797649, 
    0.04118904, 0.04250128, 0.03052695, 2.575538e-05, 7.310978e-05, 
    5.897043e-08, 0.0002337622, 4.02459e-05, 0.000108308, 0.001601278, 
    -6.365005e-07, 4.131868e-06, 5.509703e-05, 7.31947e-06,
  7.297304e-05, 0.0008289573, 1.463057e-05, -0.000101428, 0.01086299, 
    0.0581232, 0.04449405, 0.1767037, 0.01631886, 0.0191326, 0.01523838, 
    0.08801757, 0.01269966, 0.04526945, 0.02812802, 0.04084674, 0.001071775, 
    0.0003919274, 9.236447e-07, -8.071941e-09, 0.0005234284, 0.0009167605, 
    0.01624439, 0.03474087, 0.008019203, 0.0003245211, 0.00342021, 
    0.006366912, 3.327438e-06,
  0.008442303, 0.3320995, 0.328528, 0.000168742, 0.005398937, 0.1528354, 
    0.2819017, 0.2695789, 0.3529666, 0.2743067, 0.1901028, 0.1745433, 
    0.1739926, 0.07411188, 0.036632, 0.005885332, 0.0001626512, 3.165219e-05, 
    5.265436e-06, 0.01090267, 0.06348527, 0.01338306, 0.06039013, 0.1573791, 
    0.0444856, 0.01659343, 0.05058803, 0.08394339, 0.0354277,
  0.211665, 0.4205181, 0.4222841, 0.05309059, 0.02322962, 0.03654626, 
    0.3013255, 0.4393881, 0.2894511, 0.1543929, 0.228615, 0.2210441, 
    0.3263656, 0.1108465, 0.138879, 0.1484676, 0.1329019, 0.1356956, 
    0.09873941, 0.1307804, 0.220635, 0.1766838, 0.3902481, 0.1523485, 
    0.0926511, 0.1198829, 0.09348892, 0.2173419, 0.3429205,
  4.205725e-06, 0.003898357, 0.01825221, 0.1341179, 0.2279262, 0.2077232, 
    0.326694, 0.1093261, 0.2873946, 0.1296179, 0.2448447, 0.2791544, 
    0.2367147, 0.2795453, 0.19504, 0.05856578, 0.002667439, 1.523504e-05, 
    8.893556e-06, 0.01477476, 0.08200192, 0.2012077, 0.09964041, 0.07493433, 
    0.09109473, 0.03612755, 0.008131608, 0.002438669, 0.0003532503,
  8.902103e-07, 0, -9.063096e-08, 0.002198881, 0.01429288, 0.02308769, 
    0.09254354, 0.05759931, 0.05775576, 0.1731088, 0.136361, 0.1040465, 
    0.07698993, 0.1539898, 0.1899142, 0.01691324, 0.0469049, 0.0005805019, 
    0.0009451111, 0.01937726, 0.09188455, 0.0931344, 0.2269884, 0.1774219, 
    0.09954004, 0.04844669, 0.0005506795, -5.751729e-08, 2.699145e-07,
  0.001975898, -8.023259e-06, 0.006341112, 1.067748e-05, 0.002504905, 
    0.006505453, 0.0003479637, 0.01516532, 0.1022673, 0.08055302, 0.1664975, 
    0.1584308, 0.1355815, 0.2066379, 0.3075671, 0.1693322, 0.1014325, 
    0.07444192, 0.01650278, -8.347249e-05, 0.002715347, 0.06103664, 
    0.09836743, 0.1336102, 0.2009118, 0.05055862, 0.03866884, 0.02878023, 
    0.003627158,
  0.01009958, 0.008452129, 0.0006025832, 0.0006832677, 0.007528414, 
    0.002825367, -0.0001944617, 0.002691806, 0.02483595, 0.0660818, 
    0.1285147, 0.1478295, 0.1809107, 0.1569439, 0.06222009, 0.08917911, 
    0.07676138, 0.03029687, 0.01018143, 0, 0.00146341, 0.03106683, 0.1015809, 
    0.06725632, 0.06254834, 0.06220044, 0.05606576, 0.04146853, 0.02978335,
  0.01310684, 0.006985913, 0.01013401, 0.01031807, 0.004994457, 
    -6.021211e-05, 0.01144277, 0.0009240804, 0.01102135, 0.0119643, 
    0.01847429, 0.03550302, -0.0002473245, 0.009894027, 0.002877005, 
    0.01098506, -0.000475113, 0.008959194, 2.763839e-05, 0.0004375154, 
    -2.785827e-05, 0.009432598, 0.0405335, 0.000184797, 0.02708986, 
    0.01590816, 0.03134086, 0.004311363, 0.007461223,
  -5.374662e-05, 0, 0, 0, 0, 0.005017903, 0.001773867, 0.01072854, 
    -7.609918e-05, -3.219857e-05, 0.002170677, 0.0001622772, -0.0001684, 0, 
    -0.0001411295, 0, -6.324724e-06, 0, 0, 0.002379849, -0.0003697446, 
    0.006111198, 0, 0, 0, 0, -2.867993e-06, -2.378671e-05, 0.004411216,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2.896199e-05, 
    -7.840405e-05, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, -6.461369e-05, -2.766618e-06, 0, 0, -1.26121e-06, -1.350264e-05, 0, 
    0.000664924, 0.0007587769, 0, 0.0012184, 0.000877191, 6.173454e-05, 
    -1.035063e-06, 0, -1.24738e-05, 0.0005418938, 0, 0, 0.0002894463, 0, 
    -6.437507e-06, -1.920281e-05, -3.742266e-06, 0, 0, 0, 0,
  0.01264456, 0.005161592, 0.003992944, 0.002207126, 0.01465311, 0.009632178, 
    0.008795415, 0.005331158, 0.003352239, 0.001099193, -6.433447e-05, 
    0.003226266, -2.538195e-05, 0.004317432, 0.01415937, 7.326467e-05, 
    0.003610595, 0.003704811, -8.829522e-05, -0.0005288691, 0.01718705, 
    0.007955776, 0.02594117, 0.006593603, 0.0003821079, 0.0009722352, 
    0.01020145, 0.005025689, 0.0006032966,
  0.001671631, 0.0001806622, -8.914872e-06, 0.0250677, 0.02433424, 
    0.02309037, 0.01804807, -5.133555e-05, -2.634836e-05, 6.673863e-06, 
    2.960534e-08, -4.591169e-05, -9.449531e-11, 0.001959258, 0.01243902, 
    0.03215602, 0.008782187, 0.06159624, 0.05182283, 0.08694733, 0.08718526, 
    0.04034238, 0.01155197, 0.01699823, 0.005455712, 0.03211223, 0.05121338, 
    0.03361904, 0.01129132,
  0.008774184, 0.008805302, 4.134463e-07, -2.237216e-05, 2.605181e-06, 
    -9.574696e-06, 0.006451028, -3.791903e-10, -3.917083e-07, 0.006708085, 
    0.006173063, -1.648794e-05, 0.0003881025, 0.002447838, 0.0118096, 
    0.03054653, 0.08273978, 0.09261844, 0.07533646, 0.03981704, 0.04892259, 
    0.01506307, 0.004292681, 0.002768284, 0.02794599, 0.1015416, 0.02776252, 
    0.002781242, 0.007853653,
  2.426839e-06, 1.066042e-06, 1.735817e-07, 4.64421e-11, -6.034588e-11, 
    -5.617719e-09, -8.073338e-07, 1.695479e-06, 5.214083e-06, 1.031165e-07, 
    2.570432e-06, 7.122892e-07, -5.779594e-05, 0.004612892, 0.01776074, 
    0.04882551, 0.04419918, 0.02366495, 0.008800207, 0.0001502782, 
    -1.737917e-08, 2.265096e-05, 5.683296e-06, 6.347236e-06, 0.004608944, 
    0.01819702, 0.0009022886, 2.977844e-06, 1.850832e-06,
  2.942389e-05, 2.126291e-05, 5.677341e-05, -1.626392e-05, 0.001876207, 
    0.02334765, 0.04254746, 0.1522897, 0.003600392, 0.005898528, 0.01290391, 
    0.06731696, 0.01497615, 0.04016753, 0.01985886, 0.0285126, 0.0002005328, 
    0.0004568421, 1.233981e-07, 0, 8.067088e-05, 0.0001125408, 0.005596113, 
    0.004070726, 0.005224504, 2.121604e-05, 4.556189e-05, 0.000111646, 
    3.552267e-07,
  0.0001911254, 0.2264563, 0.2061397, 0.001370451, 0.001533596, 0.1176308, 
    0.180062, 0.2087511, 0.2918726, 0.2426882, 0.1417671, 0.1366654, 
    0.1676837, 0.06937612, 0.02294717, 0.004224653, 3.353776e-05, 
    4.314795e-06, 7.003222e-06, 0.001649566, 0.01129091, 0.014418, 
    0.03241739, 0.1173146, 0.02672143, 0.007672106, 0.02972401, 0.05257113, 
    0.01745847,
  0.1732695, 0.382699, 0.3567064, 0.2092224, 0.01084308, 0.008021884, 
    0.1644104, 0.3553742, 0.2078435, 0.08199296, 0.1359265, 0.1786952, 
    0.281673, 0.08568212, 0.1039738, 0.1154698, 0.08989111, 0.09127019, 
    0.05718389, 0.07111257, 0.1613243, 0.1446461, 0.3351971, 0.09219618, 
    0.05519422, 0.08234424, 0.06672814, 0.1742807, 0.2895563,
  4.597904e-05, 0.002330364, 0.01208668, 0.1330671, 0.244671, 0.1742809, 
    0.2861131, 0.09717894, 0.2616105, 0.1086609, 0.2145995, 0.2644814, 
    0.1865266, 0.1878921, 0.1382204, 0.02892573, -2.169369e-05, 4.320038e-06, 
    -5.335952e-05, 0.009458093, 0.05928129, 0.1488449, 0.06709088, 
    0.04316212, 0.05791922, 0.019192, 0.01009241, 0.0003469334, 0.0009233612,
  3.696869e-08, 0, -7.512905e-09, 0.002058587, 0.01221702, 0.01715513, 
    0.07234675, 0.1263663, 0.1139731, 0.1563251, 0.1318544, 0.07744718, 
    0.05362936, 0.1253518, 0.1768816, 0.02600947, 0.09302128, 0.01132354, 
    2.244751e-05, 0.009431764, 0.1682392, 0.04769998, 0.1494846, 0.1379976, 
    0.06941971, 0.03553664, -3.746981e-05, 3.157342e-05, -9.010663e-09,
  0.05381472, 0.007781905, 0.009336654, -9.676398e-07, 0.005348106, 
    0.01915126, 0.002342529, 0.02664643, 0.1482018, 0.1223668, 0.1710573, 
    0.1615153, 0.1332746, 0.1789322, 0.3084446, 0.2957106, 0.1838232, 
    0.1597311, 0.03398314, 0.002873673, 0.06135536, 0.09355511, 0.1480793, 
    0.09616158, 0.1883273, 0.06263497, 0.07555661, 0.07411315, 0.03573659,
  0.1383031, 0.04138316, 0.01824025, 0.009633479, 0.03538284, 0.02539278, 
    0.02302549, 0.004160226, 0.04495029, 0.1187644, 0.2118097, 0.2138588, 
    0.2130387, 0.2057588, 0.1804694, 0.1246501, 0.1200245, 0.127795, 
    0.06554785, -1.504322e-05, 0.02405509, 0.1175351, 0.1293734, 0.1613106, 
    0.1401082, 0.1558517, 0.1396035, 0.1728782, 0.1366463,
  0.08943018, 0.01714385, 0.01474307, 0.01473286, 0.007348871, 0.01475403, 
    0.03361514, 0.008967564, 0.0205135, 0.08328464, 0.1121339, 0.09870166, 
    0.01496268, 0.08389761, 0.109511, 0.1390043, 0.03652163, 0.05067529, 
    0.000392566, 0.0155328, 0.003673234, 0.03541997, 0.07294191, 0.005729061, 
    0.06678391, 0.05123838, 0.0530262, 0.0413284, 0.03804258,
  -0.0003269112, -2.872435e-05, 2.467658e-06, -8.961887e-07, 0, 0.008891834, 
    0.01633499, 0.01799048, 0.0026813, 0.01721523, 0.04350627, 0.002148446, 
    0.01444318, 0.005712075, 0.001086151, 0.0005054316, 0.002038043, 
    -1.477447e-05, -0.0001927184, 0.007376777, 0.004066667, 0.01097867, 0, 0, 
    -6.240435e-08, -6.945442e-09, -5.436686e-05, 0.005822722, 0.01115979,
  0, 0, -5.801114e-07, 0.0001768057, 2.011526e-07, 0, 0, 0, -5.0621e-07, 0, 
    3.295087e-07, 8.37147e-08, 0, 0, 0, 0, 0, 0, 0, 0, 0.0003950524, 
    0.003436489, -1.268036e-05, -1.189288e-07, -8.462742e-06, -1.915525e-06, 
    0, -5.665139e-08, 3.571549e-08,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0001804234, -6.55346e-05, 0, 
    -4.404556e-05, 0, -5.209668e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0.002316408, -5.245512e-06, 0, 0, 3.572686e-05, 0.0003282294, 
    5.688963e-05, 0.001654798, 0.003683367, -7.973632e-05, 0.001441767, 
    0.001207465, 0.006152862, 0.002098015, 0.0005458244, -7.208662e-05, 
    0.003158644, 0, 0, 0.004824418, 6.87101e-05, -4.992927e-05, 0.0003437722, 
    0.001102487, 0.0005557665, -2.468856e-05, -2.335484e-06, 0,
  0.02267619, 0.008873777, 0.02257149, 0.00622442, 0.02435272, 0.02415805, 
    0.01492906, 0.009199358, 0.008130791, 0.005700244, 0.007491674, 
    0.008787801, 0.004060952, 0.02348227, 0.04670573, 0.004902948, 0.0106774, 
    0.01328028, 0.005996025, 0.00124127, 0.02981902, 0.02198402, 0.05369898, 
    0.03169488, 0.00862345, 0.02108941, 0.01549604, 0.01174951, 0.01184588,
  0.01026356, 0.03711029, 0.02411394, 0.06949598, 0.04721304, 0.04399623, 
    0.04585201, 0.01035937, 0.003004199, 0.000113897, 0.0001991479, 
    0.0007399236, -6.590357e-05, 0.01097842, 0.02546653, 0.07006702, 
    0.04698132, 0.1080118, 0.07574487, 0.1303558, 0.1414009, 0.1082064, 
    0.07199633, 0.03783127, 0.05045009, 0.1083651, 0.1403203, 0.1108044, 
    0.04275927,
  0.005030856, 0.003765854, -4.008392e-05, -5.337547e-06, 0.0007058599, 
    0.006976208, 0.01357785, -3.808444e-12, 0.0001684034, 0.01138253, 
    0.009374458, 0.01062665, 0.01148739, 0.001901538, 0.01806493, 0.04493793, 
    0.1183546, 0.1359978, 0.08940306, 0.08304028, 0.06478469, 0.05179851, 
    0.03261172, 0.01117255, 0.03882782, 0.1157856, 0.04649676, 0.01693412, 
    0.008406741,
  1.049179e-06, 1.825549e-06, 1.194008e-07, 3.537627e-11, -3.037183e-09, 
    3.256019e-08, 5.550985e-08, -2.548036e-06, 0.00110135, 4.449758e-08, 
    4.729021e-06, 5.228126e-07, 1.47677e-07, 0.005610768, 0.01580891, 
    0.03794141, 0.03343572, 0.01714161, 0.008912717, 1.913959e-05, 
    -2.24828e-09, 1.566271e-06, 1.817927e-06, 1.243083e-06, 0.007770999, 
    0.03979573, 3.698467e-05, 5.075859e-07, 2.191856e-07,
  1.344433e-05, 9.523089e-06, 4.532987e-06, 1.103685e-05, 7.983879e-06, 
    0.007146444, 0.03005011, 0.1363533, 0.003173212, 0.001937995, 
    0.008693069, 0.07010857, 0.02184555, 0.03780043, 0.0204762, 0.02616305, 
    0.0008803117, 0.0001403902, -2.08535e-09, 0, 2.058757e-05, 3.684392e-06, 
    9.205836e-05, 0.0005290679, -3.128091e-05, 3.265978e-06, 1.145835e-06, 
    4.708627e-06, 1.840792e-07,
  -0.0001474207, 0.1222466, 0.1082582, 0.003162676, 0.000502116, 0.08809459, 
    0.1081977, 0.1650769, 0.2544084, 0.2179834, 0.09808957, 0.1403575, 
    0.1718059, 0.0731927, 0.01983079, 0.004233434, 3.541177e-05, 
    2.139094e-06, 4.192311e-06, 2.298989e-05, 0.0002566967, 0.005050411, 
    0.02778043, 0.0794395, 0.02278621, 0.003862977, 0.001840231, 0.03251898, 
    0.013701,
  0.1699101, 0.3827646, 0.3291216, 0.1830905, 0.001567189, 0.0006911115, 
    0.1068706, 0.208278, 0.1735485, 0.04919092, 0.09013875, 0.1630173, 
    0.2714438, 0.09763472, 0.09447426, 0.1111001, 0.08702082, 0.07826279, 
    0.04780573, 0.04694624, 0.1429475, 0.1349684, 0.2928866, 0.07240205, 
    0.05719548, 0.07070541, 0.06304664, 0.1588722, 0.2653473,
  4.088998e-05, 0.00227904, 0.01507062, 0.132187, 0.2222642, 0.1810299, 
    0.2681352, 0.07231269, 0.2587953, 0.07825901, 0.1951712, 0.2537754, 
    0.1616334, 0.1503794, 0.108129, 0.02237426, -9.409197e-06, 1.742262e-06, 
    -1.703709e-05, 0.007875706, 0.05151907, 0.1180079, 0.05405362, 
    0.03075598, 0.04110308, 0.01288337, 0.009672662, 0.0002139807, 0.001111827,
  5.976357e-08, 0, -4.324558e-08, 0.002082259, 0.01116804, 0.01742044, 
    0.05786711, 0.1974323, 0.1131059, 0.1261782, 0.1341943, 0.04604099, 
    0.04802599, 0.1085154, 0.1434345, 0.01593544, 0.05588474, 0.002571922, 
    1.423255e-05, 0.008597208, 0.1097629, 0.0268247, 0.1205728, 0.133154, 
    0.06541528, 0.02283954, 1.725404e-05, 7.378468e-06, -1.639471e-06,
  0.05370581, 0.0181102, 0.02272999, 5.521185e-05, 0.006887858, 0.02007012, 
    0.01727391, 0.04076009, 0.1672064, 0.1401149, 0.1769012, 0.1334062, 
    0.1219474, 0.1659556, 0.270867, 0.2776218, 0.1762581, 0.146206, 
    0.02980513, 0.006296778, 0.06689687, 0.08365438, 0.1206985, 0.06743313, 
    0.1394269, 0.04950526, 0.05857348, 0.06590894, 0.03206357,
  0.2021183, 0.1347843, 0.127382, 0.09259865, 0.1402698, 0.1239371, 
    0.08354816, 0.02474497, 0.09491029, 0.231783, 0.2192335, 0.1593749, 
    0.1906894, 0.1878914, 0.1822441, 0.1240382, 0.1169085, 0.1385633, 
    0.080474, 0.0409563, 0.08505818, 0.1364218, 0.1387773, 0.1386377, 
    0.1281808, 0.1590749, 0.1430725, 0.2178908, 0.2011036,
  0.2316586, 0.1984161, 0.1548237, 0.09185632, 0.08256169, 0.1004393, 
    0.1279729, 0.1177488, 0.1134266, 0.145088, 0.1512825, 0.1534044, 
    0.04603515, 0.2402056, 0.1491225, 0.195837, 0.1227374, 0.1628303, 
    0.02448875, 0.09526853, 0.05845111, 0.1074726, 0.1272367, 0.05952777, 
    0.1651066, 0.1092052, 0.1336941, 0.06526686, 0.1152689,
  0.07871147, 0.06777018, 0.01247534, 0.003955528, -0.0003409458, 0.02195058, 
    0.03652325, 0.08113052, 0.07861116, 0.07753536, 0.1475451, 0.0596425, 
    0.1650666, 0.114122, 0.1135478, 0.08125664, 0.04765154, 0.00713715, 
    0.007902524, 0.07694335, 0.0465367, 0.09181678, 0.03728562, -0.002792397, 
    0.05365312, -0.0001043684, 0.001300607, 0.1393825, 0.1261836,
  0.004561929, 0.02015896, 0.02541464, 0.04599505, 0.03768561, 0.03721803, 
    0.02912603, 0.03425574, 0.03789644, 0.0349574, 0.02617661, 0.009961677, 
    -0.0007381635, 0.0001536841, -4.262011e-05, 2.558602e-06, -2.382136e-06, 
    0, -1.180102e-08, 6.206989e-07, 0.0003184838, 0.01165081, 0.000972409, 
    -0.0004364192, -0.001173078, 7.962295e-05, -0.0006939247, 0.005882825, 
    0.0005861109,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.00149894, 0.00114733, 0, 
    -0.000256196, 0.003524523, 0.0007413218, 0.0008461887, 0, 0.0006636583, 
    -0.0003138113, 0, 0, 0, 0, 0,
  0.006602264, 0.004946789, 5.754493e-05, -1.719199e-07, 0, 0.0008873526, 
    0.007441835, 0.002463446, 0.004493315, 0.004543996, 0.005551777, 
    0.005376486, 0.00356446, 0.01544206, 0.02596588, 0.04156218, 0.01941897, 
    0.008639846, 0.01032458, 0.01791432, 0.03348422, 0.02232699, 0.004868253, 
    0.004839777, 0.01433505, 0.01436438, 1.977622e-05, 0.003585586, 
    0.0002029029,
  0.03041862, 0.01109526, 0.03905138, 0.02740286, 0.05458903, 0.07235049, 
    0.06514928, 0.03101253, 0.03895206, 0.02119432, 0.0354449, 0.02148322, 
    0.01559435, 0.04006399, 0.107534, 0.0353501, 0.034176, 0.02222819, 
    0.05119074, 0.01323819, 0.04907969, 0.04613118, 0.09491412, 0.06716992, 
    0.06876986, 0.09110051, 0.07146201, 0.04434795, 0.0340451,
  0.1193919, 0.1095709, 0.07547615, 0.1679234, 0.07375581, 0.06831553, 
    0.08562801, 0.03191721, 0.02442511, 0.007535968, 0.01599036, 0.05075981, 
    0.02413048, 0.05607882, 0.03803095, 0.1320176, 0.06205625, 0.1415546, 
    0.1416471, 0.2075709, 0.1702217, 0.1759039, 0.135374, 0.0603492, 
    0.1470067, 0.1121835, 0.1962979, 0.1620112, 0.1436657,
  8.583449e-05, 0.000219277, -1.763912e-05, 0.000367426, 0.001495171, 
    0.01369044, 0.01130163, -6.97324e-10, 0.001214282, 0.0226032, 0.01675061, 
    0.009767241, 0.01382617, 0.003285612, 0.02210527, 0.04028103, 0.1201856, 
    0.1209103, 0.07744456, 0.09354934, 0.06784572, 0.04545465, 0.01486027, 
    0.009012531, 0.0374728, 0.1106114, 0.06416894, 0.01571082, 0.00280101,
  1.298544e-07, 6.419215e-07, 6.65658e-08, 0, 5.70899e-08, 1.587483e-07, 
    1.080006e-06, 0.001945978, 0.01072705, -4.604987e-07, 7.04226e-05, 
    6.286486e-07, -2.433948e-06, 0.01345685, 0.01508851, 0.03287906, 
    0.02258548, 0.0103345, 0.008837378, 1.931163e-06, -3.550132e-10, 
    -5.101419e-07, 1.758346e-07, 1.446033e-07, 0.008786426, 0.01543059, 
    1.239695e-06, 2.039782e-07, 2.50663e-07,
  6.906959e-06, 5.568785e-06, 3.437079e-06, 1.257357e-05, -0.0001598029, 
    0.004712599, 0.03951912, 0.1394811, 0.002833621, 0.001875271, 
    0.006245975, 0.06719757, 0.04003806, 0.03991928, 0.02509161, 0.02132364, 
    0.0003636088, 4.545419e-05, 1.303546e-09, 0, 2.948222e-06, 4.015291e-07, 
    7.633224e-07, 0.001010913, -7.407285e-05, 2.133329e-07, 1.006012e-07, 
    3.306888e-08, 2.696252e-07,
  0.00209728, 0.04278641, 0.06164714, 0.001634743, 0.001084025, 0.06487358, 
    0.07459801, 0.1139012, 0.2123403, 0.2044888, 0.06504448, 0.1396266, 
    0.1775704, 0.06970911, 0.02206597, 0.002670377, 8.425654e-05, 
    1.363512e-07, 2.605001e-06, 7.35199e-06, 2.324168e-05, 0.002398244, 
    0.012066, 0.04969976, 0.01310007, 0.002876984, -4.555031e-05, 
    0.008430369, 0.02263236,
  0.1552123, 0.3426814, 0.2720778, 0.173484, 0.0002075568, 0.0006826747, 
    0.08187136, 0.09955608, 0.1562959, 0.03887749, 0.06621521, 0.1324169, 
    0.2495963, 0.08904381, 0.06943568, 0.1018767, 0.07827293, 0.05759596, 
    0.05016294, 0.03154838, 0.1484783, 0.1163419, 0.2165866, 0.04647464, 
    0.04634771, 0.05588467, 0.06357501, 0.1397387, 0.2407334,
  0.0001538979, 0.004671345, 0.01416242, 0.1334376, 0.1913306, 0.1801573, 
    0.2585048, 0.04960376, 0.2491753, 0.05592963, 0.1775862, 0.2256352, 
    0.1416189, 0.1192568, 0.08436357, 0.01241498, 2.479436e-06, 1.300717e-06, 
    -7.373803e-06, 0.008693366, 0.04451852, 0.09472102, 0.03409306, 
    0.01645552, 0.0257457, 0.01033813, 0.00343797, 9.764456e-05, 0.001929521,
  -2.978344e-11, -5.085902e-12, -3.986597e-09, 0.004162814, 0.006790408, 
    0.02196339, 0.04787157, 0.1942314, 0.1188506, 0.09149717, 0.1214316, 
    0.03157194, 0.0449692, 0.09015486, 0.1335222, 0.01137371, 0.04107183, 
    0.002002652, 5.975338e-06, 0.01334412, 0.07844808, 0.01278829, 
    0.08373401, 0.1292623, 0.05099702, 0.01764034, 6.04786e-06, 7.726823e-07, 
    -4.591041e-06,
  0.04282233, 0.02488986, 0.01991583, 0.0001836464, 0.008317111, 0.02576971, 
    0.02298097, 0.04888284, 0.1769447, 0.1407566, 0.1939425, 0.1098953, 
    0.1416052, 0.1589055, 0.2476894, 0.2678388, 0.1567119, 0.1244029, 
    0.03009043, 0.005824932, 0.04365207, 0.08466711, 0.09478379, 0.05625524, 
    0.1149527, 0.0399229, 0.05044799, 0.05864089, 0.01990373,
  0.1842589, 0.1038859, 0.1002816, 0.09498417, 0.1319938, 0.1210963, 
    0.09305994, 0.06637594, 0.1657708, 0.2399288, 0.1978961, 0.1322158, 
    0.1681932, 0.1695124, 0.1578025, 0.1184658, 0.1143797, 0.1309269, 
    0.07551839, 0.07349315, 0.09038097, 0.1370094, 0.1289589, 0.1251425, 
    0.1037073, 0.1321386, 0.137197, 0.196924, 0.1817441,
  0.2338909, 0.1854222, 0.181666, 0.1641048, 0.1275974, 0.1320459, 0.2670952, 
    0.1735425, 0.1715162, 0.2180247, 0.1968277, 0.1776952, 0.1078471, 
    0.2314032, 0.1376896, 0.2255288, 0.09810455, 0.2087765, 0.1771811, 
    0.1951746, 0.0825704, 0.1443931, 0.1286594, 0.09371319, 0.2357979, 
    0.1877674, 0.146121, 0.1451917, 0.1877698,
  0.1397152, 0.124821, 0.09808719, 0.1119033, 0.1484581, 0.1275488, 
    0.1258121, 0.2572165, 0.1833223, 0.1104434, 0.1482085, 0.09969529, 
    0.2139917, 0.2104435, 0.2083569, 0.1046423, 0.1018132, 0.1264224, 
    0.1533302, 0.2462898, 0.1591989, 0.1407138, 0.0581907, 0.01684675, 
    0.1434581, 0.003487744, 0.0003286455, 0.2395992, 0.1892594,
  0.1379999, 0.129527, 0.07513979, 0.09512176, 0.1163069, 0.08890437, 
    0.09076887, 0.1066319, 0.1046938, 0.1212454, 0.2071691, 0.1581107, 
    0.09074189, 0.07888147, 0.06848321, 0.05024159, 0.09048202, 0.1156144, 
    0.1567301, 0.1521342, 0.07417728, 0.07650913, 0.0542562, 0.03553874, 
    0.03798639, 0.00222929, 0.0002679068, 0.006467341, 0.08203717,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0.0001467839, 
    0.003434793, -4.004327e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, -0.0002450999, 0.008814868, 0.0009044587, 0, 0, 0, 0, 0, 0, 0, 
    0.0003227606, -0.0001453978, 0.0001001532, 0.001666013, 0.00517986, 
    0.01044169, 0.003646134, 0.01229674, 0.01536794, 0.008399932, 
    0.004350817, 0.01638816, -5.767979e-05, 0, 0, 0, -5.499584e-07, 0,
  0.01073778, 0.011346, 0.01319823, 0.01693629, 0.00253394, 0.0194757, 
    0.03488883, 0.04797737, 0.03988455, 0.01640558, 0.03717517, 0.03136328, 
    0.03999097, 0.06693851, 0.1009143, 0.1138236, 0.07580098, 0.08145902, 
    0.03524875, 0.04559362, 0.04842208, 0.02144331, 0.013982, 0.02729307, 
    0.04394176, 0.06680026, 0.04172774, 0.02151729, 0.004048311,
  0.08692296, 0.0592456, 0.160204, 0.1856715, 0.179036, 0.1859409, 0.128951, 
    0.1000954, 0.110063, 0.08380237, 0.09344611, 0.101322, 0.07333874, 
    0.09248831, 0.2508256, 0.1142436, 0.0878424, 0.08747791, 0.1090578, 
    0.06553509, 0.09930393, 0.08004526, 0.1133558, 0.1003757, 0.1228047, 
    0.2177241, 0.1121105, 0.08827565, 0.07571928,
  0.1913509, 0.1023486, 0.07126449, 0.1661589, 0.08023772, 0.07821978, 
    0.09398672, 0.02658193, 0.03647986, 0.03026316, 0.04951619, 0.09359469, 
    0.03770154, 0.09857953, 0.09154774, 0.1826977, 0.09594861, 0.1956932, 
    0.178644, 0.2455024, 0.2089833, 0.2071711, 0.1575143, 0.1119535, 
    0.1408395, 0.1078915, 0.1915054, 0.1781139, 0.1739547,
  0.0001162709, 5.336315e-06, -2.992513e-05, 0.0002195427, 0.008049021, 
    0.01628278, 0.005909942, -7.75959e-10, -3.537253e-05, 0.02662181, 
    0.01939204, 0.006626665, 0.007640487, 0.001820374, 0.01935898, 
    0.04439937, 0.1192035, 0.1083815, 0.06894019, 0.08981813, 0.05265288, 
    0.01930336, 0.00543895, 0.00699199, 0.03525908, 0.1158427, 0.06547774, 
    0.01081026, 0.002052214,
  7.897837e-09, 3.40905e-08, 4.363569e-08, -5.737744e-11, -1.47985e-07, 
    -5.442145e-05, 2.195547e-06, 0.02968305, 0.002425595, -3.857134e-05, 
    0.003918425, 1.208793e-06, 9.515114e-07, 0.03058092, 0.01343806, 
    0.03539916, 0.0202498, 0.002342488, 0.004359995, 3.986368e-06, 
    -3.121195e-10, -6.184413e-06, 1.266172e-08, -1.536125e-08, 0.01130945, 
    0.0007004798, 1.647289e-07, 1.732059e-07, 2.096105e-07,
  1.992496e-06, 1.491873e-06, 5.032917e-07, 2.029422e-05, 0.003339713, 
    0.005896761, 0.04495624, 0.1264515, 0.003639145, 0.003173684, 
    0.004184491, 0.05755537, 0.06074029, 0.03669946, 0.0161546, 0.01750577, 
    0.0004161935, 7.511389e-06, 0, 0, 6.841219e-07, 4.441322e-08, 
    1.211371e-06, 0.001693275, -1.285724e-05, 3.847252e-07, -2.275998e-08, 
    -9.862041e-10, 2.13525e-07,
  0.003406969, 0.01783264, 0.04697638, 0.008470767, 0.00157098, 0.06218614, 
    0.04332845, 0.04844843, 0.1394393, 0.195946, 0.04315083, 0.1257366, 
    0.1720953, 0.06524555, 0.02260691, 0.001749267, 6.506954e-05, 
    -4.817954e-10, 1.651549e-07, 1.040938e-06, 2.476043e-06, 6.507204e-06, 
    0.005367931, 0.02463242, 0.008642971, 0.001914836, -6.314734e-05, 
    0.0002033648, 0.01844246,
  0.1575838, 0.2934704, 0.2376687, 0.1672594, 0.0001641572, 0.001729423, 
    0.06019455, 0.03902426, 0.1459072, 0.0243057, 0.04600811, 0.09803944, 
    0.2285363, 0.0736656, 0.05567566, 0.1039758, 0.06784786, 0.04812158, 
    0.0563798, 0.03514275, 0.14177, 0.123916, 0.1600436, 0.03254435, 
    0.04144698, 0.03993921, 0.05504829, 0.1352172, 0.2368296,
  0.0001243314, 0.003617896, 0.01312159, 0.1399802, 0.2288355, 0.2369779, 
    0.2388003, 0.03428193, 0.2503525, 0.04082474, 0.1716874, 0.2025685, 
    0.1018494, 0.08487922, 0.05965241, 0.006100872, 2.450689e-07, 
    4.953638e-07, -1.948175e-05, 0.009091262, 0.04254455, 0.06744, 0.0221461, 
    0.009717618, 0.01857114, 0.006368086, 9.275856e-05, 6.949089e-05, 
    0.001803497,
  -1.138775e-08, -4.125506e-08, 0, 0.01943048, 0.008308095, 0.01976997, 
    0.04779878, 0.1734972, 0.1214309, 0.07149888, 0.101753, 0.02325816, 
    0.03963491, 0.0770653, 0.1169742, 0.009423207, 0.03372037, 0.00347203, 
    3.19324e-05, 0.01053094, 0.05325282, 0.009407125, 0.05486698, 0.1069082, 
    0.03545661, 0.01201034, 3.542199e-06, 7.250405e-08, 1.687061e-05,
  0.03731913, 0.02961019, 0.01966986, 0.0001865757, 0.0146203, 0.02960124, 
    0.03711442, 0.0652743, 0.1820347, 0.1204354, 0.2207572, 0.1181624, 
    0.1378978, 0.1385966, 0.2594764, 0.2421644, 0.1471057, 0.1253536, 
    0.03562208, 0.01279142, 0.0378967, 0.08466574, 0.06925256, 0.05068178, 
    0.08532778, 0.04225387, 0.03920965, 0.05325671, 0.02383532,
  0.1670642, 0.07827021, 0.08063293, 0.08237091, 0.1185502, 0.1108312, 
    0.09294651, 0.0872043, 0.1861701, 0.221557, 0.1796315, 0.115462, 
    0.1366171, 0.1643277, 0.1445515, 0.1126236, 0.1149168, 0.12244, 
    0.06924616, 0.06983155, 0.07043973, 0.1338872, 0.1214591, 0.1153009, 
    0.08993003, 0.1116638, 0.1459583, 0.1807162, 0.1577324,
  0.1972777, 0.15845, 0.1571281, 0.1820389, 0.16104, 0.1574281, 0.3271778, 
    0.2213805, 0.1880147, 0.2073613, 0.1716102, 0.177384, 0.1082435, 
    0.2227944, 0.1294597, 0.2059791, 0.1594493, 0.1994628, 0.2454209, 
    0.1906843, 0.1075619, 0.1346405, 0.1197666, 0.07690407, 0.2441681, 
    0.2094511, 0.144887, 0.1538981, 0.1968267,
  0.143158, 0.157228, 0.221137, 0.1681278, 0.2053323, 0.2049912, 0.1616925, 
    0.3234056, 0.2138745, 0.1225921, 0.1719179, 0.1524162, 0.1995557, 
    0.1889976, 0.2167278, 0.08909481, 0.1262663, 0.1664585, 0.1604, 
    0.2977226, 0.2475149, 0.1423507, 0.07048564, 0.09951791, 0.1719534, 
    0.0667285, 0.007360405, 0.3283008, 0.2102892,
  0.2616034, 0.2707604, 0.1757071, 0.1515462, 0.1372812, 0.125373, 0.1163189, 
    0.1403447, 0.1264116, 0.1146888, 0.1714921, 0.1488627, 0.1040724, 
    0.1175049, 0.1168731, 0.1579455, 0.1837811, 0.2094088, 0.2424776, 
    0.2454866, 0.1136743, 0.09565301, 0.09441605, 0.07125429, 0.09819949, 
    0.03502032, 0.008357204, 0.07184609, 0.1905274,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0.0003029114, -0.0001421515, 0, 
    -6.833993e-05, 0.01560512, 0.001995915, 0, 0, 3.843055e-05, 
    -1.968563e-05, 0, 0, 0, 0, 0,
  3.03774e-05, 0.01138644, 0.0666557, 0.04019859, -1.704475e-08, 0, 
    -2.905228e-05, -6.883677e-06, 0, -3.971417e-05, 0, 0.0007719947, 
    0.0007529307, 0.04525954, 0.04173731, 0.03961547, 0.03300515, 0.03138437, 
    0.0727826, 0.07503721, 0.03545958, 0.02553932, 0.04503911, 0.01407169, 
    0.01139057, 0.02884607, 0.005611651, 9.370944e-05, 7.10229e-06,
  0.03274067, 0.02351247, 0.04691754, 0.06126364, 0.08105376, 0.1065431, 
    0.1076853, 0.1023843, 0.08717668, 0.05913474, 0.07263926, 0.06851593, 
    0.1352728, 0.2116065, 0.2246, 0.2209445, 0.1626866, 0.1731945, 
    0.09624291, 0.08044552, 0.07433106, 0.03091559, 0.03775385, 0.06982788, 
    0.105391, 0.171809, 0.08164372, 0.05687328, 0.03155478,
  0.1274569, 0.1251312, 0.2465125, 0.2691723, 0.2148216, 0.2112358, 
    0.1304585, 0.1357783, 0.1450408, 0.1151271, 0.1669571, 0.1739224, 
    0.2102877, 0.2015448, 0.3043264, 0.1181271, 0.1341427, 0.1594637, 
    0.2047445, 0.1232866, 0.209056, 0.1823833, 0.1960318, 0.1629883, 
    0.152636, 0.2369135, 0.1835911, 0.1243033, 0.1082025,
  0.1610774, 0.09054825, 0.08656057, 0.1513142, 0.08075205, 0.08504158, 
    0.09938697, 0.04617272, 0.05654541, 0.06051062, 0.09107191, 0.1309518, 
    0.08338665, 0.1408715, 0.1229623, 0.1952758, 0.1049693, 0.2073549, 
    0.1676252, 0.2070052, 0.2016043, 0.2059246, 0.1783959, 0.1550071, 
    0.1236471, 0.09603681, 0.1480851, 0.1836794, 0.157277,
  2.877401e-05, 8.530792e-06, -8.438777e-06, 0.0003184245, 0.01023864, 
    0.02216941, 0.001318175, -8.403173e-11, -7.180676e-05, 0.01039987, 
    0.02466851, 0.006598706, 0.01154517, 0.003191082, 0.01843591, 0.05507009, 
    0.1092785, 0.1019171, 0.06447251, 0.1035253, 0.04232614, 0.004384562, 
    0.0003824683, 0.002873839, 0.03642337, 0.1192761, 0.07088748, 0.00765608, 
    0.0007749065,
  -1.401197e-10, 1.058022e-09, 3.752188e-08, 2.504206e-08, -7.631203e-06, 
    0.002134313, 8.778807e-07, 0.05005971, 7.152594e-05, -2.749465e-05, 
    0.000648654, 1.132883e-06, -2.050238e-05, 0.03167841, 0.01500802, 
    0.04509831, 0.009857076, -4.050063e-05, 0.003859381, 3.620987e-06, 
    3.698651e-08, -5.609208e-06, 3.235823e-09, -1.825651e-08, 0.0189792, 
    5.174744e-05, 6.303769e-08, 6.123456e-08, 7.254437e-09,
  3.872164e-07, 1.43841e-06, -2.594331e-09, 2.428688e-05, 0.005841927, 
    0.007588019, 0.05449225, 0.1135329, 0.003899551, 0.00640116, 0.004010934, 
    0.03691787, 0.06935739, 0.03435043, 0.01346296, 0.01773581, 0.0005137763, 
    -5.198792e-05, 0, 0, 5.462868e-09, -2.045805e-09, 2.625098e-06, 
    0.001140884, 5.168105e-06, 2.403078e-07, -1.623724e-08, 1.38917e-07, 
    9.591586e-08,
  0.02612831, 0.01367745, 0.03619001, 0.01206575, 0.002573241, 0.04905277, 
    0.02503162, 0.02225017, 0.08571941, 0.2095616, 0.03368194, 0.1323861, 
    0.1722232, 0.06796981, 0.01572539, 0.001640778, 0.0001804598, 
    1.191515e-08, -1.608512e-08, 1.456769e-07, 6.909948e-06, 6.825535e-07, 
    0.001295916, 0.01336316, 0.008714245, 0.002245198, -2.144384e-05, 
    8.470141e-05, 0.007335397,
  0.1463367, 0.2493357, 0.2260398, 0.1739517, 0.0003967571, 0.003249385, 
    0.0532526, 0.01932364, 0.1241159, 0.01610953, 0.03507132, 0.07304256, 
    0.2013954, 0.05797932, 0.05064682, 0.1075189, 0.06116861, 0.04867642, 
    0.07238518, 0.04852499, 0.1547156, 0.1305699, 0.1284797, 0.02277783, 
    0.03661292, 0.0284345, 0.05228389, 0.1664805, 0.2396293,
  0.0001413524, 0.004329055, 0.02311779, 0.1807219, 0.2115087, 0.1698453, 
    0.2392283, 0.02959323, 0.2362214, 0.0324899, 0.1730094, 0.1820974, 
    0.07786976, 0.06258778, 0.03680436, 0.004201292, 1.31202e-06, 
    4.712876e-07, 2.657418e-05, 0.01201181, 0.041196, 0.05202866, 0.01456588, 
    0.006765045, 0.01404194, 0.003755343, 2.454625e-05, 3.300456e-05, 
    0.001582675,
  0.000247558, -9.127724e-05, 0, 0.03574832, 0.006416891, 0.01464433, 
    0.04574297, 0.1709134, 0.1247656, 0.0613163, 0.08098398, 0.02743375, 
    0.03853012, 0.08219284, 0.1032635, 0.005449285, 0.03267299, 0.006940539, 
    4.579035e-05, 0.001795672, 0.04007816, 0.009682511, 0.03557451, 
    0.07596026, 0.02072556, 0.005779415, 3.215308e-06, 2.722876e-07, 
    0.0004359905,
  0.02659426, 0.03065672, 0.01914695, 0.0002282884, 0.02460257, 0.02539295, 
    0.04186892, 0.06256264, 0.1674297, 0.105562, 0.2221198, 0.09595359, 
    0.1168448, 0.1114326, 0.2327962, 0.2260077, 0.1546129, 0.1059998, 
    0.028972, 0.02064166, 0.02881202, 0.1066192, 0.056766, 0.04053114, 
    0.05825964, 0.04276221, 0.03131137, 0.0451501, 0.01775054,
  0.1455986, 0.07207976, 0.06121033, 0.07373175, 0.1134943, 0.1105745, 
    0.09787337, 0.06601819, 0.1923809, 0.207705, 0.1666456, 0.1009676, 
    0.1176463, 0.1337538, 0.1315787, 0.1042575, 0.1127915, 0.1205518, 
    0.0699345, 0.05814324, 0.05953065, 0.1372957, 0.1171612, 0.1122129, 
    0.08480164, 0.1074021, 0.1400179, 0.1588226, 0.1401995,
  0.1647752, 0.1428271, 0.1418345, 0.1743121, 0.1539193, 0.166846, 0.30239, 
    0.2039887, 0.167026, 0.1876981, 0.1475248, 0.1582145, 0.1052415, 
    0.2160591, 0.1323943, 0.1864069, 0.1569033, 0.1887847, 0.2624992, 
    0.1842693, 0.09805962, 0.1256615, 0.1161312, 0.07407006, 0.2340181, 
    0.2128527, 0.1514021, 0.1435307, 0.2057797,
  0.1428544, 0.1498357, 0.2457849, 0.1423524, 0.1946169, 0.192527, 0.1591201, 
    0.2780103, 0.1946613, 0.1196637, 0.1545305, 0.1524559, 0.1794156, 
    0.1861257, 0.2111993, 0.08595295, 0.1328021, 0.1649043, 0.1407698, 
    0.2908074, 0.2864408, 0.1652907, 0.06963598, 0.1189824, 0.2188024, 
    0.1188931, 0.04596858, 0.3131129, 0.2039909,
  0.2716673, 0.2783401, 0.188041, 0.1601328, 0.141531, 0.1197065, 0.1010083, 
    0.1433154, 0.1113634, 0.09344418, 0.1343369, 0.1104266, 0.1166863, 
    0.1648345, 0.1649262, 0.1754477, 0.1680975, 0.1881661, 0.2372162, 
    0.2387904, 0.1224754, 0.120258, 0.1219219, 0.0858141, 0.1365777, 
    0.04517908, 0.01774105, 0.1218399, 0.1934728,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01366269, 0.01396733, 0.007026013, 
    -0.0007409184, 0.005490471, 0.02095601, 0.00645804, 8.350571e-05, 0, 
    0.0003058634, 0.03078592, 0.04248163, -0.007082462, -0.0007087471, 0, 0,
  0.02879474, 0.06984443, 0.08735111, 0.06322122, -1.375673e-05, 0, 
    0.0007306271, 0, -9.190896e-05, 0.0004838125, -1.730339e-05, 0.00227, 
    0.04078948, 0.179146, 0.1680471, 0.1883644, 0.1851048, 0.1683914, 
    0.1555334, 0.1488048, 0.1019121, 0.07815517, 0.1027571, 0.05241512, 
    0.1579693, 0.1014396, 0.04272728, 0.01172311, 0.01553761,
  0.05823674, 0.0479998, 0.06215607, 0.1055584, 0.1947694, 0.1721974, 
    0.1611732, 0.1685799, 0.1271324, 0.1401003, 0.1859465, 0.2286259, 
    0.2384826, 0.2878287, 0.2627367, 0.2222821, 0.2058531, 0.1861965, 
    0.1381969, 0.1039167, 0.09848084, 0.07958257, 0.1407242, 0.1487596, 
    0.1911429, 0.2408066, 0.1833065, 0.1539862, 0.1040555,
  0.1241985, 0.126264, 0.2447096, 0.2659116, 0.2046902, 0.1889358, 0.1406687, 
    0.1570656, 0.1680078, 0.1658915, 0.1968377, 0.2154564, 0.244589, 
    0.2037183, 0.3209486, 0.1074487, 0.1443808, 0.1414331, 0.2144566, 
    0.1518561, 0.234091, 0.197081, 0.2137986, 0.2105931, 0.1622399, 
    0.2097072, 0.1755432, 0.1179118, 0.1262908,
  0.1523011, 0.08984277, 0.07177053, 0.1373021, 0.08094306, 0.08321516, 
    0.09712725, 0.06053023, 0.07606703, 0.05887031, 0.09026416, 0.1190385, 
    0.0839363, 0.1307362, 0.108395, 0.1797418, 0.09908079, 0.2027502, 
    0.1551547, 0.1672796, 0.2072417, 0.2133538, 0.1789097, 0.1585953, 
    0.1151458, 0.08768567, 0.1318739, 0.1752764, 0.1500872,
  0.0001239736, 3.292759e-06, -3.826454e-05, 0.0004517021, 0.005384219, 
    0.04843592, -3.781006e-05, -4.631096e-06, -1.347455e-05, 0.004323506, 
    0.01211564, 0.005599839, 0.01516818, 0.004173186, 0.02717216, 0.06552855, 
    0.1151143, 0.1155906, 0.06648261, 0.0773432, 0.02225837, 0.00565945, 
    0.0001697036, 0.005109615, 0.03917288, 0.1241111, 0.06887393, 0.0041301, 
    0.001149137,
  -4.669421e-10, -1.562843e-10, 1.934359e-08, 3.869963e-06, -4.972166e-05, 
    0.0009916734, 8.940367e-08, 0.06396245, 0.002973568, -2.389027e-06, 
    9.043953e-06, 7.772671e-07, -3.326252e-08, 0.03236575, 0.01236056, 
    0.03734693, 0.007548612, 1.91592e-05, 0.01383935, 4.704465e-06, 
    -4.569238e-08, -3.386239e-07, 0, -7.65422e-09, 0.01349091, 5.221432e-07, 
    3.024712e-09, -3.089304e-10, 1.269203e-08,
  6.581656e-07, 2.661223e-07, 5.803834e-08, 0.001318414, 0.01654358, 
    0.009773995, 0.03535593, 0.09580643, 0.00314854, 0.0112335, 0.003189638, 
    0.02022265, 0.09170692, 0.04000657, 0.01980027, 0.01399059, 0.001037378, 
    -4.269305e-05, 0, 0, 1.123572e-08, -1.922798e-09, 1.775296e-06, 
    0.001041019, 8.559682e-06, 4.195269e-07, 3.528214e-12, 3.125689e-08, 
    2.033365e-09,
  0.02154732, 0.02303097, 0.03275067, 0.01759093, 0.01264894, 0.05103735, 
    0.0165669, 0.01389623, 0.06804775, 0.1942673, 0.03500922, 0.1366025, 
    0.1817656, 0.06989999, 0.0122377, 0.00259798, 0.0003579782, 4.638674e-08, 
    -2.409248e-08, -4.342403e-05, 7.3377e-06, 1.496361e-06, 0.0001448288, 
    0.0132296, 0.01012631, 0.004306783, 9.374969e-06, 0.002198341, 0.001549692,
  0.1480555, 0.2259559, 0.2301411, 0.1945084, 0.006629851, 0.004533183, 
    0.06101679, 0.0107352, 0.1074801, 0.01606675, 0.02760614, 0.05400012, 
    0.1968296, 0.05145524, 0.04616928, 0.1028515, 0.06974766, 0.05831321, 
    0.1239092, 0.04620842, 0.1515596, 0.1339412, 0.107762, 0.01979266, 
    0.03233651, 0.02313897, 0.04791305, 0.1885829, 0.2524682,
  0.0003622167, 0.005358886, 0.04940079, 0.1586279, 0.2017498, 0.1631251, 
    0.260373, 0.04080392, 0.2386929, 0.03050121, 0.1617243, 0.1691035, 
    0.06736483, 0.05532945, 0.02261733, 0.003483581, 3.591288e-06, 
    4.317681e-07, 0.001749547, 0.01199865, 0.04183745, 0.04284047, 
    0.01225076, 0.005466507, 0.01089162, 0.002543352, 1.598248e-05, 
    5.305271e-05, 0.003125106,
  0.006470475, 0.002781572, -5.621094e-10, 0.05755918, 0.0090109, 
    0.009763409, 0.04633947, 0.1777373, 0.1372424, 0.06479598, 0.07497575, 
    0.03156123, 0.03945996, 0.06243381, 0.0979225, 0.002653999, 0.03271933, 
    0.01013347, -8.316107e-05, 0.001872966, 0.0263383, 0.01306015, 
    0.02421701, 0.0573033, 0.01648464, 0.003063227, 2.416107e-06, 
    5.987201e-08, 0.001054289,
  0.01965814, 0.02930084, 0.02072123, 0.0003329388, 0.05845809, 0.01519642, 
    0.04004256, 0.04376287, 0.133743, 0.1066979, 0.2178658, 0.08129071, 
    0.09513474, 0.08904359, 0.227976, 0.204926, 0.1420738, 0.1014554, 
    0.02234116, 0.004135725, 0.037204, 0.1105561, 0.03961646, 0.03483496, 
    0.04585838, 0.03686603, 0.03721248, 0.05772712, 0.007522576,
  0.1181448, 0.05832636, 0.04984186, 0.06446771, 0.1068567, 0.1149429, 
    0.08852787, 0.06830098, 0.1667937, 0.196631, 0.1568605, 0.08747781, 
    0.1095046, 0.1162066, 0.1346934, 0.07341041, 0.1018187, 0.120163, 
    0.06385616, 0.0483222, 0.05254448, 0.1478757, 0.1186238, 0.1175261, 
    0.08505385, 0.1162627, 0.1450078, 0.1479852, 0.1362247,
  0.1485546, 0.1235635, 0.1386827, 0.1638289, 0.1493508, 0.1550179, 
    0.2718717, 0.1787711, 0.1437259, 0.1738296, 0.140301, 0.1412232, 
    0.1058259, 0.2135751, 0.1418138, 0.1787357, 0.1622417, 0.1777595, 
    0.2542542, 0.1854199, 0.0883605, 0.1211114, 0.1156393, 0.07320244, 
    0.2258881, 0.2371807, 0.1615109, 0.1488325, 0.1882213,
  0.1677154, 0.144322, 0.2496384, 0.1326146, 0.1951129, 0.1672886, 0.1469417, 
    0.2510099, 0.1704456, 0.1189328, 0.1482176, 0.1512467, 0.1666815, 
    0.1908303, 0.2058307, 0.07825311, 0.1239485, 0.1549218, 0.1300869, 
    0.2731408, 0.2748938, 0.167066, 0.1302302, 0.1007471, 0.2214924, 
    0.1977842, 0.1142908, 0.3166901, 0.2179356,
  0.2683283, 0.2815573, 0.1713804, 0.1313583, 0.1354696, 0.1149362, 
    0.08692957, 0.1344767, 0.08914579, 0.08292567, 0.1158501, 0.0858206, 
    0.1112605, 0.1812538, 0.1941809, 0.1801623, 0.1581066, 0.174153, 
    0.2258739, 0.2188892, 0.1185147, 0.1188655, 0.1620882, 0.09071561, 
    0.1728218, 0.05021604, 0.04911159, 0.1153651, 0.1705852,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  -4.035057e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0509408, 0.0228537, 
    0.04402156, 0.05806921, 0.03157753, 0.04614952, 0.02773069, 0.0002656264, 
    -7.630673e-05, 0.01510427, 0.206903, 0.1704156, 0.06014221, 0.02426377, 
    -0.001015873, 0.0005469737,
  0.08213054, 0.1244852, 0.1438944, 0.0608713, -0.0005305075, -0.0006452381, 
    0.03123326, 9.084973e-05, -0.0007203799, 0.00403675, -0.0001100432, 
    0.007440723, 0.1746401, 0.2253044, 0.1722584, 0.2294954, 0.2452578, 
    0.1958585, 0.1989774, 0.2026027, 0.1360651, 0.1208476, 0.2165643, 
    0.1665537, 0.2598155, 0.1606345, 0.1114338, 0.06048336, 0.09225701,
  0.1221141, 0.1030714, 0.109777, 0.1579942, 0.2232031, 0.2317366, 0.1873118, 
    0.1953694, 0.1543062, 0.1770566, 0.3181901, 0.2995245, 0.2821121, 
    0.28768, 0.2573518, 0.2058978, 0.1956348, 0.1704139, 0.1300958, 
    0.09451527, 0.1112159, 0.116746, 0.2344672, 0.2089381, 0.2200945, 
    0.2884196, 0.2278255, 0.2348204, 0.1798148,
  0.1351132, 0.1432109, 0.2536233, 0.2816653, 0.2077775, 0.1770857, 
    0.1404024, 0.1728431, 0.162449, 0.2042319, 0.2124478, 0.2155956, 
    0.2264242, 0.1798917, 0.2894022, 0.1166152, 0.1332755, 0.1224423, 
    0.2024416, 0.1529135, 0.2247878, 0.1831026, 0.1995074, 0.245955, 
    0.1635354, 0.199286, 0.171442, 0.1147226, 0.1348047,
  0.1421663, 0.0928788, 0.0704551, 0.1387095, 0.0770135, 0.07926746, 
    0.117786, 0.07047149, 0.07645974, 0.05875219, 0.07713881, 0.09838737, 
    0.08839101, 0.1200835, 0.1126537, 0.1785452, 0.1038408, 0.198577, 
    0.1393449, 0.1529064, 0.2059456, 0.2149425, 0.1670617, 0.1556142, 
    0.1022871, 0.08609062, 0.1212582, 0.160345, 0.1315372,
  0.000198406, 1.102963e-06, 6.337311e-05, 0.001076503, 0.003068913, 
    0.0590106, -0.0001036839, 5.167338e-05, -1.865507e-06, 6.479955e-05, 
    0.001165684, 0.001550418, 0.02108009, 0.005620479, 0.0348824, 0.06861673, 
    0.103991, 0.1232333, 0.06860106, 0.07285856, 0.02392289, 0.006743616, 
    -9.083038e-05, 0.005445504, 0.04112147, 0.1208388, 0.07145035, 
    0.004832751, 0.001298956,
  -5.990461e-10, 3.331694e-09, 1.316657e-08, 0.0002026404, -0.0001185399, 
    0.001286156, 1.962557e-07, 0.06179791, 0.001095468, 8.304957e-07, 
    0.0001308011, 1.778076e-06, -7.145701e-08, 0.03727785, 0.01688417, 
    0.0312159, 0.01032874, 4.535209e-05, 0.02610687, 6.590495e-06, 
    -5.342342e-07, 1.604554e-07, 0, 6.303989e-09, 0.009057747, -6.041526e-06, 
    -1.512191e-09, 7.367096e-10, 0,
  3.941187e-07, 3.749657e-06, 2.862785e-07, 0.0008774832, 0.02350087, 
    0.01062312, 0.0372172, 0.08454297, 0.003666813, 0.0189493, 0.001972664, 
    0.01329, 0.104075, 0.04780095, 0.02335495, 0.01787293, 0.00305785, 
    -9.975886e-05, 0, 0, 7.797147e-09, -1.947718e-09, 2.29726e-06, 
    0.001713571, 5.812907e-06, 9.483169e-08, 1.665242e-11, 1.109105e-09, 
    -2.980223e-10,
  0.0208918, 0.05234817, 0.0505395, 0.0346492, 0.03113537, 0.04830549, 
    0.01771414, 0.01083559, 0.0575595, 0.1795178, 0.04104977, 0.1382169, 
    0.1859754, 0.07273082, 0.01183359, 0.004491395, 0.0005628824, 
    7.019184e-08, -7.767903e-09, 0.007290197, 0.0005944504, 5.790919e-07, 
    9.701229e-05, 0.01051119, 0.008151162, 0.007912118, 0.000243028, 
    0.009291415, -0.0003992162,
  0.1575951, 0.2193193, 0.219043, 0.2142294, 0.03053524, 0.003597782, 
    0.06984329, 0.007941989, 0.1068696, 0.01916059, 0.02857005, 0.04418356, 
    0.1762351, 0.04535003, 0.04421703, 0.119648, 0.07620322, 0.06955903, 
    0.1317403, 0.08971852, 0.1410623, 0.1545694, 0.1049788, 0.02105297, 
    0.02859294, 0.02198075, 0.04242102, 0.204049, 0.2826895,
  0.003957652, 0.008931569, 0.04820055, 0.1455595, 0.1699393, 0.1471654, 
    0.2774666, 0.05433707, 0.2475978, 0.03046984, 0.1574729, 0.1689119, 
    0.06943378, 0.05156625, 0.01389789, 0.00466844, -3.420754e-07, 
    -8.367732e-07, 0.002208218, 0.008294689, 0.04682069, 0.0326564, 
    0.009675209, 0.004842999, 0.007943491, 0.001714807, 4.170771e-05, 
    8.586248e-05, 0.02061402,
  0.03337893, 0.001971602, -2.897834e-07, 0.0910781, 0.01798366, 0.005043569, 
    0.04558599, 0.1923881, 0.1698375, 0.07590758, 0.0755607, 0.03506172, 
    0.04296748, 0.05543273, 0.07583921, 0.002146889, 0.04196946, 0.009777093, 
    1.326166e-05, 0.04308341, 0.02003653, 0.01905377, 0.0232858, 0.04198025, 
    0.02219776, 0.002426855, 1.163886e-06, 2.259616e-09, 0.006525431,
  0.01473245, 0.02033623, 0.02384268, 0.00047647, 0.05797435, 0.009772656, 
    0.04851342, 0.01695271, 0.09479163, 0.08868651, 0.2230936, 0.07854252, 
    0.09107957, 0.07259414, 0.2099478, 0.1862085, 0.1417877, 0.09585603, 
    0.01580063, 0.0008569849, 0.0823788, 0.1214338, 0.03095808, 0.03578651, 
    0.04161178, 0.03936501, 0.03113418, 0.03144067, 0.008784105,
  0.09738656, 0.05270083, 0.03733096, 0.06299215, 0.09403466, 0.1200053, 
    0.07472077, 0.07495644, 0.1498202, 0.1894138, 0.147611, 0.09544206, 
    0.09238015, 0.1068822, 0.130057, 0.09411322, 0.1152625, 0.1236318, 
    0.04387158, 0.03261879, 0.05511381, 0.1440084, 0.1323326, 0.1056826, 
    0.08681285, 0.1023605, 0.1482298, 0.1411055, 0.1384374,
  0.1478382, 0.1128654, 0.1461018, 0.1583602, 0.1565267, 0.1555635, 
    0.2508396, 0.1848412, 0.1176954, 0.1480476, 0.1258711, 0.1249018, 
    0.1119649, 0.225954, 0.1643513, 0.1619974, 0.1759686, 0.1713617, 
    0.2702185, 0.1751688, 0.08428188, 0.1381616, 0.1176929, 0.1220507, 
    0.2336856, 0.2573913, 0.1571319, 0.1639348, 0.1993706,
  0.1772387, 0.185243, 0.317446, 0.1297695, 0.1863343, 0.1392401, 0.1423495, 
    0.2442695, 0.1560552, 0.1149642, 0.1367753, 0.1486433, 0.1800684, 
    0.20247, 0.203283, 0.07098225, 0.1283239, 0.1549778, 0.1148835, 
    0.2551982, 0.2697471, 0.1896952, 0.1310437, 0.1179685, 0.2168119, 
    0.281137, 0.1999524, 0.3235066, 0.2249124,
  0.2529149, 0.2784873, 0.159567, 0.1242108, 0.1196341, 0.1080434, 
    0.08249618, 0.1393524, 0.07906016, 0.07577309, 0.1049325, 0.07988169, 
    0.1155356, 0.2181282, 0.2331613, 0.2034427, 0.1791282, 0.1730888, 
    0.2332181, 0.207707, 0.1195456, 0.1270901, 0.1597183, 0.08883705, 
    0.1934029, 0.08326961, 0.08082402, 0.0992576, 0.1436497,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  -0.0002515528, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0009034434, 0.06832854, 
    0.04203538, 0.1009999, 0.1174138, 0.08557181, 0.07345543, 0.05485596, 
    0.006326297, 0.002393352, 0.05742186, 0.2594861, 0.1922435, 0.1420022, 
    0.0977684, 0.004733373, 0.003789161,
  0.2477987, 0.2637111, 0.1914305, 0.08777636, -0.0009296751, -0.0009661821, 
    0.1021765, -0.001719399, -0.0005040343, 0.004507273, 0.0005574768, 
    0.004117281, 0.3019842, 0.2555603, 0.1808702, 0.2675939, 0.2746139, 
    0.1963136, 0.1923086, 0.2151263, 0.195111, 0.1696707, 0.2572669, 
    0.2537647, 0.3092633, 0.1732765, 0.1148931, 0.09171341, 0.1550966,
  0.1782473, 0.1670119, 0.2028098, 0.2204131, 0.2526025, 0.2395854, 0.208076, 
    0.2179353, 0.1727658, 0.2362003, 0.4052314, 0.3251103, 0.2868378, 
    0.2822884, 0.2607387, 0.2083651, 0.1962385, 0.1582439, 0.133449, 
    0.09416206, 0.1178071, 0.1535371, 0.2635664, 0.2149153, 0.2161424, 
    0.2758423, 0.2113163, 0.2319951, 0.1882611,
  0.1758243, 0.1728923, 0.2362681, 0.2737133, 0.2057661, 0.1759146, 
    0.1481549, 0.1838042, 0.1676976, 0.2144655, 0.2135647, 0.2043574, 
    0.2253273, 0.1624977, 0.2809778, 0.1262154, 0.1300936, 0.1121768, 
    0.209279, 0.1462327, 0.2209189, 0.175475, 0.1928111, 0.251437, 0.165758, 
    0.1848129, 0.1266005, 0.1008407, 0.1271293,
  0.1448183, 0.1065684, 0.06815793, 0.1293372, 0.08037198, 0.08052698, 
    0.1063466, 0.06305989, 0.09084527, 0.04907245, 0.07338452, 0.09332551, 
    0.09095768, 0.1204012, 0.1194036, 0.1826629, 0.1066295, 0.1959441, 
    0.1264048, 0.1506844, 0.1792743, 0.2188748, 0.1827087, 0.1548597, 
    0.08996133, 0.08156312, 0.1070428, 0.1703204, 0.1506456,
  0.000113951, -2.959241e-06, 0.0005576852, 0.002928428, 0.004161733, 
    0.05745424, -0.0001092969, 3.560014e-05, -2.078727e-05, -0.000278865, 
    -0.0001204352, 0.001198504, 0.0336758, 0.01068376, 0.04676153, 
    0.08532908, 0.1126227, 0.1255562, 0.0693797, 0.06851009, 0.02231826, 
    0.003758715, 0.0001067377, 0.01120336, 0.04884546, 0.1221633, 0.07477511, 
    0.004186378, 0.0001289641,
  5.632615e-08, 1.756625e-08, 4.198063e-09, 0.0002732246, 6.838533e-05, 
    2.000583e-05, -1.031319e-07, 0.04266144, 0.002799115, 0.0003353648, 
    0.03211048, 4.0786e-05, -5.675363e-08, 0.04117239, 0.005829241, 
    0.0266513, 0.01276938, 6.020875e-05, 0.03876195, 4.154477e-05, 
    -3.709374e-07, -9.576257e-08, 3.230783e-10, 5.96653e-08, 0.006537601, 
    3.528984e-05, 8.430663e-07, 4.299086e-09, 1.1515e-09,
  4.873543e-07, 7.826131e-05, 1.929129e-06, 0.01373859, 0.03558721, 
    0.01400654, 0.04825616, 0.07898185, 0.004775522, 0.03058318, 0.004846714, 
    0.01263234, 0.1278781, 0.06425925, 0.03250711, 0.02546035, 0.002871671, 
    -4.195145e-05, 2.164408e-10, -2.284341e-13, 4.623285e-09, 1.605842e-08, 
    4.472804e-06, 0.002030666, 2.371325e-05, 6.934937e-08, 7.544549e-09, 
    1.87992e-08, 2.138245e-08,
  0.01636745, 0.04552457, 0.1067197, 0.04775908, 0.01183248, 0.04996987, 
    0.01832589, 0.01101632, 0.0450298, 0.183003, 0.03868813, 0.1346551, 
    0.2101833, 0.06733326, 0.012851, 0.004545246, 0.001816829, -5.943477e-07, 
    1.379854e-05, 0.02378433, 0.002073931, -3.684536e-06, 0.0001427005, 
    0.01257636, 0.02019898, 0.01197995, 0.006786444, 0.003948479, 0.007956712,
  0.1699075, 0.2245108, 0.2248426, 0.2557912, 0.07813334, 0.01219707, 
    0.07491283, 0.008595733, 0.131175, 0.03800715, 0.03223127, 0.04779757, 
    0.1880267, 0.05006927, 0.05579507, 0.135552, 0.08943017, 0.08180333, 
    0.1684664, 0.1310135, 0.1524758, 0.1525982, 0.1177791, 0.02998321, 
    0.02766779, 0.02322442, 0.06044012, 0.1991149, 0.3266335,
  0.005959403, 0.01015083, 0.0324637, 0.1727744, 0.1503747, 0.160673, 
    0.3025871, 0.06686523, 0.2877653, 0.03335298, 0.1692401, 0.1674615, 
    0.07208024, 0.05824168, 0.01173269, 0.006475373, 1.32738e-05, 
    8.535368e-05, 0.01381755, 0.009534426, 0.05955734, 0.03511094, 
    0.01019543, 0.005143122, 0.007534364, 0.00124974, 2.824417e-05, 
    0.004778479, 0.009849418,
  0.002876291, 8.345352e-05, -1.283233e-06, 0.08542853, 0.02776034, 
    0.00236222, 0.05152204, 0.1896116, 0.1919386, 0.09438694, 0.08030197, 
    0.05067946, 0.05175562, 0.05674281, 0.1009118, 0.002050562, 0.0389596, 
    0.01210619, 6.374998e-05, 0.0366267, 0.04046411, 0.01948223, 0.0236324, 
    0.03584173, 0.02576561, 0.002329127, 5.058401e-06, -2.83932e-07, 
    0.02658169,
  0.01099704, 0.008782538, 0.02910977, 0.0008455216, 0.03376943, 0.004442804, 
    0.05707149, 0.005594297, 0.05546027, 0.08003798, 0.2101614, 0.07510781, 
    0.09167004, 0.06300367, 0.1794167, 0.2007289, 0.1354716, 0.09940427, 
    0.01561523, 0.001164239, 0.1195297, 0.1202524, 0.03333551, 0.03640782, 
    0.03851717, 0.04228512, 0.02543506, 0.03634621, 0.006711773,
  0.07038511, 0.06944694, 0.03943682, 0.05416522, 0.08352739, 0.1168803, 
    0.06974167, 0.08409066, 0.1364879, 0.1850044, 0.1400391, 0.08125848, 
    0.09841142, 0.09981121, 0.1228303, 0.07959299, 0.1085484, 0.111145, 
    0.04437757, 0.02803219, 0.06115218, 0.1332012, 0.1360456, 0.1074152, 
    0.08861802, 0.09152906, 0.1538983, 0.150227, 0.1114905,
  0.1196626, 0.09994389, 0.1372142, 0.1618911, 0.1752985, 0.1660986, 
    0.2432794, 0.2077393, 0.1176468, 0.119909, 0.1126311, 0.1161468, 
    0.1238445, 0.2409273, 0.1499474, 0.1578377, 0.1624788, 0.1698197, 
    0.2833977, 0.1680084, 0.07047643, 0.1473477, 0.1171552, 0.1098164, 
    0.2446848, 0.2885795, 0.2002605, 0.1898339, 0.1770443,
  0.1359247, 0.1758057, 0.3063154, 0.1328332, 0.190014, 0.1242591, 0.150484, 
    0.2608961, 0.1553403, 0.112115, 0.1183914, 0.138282, 0.1922258, 
    0.1917619, 0.1982123, 0.08195152, 0.1396394, 0.1684555, 0.09779896, 
    0.2412722, 0.2589593, 0.1927038, 0.1467027, 0.1015607, 0.1735001, 
    0.3302425, 0.2400304, 0.3211034, 0.2220302,
  0.226204, 0.2739874, 0.135381, 0.1009139, 0.1169248, 0.1054801, 0.08770832, 
    0.1282004, 0.08677221, 0.06802264, 0.08922929, 0.0821528, 0.1272208, 
    0.2356489, 0.2483654, 0.248756, 0.2369418, 0.2495137, 0.2827789, 
    0.2413777, 0.1365367, 0.163475, 0.1484139, 0.07480358, 0.1877999, 
    0.1134318, 0.0985948, 0.1145776, 0.1506981,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2.122149e-05, -2.122149e-05, 
    -2.122149e-05, -2.122149e-05, -2.122149e-05, -2.122149e-05, 
    -2.122149e-05, 0, 0, 0, 0, 0, 0, 0, 0,
  0.002864336, -5.411986e-05, 0.0006163999, 0, 0, 0, 0, 0, 0, 0, 0, 
    4.127609e-05, 0.01507585, 0.08789463, 0.07649902, 0.1405777, 0.1727097, 
    0.1432603, 0.1150908, 0.1390288, 0.05458417, 0.01934957, 0.1259264, 
    0.2437669, 0.1554793, 0.1266943, 0.09098063, 0.06266368, 0.005449696,
  0.3502121, 0.2928003, 0.2360989, 0.1000293, 2.984597e-05, 0.007744621, 
    0.1346708, -0.003016836, 0.0005443528, 0.02474459, 0.01711554, 
    0.09206583, 0.3539717, 0.2497471, 0.183408, 0.2806445, 0.2710476, 
    0.1920661, 0.1888285, 0.2428574, 0.2361455, 0.3008249, 0.3600188, 
    0.2649031, 0.3008, 0.157626, 0.1014489, 0.1055514, 0.1802387,
  0.2356213, 0.265961, 0.2433239, 0.2447322, 0.2600762, 0.2362113, 0.2050435, 
    0.2282124, 0.1710391, 0.2274534, 0.3812766, 0.3011456, 0.2798169, 
    0.2815525, 0.2530886, 0.1998545, 0.1957291, 0.1522155, 0.1228451, 
    0.09607312, 0.1162422, 0.1315707, 0.2688324, 0.2160765, 0.2261096, 
    0.2675793, 0.2203803, 0.2390924, 0.2145797,
  0.170805, 0.1728558, 0.2183399, 0.2670997, 0.2157427, 0.1696325, 0.1577267, 
    0.1977368, 0.1737853, 0.2025647, 0.1919037, 0.2068364, 0.213438, 
    0.1556037, 0.2689858, 0.1292281, 0.1362744, 0.1244675, 0.2340028, 
    0.150659, 0.2253415, 0.1760395, 0.1913918, 0.2339713, 0.1419247, 
    0.1697063, 0.1103463, 0.0888292, 0.1228427,
  0.1439348, 0.1057419, 0.06280607, 0.1252153, 0.08714741, 0.08846568, 
    0.1047599, 0.0622552, 0.08666924, 0.06218131, 0.08673678, 0.1111608, 
    0.1045849, 0.1318784, 0.1142569, 0.1772851, 0.1055048, 0.1990719, 
    0.1255426, 0.1531927, 0.1720339, 0.2055496, 0.1617654, 0.146824, 
    0.07565296, 0.0735372, 0.0939616, 0.1543704, 0.135399,
  0.0003474107, -4.255482e-05, 0.004301418, 0.006634905, 0.009698646, 
    0.0619898, 7.473366e-05, 5.808075e-05, 4.223271e-05, 0.002577025, 
    9.977251e-05, 0.008866172, 0.04551034, 0.01549555, 0.06750913, 
    0.08743899, 0.1254271, 0.1461667, 0.06949694, 0.07020997, 0.02300895, 
    0.00314377, 0.0001949817, 0.0129384, 0.04862985, 0.1290475, 0.07114551, 
    0.007915177, -0.0002807267,
  4.972042e-07, 6.982183e-08, -2.215908e-08, 1.93134e-06, 0.0004301668, 
    -6.006074e-08, -1.078165e-05, 0.0125307, 0.001697348, 0.0006824709, 
    0.04991068, 1.178452e-06, 2.997924e-08, 0.04542406, 0.004919831, 
    0.0268072, 0.02237358, 8.47616e-05, 0.05038626, 1.146921e-05, 
    -1.31092e-05, -1.049736e-06, 8.733735e-09, 1.972587e-07, 0.004985851, 
    4.293918e-05, 4.29546e-07, 6.838089e-09, 2.717659e-08,
  1.156713e-06, 0.001748136, 7.703568e-05, 0.01652159, 0.04358797, 
    0.02276007, 0.04776509, 0.07494517, 0.008876481, 0.03703106, 0.005568957, 
    0.0172966, 0.1351424, 0.07804468, 0.04384785, 0.0360622, 0.01015057, 
    0.0004154796, 9.827611e-09, 1.523742e-09, 1.476664e-07, 2.026908e-07, 
    5.048565e-06, 0.00261559, 8.072234e-05, 5.053066e-07, 1.012188e-07, 
    8.004062e-08, 1.297153e-07,
  0.01366004, 0.04320209, 0.1788616, 0.05426845, 0.005659739, 0.05379025, 
    0.01989374, 0.02232529, 0.05346523, 0.21136, 0.05415451, 0.1363653, 
    0.2124591, 0.07054688, 0.01295348, 0.003959924, 0.001923875, 
    0.0001595502, 0.0009008232, 0.00061302, -0.0001526137, 3.265978e-05, 
    0.001825906, 0.01065315, 0.01973156, 0.02714767, 0.02676378, 
    0.0002855081, 0.005105345,
  0.1703486, 0.2658535, 0.2606723, 0.3231689, 0.1351719, 0.0164012, 
    0.09057622, 0.0290916, 0.1645153, 0.06976338, 0.05321886, 0.07104712, 
    0.2148893, 0.06039747, 0.07034826, 0.1659178, 0.1107595, 0.1071787, 
    0.2188423, 0.2096466, 0.1766791, 0.1818256, 0.1511808, 0.04615366, 
    0.03461207, 0.03493997, 0.09333466, 0.253256, 0.3632873,
  0.03089315, 0.003373252, 0.02235122, 0.1528544, 0.1401345, 0.2168448, 
    0.3513572, 0.09439946, 0.3528455, 0.05217202, 0.2041321, 0.1954561, 
    0.08997141, 0.07335733, 0.01519201, 0.007128788, 0.001400369, 
    0.004575601, 0.01511092, 0.01387605, 0.08919249, 0.04646232, 0.0131287, 
    0.007637307, 0.01096069, 0.002006242, 0.001605035, 0.00588234, 0.01015136,
  6.367167e-05, 0.0001359357, 2.600233e-08, 0.04150409, 0.02061565, 
    0.005547951, 0.05965972, 0.2074404, 0.2248264, 0.1230718, 0.09880245, 
    0.07379328, 0.05992309, 0.06396652, 0.1086514, 0.003156027, 0.03440985, 
    0.003747318, 1.385438e-05, 0.007262834, 0.06462736, 0.02499012, 
    0.03584968, 0.03983309, 0.03456986, 0.003012948, 6.272759e-05, 
    7.85068e-08, 0.01497866,
  0.006593845, 0.002654359, 0.02842728, 0.001782379, 0.01433796, 0.007228737, 
    0.06038081, 0.00128195, 0.03706125, 0.07469352, 0.1912841, 0.06618225, 
    0.09576443, 0.07031568, 0.1854481, 0.2037815, 0.109586, 0.07641549, 
    0.01869581, 0.0007193777, 0.06621537, 0.1092914, 0.03555104, 0.04583302, 
    0.03743823, 0.04046315, 0.02858839, 0.03137228, 0.003784642,
  0.05482102, 0.05395301, 0.03898199, 0.06410441, 0.07848052, 0.1101927, 
    0.06923179, 0.0879604, 0.1342574, 0.1997278, 0.1354321, 0.09811264, 
    0.1063577, 0.1024702, 0.1144677, 0.0721039, 0.1278057, 0.1245315, 
    0.04251774, 0.02449919, 0.08015813, 0.1101783, 0.1367633, 0.1239176, 
    0.09927426, 0.09328858, 0.1580073, 0.1452322, 0.0999645,
  0.09788709, 0.08964894, 0.134318, 0.1372963, 0.183779, 0.200923, 0.2430956, 
    0.2403798, 0.1217242, 0.1088907, 0.1026455, 0.1126023, 0.1394391, 
    0.2557585, 0.1305227, 0.1531968, 0.1705915, 0.1613703, 0.312991, 
    0.1532686, 0.08289011, 0.1418052, 0.1399839, 0.1129543, 0.2627062, 
    0.3027266, 0.1765802, 0.1921064, 0.1881066,
  0.1702631, 0.1342987, 0.3252286, 0.100347, 0.2030649, 0.1064671, 0.1420714, 
    0.2555466, 0.1505719, 0.1103683, 0.1116084, 0.1478613, 0.162585, 
    0.1936792, 0.1909576, 0.1007884, 0.1543175, 0.1870615, 0.1042299, 
    0.2705339, 0.2707434, 0.264346, 0.2014513, 0.09724931, 0.1683679, 
    0.3406838, 0.2571258, 0.2968313, 0.2262338,
  0.2202127, 0.2758557, 0.13992, 0.1139972, 0.1088256, 0.1054207, 0.08883227, 
    0.1279634, 0.1240732, 0.07979523, 0.08292256, 0.09734032, 0.1687193, 
    0.2693931, 0.3315854, 0.3443924, 0.2920699, 0.2762321, 0.3090123, 
    0.300945, 0.1760599, 0.1736212, 0.1666088, 0.07468749, 0.1861213, 
    0.137607, 0.1139003, 0.1331123, 0.1340028,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2.122149e-05, -2.122149e-05, 
    -2.122149e-05, -2.122149e-05, -2.122149e-05, -2.122149e-05, 
    -2.122149e-05, 0, 0, 0, 0, 0, 0, 0, 0,
  0.008581975, 0.004736247, 0.009372956, 0.003449697, -2.783438e-05, 
    -3.70361e-07, 0, 0, 0, 0, -0.0003125104, 0.01956285, 0.04038547, 
    0.1264906, 0.08138669, 0.1295713, 0.1800518, 0.1952024, 0.186343, 
    0.1933907, 0.1437918, 0.1445334, 0.2151336, 0.2319521, 0.1297094, 
    0.09590606, 0.08714149, 0.119272, 0.0155916,
  0.3630623, 0.2961735, 0.2361678, 0.0951161, 0.004459579, 0.01427826, 
    0.1479446, 0.02608733, 0.02136417, 0.1325832, 0.1332613, 0.3109057, 
    0.3652345, 0.2421173, 0.1767805, 0.2857167, 0.2593951, 0.1955888, 
    0.1818519, 0.2569855, 0.2620791, 0.3494367, 0.3978615, 0.280011, 
    0.2877428, 0.149317, 0.09143606, 0.09931839, 0.2023861,
  0.2514773, 0.2676332, 0.2275737, 0.2355795, 0.2388794, 0.2301747, 
    0.2119848, 0.2345359, 0.1682324, 0.2517064, 0.3906085, 0.2728301, 
    0.2750482, 0.2800573, 0.2668841, 0.1906954, 0.1870843, 0.1734706, 
    0.1263927, 0.115844, 0.13243, 0.1461736, 0.3002343, 0.2006311, 0.2361156, 
    0.2623185, 0.2126961, 0.2307685, 0.2226322,
  0.1893242, 0.1674129, 0.1953231, 0.2476763, 0.2243993, 0.1773802, 
    0.1498241, 0.1966453, 0.1679401, 0.1827071, 0.198352, 0.2113919, 
    0.2356671, 0.1613904, 0.2718088, 0.1404236, 0.1370101, 0.1240519, 
    0.2072732, 0.1442791, 0.2274639, 0.1803055, 0.1727691, 0.2244337, 
    0.1488079, 0.1556129, 0.1124262, 0.09481361, 0.1227676,
  0.1361669, 0.1012522, 0.06689687, 0.1144674, 0.08507682, 0.08372973, 
    0.1075917, 0.07200148, 0.09564751, 0.0765323, 0.09197492, 0.1102998, 
    0.1022397, 0.127937, 0.09868452, 0.1702926, 0.1061806, 0.1997163, 
    0.1186242, 0.1595163, 0.154769, 0.1808126, 0.1436922, 0.141836, 
    0.06293973, 0.06670056, 0.08408672, 0.1574143, 0.1341516,
  0.000446211, 0.0003050867, 0.02905885, 0.01925506, 0.01363701, 0.08283595, 
    0.002843075, 8.404123e-05, 0.001236605, 0.01212575, 0.003002369, 
    0.04099017, 0.06219271, 0.02592847, 0.06795673, 0.09170081, 0.1356008, 
    0.126074, 0.06294768, 0.06780645, 0.03300377, 0.005757993, 0.001493099, 
    0.0126832, 0.04467471, 0.1393647, 0.07063989, 0.0199308, 0.004011128,
  5.975299e-07, 1.010609e-07, -3.225792e-06, 8.938559e-06, 0.003133414, 
    7.672948e-05, 0.005377081, 0.0006766794, 0.0009305206, 0.004575594, 
    0.04333902, 1.604208e-05, 1.3098e-08, 0.04888121, 0.003620941, 
    0.02773508, 0.02938428, 0.0002385124, 0.07624096, 0.000112501, 
    -8.403774e-05, -2.1852e-06, 1.239497e-08, 1.117861e-07, 0.009513431, 
    0.0001570873, 3.334671e-07, 2.35834e-08, 2.088773e-08,
  1.016857e-06, 0.005457866, 0.004049068, 0.01443008, 0.04780391, 0.03430662, 
    0.0549742, 0.08155693, 0.01072595, 0.0325927, 0.007571522, 0.011774, 
    0.144985, 0.09019772, 0.05943983, 0.04221937, 0.0180951, 0.0007299868, 
    7.508239e-08, 1.29563e-08, 2.487582e-07, 2.74435e-07, 6.180358e-06, 
    0.007870121, 0.0009336591, 1.958167e-05, -3.367627e-07, 9.34037e-08, 
    1.50116e-07,
  0.004651698, 0.03851727, 0.2442778, 0.04415279, 0.009609157, 0.07330655, 
    0.02047088, 0.02848397, 0.08055305, 0.2548797, 0.06662777, 0.1419168, 
    0.2088379, 0.08530588, 0.0121998, 0.005800809, 0.001771245, 0.007674193, 
    0.004011663, 0.0002112546, 0.004702571, 3.011592e-05, 0.01713772, 
    0.02025658, 0.03595132, 0.03399127, 0.04063417, 0.002585485, 0.007288917,
  0.216576, 0.3304771, 0.3082724, 0.4059727, 0.1738117, 0.02281885, 
    0.09979704, 0.06473114, 0.1812496, 0.07645749, 0.07740053, 0.09232993, 
    0.2365261, 0.07549044, 0.08029922, 0.1948462, 0.1215519, 0.1289074, 
    0.2480014, 0.2955033, 0.1825256, 0.2140055, 0.173333, 0.07211751, 
    0.03739349, 0.04377564, 0.1092348, 0.265676, 0.3858463,
  0.05794172, 0.003170505, 0.006646803, 0.1091928, 0.1107552, 0.1731123, 
    0.4341729, 0.1003052, 0.425229, 0.06175625, 0.2100932, 0.2026722, 
    0.09029426, 0.07707746, 0.01655513, 0.008788486, 0.001084065, 
    0.0005993504, 0.004625094, 0.01321903, 0.1104364, 0.05683387, 0.01490729, 
    0.01034933, 0.01294684, 0.002799537, 0.0006218597, 0.002165962, 
    0.004874295,
  1.388553e-05, 0.0007241213, 1.330285e-07, 0.01573533, 0.01202271, 
    0.006673319, 0.06054241, 0.2000851, 0.2409687, 0.1252339, 0.1003562, 
    0.07799821, 0.06151383, 0.06683602, 0.1183986, 0.005130841, 0.03342887, 
    -0.0004949959, 0.005272713, 0.0005471862, 0.06775863, 0.02322692, 
    0.0431231, 0.05301664, 0.03814179, 0.004194532, 0.0001486713, 
    8.796587e-08, 0.004721072,
  0.003071592, 0.001475242, 0.02840187, 0.004131869, 0.01072638, 0.009553456, 
    0.04613403, -0.0005161111, 0.02658295, 0.08242188, 0.1811213, 0.06602245, 
    0.09992206, 0.07688396, 0.1971184, 0.22157, 0.1081105, 0.07355653, 
    0.0184648, 0.001431888, 0.02651387, 0.07202185, 0.04511421, 0.05872691, 
    0.04808603, 0.04543716, 0.04036544, 0.03353407, 0.001288081,
  0.04866838, 0.07463189, 0.0485547, 0.06350186, 0.07781328, 0.1112359, 
    0.08414307, 0.08719342, 0.1303092, 0.1779458, 0.136253, 0.1149488, 
    0.1004688, 0.1054452, 0.108515, 0.07772178, 0.1254104, 0.1301397, 
    0.06860746, 0.02170912, 0.1003211, 0.09612214, 0.1403007, 0.1350246, 
    0.1031393, 0.1182577, 0.1649695, 0.1532936, 0.1116387,
  0.092734, 0.08003131, 0.1160924, 0.1262169, 0.1724245, 0.2298184, 
    0.2466433, 0.1892672, 0.1173463, 0.1101713, 0.1091689, 0.1275089, 
    0.1568032, 0.2758159, 0.1656369, 0.1698865, 0.1647543, 0.1617895, 
    0.3201251, 0.1589102, 0.08998209, 0.1590599, 0.166951, 0.1587791, 
    0.2850837, 0.3258707, 0.2174416, 0.1595591, 0.1832345,
  0.1462699, 0.1250435, 0.3124655, 0.1109451, 0.2449789, 0.1165395, 
    0.1663456, 0.2915609, 0.2305179, 0.1058064, 0.1165668, 0.1940584, 
    0.1948153, 0.1522707, 0.172741, 0.08669055, 0.1714315, 0.2412633, 
    0.1011914, 0.2844991, 0.2719873, 0.2655247, 0.1727753, 0.08036873, 
    0.1443369, 0.37167, 0.2708496, 0.2962018, 0.2036995,
  0.2236635, 0.3041916, 0.1394695, 0.08166894, 0.1177307, 0.1170351, 
    0.1242088, 0.1335492, 0.1339038, 0.1041007, 0.09829774, 0.06575613, 
    0.151371, 0.2900107, 0.3340359, 0.291611, 0.2232767, 0.2963153, 
    0.2674635, 0.1948546, 0.1565649, 0.177225, 0.1505037, 0.07895635, 
    0.1572614, 0.183345, 0.1388197, 0.1648755, 0.1391434,
  0.0002160266, 2.046304e-05, -0.0001751006, -0.0003706642, -0.0005662278, 
    -0.0007617914, -0.000957355, 0, 0, 0, 0, 0, 0, 0, -3.41448e-05, 
    -3.41448e-05, -3.41448e-05, -3.41448e-05, -3.41448e-05, -3.41448e-05, 
    -3.41448e-05, -0.0009311023, -0.0007355387, -0.0005399751, -0.0003444115, 
    -0.0001488479, 4.671573e-05, 0.0002422793, 0.0003724775,
  0.009659011, 0.02200538, 0.03799501, 0.01388146, -0.0006149547, 
    2.175257e-06, 1.048697e-06, 0, 0, 0, 0.00355367, 0.03901902, 0.03864556, 
    0.1438436, 0.08203135, 0.1383915, 0.2032284, 0.2093201, 0.2440344, 
    0.2540107, 0.2638932, 0.2171572, 0.23303, 0.2246029, 0.1238158, 
    0.08516933, 0.06948637, 0.1343175, 0.03942403,
  0.3662991, 0.3055154, 0.2474912, 0.08001627, 0.01053668, 0.0771267, 
    0.1488373, 0.08901737, 0.0895321, 0.2207804, 0.2169983, 0.3573767, 
    0.3746889, 0.2626406, 0.2219917, 0.306961, 0.2669072, 0.2190168, 
    0.179698, 0.3161855, 0.2534104, 0.3523653, 0.397757, 0.2956029, 
    0.2830876, 0.131627, 0.08922514, 0.1120253, 0.224586,
  0.2871516, 0.2674278, 0.2479399, 0.2595322, 0.2306748, 0.2175834, 
    0.2238491, 0.2692582, 0.181176, 0.2724109, 0.3915693, 0.2714758, 
    0.2837265, 0.2689973, 0.2621654, 0.1792688, 0.191057, 0.1935868, 
    0.1279541, 0.1346267, 0.1504773, 0.1548543, 0.2949968, 0.225165, 
    0.2282203, 0.2601564, 0.197869, 0.2257214, 0.2488199,
  0.1877085, 0.1727679, 0.212078, 0.2472014, 0.2189814, 0.1799169, 0.1632829, 
    0.210229, 0.1574577, 0.2023034, 0.230593, 0.2311014, 0.2350474, 
    0.1691316, 0.251052, 0.1455118, 0.1333557, 0.1318848, 0.214728, 
    0.1720855, 0.2382906, 0.1699739, 0.162859, 0.2288354, 0.1348145, 
    0.1502476, 0.113709, 0.1040927, 0.1335342,
  0.1464161, 0.1110348, 0.08083542, 0.09823814, 0.08440259, 0.0733582, 
    0.1024743, 0.09073792, 0.1019854, 0.0833921, 0.09286822, 0.1148019, 
    0.1005283, 0.1286055, 0.1040037, 0.1766791, 0.1211773, 0.1967046, 
    0.1077269, 0.1547504, 0.1534758, 0.1767443, 0.1327085, 0.141939, 
    0.06137584, 0.06041892, 0.08256654, 0.147819, 0.1300081,
  0.002202467, 0.0007041676, 0.03720996, 0.01235937, 0.01928922, 0.0749827, 
    0.009031932, 0.0006505277, 0.002761487, 0.01083804, 9.878572e-05, 
    0.0550531, 0.08015395, 0.03216868, 0.06936233, 0.1022554, 0.1391003, 
    0.1162987, 0.06757456, 0.07433644, 0.02924574, 0.01215603, 0.001928701, 
    0.01245362, 0.04673524, 0.1385873, 0.06886294, 0.02366248, 0.0155396,
  1.841043e-07, 3.103283e-08, 2.158388e-05, 0.0008026019, 0.008024446, 
    0.001883353, 0.00532094, 0.0006379407, -0.0002906185, 0.001938547, 
    0.04052252, 6.188938e-05, 2.453156e-05, 0.0515537, 0.002238727, 
    0.02581087, 0.02699671, 0.001443053, 0.08933548, 0.003756719, 
    -0.0001185769, -5.878827e-06, 7.324424e-09, 4.184187e-08, 0.0125227, 
    0.0031469, -7.865179e-06, 9.497981e-08, 1.107804e-08,
  5.364617e-06, 0.0009155684, 0.02546099, 0.004927923, 0.04969321, 
    0.02911838, 0.07688637, 0.07221089, 0.00841827, 0.02367018, 0.008163699, 
    0.008235902, 0.144428, 0.1014906, 0.06365613, 0.04660812, 0.02284284, 
    0.0009015898, 5.433705e-05, 5.349623e-08, 2.105152e-07, 1.296527e-07, 
    7.332248e-06, 0.01499765, 0.00899566, 0.005532445, 7.268584e-05, 
    1.918547e-07, 1.6048e-07,
  0.008861004, 0.04844573, 0.2661526, 0.04280498, 0.003999819, 0.06877942, 
    0.02179377, 0.03017761, 0.09359817, 0.2779329, 0.04283734, 0.093365, 
    0.1844024, 0.08093487, 0.01494578, 0.00943407, 0.002819574, 0.004156274, 
    0.0005954186, 0.0164536, 0.01040076, 0.001406546, 0.02759232, 0.04561815, 
    0.04146102, 0.02148239, 0.01567715, 0.007389848, 0.001568671,
  0.2359938, 0.3493273, 0.3444256, 0.4635637, 0.13016, 0.04829558, 0.1035184, 
    0.0584199, 0.09875801, 0.06974892, 0.04915246, 0.05302026, 0.1771875, 
    0.06528988, 0.06523908, 0.1950931, 0.138215, 0.144592, 0.2554137, 
    0.306582, 0.1478783, 0.1899952, 0.1887927, 0.08417369, 0.03332249, 
    0.04135957, 0.09532136, 0.2303739, 0.4200923,
  0.02126652, 0.01276132, 0.0003209597, 0.05141533, 0.05915979, 0.09630986, 
    0.3531917, 0.09132387, 0.4548085, 0.0533843, 0.1631467, 0.1348851, 
    0.06340352, 0.06060844, 0.01523208, 0.01193471, 0.0008714569, 
    1.141553e-05, 0.003233182, 0.008402112, 0.08071035, 0.06400845, 
    0.01354398, 0.008367361, 0.01305964, 0.001799819, 9.097949e-05, 
    0.001165606, 0.003827391,
  5.251408e-06, 0.003036458, 3.984834e-09, 0.004205873, 0.005903838, 
    0.004436262, 0.06154281, 0.2414581, 0.2484395, 0.09694804, 0.07698339, 
    0.05602558, 0.05047451, 0.06312117, 0.1105074, 0.006110695, 0.02698265, 
    -0.0004578349, 0.001320858, 2.526728e-05, 0.07443769, 0.01799207, 
    0.03194847, 0.05191237, 0.02323613, 0.005738589, 0.0001516943, 
    2.690901e-08, 0.0004397069,
  0.0005210851, 0.0009528745, 0.03448955, 0.007348468, 0.007269109, 
    0.006641608, 0.0236927, -0.000121558, 0.02199009, 0.09441464, 0.1750838, 
    0.06371142, 0.09907165, 0.07175077, 0.2349515, 0.2833907, 0.107396, 
    0.1064755, 0.02518843, 0.0006222734, 0.008216185, 0.03497785, 0.04989669, 
    0.06224768, 0.0526721, 0.05396114, 0.05461737, 0.0301649, 0.001556679,
  0.05593982, 0.0801831, 0.06941134, 0.1086893, 0.09840747, 0.08242191, 
    0.1005339, 0.0756965, 0.1194215, 0.1645613, 0.1436504, 0.1236038, 
    0.1206387, 0.137923, 0.1282842, 0.08398402, 0.1382466, 0.1412368, 
    0.08722869, 0.03660894, 0.1159859, 0.07304494, 0.1286829, 0.1382052, 
    0.1237132, 0.1296105, 0.1714392, 0.1594155, 0.1793287,
  0.0970649, 0.08222543, 0.1217577, 0.1427522, 0.178034, 0.2687149, 
    0.2370709, 0.2013339, 0.1340692, 0.1259226, 0.1118696, 0.145699, 
    0.1767967, 0.2978386, 0.1616209, 0.1591394, 0.1492061, 0.1865375, 
    0.3397966, 0.188691, 0.1079689, 0.1862734, 0.1942097, 0.1613032, 
    0.3240142, 0.3213689, 0.2404486, 0.1610533, 0.1683692,
  0.1526096, 0.1316918, 0.3506891, 0.1331602, 0.181215, 0.1226445, 0.1414853, 
    0.2911505, 0.179021, 0.1503866, 0.1285121, 0.2220692, 0.2250949, 
    0.2006544, 0.1965948, 0.1221457, 0.1566056, 0.2344848, 0.1164523, 
    0.294244, 0.2481014, 0.2251818, 0.1577379, 0.1171711, 0.1492326, 
    0.4000941, 0.2906454, 0.2977739, 0.2396523,
  0.2352769, 0.2779741, 0.1426803, 0.08663887, 0.0937534, 0.1105982, 
    0.1015109, 0.1334533, 0.1182741, 0.101809, 0.09181442, 0.1088475, 
    0.1923178, 0.2607903, 0.2587618, 0.2340647, 0.2111645, 0.2176936, 
    0.2414672, 0.2309574, 0.1599672, 0.1787379, 0.1846343, 0.08978356, 
    0.1587489, 0.208473, 0.1603705, 0.187171, 0.1635707,
  0.007446679, 0.006876235, 0.006305791, 0.005735346, 0.005164901, 
    0.004594456, 0.004024012, 0.005674387, 0.005326509, 0.004978631, 
    0.004630753, 0.004282875, 0.003934996, 0.003587118, -0.002535401, 
    -0.001098761, 0.0003378779, 0.001774517, 0.003211156, 0.004647796, 
    0.006084435, 0.00437469, 0.003856373, 0.003338057, 0.00281974, 
    0.002301424, 0.001783107, 0.001264791, 0.007903035,
  0.02753555, 0.03381344, 0.06471913, 0.05270502, 0.003969874, 0.0003586576, 
    0.0009119067, 0, 0, 5.289384e-05, 0.02527548, 0.04708225, 0.03206347, 
    0.1476341, 0.08034614, 0.1655616, 0.2798175, 0.2280052, 0.2804354, 
    0.2796884, 0.3241523, 0.2820588, 0.2224746, 0.2104045, 0.1165396, 
    0.08504811, 0.06953531, 0.1252354, 0.0572795,
  0.3520279, 0.3045838, 0.2866009, 0.07790297, 0.02507767, 0.1537106, 
    0.1522574, 0.1169422, 0.1883157, 0.284062, 0.2642897, 0.3738377, 
    0.3849139, 0.2862764, 0.2419104, 0.3342501, 0.3035451, 0.2395589, 
    0.1868338, 0.3143756, 0.3155802, 0.3600806, 0.4058398, 0.328081, 
    0.2963653, 0.1252472, 0.1249748, 0.09880415, 0.2322615,
  0.3278791, 0.3285492, 0.2922274, 0.2993289, 0.2617804, 0.2270751, 
    0.2510833, 0.3227143, 0.2555157, 0.297547, 0.3959925, 0.2609758, 
    0.269019, 0.2691243, 0.2806783, 0.1974222, 0.2213532, 0.2194712, 
    0.1447349, 0.1559801, 0.190505, 0.212041, 0.3157274, 0.2346254, 
    0.2163913, 0.2366006, 0.2040284, 0.2293249, 0.2728827,
  0.2151277, 0.1959487, 0.25281, 0.2463407, 0.2185485, 0.2085896, 0.1849637, 
    0.2487547, 0.1871002, 0.2037991, 0.2224955, 0.2369622, 0.2421265, 
    0.1737258, 0.267481, 0.1570271, 0.1179641, 0.1823931, 0.229157, 0.208027, 
    0.2461131, 0.2007915, 0.168769, 0.2311446, 0.1507008, 0.1492471, 
    0.1249687, 0.1174024, 0.144867,
  0.1660766, 0.148093, 0.08945387, 0.086315, 0.09022973, 0.08851296, 
    0.1093056, 0.09666105, 0.1060141, 0.1070462, 0.09617782, 0.1198453, 
    0.09998485, 0.125545, 0.1132138, 0.1670945, 0.1181446, 0.1907783, 
    0.1037025, 0.1544514, 0.1657713, 0.2012004, 0.1329769, 0.1454429, 
    0.04977306, 0.05578747, 0.08410471, 0.144718, 0.1478928,
  0.006478109, 0.00103988, 0.02700056, 0.01337612, 0.03381035, 0.08623219, 
    0.01698372, 0.003675241, 0.004572575, 0.01292791, 0.0002678841, 
    0.03219207, 0.06939917, 0.03437105, 0.07100168, 0.1166232, 0.1502881, 
    0.1200595, 0.08246814, 0.08440378, 0.03918139, 0.01989817, 0.003938888, 
    0.01383989, 0.05159621, 0.1323656, 0.07264505, 0.03987161, 0.0188742,
  5.277053e-08, 8.996783e-09, 0.0006173121, 0.002319402, 0.01419859, 
    0.00800237, 0.008764798, 0.003467178, -0.0001924508, 2.762961e-05, 
    0.02317826, 5.961687e-06, 0.0003801683, 0.05246842, 0.002619538, 
    0.02465694, 0.04286114, 0.00457586, 0.08090785, 0.02922108, 
    -8.567417e-05, -8.463796e-05, 2.444562e-09, 3.237396e-07, 0.009772203, 
    0.006855498, 0.0007843555, 2.675988e-07, 2.810314e-08,
  3.605948e-07, 6.708274e-05, 0.03730487, 0.03695528, 0.04530168, 0.03140326, 
    0.06137012, 0.06857453, 0.01354042, 0.01298428, 0.009336036, 0.005407819, 
    0.1540115, 0.1056107, 0.06005166, 0.05169404, 0.02988641, 0.003280184, 
    0.0001173711, 7.523177e-08, 1.261335e-07, 3.44943e-08, 3.730959e-06, 
    0.01674975, 0.07868638, 0.002819114, 0.006993998, 1.727003e-05, 
    1.197349e-07,
  0.001640152, 0.04080557, 0.2229552, 0.03465711, 0.001641296, 0.05877846, 
    0.01600134, 0.03359307, 0.06554704, 0.2394024, 0.03279354, 0.05674176, 
    0.1688238, 0.07565685, 0.01614862, 0.009418802, 0.006206684, 
    0.0007849837, 1.708104e-07, 0.0123019, 0.000789581, 0.00222591, 
    0.04101717, 0.06307165, 0.03417126, 0.01720216, 0.006512888, 0.01215071, 
    0.002399696,
  0.1399122, 0.2406994, 0.2628643, 0.5387151, 0.1242291, 0.03969803, 
    0.1214255, 0.05755027, 0.05697554, 0.05850575, 0.03652411, 0.03254685, 
    0.1369539, 0.05785963, 0.05821141, 0.192712, 0.1392873, 0.1638911, 
    0.2475053, 0.2922994, 0.1264989, 0.172964, 0.1678219, 0.08630197, 
    0.03159443, 0.04159493, 0.09123313, 0.2034004, 0.3362571,
  0.003706636, 0.008245965, -8.327462e-05, 0.05067242, 0.04000716, 
    0.06333319, 0.2985103, 0.08704837, 0.4430455, 0.04505696, 0.1451905, 
    0.09297428, 0.04944685, 0.05067903, 0.01503419, 0.01973537, 0.0002698434, 
    2.822398e-07, 0.003020688, 0.005100944, 0.05952537, 0.06267332, 
    0.01208676, 0.007947841, 0.01119613, 0.001647629, 9.161116e-06, 
    5.652536e-05, 0.001880187,
  3.331291e-06, 0.00690059, -2.165605e-11, 0.0002452436, 0.001333862, 
    0.00284172, 0.05839005, 0.2632409, 0.3032062, 0.09502304, 0.06095457, 
    0.04851776, 0.0395708, 0.03585789, 0.08132922, 0.004817754, 0.02339923, 
    0.007937218, 0.001048091, 1.212117e-05, 0.050478, 0.0196799, 0.02616686, 
    0.02483825, 0.01858586, 0.006346185, 0.0002196035, 2.015847e-08, 
    7.577571e-05,
  0.0009345433, 0.0008368084, 0.025664, 0.01137691, 0.001235611, 0.004615435, 
    0.008648489, -4.731078e-05, 0.0243552, 0.1044956, 0.1543247, 0.0461311, 
    0.1046357, 0.07032453, 0.1563414, 0.2980884, 0.1771372, 0.1046172, 
    0.03583907, 0.001204253, 0.006752549, 0.01124189, 0.03346475, 0.04762203, 
    0.04073277, 0.05943602, 0.05554745, 0.03000415, 0.001935574,
  0.04935245, 0.08977979, 0.07492485, 0.119269, 0.09412164, 0.06115909, 
    0.07463758, 0.0748265, 0.1271442, 0.1647557, 0.148904, 0.135815, 
    0.1137635, 0.1489978, 0.133591, 0.09989519, 0.1501939, 0.1471167, 
    0.1039466, 0.05801129, 0.1256765, 0.05052971, 0.1129537, 0.1661222, 
    0.1283984, 0.1396461, 0.193854, 0.1681922, 0.1659021,
  0.1328887, 0.08745764, 0.1201086, 0.1800377, 0.207279, 0.2753338, 
    0.2669611, 0.2306295, 0.173857, 0.1368171, 0.1211268, 0.1692614, 
    0.2046065, 0.3436145, 0.1807798, 0.1785908, 0.1917473, 0.2217276, 
    0.3465284, 0.2282895, 0.1069158, 0.1712149, 0.1937553, 0.1645296, 
    0.2868632, 0.3132321, 0.200136, 0.1591856, 0.1826398,
  0.1951889, 0.1261128, 0.3152251, 0.1524531, 0.1619634, 0.09198822, 
    0.1638906, 0.2740785, 0.1662812, 0.128151, 0.1020246, 0.1723084, 
    0.2058629, 0.2010746, 0.2000567, 0.1227812, 0.1677077, 0.2794488, 
    0.1093481, 0.348516, 0.2406428, 0.2923601, 0.1801575, 0.1013818, 
    0.1226011, 0.4216659, 0.314199, 0.3265671, 0.2687334,
  0.170162, 0.2548504, 0.1245647, 0.08873423, 0.08206794, 0.07243149, 
    0.08657739, 0.1424977, 0.06683684, 0.07691626, 0.08947096, 0.1273802, 
    0.1808425, 0.2886068, 0.3754984, 0.2579809, 0.2865242, 0.301021, 
    0.2240901, 0.1972514, 0.1544182, 0.1490048, 0.1730529, 0.1052154, 
    0.1346047, 0.176685, 0.156545, 0.1483037, 0.1871689,
  0.0214645, 0.01854335, 0.0156222, 0.01270105, 0.009779899, 0.006858748, 
    0.003937596, 0.0102434, 0.01133181, 0.01242022, 0.01350862, 0.01459703, 
    0.01568544, 0.01677385, -0.003368629, 0.00469959, 0.01276781, 0.02083603, 
    0.02890425, 0.03697247, 0.04504069, 0.06506079, 0.05882531, 0.05258983, 
    0.04635435, 0.04011888, 0.0338834, 0.02764792, 0.02380143,
  0.03801402, 0.03988358, 0.07253133, 0.07502115, 0.009713073, 0.0003445596, 
    0.00253253, -1.635311e-05, 1.459674e-05, 0.008146267, 0.04006093, 
    0.05536216, 0.05350034, 0.1480842, 0.08555431, 0.168799, 0.2612193, 
    0.2490354, 0.2810768, 0.3060003, 0.3813677, 0.2858297, 0.218819, 
    0.2073539, 0.1147407, 0.08852205, 0.06328828, 0.1245378, 0.08646769,
  0.3313092, 0.3034964, 0.3328121, 0.08171584, 0.06069085, 0.1946555, 
    0.184783, 0.1513309, 0.2517195, 0.3100781, 0.2950333, 0.3978636, 
    0.3771542, 0.2785131, 0.2425836, 0.3636195, 0.3351983, 0.2599477, 
    0.2221985, 0.3448736, 0.3228864, 0.357623, 0.4413357, 0.332792, 
    0.3138176, 0.1879509, 0.1654229, 0.1161887, 0.2534183,
  0.4116372, 0.3115891, 0.3158741, 0.3090705, 0.2811662, 0.2628791, 
    0.2757737, 0.3408986, 0.3491584, 0.3321744, 0.4361362, 0.2835524, 
    0.3441175, 0.3263256, 0.3504687, 0.2405011, 0.2770524, 0.2500876, 
    0.1828105, 0.1753143, 0.2222264, 0.2384001, 0.3239408, 0.2831055, 
    0.2611052, 0.2755351, 0.2709572, 0.2854628, 0.3501344,
  0.2371384, 0.2527591, 0.2600235, 0.2623598, 0.2491352, 0.2253661, 
    0.2213743, 0.2723992, 0.2227689, 0.2346795, 0.2669753, 0.2454545, 
    0.2492279, 0.2177464, 0.2578896, 0.1624601, 0.1281829, 0.1903145, 
    0.2183298, 0.222611, 0.2692582, 0.206064, 0.2017066, 0.2395732, 
    0.1431564, 0.1563088, 0.1322775, 0.139061, 0.1766867,
  0.2076546, 0.1773591, 0.1001973, 0.08486674, 0.1233783, 0.09699183, 
    0.1284655, 0.1093627, 0.1079763, 0.113998, 0.09909098, 0.1385694, 
    0.1132242, 0.1289465, 0.1233922, 0.1848167, 0.1248534, 0.198874, 
    0.1158272, 0.159564, 0.1850305, 0.220798, 0.1468169, 0.1490615, 
    0.0331898, 0.05672566, 0.09227045, 0.1573913, 0.1747219,
  0.01937838, 0.00190254, 0.00999776, 0.01309239, 0.03442447, 0.1006516, 
    0.02761501, 0.01251007, 0.01110511, 0.01906921, 0.004706616, 0.02024549, 
    0.04126866, 0.0411063, 0.07793806, 0.1435885, 0.1608663, 0.1189326, 
    0.113832, 0.1013567, 0.04421102, 0.04607138, 0.004155643, 0.0142498, 
    0.04075878, 0.128041, 0.08074683, 0.05311292, 0.03045644,
  4.710839e-08, 4.337051e-09, 0.006138586, 0.001271161, 0.03582112, 
    0.01244703, 0.01418203, 0.007911826, 0.002515808, 0.006956316, 
    0.005517318, -4.911795e-07, 0.001798651, 0.05249272, 0.00871001, 
    0.01938127, 0.06690355, 0.007558979, 0.080226, 0.04389644, 0.0001938682, 
    -2.39536e-05, 5.962001e-09, 4.269728e-06, 0.004112854, 0.00575214, 
    0.008759835, 0.0006437512, 1.854542e-07,
  1.805172e-07, -4.498875e-05, 0.01262338, 0.1336405, 0.04119954, 0.03397162, 
    0.05200658, 0.06441401, 0.01523258, 0.008636901, 0.009080421, 
    0.005831506, 0.179987, 0.1117443, 0.06482601, 0.05923598, 0.0343327, 
    0.005490074, 0.0003302635, 4.155022e-06, 3.865699e-07, 2.880479e-08, 
    1.015799e-06, 0.01771528, 0.03033252, 0.0130946, 0.02571581, 0.001263795, 
    6.712303e-08,
  8.999357e-06, 0.03106728, 0.1071231, 0.03554917, 0.002082553, 0.04503797, 
    0.01277405, 0.03423392, 0.05881013, 0.2072962, 0.03025882, 0.03961121, 
    0.1445707, 0.07349656, 0.0227361, 0.01531252, 0.01252067, 0.0004406608, 
    0.0001728048, 0.008360758, 9.999018e-06, 0.003422456, 0.0399667, 
    0.05619401, 0.02785633, 0.01236006, 0.008462358, 0.001272903, 0.002745445,
  0.1068956, 0.1689167, 0.20476, 0.5947308, 0.08638574, 0.02061655, 
    0.1356882, 0.06414133, 0.04147164, 0.04056345, 0.02991371, 0.02618135, 
    0.1198514, 0.05470121, 0.05906352, 0.1887504, 0.1517532, 0.1755339, 
    0.2403983, 0.286971, 0.1138851, 0.1595929, 0.1553764, 0.0821397, 
    0.02942746, 0.04394906, 0.09634446, 0.1875186, 0.268353,
  0.0005077532, 0.0006740707, -1.078793e-06, 0.05717322, 0.01516546, 
    0.05137583, 0.3014825, 0.08529998, 0.4371038, 0.0409099, 0.1389716, 
    0.08127527, 0.04364617, 0.04676856, 0.02004982, 0.02634264, 0.0007707095, 
    2.398584e-07, 0.003930582, 0.004038509, 0.04471734, 0.06358954, 
    0.01193017, 0.007503855, 0.01609823, 0.002256159, -2.116169e-06, 
    7.130157e-06, 0.0005462123,
  2.733075e-06, 0.003565565, -5.294436e-10, 1.300797e-05, 0.0005172199, 
    0.001128649, 0.0511422, 0.2600944, 0.3208728, 0.09732217, 0.05521822, 
    0.05010005, 0.03514655, 0.03051655, 0.07049756, 0.006664349, 0.02183319, 
    0.001242186, 0.0003175929, 4.545547e-06, 0.01647763, 0.03372732, 
    0.02336626, 0.01748782, 0.0197688, 0.006894469, 0.0007368159, 
    7.862925e-09, 1.548207e-05,
  0.004014733, 0.001098043, 0.01587601, 0.01414259, 2.634356e-05, 
    0.0007056849, 0.00255935, -7.370332e-06, 0.02458708, 0.09841986, 
    0.1437918, 0.04544626, 0.1056794, 0.07874523, 0.1256498, 0.2278704, 
    0.1447411, 0.1010788, 0.05302984, 0.001676257, 0.008102271, 0.00295708, 
    0.03262816, 0.04136164, 0.03514219, 0.04772284, 0.0646797, 0.02914645, 
    0.003513813,
  0.06590537, 0.10373, 0.09754603, 0.1174887, 0.09500784, 0.06248887, 
    0.08044909, 0.07209801, 0.1299761, 0.1642603, 0.1323573, 0.1263177, 
    0.1382752, 0.1673578, 0.1101838, 0.1102874, 0.1498691, 0.1852982, 
    0.1082614, 0.07148769, 0.1293362, 0.03047523, 0.1038256, 0.163282, 
    0.1399423, 0.1406575, 0.1996326, 0.1800523, 0.1661431,
  0.1388027, 0.08884991, 0.1547857, 0.2244467, 0.2548898, 0.3141624, 
    0.2854793, 0.2350094, 0.1789672, 0.1638459, 0.1433338, 0.1680503, 
    0.2176377, 0.3759401, 0.2140106, 0.1942635, 0.2256726, 0.2534429, 
    0.3821061, 0.2281339, 0.1149969, 0.1637171, 0.1989089, 0.1825024, 
    0.2673364, 0.3158445, 0.2415775, 0.1863206, 0.2032218,
  0.2006444, 0.1780885, 0.2947546, 0.174687, 0.1573074, 0.1673074, 0.2297425, 
    0.3471644, 0.2726726, 0.138968, 0.111079, 0.1864855, 0.2174225, 
    0.1625804, 0.2115618, 0.1447582, 0.2392364, 0.2751595, 0.1414892, 
    0.3248926, 0.2385359, 0.3065145, 0.1490997, 0.07933483, 0.09252831, 
    0.4263285, 0.3850394, 0.3056087, 0.2625019,
  0.2082907, 0.210201, 0.1485777, 0.05954123, 0.09981228, 0.08092728, 
    0.09092939, 0.1663329, 0.2070729, 0.1229575, 0.1208812, 0.1180954, 
    0.1258382, 0.2659554, 0.3228038, 0.2419979, 0.2460053, 0.3053469, 
    0.2474595, 0.2465396, 0.1635512, 0.1224859, 0.1438456, 0.1099572, 
    0.1280974, 0.1086481, 0.171245, 0.1099749, 0.2075071,
  0.06314979, 0.05838, 0.05361022, 0.04884044, 0.04407066, 0.03930087, 
    0.03453109, 0.05429926, 0.06094954, 0.06759981, 0.07425009, 0.08090036, 
    0.08755063, 0.09420091, 0.1155173, 0.1254907, 0.1354641, 0.1454375, 
    0.1554109, 0.1653843, 0.1753577, 0.13674, 0.1248861, 0.1130322, 
    0.1011783, 0.08932444, 0.07747055, 0.06561666, 0.06696561,
  0.05340203, 0.05676458, 0.07006292, 0.08341534, 0.01583333, 0.0004155693, 
    0.002751961, -0.0007635042, 0.009535271, 0.06986234, 0.04940925, 
    0.08943167, 0.06190413, 0.1395415, 0.0743154, 0.1729099, 0.2812741, 
    0.26556, 0.3013883, 0.2533722, 0.4060037, 0.3050542, 0.2501278, 
    0.2083406, 0.1132702, 0.08104965, 0.08136591, 0.1518598, 0.1107863,
  0.3396248, 0.3004176, 0.2895315, 0.06955546, 0.1040268, 0.1896671, 
    0.2238977, 0.2075007, 0.3000446, 0.3092583, 0.3242482, 0.4142685, 
    0.3512489, 0.2417437, 0.2271174, 0.3258208, 0.2750667, 0.2242774, 
    0.1853016, 0.3181148, 0.3438531, 0.3525455, 0.4214818, 0.2936136, 
    0.3464443, 0.198286, 0.1403069, 0.1150385, 0.2543606,
  0.3815583, 0.2541888, 0.3301298, 0.3126169, 0.3180368, 0.2667222, 
    0.2556149, 0.310994, 0.2914772, 0.3161277, 0.4131176, 0.2958963, 
    0.3183874, 0.3437201, 0.3298683, 0.23735, 0.2521194, 0.3161839, 0.220725, 
    0.1651533, 0.3059164, 0.2598308, 0.294972, 0.2743116, 0.2481977, 
    0.2972296, 0.2431328, 0.2465419, 0.3275435,
  0.2797801, 0.2569502, 0.270728, 0.2727881, 0.267185, 0.2751038, 0.2664361, 
    0.289491, 0.2364515, 0.2344386, 0.2708421, 0.2566188, 0.2767371, 
    0.2045767, 0.2719885, 0.1966489, 0.1356105, 0.1956227, 0.2393567, 
    0.2512739, 0.2828704, 0.227606, 0.19904, 0.2465705, 0.1393301, 0.1657481, 
    0.1520247, 0.1530002, 0.2056339,
  0.2351689, 0.1935377, 0.1172689, 0.1076892, 0.1333278, 0.1009785, 
    0.1501219, 0.1287977, 0.1471617, 0.1313668, 0.1198168, 0.1529619, 
    0.1037945, 0.1270828, 0.1468637, 0.2315619, 0.141748, 0.2117028, 
    0.1508222, 0.1749804, 0.2241595, 0.239014, 0.1566486, 0.1533073, 
    0.02658811, 0.07630404, 0.1112912, 0.164125, 0.2174814,
  0.03608857, 0.002882919, 0.002168935, 0.01818296, 0.03340066, 0.1042663, 
    0.03196708, 0.01428235, 0.02129766, 0.03558568, 0.01073354, 0.007564717, 
    0.03018554, 0.04490577, 0.09023865, 0.1608208, 0.1538836, 0.1157461, 
    0.1148808, 0.1143851, 0.05588426, 0.05781673, 0.009721396, 0.01905007, 
    0.03043533, 0.1314241, 0.08437399, 0.06744844, 0.04484176,
  -4.53981e-07, 4.370483e-09, 0.000256247, 0.001185561, 0.04759151, 
    0.02080715, 0.01341169, 0.0105939, 0.01778074, 0.007503403, 0.0001085006, 
    0.0004587255, 0.009684579, 0.05912333, 0.01838236, 0.008442435, 
    0.08238638, 0.01611586, 0.1026733, 0.04557153, 0.01049913, -2.595707e-05, 
    1.512484e-08, 6.55347e-05, 0.002897047, 0.003174909, 0.02680102, 
    0.01448445, 0.0005271586,
  1.690597e-07, -6.300433e-07, 0.001621747, 0.1838679, 0.04184924, 
    0.03846808, 0.03237753, 0.07341969, 0.02465911, 0.009201051, 0.01288477, 
    0.0104111, 0.1894361, 0.1147739, 0.07129971, 0.0600481, 0.03637385, 
    0.01550043, 0.00163903, 0.0007827119, 7.030671e-07, 6.183531e-08, 
    4.422374e-07, 0.01740231, 0.00437141, 0.001968016, 0.04789905, 
    0.002996284, 1.070823e-07,
  3.839995e-06, 0.03475593, 0.04756612, 0.05006875, 0.007755585, 0.0378422, 
    0.01290257, 0.03418205, 0.05902782, 0.1881762, 0.03278944, 0.03024673, 
    0.133431, 0.05807595, 0.02718121, 0.03175658, 0.02190942, 0.002686531, 
    0.0002444456, 0.001444958, 1.509816e-05, 0.002185303, 0.03189052, 
    0.04094713, 0.02423472, 0.009379954, 0.009094382, 0.002649877, 
    0.0004355467,
  0.08789521, 0.144727, 0.1757112, 0.5715674, 0.05297252, 0.006341144, 
    0.141837, 0.05466149, 0.03522527, 0.03119845, 0.02588642, 0.02426936, 
    0.1061348, 0.05427707, 0.05946488, 0.175809, 0.1518278, 0.1705274, 
    0.2383989, 0.2587725, 0.1106146, 0.1493134, 0.176091, 0.07625719, 
    0.02920389, 0.04255888, 0.103169, 0.1913189, 0.2436212,
  0.0001203896, 0.0005431662, 1.054303e-06, 0.05465809, 0.008025489, 
    0.04167806, 0.2932728, 0.1068806, 0.4391718, 0.03838855, 0.1271495, 
    0.07934279, 0.0398337, 0.04050243, 0.02295126, 0.02438636, 0.005209556, 
    0.0001011331, 0.00756303, 0.003641269, 0.03168553, 0.06545778, 
    0.01248182, 0.007303797, 0.02166202, 0.009776046, -1.533584e-05, 
    1.492925e-06, 0.0001666207,
  2.119868e-06, 0.0003951292, -8.230479e-08, 6.343698e-06, 0.0002962912, 
    0.0002623703, 0.04685929, 0.2866252, 0.3015162, 0.126829, 0.05330433, 
    0.0523644, 0.02983207, 0.02998496, 0.06639704, 0.01213529, 0.02451402, 
    0.006589624, 1.120956e-05, 1.936326e-06, 0.004234998, 0.01636719, 
    0.02426459, 0.01537387, 0.02693162, 0.009503039, 0.001336489, 
    2.587803e-07, 6.15116e-06,
  0.001026059, 0.00121371, 0.01419896, 0.0161424, -8.741033e-05, 1.01283e-05, 
    1.928886e-05, 4.28247e-07, 0.01698082, 0.08953469, 0.1413596, 0.06347726, 
    0.1177309, 0.08402803, 0.1214764, 0.2109127, 0.09349647, 0.1146524, 
    0.05180494, 0.0006890266, 0.006798355, 0.0005473556, 0.02725325, 
    0.039416, 0.03578089, 0.04496579, 0.06951976, 0.04120534, 0.003495508,
  0.05359575, 0.105758, 0.08978193, 0.1309123, 0.08141571, 0.03190606, 
    0.07313658, 0.0682625, 0.1356939, 0.1636847, 0.127671, 0.1181653, 
    0.1134142, 0.1630099, 0.1328178, 0.1223258, 0.1431821, 0.195841, 
    0.1300224, 0.08257548, 0.09369187, 0.02076514, 0.09551562, 0.1365849, 
    0.1349763, 0.1504589, 0.1950771, 0.1744974, 0.1588905,
  0.1663986, 0.09099815, 0.1934458, 0.2324531, 0.3248321, 0.308166, 
    0.2888796, 0.2900599, 0.1908412, 0.1898019, 0.2073118, 0.2030379, 
    0.2443239, 0.4063522, 0.2175968, 0.2101688, 0.2501895, 0.2679842, 
    0.3917858, 0.2786627, 0.1066356, 0.1622901, 0.1772232, 0.2119788, 
    0.2525946, 0.3091679, 0.2747456, 0.2373682, 0.2390236,
  0.2396239, 0.198552, 0.359724, 0.2287095, 0.2703872, 0.1976201, 0.2789714, 
    0.362149, 0.2467112, 0.1976573, 0.08905097, 0.2065463, 0.237152, 
    0.2061242, 0.2599405, 0.1467917, 0.2812458, 0.3129689, 0.1647381, 
    0.3209449, 0.2748538, 0.3263509, 0.2099526, 0.06558834, 0.1197799, 
    0.4149279, 0.3106381, 0.3298766, 0.277487,
  0.2419476, 0.271347, 0.1750976, 0.06401429, 0.1027072, 0.1225685, 
    0.09450018, 0.1704559, 0.1551043, 0.1916475, 0.2142574, 0.1630323, 
    0.1631553, 0.2909999, 0.2878424, 0.2776053, 0.3287221, 0.2720599, 
    0.2316363, 0.3081598, 0.2020005, 0.1407718, 0.1049603, 0.1445977, 
    0.1115404, 0.0716546, 0.1287548, 0.1242414, 0.2791852,
  0.1342186, 0.1304251, 0.1266316, 0.1228381, 0.1190445, 0.115251, 0.1114575, 
    0.1663201, 0.1777494, 0.1891787, 0.2006079, 0.2120372, 0.2234665, 
    0.2348958, 0.2365174, 0.2434325, 0.2503477, 0.2572629, 0.264178, 
    0.2710932, 0.2780083, 0.2153808, 0.2008298, 0.1862789, 0.171728, 
    0.1571771, 0.1426262, 0.1280753, 0.1372534,
  0.0712808, 0.07508865, 0.09017976, 0.08627804, 0.02635114, 0.00301721, 
    0.00527258, 0.001867392, 0.05636868, 0.09020048, 0.08217612, 0.09332283, 
    0.09142008, 0.1393723, 0.07190426, 0.1845375, 0.2852411, 0.2849573, 
    0.2903343, 0.227829, 0.4417018, 0.3356352, 0.2865046, 0.2219317, 
    0.1158931, 0.09146987, 0.09277428, 0.1561879, 0.1086293,
  0.3198772, 0.2948547, 0.2912145, 0.05993674, 0.1407664, 0.1826242, 
    0.2744268, 0.2544754, 0.3232637, 0.3262052, 0.3548848, 0.4473639, 
    0.3196267, 0.2489998, 0.2017588, 0.2961356, 0.210161, 0.1877657, 
    0.1696519, 0.3283329, 0.2845413, 0.3685673, 0.3279666, 0.2842376, 
    0.3463817, 0.1476292, 0.1078126, 0.1757858, 0.2581936,
  0.2863515, 0.2450706, 0.292331, 0.286041, 0.2979868, 0.2903906, 0.3089789, 
    0.3440546, 0.2681619, 0.2939469, 0.3933404, 0.2750254, 0.3174405, 
    0.2694504, 0.2675053, 0.2074211, 0.2243441, 0.2684382, 0.2268279, 
    0.275408, 0.3199635, 0.2543034, 0.2849715, 0.2333157, 0.249261, 
    0.2536312, 0.2388917, 0.2228034, 0.2882378,
  0.3178728, 0.2495639, 0.2823265, 0.3051242, 0.2948323, 0.3132006, 
    0.2675509, 0.3105143, 0.2450815, 0.2431469, 0.2808087, 0.2528005, 
    0.3143277, 0.1763719, 0.2807835, 0.1973166, 0.1476277, 0.2489421, 
    0.2468517, 0.268102, 0.2638788, 0.2325201, 0.2008921, 0.2502153, 
    0.1240043, 0.1759148, 0.1640976, 0.1725988, 0.2444233,
  0.2557767, 0.2266233, 0.1402048, 0.1610479, 0.1641939, 0.1385023, 0.173807, 
    0.1438241, 0.1679214, 0.146587, 0.1299327, 0.1651399, 0.08772518, 
    0.1279675, 0.1746223, 0.2368531, 0.1567171, 0.2378125, 0.1643003, 
    0.1722519, 0.2510127, 0.2457501, 0.1895303, 0.1571799, 0.03087723, 
    0.09366576, 0.1444155, 0.2035529, 0.2583374,
  0.04472141, 0.009064987, 0.0009593302, 0.02131135, 0.02974446, 0.07664558, 
    0.05069601, 0.03023242, 0.04356996, 0.068524, 0.002844721, 0.001036686, 
    0.03018887, 0.05650691, 0.08550255, 0.1565283, 0.1504181, 0.1279127, 
    0.1052124, 0.1309997, 0.08016549, 0.05669371, 0.01739224, 0.01538327, 
    0.0310665, 0.1333563, 0.1034388, 0.07104891, 0.0631846,
  2.444057e-05, 5.213523e-09, -3.894589e-05, 0.004495005, 0.05860791, 
    0.02810607, 0.03720134, 0.01852377, 0.01354008, 0.002019476, 
    3.112232e-06, 9.207248e-06, 0.02975223, 0.06272616, 0.02413063, 
    0.01095826, 0.1150435, 0.03145799, 0.1076505, 0.0564822, 0.05577606, 
    0.001597212, 1.824762e-06, 0.0003237851, 0.002373047, 0.005937437, 
    0.05309101, 0.05118385, 0.01539217,
  3.700059e-07, 6.473929e-07, 0.0002021888, 0.12887, 0.04263043, 0.04917568, 
    0.04744345, 0.07609729, 0.04611778, 0.01719037, 0.01738703, 0.02022122, 
    0.1873433, 0.1084062, 0.07644475, 0.04821117, 0.03596679, 0.01748822, 
    0.008221581, 0.008850987, 0.0001223269, 7.15111e-07, 3.43869e-07, 
    0.01615565, 0.000757842, -1.026642e-05, 0.04614817, 0.006618615, 
    6.319534e-05,
  9.093983e-06, 0.04700384, 0.02140508, 0.04951011, 0.02297786, 0.03375065, 
    0.01247046, 0.03373182, 0.06110634, 0.1657875, 0.03538435, 0.02472793, 
    0.1209379, 0.04389954, 0.02366083, 0.03137815, 0.02397347, 0.008877786, 
    0.003168387, 0.0008245771, 0.0001426345, 0.002402568, 0.02409528, 
    0.03468252, 0.02353899, 0.008346973, 0.01216512, 0.003535288, 0.000121668,
  0.09360344, 0.121434, 0.1494053, 0.5103624, 0.01440822, 0.002655181, 
    0.116506, 0.04465931, 0.0241325, 0.02509554, 0.02187876, 0.02214887, 
    0.08592492, 0.04755, 0.05620164, 0.1555692, 0.1401654, 0.1564773, 
    0.2297099, 0.2214804, 0.1147882, 0.1352637, 0.1926076, 0.07689819, 
    0.02670129, 0.04481631, 0.09664709, 0.2065616, 0.2287297,
  4.370584e-05, 0.0001239991, 1.853994e-07, 0.04331736, 0.005353959, 
    0.02180435, 0.2730501, 0.1222666, 0.4158033, 0.03723255, 0.1087651, 
    0.07377833, 0.03208279, 0.03403243, 0.02013978, 0.02747439, 0.010538, 
    0.002797632, 0.01725696, 0.007929699, 0.02070923, 0.06200601, 0.01177301, 
    0.007109323, 0.02944078, 0.03192951, -8.158109e-05, 8.023191e-07, 
    5.898886e-05,
  1.748188e-06, 7.95521e-05, 7.251871e-05, 2.974701e-06, 0.000242558, 
    5.955664e-05, 0.03912271, 0.2875643, 0.298427, 0.1380702, 0.04974111, 
    0.05457314, 0.02804822, 0.02872448, 0.05965412, 0.02158966, 0.03301325, 
    0.02162733, 1.080048e-05, 1.010038e-06, 0.001260877, 0.0061426, 
    0.02761705, 0.01351041, 0.0305935, 0.0287404, 0.003848872, 9.138794e-06, 
    2.778269e-06,
  0.000429887, 0.0006079909, 0.01295487, 0.03358236, -6.655246e-05, 
    4.631254e-07, -3.413072e-05, 4.569365e-07, 0.01259538, 0.08408369, 
    0.1505588, 0.0769262, 0.1243407, 0.09819002, 0.131549, 0.2117161, 
    0.08051648, 0.0956331, 0.0539213, 6.011417e-05, 0.003371964, 
    0.0002663335, 0.02105867, 0.04378808, 0.03749653, 0.04950252, 0.0754793, 
    0.05990358, 0.005350763,
  0.04285323, 0.08713896, 0.07686506, 0.1185513, 0.04386221, 0.01751729, 
    0.04482519, 0.06516504, 0.1403266, 0.152209, 0.1004653, 0.1178706, 
    0.1019595, 0.1728064, 0.1693928, 0.1545098, 0.1463452, 0.1779698, 
    0.1268081, 0.08481475, 0.05767938, 0.01401897, 0.09053945, 0.1345523, 
    0.1484703, 0.1603312, 0.2149495, 0.1731029, 0.1453779,
  0.1753576, 0.09823967, 0.2083788, 0.2233125, 0.3027179, 0.292627, 0.278089, 
    0.3013885, 0.1756976, 0.1645606, 0.1940332, 0.1998822, 0.2526547, 
    0.4385566, 0.2052368, 0.2058713, 0.2544945, 0.2633857, 0.3798257, 
    0.2437487, 0.1475948, 0.1419974, 0.1646072, 0.2374474, 0.2505085, 
    0.3154736, 0.2928056, 0.2475042, 0.2350677,
  0.2425976, 0.1623146, 0.452762, 0.2495054, 0.3833849, 0.1763407, 0.2691121, 
    0.3236094, 0.2578969, 0.1382182, 0.1228501, 0.2248386, 0.2085948, 
    0.1534574, 0.246217, 0.1400691, 0.2739806, 0.364988, 0.1441436, 
    0.3282321, 0.303126, 0.3043588, 0.2602482, 0.1169707, 0.122616, 0.408255, 
    0.348652, 0.3349984, 0.3046175,
  0.293837, 0.3322507, 0.2293331, 0.09673965, 0.1262362, 0.1629551, 
    0.1591236, 0.1516425, 0.1257854, 0.2135779, 0.1679524, 0.224553, 
    0.2419288, 0.2855199, 0.2523985, 0.2827301, 0.2925228, 0.2596511, 
    0.2096046, 0.2598795, 0.20816, 0.1589552, 0.1188307, 0.1478063, 
    0.09166197, 0.08040835, 0.1043485, 0.1789563, 0.3375504,
  0.1592852, 0.1587761, 0.158267, 0.1577579, 0.1572489, 0.1567398, 0.1562307, 
    0.1805606, 0.1966947, 0.2128287, 0.2289627, 0.2450967, 0.2612307, 
    0.2773647, 0.3243211, 0.3261608, 0.3280006, 0.3298404, 0.3316802, 
    0.3335199, 0.3353597, 0.2369409, 0.2194762, 0.2020115, 0.1845468, 
    0.167082, 0.1496173, 0.1321526, 0.1596925,
  0.07618497, 0.07596207, 0.09071589, 0.08780678, 0.05200276, 0.03786549, 
    0.02833865, 0.03140046, 0.08548263, 0.09370319, 0.1045043, 0.1095205, 
    0.1200909, 0.1370653, 0.06660247, 0.1984944, 0.2788662, 0.2958152, 
    0.2756163, 0.2305274, 0.4636271, 0.3580842, 0.3040294, 0.2392144, 
    0.1174693, 0.09508719, 0.1093741, 0.1626102, 0.09748238,
  0.2930869, 0.2709732, 0.2759939, 0.05134571, 0.1516754, 0.1939054, 
    0.3004006, 0.2884204, 0.3221162, 0.3401144, 0.3786857, 0.462667, 
    0.3078805, 0.2567413, 0.2043259, 0.2837394, 0.2119089, 0.2075848, 
    0.1673197, 0.3825119, 0.3320531, 0.350307, 0.2815689, 0.2858258, 
    0.3446551, 0.1158974, 0.105072, 0.1736175, 0.3199679,
  0.3047284, 0.2707191, 0.314294, 0.3586163, 0.3490745, 0.3199688, 0.3222653, 
    0.3946178, 0.2688271, 0.3690541, 0.3994727, 0.3050027, 0.3362154, 
    0.2537308, 0.3183853, 0.2621451, 0.2349757, 0.2616402, 0.2354596, 
    0.3339474, 0.3122896, 0.2532593, 0.3023876, 0.2277284, 0.2855189, 
    0.2614491, 0.2906407, 0.2462773, 0.320906,
  0.3388169, 0.2907534, 0.2963921, 0.321927, 0.3312503, 0.3314441, 0.287439, 
    0.3436204, 0.2951066, 0.2798349, 0.3046473, 0.2704033, 0.2814198, 
    0.2185837, 0.2801888, 0.2081663, 0.2178241, 0.243346, 0.2607603, 
    0.3186656, 0.2922147, 0.2863975, 0.2197035, 0.2605596, 0.1247852, 
    0.1942701, 0.2073374, 0.2869006, 0.3190905,
  0.2965122, 0.2744955, 0.2091085, 0.2568475, 0.2166381, 0.1991876, 
    0.1855227, 0.1511774, 0.1849861, 0.1707039, 0.1900466, 0.1888736, 
    0.09558254, 0.14879, 0.1889932, 0.2587595, 0.1918708, 0.2494155, 
    0.1977357, 0.1960324, 0.2636363, 0.2725899, 0.1978341, 0.1655923, 
    0.04152941, 0.1161317, 0.2142741, 0.3072173, 0.3307005,
  0.061173, 0.02754022, 0.0002332215, 0.03178235, 0.04711728, 0.08028948, 
    0.07146133, 0.07620514, 0.09662422, 0.1324147, 0.000460525, 1.017582e-05, 
    0.02614455, 0.1458672, 0.1091344, 0.1591518, 0.149475, 0.1377707, 
    0.1668051, 0.1406872, 0.09062269, 0.08181216, 0.05739446, 0.01702402, 
    0.0313907, 0.1345741, 0.1343474, 0.1073391, 0.08477859,
  0.0006307834, 5.303095e-09, -3.571974e-05, 0.005814321, 0.05501902, 
    0.0377283, 0.09296606, 0.1391459, 0.1658697, 0.006301678, 3.920962e-08, 
    2.488724e-08, 0.02271358, 0.06961032, 0.05726441, 0.01732509, 0.1052874, 
    0.03764132, 0.1013552, 0.0863437, 0.09367665, 0.02498443, 0.00536391, 
    0.0004127602, 0.001068673, 0.03443292, 0.05360417, 0.1336788, 0.05003422,
  4.312892e-06, 5.837049e-06, 6.402964e-05, 0.05369364, 0.04760396, 
    0.05823007, 0.06933107, 0.08411618, 0.04957619, 0.03460601, 0.0177358, 
    0.02787969, 0.2003965, 0.09904063, 0.079065, 0.03799313, 0.03251395, 
    0.02000671, 0.0152907, 0.0226136, 0.003425331, 0.0001131168, 
    1.666698e-07, 0.01853858, 0.0001263019, -4.243816e-06, 0.04318836, 
    0.01833214, 0.001844908,
  0.001462281, 0.05958731, 0.01489566, 0.03148524, 0.03337872, 0.03956139, 
    0.01267484, 0.0300403, 0.05889635, 0.1557634, 0.03493551, 0.02170999, 
    0.1047611, 0.03518454, 0.02200239, 0.02485449, 0.02125967, 0.01940115, 
    0.01282391, 0.008712421, 0.0009506488, 0.002189543, 0.01156321, 
    0.04021746, 0.02503577, 0.007179108, 0.01635111, 0.008817083, 0.001907357,
  0.110934, 0.1076327, 0.1343116, 0.4420601, 0.001713521, 0.005031927, 
    0.08345053, 0.03695064, 0.01627813, 0.02207241, 0.01945384, 0.01946424, 
    0.06896959, 0.04015234, 0.04659612, 0.1316298, 0.1213267, 0.1423489, 
    0.1996251, 0.1872363, 0.1033571, 0.1141104, 0.1916623, 0.0800509, 
    0.02504086, 0.04112037, 0.07926039, 0.1830181, 0.2074114,
  9.011597e-06, 1.73026e-05, 4.14064e-08, 0.0305468, 0.004167138, 
    0.009279437, 0.2563413, 0.1287902, 0.3903761, 0.03489736, 0.0909822, 
    0.06400787, 0.02771376, 0.02760244, 0.01889375, 0.02852137, 0.02192413, 
    0.01413877, 0.02148838, 0.02231547, 0.01420982, 0.06407991, 0.01312075, 
    0.007994494, 0.03860923, 0.05198781, 0.004611186, 2.792436e-07, 
    1.759929e-05,
  1.488526e-06, 1.866695e-05, 4.086375e-05, 1.277933e-06, 8.762677e-05, 
    7.12374e-06, 0.02773554, 0.2567676, 0.3116795, 0.1323296, 0.0480662, 
    0.05299543, 0.0259683, 0.02765756, 0.04228713, 0.02723046, 0.03209761, 
    0.08148096, 0.0003042181, 3.047718e-07, 0.0005296161, 0.003173182, 
    0.02841889, 0.01216147, 0.02865921, 0.03584332, 0.04046752, 0.0003728799, 
    1.474587e-06,
  0.0001045185, 0.0005834518, 0.00725449, 0.07845761, -4.907788e-05, 
    1.082694e-07, -1.816161e-05, 4.509777e-07, 0.01531518, 0.08266941, 
    0.1511213, 0.08699935, 0.1267367, 0.1195547, 0.1464708, 0.2102852, 
    0.0776717, 0.1179199, 0.08369935, -4.901174e-05, 0.0007374536, 
    0.0001380259, 0.02373009, 0.04979552, 0.0395553, 0.05351884, 0.1066385, 
    0.08779556, 0.009050288,
  0.07799996, 0.09212509, 0.09968976, 0.1029575, 0.03531394, 0.01458192, 
    0.03382919, 0.0648907, 0.1352848, 0.1166309, 0.09045617, 0.1073755, 
    0.133407, 0.2183645, 0.1805998, 0.160183, 0.1807491, 0.1872779, 
    0.1680666, 0.1017032, 0.03955677, 0.01216571, 0.09134822, 0.1491802, 
    0.1458468, 0.1859856, 0.272742, 0.1835607, 0.1410583,
  0.1650737, 0.1322701, 0.1983174, 0.229325, 0.2895413, 0.2765652, 0.2814663, 
    0.2569577, 0.182976, 0.1526029, 0.189784, 0.2308957, 0.2923459, 
    0.4565641, 0.2421446, 0.2297929, 0.2784806, 0.2709022, 0.4148748, 
    0.244492, 0.21067, 0.1625339, 0.1561885, 0.2975922, 0.2672586, 0.2862929, 
    0.3604952, 0.3294352, 0.2746058,
  0.2338355, 0.197515, 0.4693961, 0.3693068, 0.3142444, 0.149825, 0.2810897, 
    0.3248116, 0.2577342, 0.1540039, 0.1569857, 0.2948001, 0.2127889, 
    0.183615, 0.2497743, 0.1790338, 0.3046472, 0.3424569, 0.1981234, 
    0.3371717, 0.3398778, 0.3508301, 0.2906707, 0.1093093, 0.131161, 
    0.4487142, 0.3593158, 0.3313876, 0.302333,
  0.3828615, 0.4033649, 0.2966847, 0.1960951, 0.1406837, 0.209952, 0.2202869, 
    0.1927059, 0.1945576, 0.2314924, 0.1488042, 0.3233904, 0.2849782, 
    0.3194553, 0.2676592, 0.3195936, 0.2961008, 0.2977239, 0.2638597, 
    0.2236262, 0.1929874, 0.1498078, 0.1476891, 0.1505651, 0.100465, 
    0.1004447, 0.1217748, 0.1913524, 0.4103503,
  0.1759438, 0.1774538, 0.1789638, 0.1804739, 0.1819839, 0.1834939, 
    0.1850039, 0.2077958, 0.2253419, 0.242888, 0.2604341, 0.2779801, 
    0.2955263, 0.3130724, 0.3567401, 0.3554063, 0.3540724, 0.3527386, 
    0.3514047, 0.3500708, 0.348737, 0.2583512, 0.240629, 0.2229067, 
    0.2051845, 0.1874622, 0.16974, 0.1520177, 0.1747358,
  0.08203961, 0.06799297, 0.08251683, 0.08659883, 0.06875537, 0.07437186, 
    0.07345548, 0.06551317, 0.1282548, 0.1025442, 0.1141679, 0.1141279, 
    0.134542, 0.1183382, 0.05774022, 0.195823, 0.2924675, 0.2941795, 
    0.2543571, 0.2160921, 0.5133983, 0.380771, 0.2982916, 0.248996, 
    0.1259176, 0.0991228, 0.1201934, 0.1603016, 0.09570849,
  0.3014432, 0.2663286, 0.2513016, 0.05629902, 0.163739, 0.1997162, 0.242084, 
    0.3136636, 0.3456519, 0.3624935, 0.3978293, 0.443414, 0.3057848, 
    0.270859, 0.2517673, 0.3375781, 0.2613709, 0.2242695, 0.2039498, 
    0.4366036, 0.3998759, 0.3068892, 0.287076, 0.3047761, 0.3447757, 
    0.1616883, 0.0829335, 0.1312709, 0.3067495,
  0.3638736, 0.3284988, 0.4242383, 0.4087986, 0.3884094, 0.3326479, 
    0.3101495, 0.4221729, 0.2636665, 0.3983908, 0.3788533, 0.3197421, 
    0.3998714, 0.3072114, 0.4152443, 0.3526746, 0.3116623, 0.3218061, 
    0.308708, 0.4636244, 0.3004422, 0.2338918, 0.3274692, 0.223963, 
    0.2937298, 0.2611579, 0.3005927, 0.3125721, 0.3984076,
  0.3049237, 0.2577946, 0.2674662, 0.3052876, 0.3248911, 0.3313854, 
    0.3133547, 0.3190832, 0.2838649, 0.307907, 0.286576, 0.2872213, 
    0.3077109, 0.2494465, 0.3269478, 0.2410613, 0.3157593, 0.3033321, 
    0.2972185, 0.4356259, 0.3804087, 0.2868622, 0.2358276, 0.2686857, 
    0.1257842, 0.2197464, 0.3083215, 0.2835865, 0.3153569,
  0.3147412, 0.2560363, 0.1899468, 0.2143542, 0.2464467, 0.1698759, 0.184293, 
    0.1602298, 0.16639, 0.1572733, 0.1643088, 0.1553898, 0.07917149, 
    0.160671, 0.2276768, 0.294806, 0.2637723, 0.2728257, 0.2107789, 
    0.2246714, 0.2533109, 0.2877769, 0.2382276, 0.1784131, 0.04861082, 
    0.1586212, 0.3127484, 0.3046092, 0.3047679,
  0.1568641, 0.05676162, -3.556393e-05, 0.07434141, 0.08009174, 0.08400072, 
    0.07390482, 0.2265565, 0.1417264, 0.158109, -1.72929e-05, 2.402808e-05, 
    0.01707201, 0.1454181, 0.1365629, 0.1868445, 0.1954718, 0.1528533, 
    0.15408, 0.1792526, 0.09806459, 0.1818979, 0.08627917, 0.02228395, 
    0.03913837, 0.1496857, 0.1692128, 0.1534415, 0.1404928,
  0.07456677, -7.404271e-08, -1.697031e-05, 0.04760884, 0.0564165, 
    0.06580555, 0.1239519, 0.2298811, 0.2344232, 0.006792587, 4.686243e-08, 
    3.881086e-08, 0.07109506, 0.1999191, 0.1237953, 0.0463328, 0.08531121, 
    0.02769515, 0.11118, 0.09772803, 0.1784479, 0.2041942, 0.08322363, 
    -0.0004709911, 0.000690188, 0.01885851, 0.06540006, 0.1326355, 0.2445291,
  0.001093703, 3.587716e-05, 3.288302e-05, 0.02242344, 0.05054222, 
    0.05060461, 0.06294368, 0.08707622, 0.04937719, 0.0456269, 0.01767562, 
    0.03325573, 0.2021835, 0.1075092, 0.07984652, 0.0366155, 0.03511066, 
    0.02533735, 0.02187512, 0.03258964, 0.02837576, 0.05275864, -6.26243e-05, 
    0.0172945, 6.020489e-05, 7.092723e-07, 0.06224363, 0.02180693, 0.01611231,
  0.01573234, 0.08555542, 0.01415998, 0.02614426, 0.03704266, 0.04380819, 
    0.01622719, 0.03119703, 0.05888176, 0.1455053, 0.03318712, 0.02015977, 
    0.0820464, 0.03182547, 0.02256108, 0.0212037, 0.0174783, 0.01414017, 
    0.0134141, 0.02274843, 0.002016739, 0.001533027, 0.006143028, 0.07419441, 
    0.02553776, 0.007592671, 0.02387384, 0.03240998, 0.01782402,
  0.1251601, 0.1004003, 0.1073836, 0.3971114, -0.0004848779, 0.01474863, 
    0.0596663, 0.03060048, 0.01215909, 0.02270043, 0.01884687, 0.01929491, 
    0.05554276, 0.03596977, 0.04211761, 0.1062979, 0.09591477, 0.1214579, 
    0.1668447, 0.1627345, 0.09311395, 0.1032152, 0.1855358, 0.07344235, 
    0.02512878, 0.04177045, 0.06769036, 0.1651254, 0.190206,
  6.361122e-07, 5.350932e-07, 2.140921e-08, 0.01906074, 0.003928986, 
    0.004397914, 0.242807, 0.1287129, 0.3472699, 0.03252513, 0.07432164, 
    0.05385631, 0.02739413, 0.02698835, 0.02244844, 0.03602117, 0.07890671, 
    0.07766392, 0.0163796, 0.04599919, 0.01345136, 0.06366232, 0.01591922, 
    0.01044082, 0.04070146, 0.08567808, 0.05073491, 9.376993e-07, 6.001553e-06,
  1.304998e-06, 2.373989e-06, 0.001167762, 5.534475e-07, 8.163814e-05, 
    -5.811163e-06, 0.0170717, 0.2149164, 0.2954024, 0.1150557, 0.05221134, 
    0.04884546, 0.0252593, 0.02864267, 0.03566711, 0.0367431, 0.03737906, 
    0.1113949, 0.02142905, 4.577736e-08, 0.0003049256, 0.00185987, 0.0346514, 
    0.01332176, 0.03047636, 0.03840508, 0.07898514, 0.009337289, 8.93933e-07,
  0.001110561, 0.001223014, 0.00533763, 0.1320565, -3.37136e-05, 
    5.165495e-08, -1.580826e-06, 4.798786e-07, 0.01589886, 0.08096499, 
    0.1500922, 0.0919214, 0.1570755, 0.1445073, 0.1670927, 0.2058295, 
    0.092525, 0.168384, 0.1342094, -4.051447e-05, 2.351388e-05, 4.928145e-05, 
    0.02547498, 0.04926597, 0.0391778, 0.112425, 0.1217443, 0.1133781, 
    0.01220274,
  0.07616664, 0.1457938, 0.1237263, 0.1151405, 0.03788573, 0.01158252, 
    0.02528585, 0.07395785, 0.1423568, 0.1075738, 0.08722847, 0.1023271, 
    0.1428791, 0.2577081, 0.177729, 0.1895005, 0.199782, 0.213048, 0.2223709, 
    0.0829726, 0.03402762, 0.01535539, 0.09243704, 0.1449977, 0.1348975, 
    0.2170938, 0.3196287, 0.2114705, 0.1804466,
  0.1532152, 0.1445084, 0.1911179, 0.1956381, 0.2404798, 0.2245611, 0.309939, 
    0.2002272, 0.1737956, 0.1513908, 0.1648789, 0.2744251, 0.2888425, 
    0.4814216, 0.2776279, 0.2321593, 0.3219257, 0.25381, 0.4250508, 
    0.2241145, 0.1948303, 0.1867854, 0.1728986, 0.3143097, 0.2853727, 
    0.2466528, 0.5153209, 0.3588771, 0.3152865,
  0.2537118, 0.2766117, 0.5318269, 0.3938281, 0.3000612, 0.2037164, 
    0.3403691, 0.3502395, 0.2438213, 0.2149682, 0.2072929, 0.3097396, 
    0.292562, 0.2221637, 0.2838821, 0.2476309, 0.2800088, 0.3297847, 
    0.1696546, 0.3307047, 0.3461825, 0.3755262, 0.3187284, 0.1297562, 
    0.119537, 0.4141769, 0.3688061, 0.3242279, 0.3216553,
  0.4148746, 0.3947733, 0.2063844, 0.2348591, 0.1390782, 0.2395373, 
    0.2153922, 0.2558154, 0.2084407, 0.2753047, 0.331525, 0.3071029, 
    0.3211385, 0.3589697, 0.2717421, 0.3232224, 0.3366477, 0.3224712, 
    0.2623208, 0.2761457, 0.2759947, 0.1881519, 0.1629674, 0.1661588, 
    0.1164274, 0.1240022, 0.09975233, 0.2169119, 0.4107077,
  0.1763586, 0.1788832, 0.1814077, 0.1839323, 0.1864569, 0.1889815, 
    0.1915061, 0.2246802, 0.2425663, 0.2604525, 0.2783387, 0.2962248, 
    0.314111, 0.3319972, 0.3615003, 0.3587998, 0.3560992, 0.3533986, 
    0.350698, 0.3479975, 0.3452969, 0.2735529, 0.2558427, 0.2381325, 
    0.2204224, 0.2027122, 0.185002, 0.1672918, 0.1743389,
  0.08330896, 0.06205471, 0.07104078, 0.08360831, 0.09332044, 0.1190267, 
    0.1115231, 0.1353769, 0.1369025, 0.1047072, 0.1160468, 0.1173795, 
    0.1463819, 0.09730852, 0.05888563, 0.1999524, 0.294988, 0.2786012, 
    0.2382745, 0.2416332, 0.5433554, 0.4148774, 0.2987111, 0.223396, 
    0.1136606, 0.08964467, 0.1360068, 0.179336, 0.1048075,
  0.3214, 0.2844055, 0.2296449, 0.05638606, 0.1848701, 0.2159761, 0.1838363, 
    0.3317488, 0.3733881, 0.3903856, 0.4138238, 0.4181159, 0.2874851, 
    0.2619351, 0.2670628, 0.3632205, 0.3519754, 0.2947283, 0.2696981, 
    0.4172461, 0.3984477, 0.311615, 0.3116365, 0.3214802, 0.3845513, 
    0.1976042, 0.1326298, 0.09517792, 0.2885612,
  0.4265862, 0.3207289, 0.4175475, 0.4310397, 0.434403, 0.3669153, 0.3077672, 
    0.4189579, 0.3375817, 0.4276633, 0.4312152, 0.3380273, 0.4326022, 
    0.4037816, 0.4116656, 0.3901263, 0.337565, 0.4494316, 0.4718605, 
    0.4119092, 0.2801492, 0.2349897, 0.2928668, 0.247481, 0.330261, 
    0.3184689, 0.3154352, 0.3717213, 0.4298067,
  0.2433611, 0.2273239, 0.2261559, 0.2741545, 0.3053564, 0.3217429, 
    0.3295766, 0.2969635, 0.2696255, 0.2682657, 0.243793, 0.2808893, 
    0.2816476, 0.290884, 0.3914351, 0.3035712, 0.3877025, 0.3465868, 
    0.3759524, 0.4217923, 0.3417927, 0.3032535, 0.2729884, 0.3025985, 
    0.1420409, 0.2546976, 0.3820117, 0.2608763, 0.2548983,
  0.284082, 0.2062201, 0.113872, 0.1751954, 0.196483, 0.1673006, 0.1674025, 
    0.152216, 0.1937811, 0.182132, 0.1498037, 0.1069944, 0.04422174, 
    0.1167606, 0.2790841, 0.2766842, 0.2399255, 0.2804386, 0.1496749, 
    0.1894422, 0.2136562, 0.2696408, 0.1668102, 0.2279122, 0.04725415, 
    0.1422643, 0.2636658, 0.227293, 0.2618833,
  0.2714844, 0.147476, -5.572653e-05, 0.09965703, 0.1252294, 0.08843037, 
    0.2606451, 0.241529, 0.1905673, 0.07064289, -4.085043e-05, 0.000101651, 
    0.009526741, 0.113008, 0.09473585, 0.1596432, 0.1502409, 0.1047126, 
    0.1201989, 0.1323369, 0.08713427, 0.1581398, 0.09949489, 0.02216776, 
    0.03779055, 0.1935141, 0.1799814, 0.1526656, 0.2474778,
  0.2736689, -0.0001208469, -5.847875e-06, 0.04929538, 0.0754111, 0.06998478, 
    0.1226498, 0.2238287, 0.1990965, 0.01440808, 4.09408e-10, 4.450801e-09, 
    0.1184264, 0.2561063, 0.1183576, 0.09981892, 0.07955453, 0.0370669, 
    0.1206303, 0.1314292, 0.2191796, 0.3243612, 0.1671493, 0.00529705, 
    0.002574567, 0.01098044, 0.07741981, 0.1682706, 0.5027745,
  0.01123349, 0.00365536, 1.140384e-05, 0.01214196, 0.05253672, 0.057163, 
    0.06471141, 0.08532964, 0.07054497, 0.07100061, 0.02135189, 0.05627968, 
    0.1978747, 0.1019832, 0.07635816, 0.04927916, 0.0968876, 0.06309575, 
    0.03636681, 0.06908336, 0.1627261, 0.1512153, 0.008268531, 0.01269825, 
    2.283236e-05, 3.178619e-07, 0.09686688, 0.05186382, 0.1975255,
  0.07879589, 0.1963869, 0.01080794, 0.02189863, 0.04170938, 0.04218539, 
    0.03021268, 0.0357687, 0.05265338, 0.1335738, 0.04109748, 0.02258546, 
    0.07757128, 0.03344141, 0.03736362, 0.02139839, 0.01484026, 0.01073362, 
    0.008938954, 0.02272002, 0.0251982, 0.001533796, 0.00186945, 0.05605341, 
    0.01777319, 0.01186842, 0.04199517, 0.08287425, 0.07742352,
  0.1314692, 0.1022112, 0.07552379, 0.3739646, -0.0005927157, 0.01540824, 
    0.04013932, 0.02973633, 0.009638736, 0.02747354, 0.02186056, 0.02249755, 
    0.04999255, 0.05069313, 0.03996329, 0.09241229, 0.08859712, 0.1015832, 
    0.1392252, 0.1260341, 0.08677651, 0.09276846, 0.1646231, 0.06849863, 
    0.03013923, 0.04668197, 0.05966071, 0.1393766, 0.1819727,
  -2.124694e-07, -1.147265e-06, 1.480931e-08, 0.01570448, 0.00298712, 
    0.004074647, 0.2082229, 0.1167296, 0.3060956, 0.02434468, 0.06600805, 
    0.05657459, 0.03258007, 0.03059856, 0.0310284, 0.05066151, 0.1745837, 
    0.1660223, 0.06962329, 0.07088955, 0.01501182, 0.07114318, 0.02086409, 
    0.01214926, 0.04502227, 0.1118806, 0.09886758, -1.480114e-05, 2.997655e-06,
  1.193232e-06, -1.07482e-05, 0.003373003, 2.945689e-07, 5.562343e-06, 
    -1.678395e-06, 0.01062605, 0.2175712, 0.2767744, 0.08490705, 0.05593747, 
    0.04949982, 0.02862971, 0.03817261, 0.03959213, 0.04356652, 0.05148574, 
    0.1172609, 0.07314806, 1.614842e-07, 0.0001635221, 0.001313987, 
    0.02764335, 0.02169193, 0.03879874, 0.04568056, 0.1147666, 0.07512209, 
    -2.95691e-06,
  0.002433044, 0.002508076, 0.002070117, 0.1916235, -2.959573e-05, 
    3.358695e-08, 1.129963e-05, 4.385398e-07, 0.01295042, 0.07065592, 
    0.1532457, 0.08976341, 0.2197199, 0.1926908, 0.2057664, 0.2015604, 
    0.1670603, 0.2297229, 0.313288, -1.272011e-06, 2.109351e-06, 
    9.733132e-06, 0.0102538, 0.04418607, 0.05004732, 0.1372203, 0.1658054, 
    0.1673397, 0.02074802,
  0.08872404, 0.1290595, 0.1575623, 0.0695217, 0.03976561, 0.004385082, 
    0.0193029, 0.09010168, 0.1221589, 0.09172752, 0.07247405, 0.08377918, 
    0.1458162, 0.3048073, 0.194768, 0.3148196, 0.3433364, 0.3524158, 
    0.2179552, 0.05998161, 0.02779328, 0.01117056, 0.1008178, 0.1326682, 
    0.1136372, 0.2523538, 0.3473126, 0.2284462, 0.2390737,
  0.1449536, 0.07580628, 0.1679283, 0.1795691, 0.2015563, 0.1796456, 
    0.2574477, 0.2081422, 0.1441459, 0.1624678, 0.1448776, 0.3029846, 
    0.2691537, 0.5060894, 0.3376263, 0.2816398, 0.3528352, 0.2402374, 
    0.3986765, 0.2318985, 0.1644563, 0.1718611, 0.2074724, 0.2888751, 
    0.3151721, 0.2235364, 0.5870371, 0.3777871, 0.2993082,
  0.3637545, 0.380839, 0.5728278, 0.4027712, 0.3489835, 0.2229696, 0.3783103, 
    0.3454776, 0.2267032, 0.2921609, 0.2547744, 0.3247086, 0.3677038, 
    0.2765089, 0.2392983, 0.2829391, 0.3167826, 0.3291017, 0.2232553, 
    0.3739876, 0.3569096, 0.4258552, 0.3275711, 0.1512748, 0.1224861, 
    0.3823604, 0.377387, 0.3281539, 0.3865241,
  0.4487998, 0.428105, 0.2643251, 0.2442356, 0.2038878, 0.2288018, 0.2166498, 
    0.27961, 0.2638391, 0.3374988, 0.3977396, 0.3222591, 0.3156563, 0.383204, 
    0.3102138, 0.317788, 0.4502756, 0.4046703, 0.3275289, 0.3963339, 
    0.3194701, 0.1698889, 0.164261, 0.2178244, 0.1919537, 0.1325021, 
    0.1100376, 0.2496139, 0.4060051,
  0.1922017, 0.1938577, 0.1955137, 0.1971697, 0.1988257, 0.2004817, 
    0.2021378, 0.2230725, 0.2415055, 0.2599386, 0.2783716, 0.2968046, 
    0.3152377, 0.3336707, 0.3620894, 0.3581122, 0.3541349, 0.3501576, 
    0.3461804, 0.3422032, 0.3382259, 0.2785932, 0.2624814, 0.2463696, 
    0.2302578, 0.214146, 0.1980342, 0.1819224, 0.1908769,
  0.09728622, 0.06295542, 0.0611972, 0.07840845, 0.1084026, 0.1554109, 
    0.1681722, 0.1648664, 0.1395117, 0.1129761, 0.1151599, 0.1370627, 
    0.1666395, 0.08102035, 0.055025, 0.1695853, 0.2882846, 0.2635512, 
    0.2325062, 0.2478379, 0.5658612, 0.4720827, 0.2985639, 0.177272, 
    0.1134606, 0.09629396, 0.1677843, 0.1846892, 0.122446,
  0.3315383, 0.2972835, 0.2046876, 0.05490723, 0.1991511, 0.2359552, 
    0.1139921, 0.3426331, 0.3979037, 0.3867839, 0.4287585, 0.3898543, 
    0.2625022, 0.2585195, 0.2989006, 0.361467, 0.4097755, 0.318913, 
    0.2911327, 0.3898485, 0.4112295, 0.358268, 0.3583207, 0.3405012, 
    0.413574, 0.2415098, 0.2040716, 0.1062448, 0.2808718,
  0.3978991, 0.3564672, 0.3828109, 0.3197799, 0.3898989, 0.4977019, 
    0.3278296, 0.428818, 0.3930993, 0.3446762, 0.4105962, 0.3695578, 
    0.462116, 0.4947417, 0.4329331, 0.4191185, 0.463138, 0.4550065, 
    0.4491903, 0.2915059, 0.196286, 0.1745756, 0.2678748, 0.3058377, 
    0.3890316, 0.3839463, 0.3135659, 0.3739813, 0.4472049,
  0.1835547, 0.1830775, 0.2137364, 0.272216, 0.3121574, 0.3330002, 0.3251337, 
    0.2729465, 0.254658, 0.2262287, 0.1900761, 0.2227325, 0.2601109, 
    0.2460098, 0.336844, 0.2316584, 0.2927438, 0.3345167, 0.2998011, 
    0.3050272, 0.2935941, 0.2632061, 0.2526118, 0.3383081, 0.1257192, 
    0.2674937, 0.347839, 0.2216812, 0.1816822,
  0.2731953, 0.1426316, 0.07662715, 0.1671076, 0.171598, 0.1477372, 
    0.1213024, 0.1396241, 0.2245007, 0.1502643, 0.1537716, 0.07022617, 
    0.0209748, 0.1032302, 0.2955672, 0.207573, 0.2124131, 0.2691215, 
    0.120367, 0.1479256, 0.2143122, 0.2325245, 0.1807758, 0.2427031, 
    0.04168149, 0.09863828, 0.2174538, 0.2198402, 0.2711334,
  0.2332164, 0.1758035, 5.732075e-06, 0.07462044, 0.09845728, 0.1195986, 
    0.1495384, 0.08100181, 0.1284369, 0.01755826, -7.318069e-06, 
    8.065265e-06, 0.007111096, 0.05137775, 0.08483481, 0.1313366, 0.1087548, 
    0.08160558, 0.1196519, 0.1139574, 0.08417404, 0.1420814, 0.1047924, 
    0.02565016, 0.03508775, 0.120685, 0.09530281, 0.1628586, 0.2036506,
  0.5719216, -8.878505e-06, -4.415546e-07, 0.03231655, 0.08199596, 0.0362652, 
    0.05520987, 0.09051578, 0.1323227, 0.00397808, 1.236998e-08, 
    3.740311e-09, 0.05257892, 0.1654318, 0.07884607, 0.09206183, 0.1092734, 
    0.08195592, 0.08839708, 0.07073544, 0.1108297, 0.3191435, 0.4191681, 
    0.00649534, 0.006887213, 0.01212146, 0.03355726, 0.115631, 0.2706923,
  0.2634633, 0.05529023, 1.911769e-06, 0.009165622, 0.0464277, 0.06113408, 
    0.09505016, 0.0820729, 0.06083326, 0.09500928, 0.04578404, 0.05398129, 
    0.1871694, 0.09449632, 0.07055319, 0.04292654, 0.04458752, 0.03200384, 
    0.01844706, 0.04162484, 0.1238345, 0.3656968, 0.03160128, 0.00677513, 
    5.161632e-06, 8.728907e-08, 0.07032105, 0.0575987, 0.3397927,
  0.2720981, 0.2385009, 0.005643215, 0.02324216, 0.04717734, 0.1516787, 
    0.1205857, 0.1187301, 0.03582406, 0.1245222, 0.06389014, 0.03117246, 
    0.1091298, 0.05056293, 0.03196932, 0.02363914, 0.01886171, 0.01384422, 
    0.01292111, 0.02100227, 0.08597622, 0.02253539, 0.00360171, 0.02132403, 
    0.006694854, 0.0458906, 0.06078118, 0.1628359, 0.232838,
  0.1232634, 0.08280474, 0.0518341, 0.3346717, -0.0003714475, 0.01688465, 
    0.03426623, 0.03138477, 0.005955819, 0.03054229, 0.02199884, 0.04846367, 
    0.07308061, 0.0442865, 0.04095764, 0.07251426, 0.07590939, 0.09600443, 
    0.1410738, 0.1067338, 0.1066154, 0.08551787, 0.1442993, 0.05041735, 
    0.06142011, 0.05992213, 0.06693979, 0.1357049, 0.1694476,
  -2.803305e-07, -2.755011e-07, 1.155452e-08, 0.009604444, 0.001315454, 
    0.01414678, 0.1600204, 0.105772, 0.2516536, 0.02448, 0.0690391, 
    0.06294779, 0.03500706, 0.03195795, 0.03112164, 0.04250262, 0.1007148, 
    0.2236956, 0.3612813, 0.07860845, 0.0240253, 0.08230517, 0.06719524, 
    0.03488553, 0.04241977, 0.1065598, 0.2261422, 0.005666592, -1.104069e-06,
  1.121455e-06, -0.000124841, 0.006002349, 2.113769e-07, 7.984322e-07, 
    -2.985143e-06, 0.006888578, 0.2495899, 0.265876, 0.05517905, 0.09507485, 
    0.05661807, 0.08209601, 0.06120073, 0.08895907, 0.07308931, 0.07033686, 
    0.1421355, 0.3653249, 0.0002024623, 0.0001154501, 0.0007089571, 
    0.01715201, 0.08440508, 0.04121076, 0.09147857, 0.1149083, 0.2510894, 
    -0.0004063357,
  0.001059254, 0.002183171, 0.001012401, 0.2501248, -2.508708e-05, 
    2.449921e-08, 1.192782e-05, 3.611103e-07, 0.01068132, 0.06605004, 
    0.1476864, 0.1035195, 0.2373054, 0.2291931, 0.2568891, 0.2185068, 
    0.3520115, 0.2397023, 0.4348424, -4.473421e-06, 2.034556e-06, 
    -9.552943e-05, 0.003167439, 0.0495506, 0.09463645, 0.2841251, 0.2122388, 
    0.158361, 0.03892102,
  0.0686477, 0.1330527, 0.08814064, 0.04781751, 0.0400963, 0.001000401, 
    0.01525033, 0.08888358, 0.1043302, 0.08859308, 0.05902718, 0.07360268, 
    0.1600639, 0.3732726, 0.3240717, 0.4107186, 0.4372369, 0.469398, 
    0.2990804, 0.05702625, 0.03478351, 0.01908557, 0.1067628, 0.1265283, 
    0.1074848, 0.2783109, 0.328709, 0.2147419, 0.2692578,
  0.164496, 0.07075509, 0.1333537, 0.1560356, 0.1886341, 0.135416, 0.2128888, 
    0.1858084, 0.113198, 0.1722762, 0.1280416, 0.2759209, 0.2384436, 
    0.4380957, 0.3337866, 0.4280885, 0.3428505, 0.2225575, 0.3642511, 
    0.1911002, 0.1102616, 0.149045, 0.2702195, 0.2977901, 0.344863, 
    0.1997205, 0.5142438, 0.3815652, 0.2880194,
  0.5182992, 0.4400854, 0.5883374, 0.4223408, 0.4425892, 0.3296894, 
    0.4596061, 0.3742176, 0.2416926, 0.4038263, 0.2666487, 0.4186357, 
    0.4126573, 0.3199518, 0.2465029, 0.3778269, 0.35761, 0.3878014, 
    0.3374922, 0.4612742, 0.4552454, 0.5011159, 0.3771829, 0.2490074, 
    0.2299382, 0.3748, 0.4085608, 0.3262765, 0.4653973,
  0.5731998, 0.5152426, 0.4893726, 0.4961754, 0.4758643, 0.3258255, 
    0.2840427, 0.3692157, 0.4330096, 0.4325732, 0.4227887, 0.360719, 
    0.3738634, 0.5012763, 0.5278811, 0.5058793, 0.5958735, 0.572967, 
    0.4306061, 0.4707635, 0.4795137, 0.2447456, 0.2355799, 0.3007193, 
    0.2317791, 0.1505629, 0.1211045, 0.3050085, 0.518512,
  0.1948528, 0.1955874, 0.1963221, 0.1970567, 0.1977914, 0.198526, 0.1992607, 
    0.2117471, 0.2298008, 0.2478545, 0.2659082, 0.2839618, 0.3020155, 
    0.3200692, 0.3488154, 0.3428899, 0.3369645, 0.331039, 0.3251135, 
    0.319188, 0.3132626, 0.2668405, 0.2539777, 0.2411148, 0.228252, 
    0.2153891, 0.2025262, 0.1896634, 0.194265,
  0.151472, 0.05482477, 0.05889042, 0.06910955, 0.1174842, 0.1716924, 
    0.2059315, 0.1856968, 0.1220644, 0.1151452, 0.1112903, 0.1469263, 
    0.2123072, 0.06439742, 0.05570725, 0.1815118, 0.3120275, 0.2495791, 
    0.2180061, 0.2367573, 0.5789504, 0.4944092, 0.3034737, 0.1635034, 
    0.1162637, 0.1117811, 0.2187276, 0.1902462, 0.1511501,
  0.3207509, 0.2756155, 0.1948447, 0.02618298, 0.1896525, 0.2501747, 
    0.05170862, 0.3521373, 0.4373785, 0.3763792, 0.4126728, 0.3745924, 
    0.2183394, 0.2239273, 0.3037959, 0.3948661, 0.4246727, 0.329438, 
    0.3108859, 0.3986254, 0.4592191, 0.3500494, 0.3443791, 0.3462492, 
    0.4272231, 0.2727102, 0.2070214, 0.1436408, 0.2549107,
  0.4166008, 0.3943366, 0.289497, 0.2522808, 0.314844, 0.5367137, 0.3009505, 
    0.4369909, 0.4154646, 0.2537161, 0.3519561, 0.3285162, 0.4574956, 
    0.5286415, 0.4348383, 0.4062627, 0.5707286, 0.4715098, 0.3992496, 
    0.2044159, 0.1470059, 0.11512, 0.2233737, 0.2582149, 0.3955085, 
    0.4386395, 0.3411765, 0.3667045, 0.4861306,
  0.1419566, 0.15077, 0.2058188, 0.2694597, 0.2930774, 0.3608749, 0.3168457, 
    0.2759758, 0.2284244, 0.2003509, 0.1485031, 0.1932448, 0.2347629, 
    0.1983524, 0.2796654, 0.2019826, 0.1798033, 0.2855298, 0.262386, 
    0.2418932, 0.2541939, 0.2391946, 0.2344857, 0.3499528, 0.1400077, 
    0.267197, 0.28796, 0.2081262, 0.1358867,
  0.2462664, 0.09139904, 0.04859645, 0.1545394, 0.1717477, 0.1420598, 
    0.1259361, 0.1430962, 0.1839013, 0.07907825, 0.1121198, 0.04147402, 
    0.007885793, 0.08083565, 0.3063281, 0.195391, 0.1867336, 0.2152693, 
    0.1120596, 0.1378767, 0.2197102, 0.207667, 0.1656398, 0.2518564, 
    0.02773374, 0.08547837, 0.189188, 0.2217973, 0.2478313,
  0.08337957, 0.1331204, -0.0001207297, 0.03623012, 0.1006652, 0.07795601, 
    0.05467223, 0.02377812, 0.04001994, 0.005376615, -1.670755e-06, 
    -1.164689e-06, 0.005520649, 0.02600296, 0.0673025, 0.1139248, 0.09104127, 
    0.07535335, 0.09268355, 0.1084712, 0.09950116, 0.0870624, 0.14454, 
    0.02748151, 0.0415485, 0.08828179, 0.06270459, 0.06764948, 0.06814925,
  0.2828578, -0.0007074515, -5.958593e-08, 0.01976838, 0.02392315, 
    0.01108506, 0.01127169, 0.02658982, 0.04681809, 0.003883939, 
    1.054496e-08, 2.96755e-09, 0.01769259, 0.1207287, 0.06861106, 0.06168263, 
    0.1214444, 0.04392862, 0.04320163, 0.02628364, 0.0328479, 0.1486463, 
    0.2349551, 0.006488728, 0.009015142, 0.01288059, 0.00637976, 0.04060861, 
    0.07476919,
  0.465885, 0.1599049, 8.957132e-08, 0.01649832, 0.02744432, 0.02023157, 
    0.03485328, 0.05485233, 0.02190723, 0.04277431, 0.0239404, 0.02448548, 
    0.1486452, 0.06184954, 0.02888224, 0.01959533, 0.01013919, 0.006552672, 
    0.003083253, 0.009831758, 0.04055956, 0.2569112, 0.2069273, 0.003764657, 
    5.554497e-07, 5.473207e-08, 0.01546129, 0.009228948, 0.1295211,
  0.3359347, 0.1391686, 0.002297969, 0.02431043, 0.04887371, 0.04553749, 
    0.06791972, 0.05874753, 0.05105073, 0.0958927, 0.04165837, 0.03633947, 
    0.06502837, 0.02067134, 0.01457692, 0.01197876, 0.01444717, 0.01013147, 
    0.01221862, 0.02284369, 0.1327058, 0.2427831, 0.03792665, 0.008048793, 
    0.001793577, 0.04153723, 0.0169167, 0.03166545, 0.246604,
  0.07714098, 0.05810122, 0.03303315, 0.3156083, -0.0002155756, 0.01553931, 
    0.0382695, 0.01455699, 0.0009591303, 0.008986213, 0.009453107, 
    0.09999643, 0.04988672, 0.04459284, 0.03929109, 0.06662515, 0.06993818, 
    0.08268622, 0.1450071, 0.1353942, 0.1342257, 0.1306819, 0.1413302, 
    0.04426108, 0.02293243, 0.04433436, 0.06077238, 0.113314, 0.1314456,
  -2.117772e-07, -9.329019e-08, 1.030341e-08, 0.008866549, 0.0004280354, 
    0.05010273, 0.1527544, 0.07513566, 0.2209762, 0.04512094, 0.05585144, 
    0.05041556, 0.01690028, 0.01290351, 0.005696812, 0.008609978, 0.02593642, 
    0.08830779, 0.2907642, 0.2376665, 0.08132529, 0.08359775, 0.004776907, 
    0.006138148, 0.01583914, 0.02629235, 0.1540092, 0.1306916, -3.205393e-05,
  1.074607e-06, 5.505273e-05, 0.00291415, 1.739243e-07, 5.151651e-07, 
    -8.488718e-07, 0.0006831869, 0.2820134, 0.2631213, 0.03462398, 
    0.08683048, 0.1003125, 0.1148972, 0.07544307, 0.1277711, 0.1015642, 
    0.07643538, 0.08263135, 0.3605435, 0.036899, 6.734538e-05, 0.001414517, 
    0.008090446, 0.05017033, 0.02449385, 0.07365064, 0.1088438, 0.1417052, 
    -0.000391536,
  0.0001679652, 0.00128776, 0.000131606, 0.3014453, -4.155982e-05, 
    2.215672e-08, 1.06733e-05, 2.961769e-07, 0.008651647, 0.06001472, 
    0.1574082, 0.137916, 0.361852, 0.2078298, 0.2924715, 0.3157615, 
    0.4602533, 0.263638, 0.3778146, -0.0001020863, 1.363466e-06, 
    0.0008827558, 0.0014704, 0.1085671, 0.1726817, 0.2506618, 0.1382245, 
    0.1633007, 0.1527871,
  0.08645558, 0.0804019, 0.0502264, 0.03745959, 0.02512994, 8.593064e-05, 
    0.01479327, 0.06875179, 0.1091127, 0.1000439, 0.04747528, 0.06178712, 
    0.2544249, 0.4385315, 0.4277074, 0.5543044, 0.5643436, 0.5633941, 
    0.3067625, 0.06027294, 0.02880016, 0.02410387, 0.1158289, 0.1250017, 
    0.1030452, 0.3006313, 0.253205, 0.2544169, 0.3191301,
  0.1696512, 0.08865927, 0.1290024, 0.1285794, 0.1595968, 0.1057177, 
    0.1889887, 0.1473828, 0.0935495, 0.1482528, 0.1090742, 0.2513692, 
    0.256999, 0.4019026, 0.4005301, 0.4927758, 0.3519843, 0.2006893, 
    0.3369056, 0.1674328, 0.07687048, 0.1260891, 0.2175736, 0.2834074, 
    0.4435702, 0.1921445, 0.479993, 0.4099834, 0.3000909,
  0.4936979, 0.3637868, 0.5746059, 0.4161027, 0.4931384, 0.4137347, 
    0.4411897, 0.3666567, 0.2210015, 0.3454424, 0.2687859, 0.4750513, 
    0.4999123, 0.4596357, 0.3977863, 0.5262501, 0.5423355, 0.4287092, 
    0.3543631, 0.5385921, 0.5224198, 0.5506164, 0.3579988, 0.2934752, 
    0.2400745, 0.4049666, 0.4234225, 0.333066, 0.5808665,
  0.6789983, 0.4903946, 0.610113, 0.6501298, 0.7230231, 0.691236, 0.5472544, 
    0.6049132, 0.6622974, 0.6606581, 0.6691633, 0.6626302, 0.7440068, 
    0.829618, 0.7848232, 0.7403017, 0.7876721, 0.7865161, 0.7919394, 
    0.6809006, 0.5668297, 0.3320383, 0.1976843, 0.3741073, 0.320393, 
    0.1463208, 0.1808746, 0.4527749, 0.7183319,
  0.1568702, 0.156603, 0.1563359, 0.1560687, 0.1558015, 0.1555343, 0.1552672, 
    0.1648941, 0.181806, 0.198718, 0.2156299, 0.2325419, 0.2494538, 
    0.2663658, 0.3106571, 0.3044272, 0.2981973, 0.2919674, 0.2857375, 
    0.2795077, 0.2732778, 0.2344411, 0.2240262, 0.2136113, 0.2031965, 
    0.1927816, 0.1823667, 0.1719518, 0.1570839,
  0.1758619, 0.06834692, 0.04718192, 0.06710514, 0.08287159, 0.1537832, 
    0.1853707, 0.1565416, 0.09295134, 0.1149097, 0.07914707, 0.1210736, 
    0.2738522, 0.05655844, 0.06379407, 0.2408199, 0.3567107, 0.2683582, 
    0.2199895, 0.2062078, 0.5812964, 0.5094246, 0.3000543, 0.1617722, 
    0.1422976, 0.1158486, 0.2280562, 0.2007054, 0.1946462,
  0.2810569, 0.2399671, 0.1551634, 0.002613053, 0.1391032, 0.2279521, 
    0.01558301, 0.3415617, 0.4400302, 0.3501131, 0.3765396, 0.3737751, 
    0.1831083, 0.1830077, 0.2896765, 0.4318929, 0.4418248, 0.3587485, 
    0.3257998, 0.4234834, 0.466542, 0.3542925, 0.3078168, 0.3402171, 
    0.4220212, 0.2769518, 0.2258027, 0.1916383, 0.2692752,
  0.5005873, 0.3868446, 0.2039941, 0.1900674, 0.2559372, 0.4490071, 
    0.3568573, 0.4712854, 0.3956599, 0.1821247, 0.2919655, 0.2962492, 
    0.424319, 0.4898199, 0.4348169, 0.3955538, 0.5424349, 0.5175626, 
    0.3281546, 0.1474877, 0.1161183, 0.07602599, 0.1760948, 0.1835758, 
    0.3345734, 0.4606599, 0.3848363, 0.386744, 0.5210773,
  0.1091849, 0.130724, 0.1999369, 0.2612889, 0.3080927, 0.3576313, 0.3213765, 
    0.2673745, 0.2064272, 0.1743684, 0.1211755, 0.1648647, 0.1935679, 
    0.1882128, 0.2384153, 0.1957945, 0.1426993, 0.2495228, 0.2050723, 
    0.1983701, 0.204464, 0.2214623, 0.1991131, 0.3019018, 0.1323455, 
    0.2400292, 0.2466516, 0.1717097, 0.1137425,
  0.1968409, 0.05681221, 0.02692121, 0.1304626, 0.1400234, 0.1287282, 
    0.1066736, 0.09381744, 0.1063664, 0.03911518, 0.05826829, 0.02380493, 
    0.00185164, 0.05361634, 0.2718395, 0.1480219, 0.1279625, 0.1927662, 
    0.1126175, 0.1258248, 0.2129027, 0.197518, 0.1388404, 0.2692886, 
    0.01928471, 0.06487697, 0.1692006, 0.2031234, 0.202514,
  0.02282266, 0.05959606, 0.0002358957, 0.02227857, 0.06067599, 0.0503395, 
    0.02746588, 0.009526973, 0.01605344, 0.002546357, -4.237785e-07, 
    -7.562887e-07, 0.004402373, 0.01475515, 0.04165181, 0.09932513, 
    0.07815401, 0.09301714, 0.08405458, 0.1084908, 0.06035878, 0.0410348, 
    0.1104764, 0.01831398, 0.05792639, 0.06987045, 0.0390453, 0.02473781, 
    0.02599667,
  0.1063272, -0.0001002673, -2.30554e-08, 0.00504182, 0.0001690097, 
    0.001450194, 0.002229462, 0.007792335, 0.01447119, 0.0008273568, 
    8.405014e-09, 2.828845e-09, 0.008224263, 0.08389134, 0.04830704, 
    0.04616193, 0.05170606, 0.009212852, 0.02613202, 0.009821968, 
    0.007371245, 0.04786104, 0.1258586, 0.005710502, 0.01086775, 0.01819814, 
    0.00153729, 0.01300458, 0.02097315,
  0.2597151, 0.2999083, 2.430087e-07, 0.02853713, 0.01120433, 0.003609334, 
    0.01172202, 0.03814005, 0.007697537, 0.006314186, 0.02034635, 
    0.005369633, 0.1148657, 0.0318735, 0.007113214, 0.003759898, 0.001449671, 
    0.0006672264, 5.704183e-05, 0.001086842, 0.007740081, 0.09388878, 
    0.1819442, 0.001140585, 1.165463e-08, 4.535622e-08, -0.002248707, 
    0.001657963, 0.04469734,
  0.09813116, 0.07475897, 0.001471541, 0.01464283, 0.05146807, 0.01883575, 
    0.007447421, 0.01356072, 0.05228171, 0.06331859, 0.02646808, 0.01084189, 
    0.05789999, 0.008168408, 0.003376015, 0.0009385778, 0.003474557, 
    0.001271931, 0.006184881, 0.01326601, 0.07321888, 0.5542201, 0.3123464, 
    0.00399848, 0.0005808712, 0.004537097, 0.001788139, 0.007869572, 
    0.07410248,
  0.05763244, 0.0495728, 0.02433449, 0.3102084, -0.0001271527, 0.006347214, 
    0.05349112, 0.0028471, -0.001173316, 0.001264245, 0.004257513, 
    0.02088401, 0.03419126, 0.01759196, 0.01506142, 0.05943453, 0.04936815, 
    0.06366399, 0.08947369, 0.09289058, 0.04707957, 0.09185181, 0.20317, 
    0.03301858, 0.006632305, 0.01489893, 0.04371348, 0.08160685, 0.115598,
  -1.0142e-07, -1.499936e-08, 9.650109e-09, 0.005020908, 0.000170449, 
    0.05619903, 0.1386424, 0.02696915, 0.2285937, 0.02295723, 0.02706421, 
    0.02439615, 0.002621235, 0.003963377, 0.000761889, 0.0006757253, 
    0.006038873, 0.027133, 0.1346844, 0.4146937, 0.1886854, 0.07429373, 
    0.0004254903, -0.001223229, 0.004214784, 0.004648277, 0.06022971, 
    0.1750025, -2.079719e-05,
  1.042773e-06, 0.0005434785, 0.0009253918, 5.913201e-08, 4.281608e-07, 
    -1.127816e-07, -0.001175028, 0.2861376, 0.2588388, 0.0246408, 0.04436732, 
    0.1092578, 0.03014897, 0.01537173, 0.05586575, 0.01979173, 0.01484316, 
    0.01718007, 0.1663795, 0.130464, 2.863987e-05, 0.0008993449, 0.002807171, 
    0.006969507, 0.002695472, 0.007196472, 0.02594725, 0.06997573, 
    -0.0006208146,
  -0.0003001762, 0.0003053831, -0.0001721946, 0.3627845, -5.391194e-05, 
    2.018402e-08, 9.641991e-06, 2.688118e-07, 0.009572534, 0.05894575, 
    0.1795292, 0.1316436, 0.4573931, 0.2213626, 0.3166007, 0.4504717, 
    0.4344447, 0.1800726, 0.2707078, -0.000569976, 3.337926e-06, 0.009948395, 
    0.001445197, 0.1512989, 0.1644793, 0.1897012, 0.08421006, 0.1289482, 
    0.1978655,
  0.1138817, 0.05391433, 0.03726151, 0.02651612, 0.0124048, -1.882027e-05, 
    0.01198373, 0.06911759, 0.1026294, 0.09400312, 0.03999789, 0.05054571, 
    0.4319454, 0.5263203, 0.6862211, 0.652258, 0.62059, 0.582315, 0.2215389, 
    0.06172886, 0.02428118, 0.02547231, 0.1366837, 0.112805, 0.106304, 
    0.25521, 0.2183397, 0.1924611, 0.3151271,
  0.3442896, 0.1123292, 0.1032861, 0.1155539, 0.1386019, 0.07922357, 
    0.1595393, 0.1201312, 0.08942021, 0.142817, 0.09189312, 0.2535963, 
    0.2821794, 0.4451995, 0.4917199, 0.525711, 0.3460746, 0.1853674, 
    0.3152359, 0.1505351, 0.06460612, 0.08975792, 0.1544934, 0.2304569, 
    0.4520517, 0.174321, 0.4082365, 0.3760517, 0.357982,
  0.4694515, 0.3358745, 0.5297266, 0.3372689, 0.4836455, 0.4156707, 
    0.4572708, 0.3623741, 0.227707, 0.2451049, 0.259903, 0.4554838, 
    0.4505191, 0.484968, 0.4213334, 0.4476289, 0.447706, 0.3628608, 0.317798, 
    0.453874, 0.5584948, 0.5346997, 0.3191379, 0.3097863, 0.2823399, 
    0.3875195, 0.3884639, 0.3362488, 0.5793621,
  0.6735156, 0.4657592, 0.5469996, 0.5685727, 0.6399997, 0.6763134, 
    0.7088562, 0.7272457, 0.7722959, 0.8182368, 0.7310299, 0.7035984, 
    0.7676564, 0.7724437, 0.7337182, 0.7147665, 0.7223498, 0.7447305, 
    0.7564554, 0.7316545, 0.5530442, 0.4143726, 0.1764175, 0.5090266, 
    0.3339795, 0.127296, 0.1610596, 0.5099129, 0.7284623,
  0.1284978, 0.1314706, 0.1344433, 0.1374161, 0.1403888, 0.1433616, 
    0.1463344, 0.1427807, 0.1577725, 0.1727644, 0.1877562, 0.202748, 
    0.2177399, 0.2327317, 0.2363983, 0.2281164, 0.2198346, 0.2115527, 
    0.2032709, 0.194989, 0.1867071, 0.1827117, 0.173029, 0.1633462, 
    0.1536635, 0.1439808, 0.134298, 0.1246153, 0.1261196,
  0.1845847, 0.06501874, 0.04124848, 0.06716987, 0.06808913, 0.09941331, 
    0.1113235, 0.1182537, 0.0492877, 0.05554491, 0.05474397, 0.06374349, 
    0.2252508, 0.04670739, 0.09842148, 0.3221922, 0.3659617, 0.3292642, 
    0.2018663, 0.2114735, 0.5658338, 0.5380318, 0.3005307, 0.1614715, 
    0.1637844, 0.128512, 0.2433842, 0.2055509, 0.2524196,
  0.2396668, 0.1970159, 0.1331588, -0.002076382, 0.08703579, 0.2020386, 
    0.00735317, 0.3062405, 0.4392489, 0.3230649, 0.3321146, 0.3950489, 
    0.1345772, 0.1377226, 0.289425, 0.4775101, 0.4862003, 0.3747028, 
    0.3367281, 0.4676149, 0.4732859, 0.3653811, 0.2929818, 0.3035256, 
    0.4228235, 0.3165678, 0.25628, 0.2846913, 0.3058794,
  0.5612812, 0.3900776, 0.1539355, 0.1449783, 0.2036608, 0.3306946, 
    0.3853155, 0.5100023, 0.3259706, 0.1299031, 0.2347157, 0.2614949, 
    0.3865069, 0.4197726, 0.3959489, 0.4084237, 0.5003402, 0.5401309, 
    0.2601445, 0.1106306, 0.0979198, 0.05896465, 0.1407689, 0.1559489, 
    0.2690378, 0.4510759, 0.393701, 0.3854219, 0.5808198,
  0.09026996, 0.1230949, 0.1939045, 0.2463816, 0.3044255, 0.319657, 
    0.2866243, 0.2295814, 0.1758374, 0.1450764, 0.09707054, 0.1279282, 
    0.1424735, 0.168614, 0.180476, 0.1559017, 0.1244886, 0.2204838, 
    0.1461011, 0.1540326, 0.1635549, 0.1768686, 0.1442476, 0.2567277, 
    0.1044004, 0.1891218, 0.2162209, 0.1481006, 0.09574169,
  0.1424208, 0.03127898, 0.01547858, 0.1017403, 0.1024408, 0.1074743, 
    0.06451267, 0.05986921, 0.0829825, 0.02000404, 0.03514828, 0.01190163, 
    0.000644804, 0.03779735, 0.2162596, 0.1048294, 0.088888, 0.1706415, 
    0.1094354, 0.1038655, 0.1749417, 0.1680055, 0.09711567, 0.2721863, 
    0.01536792, 0.05248524, 0.1365813, 0.1501641, 0.1348931,
  0.00907144, 0.02407305, 0.0006285029, 0.00914345, 0.04277257, 0.03008873, 
    0.01771161, 0.005339608, 0.008936046, 0.001557666, -2.105369e-07, 
    -4.313866e-07, 0.003935924, 0.009586089, 0.03043782, 0.08304232, 
    0.06750544, 0.0949083, 0.07008929, 0.07573494, 0.03183659, 0.02151036, 
    0.04334149, 0.01845662, 0.05066349, 0.04481945, 0.02126676, 0.009162093, 
    0.01126105,
  0.04540529, 0.0005821273, -2.945886e-08, 0.002502748, -0.001889801, 
    0.0003659934, 0.0007536453, 0.003332828, 0.006421742, 0.0002940435, 
    5.732074e-09, 1.450926e-09, 0.00242931, 0.06694, 0.01375981, 0.01349676, 
    0.02855476, 0.002152387, 0.01695625, 0.004935286, 0.002205728, 
    0.01894292, 0.0541519, 0.01513926, 0.006148569, 0.02903773, 0.0006666686, 
    0.00496253, 0.008483893,
  0.1231533, 0.1793471, 1.866898e-07, 0.02380756, 0.00351787, 0.0004902777, 
    0.002534319, 0.02321823, 0.0009012501, -0.002167641, 0.01050413, 
    0.000622591, 0.06683268, 0.01258453, 0.001846419, 0.0005180937, 
    0.0004331036, 0.0002141065, 8.677116e-06, 0.0003750774, 0.00285405, 
    0.03469484, 0.07823324, 0.0002216727, 1.55615e-08, 4.018595e-08, 
    -0.00211201, 0.0008067553, 0.01794447,
  0.03937148, 0.05607187, 0.0007255389, 0.007794948, 0.009051945, 
    0.006759357, 0.001889911, 0.003987547, 0.04863559, 0.04407391, 
    0.003198188, 0.00655517, 0.04346251, 0.005738768, 0.0002984012, 
    4.192837e-05, 7.035666e-05, 2.389863e-05, 8.964774e-05, 0.001377237, 
    0.01355124, 0.2462744, 0.2962102, 0.001588632, 0.0001923389, 
    0.0008030977, 0.0001121013, 0.003739036, 0.02569671,
  0.04352068, 0.04702965, 0.01727971, 0.3195242, -6.589372e-05, 0.0003418633, 
    0.06423149, 0.0001531143, -0.001787656, 2.562419e-05, 0.0005618429, 
    0.004733036, 0.02382801, 0.006816289, 0.00146107, 0.03965424, 0.02338221, 
    0.0320676, 0.06153407, 0.04610131, 0.01656486, 0.04227303, 0.2449904, 
    0.01687332, 0.002263519, 0.003233098, 0.01171199, 0.04168916, 0.0928541,
  -2.620669e-08, 2.75707e-08, 9.464034e-09, 0.002892182, 5.341021e-05, 
    0.02501581, 0.08789416, 0.002403191, 0.2548555, 0.004696927, 0.009744643, 
    0.009583055, 3.353881e-05, 0.00119948, 1.67419e-05, 0.0001290104, 
    0.002008055, 0.008866213, 0.05100301, 0.2282797, 0.05250159, 0.06644987, 
    0.0001174129, -0.001776438, 0.001325297, 0.001013896, 0.02082951, 
    0.1364723, -4.058392e-06,
  1.019717e-06, 0.0009159778, 0.0004159342, -5.214942e-07, 3.792387e-07, 
    -6.90228e-09, -0.002966644, 0.2715399, 0.2603948, 0.01495397, 
    0.009789336, 0.0295297, 0.007622913, 0.002332875, 0.01051807, 0.0045423, 
    0.003635325, 0.004822348, 0.06384259, 0.09453814, 5.522367e-06, 
    0.000287375, 0.0009577625, 0.002132094, 0.0002043148, 0.001699861, 
    0.007185783, 0.02901129, 0.0004518252,
  -0.0006455004, -6.561014e-05, -7.691711e-05, 0.3767111, -5.575289e-05, 
    1.771866e-08, 8.970857e-06, 2.597025e-07, 0.01509114, 0.04833976, 
    0.1847133, 0.1426934, 0.4152979, 0.2031664, 0.301042, 0.4215336, 
    0.3728454, 0.1089234, 0.1949011, -0.001527733, 3.259735e-06, 0.02082597, 
    0.00165051, 0.1672446, 0.1133536, 0.1559265, 0.04937338, 0.09710307, 
    0.1607428,
  0.09903754, 0.04681642, 0.02647922, 0.02077976, 0.00336815, -6.233491e-06, 
    0.008399554, 0.06579655, 0.08858276, 0.09036814, 0.03654253, 0.04250879, 
    0.4617843, 0.5364229, 0.6473976, 0.6524091, 0.574407, 0.4587408, 
    0.1401289, 0.06177719, 0.02021207, 0.01935896, 0.1301349, 0.09708839, 
    0.1107756, 0.24596, 0.1859078, 0.1349495, 0.3087045,
  0.3390722, 0.1163395, 0.07906094, 0.1023859, 0.1231132, 0.06545755, 
    0.1339174, 0.09870682, 0.0862023, 0.1307755, 0.08821128, 0.2384795, 
    0.2877417, 0.4253229, 0.5354749, 0.4908079, 0.3297321, 0.1757958, 
    0.2898907, 0.1355644, 0.05660295, 0.08283329, 0.1467357, 0.1990244, 
    0.4979939, 0.1708274, 0.3437876, 0.28499, 0.4725924,
  0.4785314, 0.2929911, 0.478523, 0.2980411, 0.391381, 0.4267752, 0.3920604, 
    0.3311428, 0.1978231, 0.2053982, 0.2048319, 0.4053116, 0.4194649, 
    0.4896213, 0.3301191, 0.3561922, 0.3393258, 0.3118911, 0.259255, 
    0.3499279, 0.5304885, 0.4892305, 0.2811061, 0.2889227, 0.3025053, 
    0.3551391, 0.3317108, 0.3150065, 0.6047417,
  0.662185, 0.4054953, 0.4589642, 0.4338736, 0.5017503, 0.5811636, 0.6515051, 
    0.6536145, 0.7202498, 0.7821454, 0.6428874, 0.6821726, 0.6582134, 
    0.6588091, 0.6226616, 0.6056715, 0.5866997, 0.614947, 0.6146146, 
    0.6840222, 0.5214095, 0.388511, 0.2914492, 0.5795112, 0.2695397, 
    0.1346591, 0.1264676, 0.4995057, 0.6719211,
  0.0700592, 0.07063691, 0.07121462, 0.07179233, 0.07237004, 0.07294774, 
    0.07352545, 0.09955198, 0.1135503, 0.1275486, 0.141547, 0.1555453, 
    0.1695436, 0.183542, 0.1783181, 0.1733237, 0.1683293, 0.1633349, 
    0.1583406, 0.1533462, 0.1483518, 0.164725, 0.1551433, 0.1455617, 0.13598, 
    0.1263983, 0.1168167, 0.107235, 0.06959704,
  0.1635979, 0.05191122, 0.03725844, 0.0683798, 0.07440776, 0.04810651, 
    0.05846119, 0.06842825, 0.003048935, 0.004009211, 0.006635937, 
    0.04149742, 0.1719892, 0.03536854, 0.1463607, 0.3677615, 0.3477157, 
    0.3859498, 0.1664098, 0.2151254, 0.5502833, 0.5568498, 0.2653209, 
    0.1294992, 0.1913107, 0.1855772, 0.2475805, 0.2158878, 0.2784554,
  0.2154417, 0.1483559, 0.1183127, -0.001766584, 0.05675454, 0.1756903, 
    0.002484148, 0.2410125, 0.4383447, 0.2659083, 0.2785066, 0.411174, 
    0.09911273, 0.1020417, 0.3297589, 0.518374, 0.4735483, 0.3806971, 
    0.3213595, 0.4406885, 0.4800222, 0.3838298, 0.2752162, 0.270441, 
    0.4318581, 0.3531989, 0.2943996, 0.3512027, 0.2920791,
  0.5786644, 0.3898435, 0.1157764, 0.1054082, 0.1595979, 0.2529521, 
    0.3781774, 0.4629209, 0.2596014, 0.08604325, 0.1833192, 0.2254245, 
    0.3397321, 0.3456532, 0.3257472, 0.3467878, 0.4377888, 0.515299, 
    0.2046387, 0.08088342, 0.08688816, 0.04795132, 0.1129795, 0.1281087, 
    0.2347877, 0.4013249, 0.3853808, 0.3603276, 0.5342591,
  0.07522976, 0.1100103, 0.1686724, 0.2116542, 0.269673, 0.2575688, 
    0.2340894, 0.1801538, 0.1400877, 0.1074088, 0.07171082, 0.08929208, 
    0.09486067, 0.1151063, 0.1366006, 0.1201274, 0.1013301, 0.1801843, 
    0.09039212, 0.104717, 0.1264589, 0.1282169, 0.09825499, 0.2177595, 
    0.08275905, 0.1490074, 0.1773601, 0.1092028, 0.0802523,
  0.0969108, 0.0180153, 0.0101831, 0.07553931, 0.0653271, 0.07343207, 
    0.03571931, 0.03748116, 0.06749289, 0.009547734, 0.0146423, 0.005963818, 
    0.0003474209, 0.02540489, 0.1643984, 0.07665755, 0.06546271, 0.1318838, 
    0.08869255, 0.07088302, 0.1407414, 0.1243106, 0.06159419, 0.2499335, 
    0.01268116, 0.03849412, 0.08559027, 0.1008005, 0.08062088,
  0.005391149, 0.013802, 0.0003565093, 0.003469971, 0.01827424, 0.0194242, 
    0.01061769, 0.003579797, 0.006040455, 0.00110667, -1.689491e-07, 
    -2.67021e-07, 0.003570393, 0.00653164, 0.01931501, 0.06323352, 
    0.05448241, 0.07221162, 0.05317958, 0.04342252, 0.01667558, 0.01174505, 
    0.02289223, 0.01082357, 0.03896144, 0.02477633, 0.009971899, 0.005263375, 
    0.006201567,
  0.02472785, 0.001532098, -1.25671e-06, 0.001594752, -0.001825254, 
    0.0001760504, 0.0003774699, 0.00180353, 0.00363581, 0.000150508, 
    4.471502e-09, 1.344177e-09, 0.001300662, 0.02538566, 0.004498725, 
    0.003825113, 0.008260486, 0.0011246, 0.008990538, 0.002262962, 
    0.001093222, 0.009712229, 0.02707968, 0.01235839, 0.002167181, 
    0.04240981, 0.0003749681, 0.002464316, 0.004629469,
  0.06484129, 0.08230146, 1.42786e-07, 0.009763521, 0.0005983294, 
    0.0002180947, 0.0006266322, 0.01032077, 0.0001771239, -0.002768504, 
    0.003490747, 0.0001515018, 0.03308757, 0.004953372, 0.0005105886, 
    0.000154778, 0.0002483341, 0.0001220821, 1.442391e-06, 0.0002154355, 
    0.001496079, 0.01680302, 0.04085848, 0.0006927701, 3.507449e-08, 
    3.569624e-08, -0.001831706, 0.0005006234, 0.009593799,
  0.02162953, 0.05318834, 0.0007438284, 0.003472846, 0.001530669, 0.00337903, 
    0.0009354128, 0.001621918, 0.04365164, 0.04941144, 0.0006284533, 
    0.003025725, 0.02570529, 0.003280131, 8.599489e-05, 1.415188e-05, 
    1.982688e-05, 6.313491e-06, 1.664752e-05, 0.0001591967, 0.003366159, 
    0.1108548, 0.1473408, 0.0005894454, 7.028614e-05, 0.0003418862, 
    3.886122e-05, 0.002223235, 0.01348432,
  0.03792865, 0.04021942, 0.00704743, 0.306791, -3.063001e-05, 5.861513e-05, 
    0.05399226, 1.589456e-05, -0.001134965, 1.055331e-05, 4.116389e-05, 
    0.001963922, 0.01135088, 0.002573247, -3.58934e-05, 0.01783452, 
    0.01100455, 0.01704368, 0.03314135, 0.01773497, 0.007385311, 0.01968224, 
    0.206545, 0.01377618, 0.001036897, 0.001506236, 0.003101738, 0.01717241, 
    0.07209352,
  1.02244e-08, 1.860259e-08, 9.497556e-09, 0.001259879, 1.408857e-05, 
    0.004666796, 0.03714192, -0.0004557881, 0.2542894, 0.0004348091, 
    0.003584788, 0.003675018, -4.106382e-05, 0.0004398121, 8.262572e-06, 
    6.837906e-05, 0.0009983561, 0.00406667, 0.01990391, 0.1250525, 
    0.01542476, 0.05635059, 4.742858e-05, -0.001295559, 0.0003117414, 
    0.0004796814, 0.008621169, 0.09152549, -9.888237e-07,
  1.00266e-06, 0.0006359376, 0.0001868268, -9.026208e-07, 3.49597e-07, 
    4.027995e-10, -0.00200779, 0.2460127, 0.2477188, 0.01069644, 0.003032912, 
    0.01045955, 0.001900865, 0.0007461772, 0.004544992, 0.001797086, 
    0.001882175, 0.002477094, 0.03024894, 0.05937285, 2.56968e-06, 
    5.480801e-05, 0.0004810141, 0.001131105, 6.363571e-05, 0.0008352418, 
    0.003715388, 0.01095847, 0.0005002905,
  -0.0006617452, -9.32172e-05, -4.42957e-05, 0.3656584, -5.185092e-05, 
    1.765547e-08, 8.482953e-06, 2.554772e-07, 0.0100537, 0.03614398, 
    0.1753655, 0.1736167, 0.3399421, 0.1622923, 0.272578, 0.3139438, 
    0.2453085, 0.05289848, 0.1420312, -0.001876726, 2.833878e-06, 0.02409728, 
    0.0009135872, 0.1945083, 0.05084839, 0.08320695, 0.02274667, 0.06236001, 
    0.1638235,
  0.08411491, 0.04221055, 0.01704846, 0.01466356, 0.001171401, 3.568951e-06, 
    0.004490953, 0.06077865, 0.07353808, 0.09120362, 0.03143427, 0.03890138, 
    0.4626204, 0.4817391, 0.5438559, 0.6046128, 0.5324391, 0.3680565, 
    0.08967076, 0.05923732, 0.01634097, 0.01138612, 0.1200738, 0.08512232, 
    0.130004, 0.2483011, 0.1603232, 0.09711184, 0.2688766,
  0.3511528, 0.1075828, 0.05338072, 0.07797532, 0.1019516, 0.05764478, 
    0.1150344, 0.07436865, 0.08049466, 0.1214503, 0.07766411, 0.2201125, 
    0.2755585, 0.3645841, 0.4985292, 0.4125121, 0.2995455, 0.1686272, 
    0.2429264, 0.1222915, 0.04284919, 0.07841371, 0.1560551, 0.1662639, 
    0.4706891, 0.1594074, 0.2855357, 0.2332949, 0.4355261,
  0.4856592, 0.2325097, 0.4126404, 0.2466873, 0.2996531, 0.3880784, 
    0.3378824, 0.2765836, 0.1708814, 0.1813317, 0.1705386, 0.366988, 
    0.3726056, 0.4635521, 0.2665504, 0.3107522, 0.2748411, 0.2825834, 
    0.2365614, 0.2789935, 0.5071715, 0.4448833, 0.2478198, 0.2371508, 
    0.2703474, 0.3011689, 0.3001365, 0.3094095, 0.6114403,
  0.6418057, 0.3608042, 0.3893409, 0.3867677, 0.393964, 0.5059413, 0.5855312, 
    0.5849905, 0.638949, 0.676502, 0.589806, 0.5976524, 0.5497825, 0.5620858, 
    0.501848, 0.5051529, 0.4802448, 0.5471856, 0.5300862, 0.6038363, 
    0.4622464, 0.3043807, 0.2809014, 0.5034329, 0.2148865, 0.1261641, 
    0.1136087, 0.4396156, 0.6183649,
  0.03026015, 0.02723086, 0.02420156, 0.02117226, 0.01814296, 0.01511367, 
    0.01208437, 0.01826215, 0.02654504, 0.03482793, 0.04311081, 0.0513937, 
    0.05967659, 0.06795947, 0.08370099, 0.08631142, 0.08892185, 0.09153228, 
    0.09414271, 0.09675314, 0.09936357, 0.09856281, 0.09069879, 0.08283477, 
    0.07497075, 0.06710673, 0.05924271, 0.05137869, 0.03268359,
  0.137531, 0.02514263, 0.03225651, 0.09507416, 0.05994924, 0.01945458, 
    0.04012507, 0.02786679, 0.01440532, 0.01017361, 0.01058812, 0.01004431, 
    0.1249691, 0.02054236, 0.2189172, 0.3771136, 0.2844497, 0.3953283, 
    0.1668855, 0.2381677, 0.5164024, 0.5651529, 0.2465547, 0.1191978, 
    0.2254022, 0.240667, 0.2468019, 0.1990608, 0.2663544,
  0.1738404, 0.1087359, 0.1298583, -0.0009113225, 0.05175025, 0.1421361, 
    0.001691045, 0.1789038, 0.4287653, 0.1976484, 0.2330915, 0.4123705, 
    0.07340984, 0.08572299, 0.3585185, 0.489945, 0.4462291, 0.3681595, 
    0.302954, 0.4178764, 0.4441908, 0.3769837, 0.2674367, 0.2344683, 
    0.4003735, 0.396422, 0.353741, 0.3353191, 0.2375358,
  0.4926292, 0.3342451, 0.08364753, 0.07132013, 0.118558, 0.1938351, 
    0.3496634, 0.4022164, 0.2119393, 0.05643957, 0.13717, 0.1767253, 
    0.2845753, 0.2687251, 0.2362974, 0.2618336, 0.3555527, 0.4402909, 
    0.1576596, 0.06301466, 0.07213809, 0.03765273, 0.08837649, 0.09883601, 
    0.1891457, 0.3239457, 0.3613297, 0.3273022, 0.4506879,
  0.06020066, 0.08908387, 0.1347005, 0.1670288, 0.2218618, 0.2019603, 
    0.1836044, 0.1348145, 0.1061181, 0.07598175, 0.04906181, 0.0578695, 
    0.05452505, 0.06830198, 0.09496643, 0.08802041, 0.07589384, 0.1196715, 
    0.05332131, 0.06856392, 0.09305301, 0.08865271, 0.06508242, 0.1853525, 
    0.0568321, 0.1060276, 0.1301471, 0.08102197, 0.06156274,
  0.06099704, 0.01014755, 0.006627414, 0.04342284, 0.03758433, 0.04760003, 
    0.01962339, 0.0207231, 0.04594038, 0.004891892, 0.006692719, 0.003122213, 
    0.0002446797, 0.01749127, 0.123637, 0.04882554, 0.04264146, 0.09407109, 
    0.06276995, 0.04271853, 0.107835, 0.08361137, 0.03570497, 0.2208595, 
    0.008269561, 0.02284287, 0.05309909, 0.06957772, 0.04376669,
  0.003850205, 0.009432833, -0.0001032449, 0.001804954, 0.00645357, 
    0.009773869, 0.006628566, 0.002741918, 0.004566219, 0.0008542637, 
    -1.226081e-07, -1.847057e-07, 0.002985657, 0.004121229, 0.01202223, 
    0.04447807, 0.03567924, 0.05090211, 0.03329811, 0.02121277, 0.008636835, 
    0.00699708, 0.01527842, 0.007318375, 0.03060975, 0.01135508, 0.004923654, 
    0.003823094, 0.004058212,
  0.01610543, 0.001691538, -3.500113e-06, 0.001148929, -0.001363939, 
    0.0001123249, 0.0002309253, 0.00115164, 0.002400722, 9.452904e-05, 
    7.164727e-09, 1.33321e-09, 0.0008766084, 0.01160921, 0.002038642, 
    0.00184066, 0.003292175, 0.0007359359, 0.004361512, 0.0007822202, 
    0.0006811586, 0.006016043, 0.01768505, 0.01067432, 0.001085799, 
    0.04510019, 0.000245953, 0.001470326, 0.003011823,
  0.04150983, 0.03521562, 1.140304e-07, 0.004917676, 0.0002158841, 
    0.0001340009, 0.000295443, 0.003987311, 0.0001025137, -0.001712275, 
    0.001712619, 8.936467e-05, 0.01322206, 0.001543477, 0.0002018596, 
    7.971406e-05, 0.0001676497, 8.277241e-05, 2.773674e-07, 0.0001470552, 
    0.0009631212, 0.01025641, 0.02557189, 0.0003807685, 2.544548e-08, 
    3.471084e-08, -0.00123043, 0.0003536366, 0.006196555,
  0.01437175, 0.04396359, 0.0005823874, 0.001524606, 0.0006727932, 
    0.001822376, 0.0005924846, 0.0009610478, 0.03380376, 0.05335856, 
    0.0003088959, 0.001238543, 0.01174188, 0.00165455, 4.754822e-05, 
    7.755271e-06, 9.122368e-06, 2.917049e-06, 6.394757e-06, 7.327378e-05, 
    0.001637443, 0.06300907, 0.09882038, 0.001321694, -0.0002340331, 
    0.0001956524, 2.240567e-05, 0.001519964, 0.008838852,
  0.01999117, 0.02637942, 0.002491167, 0.2725923, -1.337103e-05, 
    2.986346e-05, 0.03326556, 8.476111e-06, -0.0004890776, 5.544728e-06, 
    -1.461411e-05, 0.001161827, 0.004795947, 0.001047925, -1.004542e-05, 
    0.007086243, 0.004754095, 0.007833209, 0.01595303, 0.007408712, 
    0.003237484, 0.00880372, 0.1652487, 0.0155558, 0.0003509828, 
    0.0007761329, 0.00113267, 0.007189163, 0.04371162,
  2.329858e-08, 3.256746e-08, 9.549616e-09, 0.0006789042, 1.918806e-06, 
    0.001649046, 0.01030086, -0.0004070209, 0.2094078, 0.000172444, 
    0.00144126, 0.001398908, -1.334553e-05, 0.0001332661, 4.337234e-06, 
    4.383182e-05, 0.0006185411, 0.002398206, 0.01086501, 0.0777852, 
    0.008230704, 0.04838206, 2.377706e-05, -0.0009381439, 9.461925e-05, 
    0.0002948704, 0.005067224, 0.04920079, -2.926317e-07,
  9.896564e-07, 0.000221122, 9.639763e-05, -1.442511e-06, 3.317178e-07, 
    5.500346e-10, -0.004411305, 0.2230837, 0.2273295, 0.005394469, 
    0.001627397, 0.005001086, 0.0009217476, 0.0003280943, 0.002726246, 
    0.001128904, 0.001243686, 0.001560756, 0.01839526, 0.04291041, 
    9.631605e-07, 2.47531e-05, 0.0009173838, 0.0007189135, 3.041661e-05, 
    0.0005231895, 0.002389233, 0.006203501, 0.0002322032,
  -0.0003711177, -0.000103183, -3.096563e-05, 0.329091, -4.969447e-05, 
    1.758558e-08, 8.103961e-06, 2.551251e-07, 0.005170337, 0.02463972, 
    0.164693, 0.1523244, 0.2627801, 0.1151923, 0.2173462, 0.2029968, 
    0.1307149, 0.02433658, 0.09938753, -0.001768771, 2.548599e-06, 
    0.02050032, 0.0007899478, 0.1654495, 0.02131846, 0.03693521, 0.007285497, 
    0.03191181, 0.1265461,
  0.05786698, 0.03778069, 0.01026542, 0.01027117, 0.0006055873, 3.003565e-06, 
    0.00243811, 0.05358332, 0.06101552, 0.08532482, 0.03084633, 0.03444763, 
    0.4337384, 0.4274294, 0.4291856, 0.5326432, 0.5138137, 0.2911961, 
    0.05672492, 0.05466264, 0.01203786, 0.006430745, 0.1128684, 0.07318874, 
    0.1252394, 0.2308254, 0.1178393, 0.06092219, 0.172046,
  0.3119053, 0.09581026, 0.03371965, 0.05100704, 0.08245726, 0.04309843, 
    0.09435336, 0.04963258, 0.07973816, 0.1118788, 0.06400566, 0.190014, 
    0.2536992, 0.291917, 0.390787, 0.3338622, 0.2679752, 0.1510242, 
    0.1812897, 0.1062615, 0.03225667, 0.07444184, 0.144218, 0.1419021, 
    0.3951676, 0.1602436, 0.2048879, 0.1811576, 0.3884591,
  0.4277725, 0.1838876, 0.3481946, 0.1781398, 0.241576, 0.3426277, 0.2877622, 
    0.2360296, 0.149483, 0.1624256, 0.1371467, 0.3251471, 0.3242564, 
    0.4539891, 0.219458, 0.2872077, 0.2290744, 0.2551198, 0.2064772, 
    0.2276087, 0.4352622, 0.4130967, 0.2208441, 0.2032852, 0.259716, 
    0.2564377, 0.2907939, 0.3024209, 0.5931555,
  0.6306549, 0.3167647, 0.3501431, 0.3549451, 0.3033126, 0.4290445, 
    0.5137381, 0.4952533, 0.5551118, 0.57412, 0.5332496, 0.4645289, 
    0.4275312, 0.4337626, 0.3796184, 0.3805573, 0.3843033, 0.4663758, 
    0.4368408, 0.4802997, 0.3901204, 0.2361192, 0.2355735, 0.4386821, 
    0.1792087, 0.0990536, 0.09075168, 0.3870497, 0.5428362,
  0.01819965, 0.01728851, 0.01637737, 0.01546622, 0.01455508, 0.01364394, 
    0.01273279, 0.01960096, 0.02411898, 0.02863699, 0.03315501, 0.03767302, 
    0.04219104, 0.04670905, 0.0525371, 0.05337297, 0.05420884, 0.05504472, 
    0.05588059, 0.05671647, 0.05755234, 0.0457851, 0.04134235, 0.03689961, 
    0.03245686, 0.02801412, 0.02357137, 0.01912862, 0.01892857,
  0.06960107, 0.03516091, 0.06850617, 0.09947531, 0.05304962, 0.03346336, 
    0.0335886, 0.005440895, 0.01532477, 0.01320067, 0.005269032, 0.00763805, 
    0.08682213, 0.01543187, 0.3392007, 0.3039553, 0.2585788, 0.4233045, 
    0.1706736, 0.3114015, 0.5089387, 0.6082933, 0.2458344, 0.1129313, 
    0.2313717, 0.2609248, 0.2578146, 0.1617857, 0.2710582,
  0.1218174, 0.09173458, 0.1194159, -0.0006789819, 0.02635951, 0.1044161, 
    0.001006061, 0.1473964, 0.3979247, 0.1748008, 0.2131043, 0.4101847, 
    0.05544093, 0.06194218, 0.3415412, 0.4586265, 0.4250912, 0.317061, 
    0.2932095, 0.3766904, 0.3849812, 0.3493571, 0.2663053, 0.2098261, 
    0.357989, 0.3902552, 0.3428388, 0.2950636, 0.183148,
  0.3886599, 0.2626729, 0.07052275, 0.05354904, 0.0907254, 0.1630552, 
    0.3233312, 0.3563901, 0.1800611, 0.04196935, 0.1069771, 0.1472759, 
    0.2341979, 0.2152414, 0.1775933, 0.1994904, 0.306209, 0.3695167, 
    0.1271532, 0.05068824, 0.05907646, 0.03039935, 0.07033113, 0.08080625, 
    0.1538961, 0.2721278, 0.3249394, 0.2976181, 0.3721658,
  0.04952171, 0.07167187, 0.1113186, 0.1414945, 0.1963311, 0.1658773, 
    0.1540294, 0.1053821, 0.0855334, 0.0571604, 0.03744159, 0.04111276, 
    0.03472256, 0.04367759, 0.06498589, 0.05752612, 0.05508486, 0.08244041, 
    0.03459389, 0.05104062, 0.07082071, 0.06350669, 0.04819838, 0.1665938, 
    0.04273712, 0.07560353, 0.09894786, 0.0634019, 0.04875526,
  0.04038524, 0.006574429, 0.005119926, 0.02555714, 0.02233977, 0.03144703, 
    0.01253051, 0.01247316, 0.0311033, 0.003022791, 0.004368943, 0.001898844, 
    0.000194562, 0.01080436, 0.09927227, 0.03328206, 0.02728557, 0.06538352, 
    0.04428257, 0.02631272, 0.08563509, 0.05037469, 0.02201156, 0.1961011, 
    0.004447956, 0.0116971, 0.03338045, 0.04834408, 0.0268912,
  0.003037544, 0.007313231, -0.0002102402, 0.001252675, 0.003758265, 
    0.005839967, 0.004524992, 0.002253173, 0.003737939, 0.0006992475, 
    -1.025876e-07, -1.275683e-07, 0.002851984, 0.00265789, 0.008040719, 
    0.0291448, 0.02309775, 0.02943762, 0.02003359, 0.01263981, 0.005219806, 
    0.004865183, 0.01172614, 0.006106337, 0.02442016, 0.005670774, 
    0.002758693, 0.00303733, 0.003056131,
  0.01193117, 0.0007346731, -4.451166e-06, 0.0009051611, -0.0008982868, 
    8.328023e-05, 0.0001640249, 0.0008408241, 0.001790021, 6.79741e-05, 
    7.092283e-09, 1.399362e-09, 0.0006773511, 0.006756092, 0.001450051, 
    0.001294194, 0.001741222, 0.000545139, 0.00233295, 0.0004579666, 
    0.000492951, 0.004304883, 0.0132088, 0.009909105, 0.0006564164, 
    0.04032856, 0.000181852, 0.001018794, 0.002224224,
  0.0303744, 0.01970896, 9.420509e-08, 0.003824725, 0.0001203308, 
    9.669257e-05, 0.0002001956, 0.001524325, 7.191647e-05, -0.0009082765, 
    0.0011635, 6.536367e-05, 0.005995339, 0.0006497351, 0.0001125222, 
    5.279764e-05, 0.0001277246, 6.332865e-05, 3.503577e-08, 0.0001129418, 
    0.0007109269, 0.00729915, 0.0185506, 0.001312097, 2.41687e-08, 
    3.374344e-08, -0.0007661426, 0.0002764741, 0.004571575,
  0.01082106, 0.03823053, 0.000316548, 0.0007205267, 0.0004344366, 
    0.001119407, 0.0004330243, 0.0006896588, 0.03202637, 0.06019191, 
    0.0002086821, 0.0005872, 0.005831015, 0.0008314417, 3.343091e-05, 
    5.553072e-06, 5.527988e-06, 1.867499e-06, 3.865963e-06, 4.583549e-05, 
    0.001052797, 0.04356652, 0.07509963, 0.004412466, -0.0002244499, 
    0.0001340587, 1.596886e-05, 0.001161048, 0.006554269,
  0.01159298, 0.01568969, 0.0009088295, 0.2235483, -6.47785e-06, 
    1.909725e-05, 0.02039087, 5.545095e-06, -0.0003253138, 3.928583e-06, 
    -2.409649e-06, 0.0008204444, 0.002197946, 0.0004961583, 5.221851e-06, 
    0.003118948, 0.002230119, 0.003373086, 0.007341073, 0.003355783, 
    0.001683239, 0.003968901, 0.1375015, 0.01983921, 0.0001391093, 
    0.0003839122, 0.0005286727, 0.003129031, 0.0270983,
  2.274609e-08, 3.25324e-08, 9.611282e-09, 0.0004299814, 1.879874e-07, 
    0.0009707732, 0.004672521, -0.0002446058, 0.1419594, 1.838198e-05, 
    0.0007082306, 0.0006807347, -1.225443e-06, 8.071311e-05, 2.948799e-06, 
    3.279344e-05, 0.0004217283, 0.001678464, 0.007454018, 0.05129585, 
    0.005599593, 0.04067175, 1.423251e-05, -0.0009717011, 4.43395e-05, 
    0.0002110233, 0.003533905, 0.02858509, -1.272929e-07,
  9.796501e-07, 0.0001104714, 6.422031e-05, -9.140434e-07, 3.179547e-07, 
    5.405683e-10, -0.005116168, 0.2084733, 0.2057733, 0.002653488, 
    0.001139013, 0.003328857, 0.000626069, 0.0001884724, 0.001953907, 
    0.0008107607, 0.0009365327, 0.001145872, 0.01301198, 0.03361657, 
    6.640955e-07, 0.0001268519, 0.007170723, 0.0005223694, 1.875581e-05, 
    0.0003778345, 0.001757918, 0.004427865, 4.266208e-05,
  -0.0003216909, -0.0001217898, -3.03964e-05, 0.2927364, -5.29305e-05, 
    1.752441e-08, 7.802682e-06, 2.537769e-07, 0.003010963, 0.0163517, 
    0.1484862, 0.1154637, 0.176878, 0.07820071, 0.1608899, 0.1233585, 
    0.06603269, 0.01102696, 0.07728302, -0.001901497, 2.482978e-06, 
    0.01662671, 0.003673556, 0.1299984, 0.01192923, 0.02075261, 0.003721796, 
    0.01934124, 0.102355,
  0.04111373, 0.03881125, 0.007342754, 0.006825244, 0.0003852355, 
    2.413732e-06, 0.001610641, 0.04865232, 0.05382321, 0.07950934, 
    0.03472765, 0.03186932, 0.3731572, 0.3684945, 0.3232263, 0.4271591, 
    0.4398433, 0.2146308, 0.03734579, 0.05214999, 0.00981951, 0.004037617, 
    0.1033848, 0.06909465, 0.1088941, 0.1903389, 0.07817137, 0.03492654, 
    0.1146104,
  0.2651533, 0.08298669, 0.02081861, 0.03943569, 0.06807432, 0.03391898, 
    0.07859844, 0.0371621, 0.08962573, 0.1011636, 0.05913972, 0.1686229, 
    0.2327188, 0.2256278, 0.2993994, 0.2319055, 0.235653, 0.1396005, 
    0.1307476, 0.09261195, 0.02568606, 0.06729385, 0.127028, 0.1137896, 
    0.3112134, 0.172707, 0.1358824, 0.1281758, 0.3446015,
  0.324662, 0.1462078, 0.2952139, 0.1191725, 0.2078142, 0.299406, 0.2465166, 
    0.2011569, 0.1317905, 0.1404374, 0.1203796, 0.2903301, 0.2841758, 
    0.4182116, 0.1986683, 0.2530291, 0.1923742, 0.2220796, 0.1854801, 
    0.1855115, 0.3745785, 0.3870451, 0.1967572, 0.1835297, 0.2249881, 
    0.2248962, 0.2806822, 0.2865295, 0.5236415,
  0.5930089, 0.3007986, 0.3021736, 0.3106067, 0.2454652, 0.3729887, 
    0.4391998, 0.4436946, 0.4674167, 0.4704157, 0.4469511, 0.3799439, 
    0.3526047, 0.3429368, 0.3061883, 0.2959377, 0.3014723, 0.3676476, 
    0.347252, 0.39959, 0.3333325, 0.193519, 0.2108373, 0.3899055, 0.151797, 
    0.08854784, 0.07357229, 0.3505169, 0.4760602,
  0.0121508, 0.01135126, 0.01055173, 0.009752188, 0.00895265, 0.008153113, 
    0.007353575, 0.007221668, 0.01027636, 0.01333106, 0.01638575, 0.01944044, 
    0.02249514, 0.02554983, 0.03916645, 0.04054419, 0.04192192, 0.04329965, 
    0.04467738, 0.04605512, 0.04743285, 0.03660311, 0.03297022, 0.02933733, 
    0.02570444, 0.02207155, 0.01843866, 0.01480578, 0.01279043,
  0.05753171, 0.04256249, 0.08711712, 0.04460485, 0.0318203, 0.01623998, 
    0.03066499, 0.0050097, 0.02365676, 0.0122306, 0.001347897, 0.005670969, 
    0.0644554, 0.01324668, 0.35833, 0.1693116, 0.1999322, 0.4611131, 
    0.1827686, 0.358369, 0.5126143, 0.6605345, 0.2388224, 0.111539, 
    0.2196888, 0.274131, 0.2748671, 0.1662011, 0.1895752,
  0.1065862, 0.08394889, 0.1060054, -0.0006579371, 0.003056939, 0.09453619, 
    0.001330432, 0.1355821, 0.3735937, 0.1691372, 0.200575, 0.4073117, 
    0.04982046, 0.05314043, 0.3162974, 0.4357972, 0.3947513, 0.3063129, 
    0.2595129, 0.348904, 0.3397274, 0.3346944, 0.248367, 0.186784, 0.3348817, 
    0.3659982, 0.313218, 0.2695975, 0.1524781,
  0.3407564, 0.2375247, 0.06210971, 0.04591633, 0.0780756, 0.1483535, 
    0.2892658, 0.3367693, 0.1646442, 0.0357881, 0.09068955, 0.1310187, 
    0.1962412, 0.1822275, 0.1485084, 0.1626739, 0.2661432, 0.316657, 
    0.1068312, 0.04368322, 0.04940806, 0.02666309, 0.06028316, 0.07081447, 
    0.1352523, 0.2436414, 0.3110915, 0.2714099, 0.3320436,
  0.04136923, 0.05954987, 0.0955269, 0.1252328, 0.1711913, 0.1472865, 
    0.1336569, 0.09056427, 0.07404116, 0.04840386, 0.03186419, 0.03323919, 
    0.02686421, 0.03122616, 0.04519005, 0.04224567, 0.04174294, 0.06365409, 
    0.02552336, 0.04042848, 0.05968792, 0.05192834, 0.04086956, 0.1842612, 
    0.03505281, 0.05985705, 0.08353434, 0.05331469, 0.04276314,
  0.03035555, 0.005174429, 0.004470988, 0.01854751, 0.01523594, 0.02343113, 
    0.009982299, 0.0092499, 0.02340205, 0.002394234, 0.003508255, 
    0.001463237, 0.0001719245, 0.007298341, 0.08831924, 0.02325669, 
    0.01946738, 0.04759247, 0.03546187, 0.01953771, 0.06737957, 0.03468246, 
    0.0162501, 0.1873233, 0.003008323, 0.007241363, 0.02424681, 0.03703766, 
    0.01989603,
  0.002617602, 0.006199855, -0.0003986501, 0.001020013, 0.002611144, 
    0.003822061, 0.003572563, 0.001993618, 0.003285915, 0.0005934744, 
    -8.416939e-08, -8.798045e-08, 0.005736274, 0.002006612, 0.005763745, 
    0.01883687, 0.01352485, 0.01660252, 0.01187576, 0.008847479, 0.003432256, 
    0.00393799, 0.009815505, 0.005442313, 0.02408074, 0.003899717, 
    0.001994443, 0.002591811, 0.002566065,
  0.009925966, 0.0005319737, -6.935134e-06, 0.0007809498, -0.0007827659, 
    7.137809e-05, 0.0001356962, 0.0007070348, 0.001510023, 5.566505e-05, 
    6.95203e-09, 1.308753e-09, 0.0005626768, 0.004688894, 0.001098282, 
    0.001055664, 0.001250785, 0.0004317756, 0.001578402, 0.0003466828, 
    0.0004053603, 0.003505157, 0.01107035, 0.009248038, 0.0004562457, 
    0.04345576, 0.0001515463, 0.0008227688, 0.001849785,
  0.02490139, 0.01324381, 7.953219e-08, 0.005943213, 8.917008e-05, 
    8.135125e-05, 0.0001870717, 0.0008000722, 6.025259e-05, -0.000712569, 
    0.0009249651, 5.398467e-05, 0.00388101, 0.0004199879, 8.146009e-05, 
    4.145824e-05, 0.0001097371, 5.428364e-05, -1.601406e-08, 9.710295e-05, 
    0.0005993701, 0.005951218, 0.01517062, 0.01526983, 4.923777e-08, 
    3.336459e-08, -0.0006343724, 0.0002379754, 0.003803961,
  0.009004345, 0.07126547, 0.003599384, 0.0004288547, 0.0003336509, 
    0.000841709, 0.0003023483, 0.0005620388, 0.04863036, 0.1052996, 
    0.0001668282, 0.0003820046, 0.003819125, 0.0005321714, 2.758942e-05, 
    4.751686e-06, 4.670841e-06, 1.803567e-06, 2.96844e-06, 3.588649e-05, 
    0.0008133493, 0.03435031, 0.06262764, 0.01364335, 0.0002263926, 
    0.0001071597, 1.323348e-05, 0.0009821001, 0.005404198,
  0.04155188, 0.02543712, 0.00119855, 0.2033871, -3.987506e-06, 1.499036e-05, 
    0.02748721, 4.657487e-06, -0.002079314, 3.292642e-06, 7.708047e-06, 
    0.0006526224, 0.001438791, 0.000325185, 8.123106e-06, 0.001944716, 
    0.001337441, 0.001881377, 0.004309152, 0.002203289, 0.001087566, 
    0.002456807, 0.2021639, 0.03698348, 8.626722e-05, 0.0002430265, 
    0.0003638494, 0.001888655, 0.0511839,
  2.16487e-08, 1.89985e-08, 9.690491e-09, 0.0003211894, 1.440779e-07, 
    0.0007294414, 0.002624191, -0.0002001177, 0.1596311, -0.0007050584, 
    0.000452469, 0.000456103, 1.768462e-06, 6.337023e-05, 2.360228e-06, 
    2.75741e-05, 0.0003468123, 0.001376233, 0.005990925, 0.03946381, 
    0.004215475, 0.03751212, 1.042492e-05, -0.001725008, 2.949069e-05, 
    0.0001745509, 0.002857928, 0.02010324, -6.435111e-08,
  9.712766e-07, 7.051775e-05, 4.812688e-05, -5.347321e-07, 3.093169e-07, 
    5.457322e-10, -0.004065198, 0.2081192, 0.2022517, 0.002198143, 
    0.0008866985, 0.002588416, 0.0005332857, 0.000135775, 0.001556308, 
    0.0006425385, 0.0007786223, 0.0009394811, 0.0105413, 0.02819451, 
    6.390174e-07, 0.008544812, 0.03701534, 0.0004226438, 1.370624e-05, 
    0.0003067122, 0.00144349, 0.003624532, -1.48028e-05,
  0.0003012783, -0.0001526675, -0.0001301185, 0.2848418, -5.505703e-05, 
    1.738059e-08, 7.562837e-06, 2.525039e-07, 0.002232063, 0.01369767, 
    0.1627296, 0.08316582, 0.1234791, 0.05101468, 0.1174067, 0.07941674, 
    0.04516828, 0.00773121, 0.04783796, -0.002160446, 2.708524e-06, 
    0.01430836, 0.02434723, 0.1014361, 0.008636427, 0.01355777, 0.002620034, 
    0.01246172, 0.08525462,
  0.03057639, 0.05074201, 0.01543186, 0.004377462, 0.0002942115, 
    2.200156e-06, 0.00133737, 0.04800153, 0.06352034, 0.08905759, 0.08834352, 
    0.05561493, 0.3099946, 0.3132563, 0.2448718, 0.3260332, 0.3284041, 
    0.1454034, 0.02645906, 0.05576526, 0.0104255, 0.003167034, 0.1112494, 
    0.1232737, 0.09823585, 0.1511585, 0.05526786, 0.02359406, 0.08644194,
  0.2374677, 0.09575307, 0.01875149, 0.03995004, 0.08368818, 0.04358585, 
    0.09166358, 0.07663622, 0.1275166, 0.1248866, 0.08664388, 0.1762416, 
    0.2326242, 0.2056535, 0.2455086, 0.1778378, 0.2275159, 0.1350854, 
    0.1209722, 0.09130193, 0.02594614, 0.07711551, 0.1023101, 0.1145331, 
    0.2514798, 0.1400785, 0.1011264, 0.09935163, 0.3017041,
  0.2615137, 0.1211483, 0.2674552, 0.08668736, 0.1792904, 0.2728664, 
    0.2360992, 0.200028, 0.1356132, 0.1358514, 0.1364985, 0.2855454, 
    0.2697304, 0.3671907, 0.187495, 0.2030177, 0.1717574, 0.1906899, 
    0.1727353, 0.1564863, 0.3290415, 0.3656254, 0.1851247, 0.1754916, 
    0.1945592, 0.2032356, 0.2864765, 0.2550341, 0.4247549,
  0.5013993, 0.2662974, 0.2684119, 0.2531662, 0.2090493, 0.33086, 0.3944924, 
    0.4091697, 0.4185853, 0.4066308, 0.3724548, 0.3138628, 0.2951699, 
    0.2852121, 0.2616006, 0.2489989, 0.2526987, 0.3066558, 0.3002006, 
    0.3554213, 0.2976957, 0.1680116, 0.1945624, 0.3562287, 0.1375932, 
    0.08623026, 0.0680086, 0.3321925, 0.4054506,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2.401027e-05, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, -2.885349e-06, 0, -4.791023e-06, 0, 0, -1.934039e-05, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 1.171923e-06, 0, 0, 0, 1.90944e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.460109e-05, 0, -5.882556e-05, 0, 0, 0, 
    0, 0, 0, -7.31438e-06, 0, 0, 2.493059e-05, 0, 0, -9.000839e-06, 0, 0,
  0, 0, 0, 0, 0, 0, -3.98339e-05, 0, -2.958632e-05, 0, 0, 0.0009410249, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, -3.528134e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 4.895271e-05, 0, 0, 0, 0.003302375, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, -8.091683e-06, 0, 0, 0, 0, 0, 0, 0, -6.682684e-06, 0, 0.0003267125, 0, 
    -0.0001037551, 0, 0.00329614, 0, 0.000786463, 0, -3.634716e-05, 
    -2.766303e-05, 0, -5.783729e-05, 2.07785e-05, -7.483203e-07, 0, 
    -6.884534e-05, -1.76848e-06, 0,
  0, 0, 0, 0, 0, 0, 0.002205595, 0, -6.356021e-05, 0, 0.0002091525, 
    0.002607881, -2.913835e-05, 0, 0, 0, 0, 0, 0, 0, 0, -8.684077e-05, 0, 0, 
    0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, -2.417854e-05, 0, 0, 0, -2.628852e-07, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, -7.056269e-05, 0, 0, 0, 0, -1.430668e-06, 0, 
    -5.198449e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 4.024574e-05, -6.447473e-06, 0, 0, 0.005779605, 0, 0.001941693, 0, 
    0.000177481, 0, 0, 3.064986e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0,
  0, 0.0001104622, 3.176574e-05, 0, 0, 0, 0, 0, 0, -4.508129e-05, 0, 
    0.002298785, 0.0002066295, -0.0001497798, 0.0006907218, 0.003648158, 
    0.0007739082, 0.0009950601, -3.793522e-05, 0.001243902, 0.002264494, 
    -0.0001268521, 0.000395122, 0.0001979397, -4.435297e-05, 0, 0.003149966, 
    0.001763256, 0,
  0, 0, 0, 0, 0, 0, 0.006621389, -1.356363e-05, -7.550472e-05, 0, 0.00286858, 
    0.006023736, 0.0003682322, 0, 0, 0, 0, 0, 0, 0, 0.0002656846, 
    -0.0002944221, 0, 0, 0.0002353721, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, -7.253564e-05, 0, 0, 0, -3.324549e-06, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.000745061, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -1.202813e-05, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0.0005246676, 0, 0, 0, 0, -2.426507e-05, 0.0002923363, 
    -0.0001065971, 0.0008979059, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0.0001743505, 0.0002899383, 0, 0, 0.01588845, 0, 0.004156548, 0, 
    0.00247393, 0, 0, -1.622574e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0,
  0, 0.0006499379, 4.764861e-05, 0, 0, 0, 0, 0, 0.002805939, 0.0008179769, 0, 
    0.008471906, 0.00170562, 0.00228957, 0.002982117, 0.008840803, 
    0.0007554617, 0.002719431, 0.000463238, 0.00400652, 0.006571392, 
    0.001274173, 0.003574144, 0.0003228875, -6.184263e-05, 0, 0.00694075, 
    0.005791075, 0,
  0, 0, 0, 0, 0, 0, 0.01716203, 0.0007721885, 0.002879558, 0.001636181, 
    0.005173641, 0.01082025, 0.002413117, 0, 0, 0, 0, 0, 0, -2.061867e-06, 
    0.0003464514, -0.000352957, -8.799553e-06, 0, 0.001237081, -2.693258e-05, 
    0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0.0002022481, 0, 0, 0, 5.555921e-05, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.003640917, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.002825432, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -3.011528e-06, 0, -8.719199e-06, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0002741901, -3.631674e-06, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0004051809, -7.005636e-06, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.180436e-05, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0.005826164, 0, 0, 0, -1.16398e-10, 0.0002071851, 
    0.0008529, -0.0001286289, 0.002572715, -0.0001181483, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0.0005745922, 0.005021226, 0, 0, 0.02942212, 0, 0.01297063, 0, 
    0.009403836, 0, -3.364201e-05, 5.038665e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.001188516, 0, 0, 0, 0, 0,
  -4.317789e-05, 0.0009528289, 0.0001396947, -4.125041e-06, 0, 0, 0, 0, 
    0.004279865, 0.003846675, 0, 0.01305194, 0.00751104, 0.004247705, 
    0.004199245, 0.01558102, 0.001429829, 0.007323119, 0.0007174498, 
    0.006575704, 0.01965022, 0.004055633, 0.01110678, 0.0006000181, 
    -3.571274e-05, 0, 0.011812, 0.00862183, 0.001829072,
  0, 0, 0, 0, 0, 0, 0.02740484, 0.001296942, 0.004044069, 0.004672985, 
    0.01099289, 0.02069816, 0.009584604, 0, 0, 0, 0, 0, 0, -1.421314e-05, 
    0.0003431737, 0.001324073, -0.0001635584, -2.025931e-05, 0.003681996, 
    9.845137e-05, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0.001250894, 0.0006807871, 0, 0, 0.0005040577, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.0002858793, 0, -7.861868e-05, 0.00599708, 
    -3.284523e-05, -7.537638e-06, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, -2.411571e-05, 0, 0, 0.007292192, -3.591214e-05, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, -5.408843e-05, -2.772307e-05, 0.0002394463, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -3.219632e-07, 0, 0, 0, 0, 0, 0, 0, 
    0, -2.924148e-05, 8.011026e-05, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -1.924857e-06, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, -2.019838e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.003093018, -2.826855e-05, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001577418, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.002022492, -0.0001513781, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -7.280593e-06, 0.003049273, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, -1.993507e-05, 0, 0.01289712, -4.707992e-05, 0, 0, 
    -6.543515e-07, 0.0008457542, 0.003707746, 0.0005946158, 0.008458326, 
    0.001169013, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0.01059624, 0.008087801, 0, 0, 0.04132331, -2.132882e-05, 0.02484639, 
    -1.126918e-05, 0.02048701, 0, 0.0001200826, 0.000949186, 2.182268e-05, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0.001635347, 0, 0, 0, 0, 0,
  -9.695714e-05, 0.004545026, 0.0008176908, 0.0003896091, 0, 0, 0, 
    -1.404509e-05, 0.00906711, 0.009577594, -2.177337e-05, 0.01850877, 
    0.0181259, 0.006558475, 0.01265545, 0.02738602, 0.003395899, 0.01489431, 
    0.002322681, 0.01060305, 0.04792868, 0.01399404, 0.01770604, 0.001846145, 
    9.072803e-05, 0, 0.01395459, 0.01908179, 0.005776669,
  0, 0, 0, 0, 0, -3.576635e-05, 0.03610258, 0.007028489, 0.006636528, 
    0.01610564, 0.02002669, 0.0352751, 0.01791885, -3.255306e-05, 0, 0, 0, 0, 
    0, -1.412524e-06, 0.0005643644, 0.006953236, -8.299501e-05, 
    -0.0001073609, 0.007427106, 0.0006338549, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0.002516205, 0.001011219, 0.00205403, 0, 0.00174323, 
    0, 0, 0, 0, 0, 0, 0, 0, 0.001285079, -1.753795e-05, -0.0001248528, 
    0.008689677, 6.816417e-05, 0.0002589766, 0, 0, 0,
  0, -4.730377e-06, 0, 0, 0, 0, 0, 0, -3.47651e-05, -4.903093e-06, 
    0.001645984, 0.01826037, 0.003183918, -5.585709e-06, -3.727152e-05, 0, 0, 
    0, 0, 0, 0, -1.595914e-07, 0.0003632332, -2.788726e-05, 0.001232861, 
    -1.16588e-06, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0006497428, 9.85459e-05, -2.486679e-05, 
    -1.174487e-05, 0, 0, -3.366158e-06, 0, 0, 0, 0, 0.0005942085, 
    0.004062762, 0.001384351, 0.001718518, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.001839791, -1.022239e-05, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0.001231963, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.0003162549, 0, 0, 0,
  0, 0, 0, 0.003548099, -4.080192e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -8.930522e-07, 0, -1.183146e-05, 0, -3.696603e-05, -3.128804e-05, 
    -1.438853e-05, 0, 0, 0, 0.003743166, 0.002892546, 0.002220919, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0002677467, -1.702051e-05, 
    0.005182554, 0, 0, 0.0008410819, 0, 0, 0, 0, 0, -1.261806e-05, 
    0.007928712, 0.001881353, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.623415e-06, 0.009881531, 
    0.008015256, -2.317509e-05, 0, 0, 0, 0, -8.247241e-06, 0, 0, 0, 0, 0, 0,
  0, 0, -2.141371e-06, 0, -3.87568e-05, 0, 0.02024536, 0.0006212561, 0, 0, 
    -7.925437e-05, 0.003531598, 0.008288936, 0.003086605, 0.01824059, 
    0.002432032, -0.0001932416, 0, 0, 0, 0, 0, 0, -1.973217e-05, 0, 0, 0, 0, 0,
  0, 0.0273324, 0.01040807, 0, 0, 0.05565038, -6.525903e-05, 0.04371369, 
    0.001856919, 0.03144366, 9.767956e-05, 0.003926091, 0.01019987, 
    0.0005490175, -4.571758e-06, 0, 0, 0, 0, 0, 0, 0, -1.010451e-05, 
    0.001651413, 0, 0, 0, 0, -2.444366e-05,
  -0.0003105918, 0.01075401, 0.001639323, 0.001743669, 0, 0, 0, -0.000120025, 
    0.01541055, 0.02331573, 0.0002597379, 0.0315127, 0.0312873, 0.01251896, 
    0.02832849, 0.04029263, 0.008215222, 0.02349936, 0.004586778, 0.02222881, 
    0.1012551, 0.03395707, 0.02629954, 0.002486237, 0.001823563, 0, 
    0.02004984, 0.03870206, 0.009706918,
  0, 0, 0, 0, -7.875715e-07, -0.0001290697, 0.0432997, 0.01601782, 
    0.01435583, 0.0257651, 0.03045842, 0.06363311, 0.02933216, 0.0001996029, 
    -9.116492e-06, 0, 0, 0, 0, -2.53458e-05, 0.006074538, 0.01581245, 
    0.0002919943, 0.0008762983, 0.01347012, 0.001975615, 0, 0, 0,
  0, 0, 0, 0, 0, 0, -1.430088e-11, 0.003542914, 0.003654773, 0.004547295, 0, 
    0.008592823, -5.685184e-06, 1.467849e-05, 0, 0, 0, 0, 0, 0, 0.001407243, 
    0.001428858, 4.053533e-05, 0.01484231, 0.0001565323, 0.0003908274, 0, 0, 0,
  0, 0.000554714, 0, 0, 0, 0, -4.438134e-06, 0, -3.473069e-05, 0.0008295217, 
    0.007025765, 0.03946252, 0.01152638, -2.543774e-05, -9.330383e-05, 
    0.0007585931, -6.857404e-06, 0, 0, 0, 0, 0.002984343, 0.003670877, 
    0.003857651, 0.005898936, 4.518249e-05, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -5.844872e-06, 0.003906639, 0.007690257, 
    -5.743422e-05, 0.006250051, 0, 8.089578e-05, 0.001036052, 0, 0, 0, 
    -6.107984e-07, 0.004726768, 0.005550263, 0.007671309, 0.006263968, 
    0.0007260338, -2.708817e-05, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.003213903, 0, 0, 0, 0, 0, 0, 
    0.004035868, -3.10107e-05, 0.002654981, -2.966249e-05, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, -1.795162e-05, 0, -4.776942e-06, 0.004333835, -1.618304e-05, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0002871542, 0, 0, 0, 0, 0, 0.001317123, 0, 
    0, 0,
  0, 0, 0, 0.007785543, 0.0008202835, 0, -1.991036e-06, 0, 0, 0, 0, 0, 0, 0, 
    0.003234434, 0, 0.002689696, 1.282078e-05, 0.00336118, 0.001430502, 
    -1.438853e-05, 0, 0, 0, 0.004775973, 0.009362582, 0.009979904, 
    -6.872343e-06, -4.036326e-05,
  0, 0, 0, -4.075883e-07, 0, 0, 0, 0, 0, 0, 0, 2.904303e-07, 0, 0.004568715, 
    -0.0001409721, 0.01146737, 0.001895441, 0.0002249151, 0.006823393, 
    0.0009143597, 0, 0, 0, 0, 0.0004021841, 0.01610726, 0.006727695, 
    2.006663e-05, 0,
  0, 0, -1.589759e-07, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0006945117, 
    -3.055199e-09, 0.01475689, 0.0303733, 0.0107807, 0.0007539515, 
    -0.0001495102, 0, -1.358706e-08, 0, -1.207367e-06, 0, 9.685131e-06, 
    0.000272576, 0, 0, 0,
  0, -8.32376e-06, -7.930318e-06, 0, -5.296262e-05, 0, 0.03634447, 
    0.004636737, 5.31793e-05, 0, 0.001510937, 0.01797972, 0.01875126, 
    0.01196172, 0.0366576, 0.007201798, -0.0002155428, 0, 0, 0, 0, 0, 
    -6.60247e-10, 0.0001401686, 0.000916532, 0, 0, 0, 0,
  2.092178e-06, 0.05216857, 0.0176887, 2.722883e-08, -1.888678e-06, 
    0.08088491, 0.0008659756, 0.07272999, 0.01097959, 0.05426104, 
    0.0005367566, 0.01196955, 0.02885321, 0.008837009, 8.429843e-06, 0, 0, 0, 
    0, -8.766196e-06, 1.937777e-06, 2.376096e-06, -0.0001407508, 0.01320954, 
    0, 0, 0, -8.831025e-11, -3.505771e-05,
  0.004096767, 0.02293777, 0.009922883, 0.002680472, 0, -5.476682e-06, 
    0.0009028681, 0.004101539, 0.0329686, 0.0502232, 0.003660451, 0.0505907, 
    0.06092082, 0.04096077, 0.04255554, 0.06143811, 0.01435886, 0.0319919, 
    0.006983162, 0.03494576, 0.1662833, 0.08050378, 0.05178137, 0.01888417, 
    0.00451941, 8.450127e-05, 0.03383452, 0.05599162, 0.01786342,
  0, 0, 0.0003753834, 0, -8.186501e-05, 0.001531759, 0.05257159, 0.05160455, 
    0.03553943, 0.04473482, 0.04354303, 0.09444265, 0.05111518, 0.004348783, 
    0.0001051538, -8.176678e-05, 0.0008122839, 0, 0, 0.0004237178, 
    0.02061464, 0.05203418, 0.003984558, 0.004894396, 0.01430768, 
    0.007696267, 0, 0, 0,
  0, 0, 0, 0, 0, 0, -1.615595e-05, 0.005724604, 0.008697526, 0.008851214, 
    -0.0001163668, 0.02487153, 7.322789e-05, 0.004950765, 0.002508576, 0, 
    7.764653e-05, 0, 0, 0, 0.007276843, 0.007667687, 0.003232101, 0.02172668, 
    0.01087171, 0.001811118, 0, 0, 0,
  0, 0.002955797, 0, -3.402787e-11, 1.203276e-12, 0, -7.055456e-05, 
    -2.969611e-08, 2.355822e-06, 0.006852121, 0.01800783, 0.06848649, 
    0.02075541, 0.009035046, 0.003290333, 0.007614471, 0.0008692407, 0, 0, 0, 
    0.0001580211, 0.004240933, 0.01323995, 0.009234586, 0.01777294, 
    0.007484361, 0, -4.838567e-05, 0,
  -1.210579e-05, 2.850951e-05, 0, 0, 0, -1.617759e-07, 0, 0, 0, 0.0009127535, 
    0.006433053, 0.008855158, 0.01800061, 0.006650765, 0.0110734, 
    0.0004654254, 0.003052743, 0.003565261, 0, 0, 0, -1.22872e-06, 0.0130164, 
    0.007563146, 0.02737029, 0.011934, 0.01393668, 0.002438306, -0.0001288479,
  0, 0, -1.824927e-05, -7.057766e-07, 0, 0.001259303, 0, 0, 0, 0, 
    -7.860235e-05, 0, 0, 0, -1.677596e-05, 0.006688788, 0, 0, 0, 0, 0, 0, 
    0.004121576, 0.002018462, 0.006432899, 0.0008186764, 0, -2.58125e-05, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  -5.144607e-05, 0, -3.403096e-05, 0, 0.001310021, 0.007141874, 0.001243485, 
    0.0005337454, 0, 0, 0, 0, 0, 0, 0, 0, 0, -4.470169e-06, -1.5639e-05, 
    0.003422877, 0.0002878328, 0, 0, 0, 0, 0.003842139, 0, 0.0001325598, 
    -1.232456e-06,
  -9.034812e-06, 0, 0, 0.01260622, 0.001874587, 0.008862468, 0.003391458, 
    -6.622807e-06, 0, 0, 0, 0, -9.925232e-05, -8.704174e-05, 0.005202365, 0, 
    0.006886694, 0.007086349, 0.01029335, 0.01293246, 0.0007078527, 
    -0.0001192278, 0.0001609344, 0.0004549661, 0.005533927, 0.01642862, 
    0.03194568, 0.0004823171, 0.003814843,
  -3.910696e-08, 0, 1.702122e-07, 2.06656e-05, 0, 0, 0, 0, 1.697556e-09, 
    -6.836057e-11, 4.008837e-12, -2.343837e-07, 0, 0.007425264, 0.002971118, 
    0.01858688, 0.009765988, 0.006378265, 0.03548193, 0.00227386, 
    0.0001115058, 1.466678e-07, 4.557826e-08, -9.238133e-08, 0.001760739, 
    0.02876441, 0.01373047, 0.001949104, -3.937268e-11,
  0, 0, -2.891937e-05, 0, 0, -5.155424e-10, -4.257189e-07, 1.192418e-06, 
    1.960487e-06, 1.307228e-06, 6.648388e-07, 2.789557e-07, 0.01207502, 
    3.076246e-05, 0.02603712, 0.06795529, 0.02059851, 0.01100557, 
    -0.0001403284, -8.46323e-06, 1.114648e-05, 4.639544e-07, 5.943124e-06, 
    0.0003039726, 0.0001568282, 0.0008474819, -2.882983e-07, 0, 0,
  -2.177232e-08, -1.498588e-05, -1.534507e-06, -6.926207e-10, 1.970371e-05, 
    1.715027e-06, 0.04419969, 0.04671891, 0.007230692, 7.832e-06, 0.02065603, 
    0.1128452, 0.09807978, 0.1130432, 0.08014221, 0.05557565, 0.001418389, 
    -2.884891e-07, 2.839801e-07, 2.687284e-06, 0.0001892844, -2.277595e-05, 
    0.0001381799, 0.004560643, 0.001638714, 0, -2.679293e-05, -1.489458e-08, 0,
  0.008869958, 0.109458, 0.05261047, 1.367972e-05, -1.701065e-05, 0.1075438, 
    0.01557438, 0.2159709, 0.09300619, 0.08761065, 0.03162543, 0.05784552, 
    0.1081422, 0.08736869, 0.005765383, 0.0004251674, 0.0003901203, 
    1.636583e-07, -1.029876e-06, 2.388869e-05, 0.01493028, 0.003583814, 
    0.01233868, 0.08971781, 0.0004520635, 0, -1.784809e-07, 0.005763104, 
    0.0001322083,
  0.03844068, 0.06685121, 0.04560157, 0.002944143, -2.004523e-06, 
    0.004188992, 0.02407544, 0.5145487, 0.4332523, 0.4157121, 0.2743606, 
    0.278168, 0.2776654, 0.2379876, 0.1692459, 0.1459754, 0.04415715, 
    0.0328822, 0.01575417, 0.1019194, 0.3631768, 0.3058417, 0.09457181, 
    0.09880007, 0.01038573, 0.006253699, 0.06014709, 0.08138933, 0.04090833,
  0.0001586392, -0.0001170466, 0.001648428, 0.0004440316, 0.007773133, 
    0.09066294, 0.3069198, 0.166392, 0.2195371, 0.1146235, 0.1436055, 
    0.263971, 0.1924345, 0.07173517, 0.007663263, -0.0002701442, 0.004220613, 
    -5.484889e-09, 4.658742e-06, 0.03054504, 0.1410614, 0.1637516, 
    0.08537691, 0.09847355, 0.0200175, 0.0106638, 0.009287824, 5.706633e-05, 
    0.002854707,
  -2.664782e-08, -3.06655e-09, 0, 1.483516e-09, 6.956132e-08, -1.632658e-06, 
    0.0001628772, 0.01359382, 0.01662112, 0.1017607, 0.08278968, 0.1017264, 
    0.05013461, 0.04948949, 0.01327616, -5.466301e-06, 0.00112292, 
    2.261294e-06, 8.741631e-10, -1.011277e-07, 0.03294909, 0.03856518, 
    0.03091458, 0.04488255, 0.02586925, 0.007819562, 2.999047e-06, 
    -9.107041e-07, 0,
  0, 0.009180635, 0, -1.281392e-09, -6.5624e-07, 0, -6.072579e-05, 
    0.001362864, 0.004075754, 0.01367426, 0.03583599, 0.1354049, 0.07490934, 
    0.03879922, 0.01400952, 0.02036911, 0.007284933, 2.180109e-06, 
    3.211857e-09, 0, 0.0012521, 0.005664492, 0.02626542, 0.02081402, 
    0.02901369, 0.0113104, 0.0002490241, -5.600277e-05, 0.0006025081,
  7.441651e-05, 0.001098133, 0, 5.351494e-06, -5.052778e-06, 1.705373e-06, 0, 
    0, -0.0001421905, 0.007565149, 0.0115982, 0.02365429, 0.05397724, 
    0.02805149, 0.01724829, 0.007223434, 0.02481448, 0.007152211, 
    0.0001935832, 0, -6.051559e-06, -3.398541e-06, 0.02489635, 0.008526746, 
    0.05076202, 0.02803661, 0.05646199, 0.009311071, 0.005591947,
  0.0008489902, -0.0001363174, 0.00742354, 0.0006561212, -0.000140217, 
    0.002495304, 0, 0, 0, 0, -0.0002105836, -1.434892e-05, 0, -6.251971e-06, 
    -0.000128086, 0.008615058, 0.004154322, 0.0002177044, 3.196634e-05, 
    0.0004922407, 0, -0.0001167661, 0.004696934, 0.004072099, 0.01518659, 
    0.007663576, 0.0008164294, 0.001338142, 0.003372651,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -3.12501e-05, 1.229202e-05, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.187913e-08, 
    0, 0, 0, 0, 0, 0, 0, 0,
  -0.0001325969, 0, 1.288059e-05, -6.83179e-05, 0.006314113, 0.01120497, 
    0.003940168, 0.001276517, 0, 0, 0, 0, 0, 0, 0, -5.302944e-06, 0, 
    -6.969212e-06, -0.0002350259, 0.00768957, 0.002498706, 0.0005029249, 0, 
    0, 0, 0.01030115, 0, 0.002207836, 8.17445e-05,
  0.0006475869, -6.370721e-08, 2.774897e-08, 0.0182349, 0.007750311, 
    0.02030145, 0.004449199, -4.369444e-05, 0, -6.348574e-11, 1.390223e-07, 
    -4.4534e-06, -0.0001950272, 0.002641438, 0.009454589, 0.0003321272, 
    0.01026345, 0.02095142, 0.02457897, 0.02925586, 0.01255388, 
    -0.0001592031, 0.001209999, 0.001249667, 0.008377478, 0.02682371, 
    0.05276891, 0.009729662, 0.01803967,
  0.0002772739, 2.133428e-06, 3.225898e-05, 0.0009694434, 3.173979e-07, 
    0.0008040505, 0, 0, 1.873999e-07, 2.302082e-06, 6.870837e-07, 
    0.0001994411, -2.025606e-08, 0.01020399, 0.01758482, 0.02646878, 
    0.03288413, 0.03071695, 0.07308685, 0.007767564, 0.001555161, 
    0.001300117, 0.001958351, 0.0005647144, 0.0162973, 0.06397191, 
    0.03928927, 0.03765384, 0.001912495,
  1.370449e-06, 2.180306e-05, -6.252283e-05, -7.419713e-11, 0, -8.782334e-11, 
    -7.541108e-07, 0.0002743935, 2.183507e-06, 1.527182e-06, 6.978579e-07, 
    1.032096e-06, 0.03245509, 0.00267597, 0.04959945, 0.1311635, 0.09554788, 
    0.05254273, 0.007264138, 0.002598544, 9.55543e-06, 1.360275e-05, 
    2.604754e-05, 0.02413991, 0.038744, 0.006914194, 0.001853655, 
    8.518954e-05, 0.006661699,
  8.6344e-06, -8.482177e-05, 0.009438254, -1.498741e-07, 0.0002579533, 
    0.01807005, 0.06628554, 0.08138935, 0.005037817, -1.034742e-05, 
    0.03125528, 0.09677937, 0.08529846, 0.1060898, 0.08254967, 0.07683841, 
    0.02171867, -5.394287e-06, 1.874802e-06, 9.876395e-06, 0.01406896, 
    0.0004193836, 0.0008624402, 0.06300855, 0.1149842, 1.095136e-06, 
    0.0002185773, 2.273719e-05, 3.34639e-06,
  0.1091818, 0.472166, 0.4190605, 0.001088966, 0.0005579419, 0.14513, 
    0.09677143, 0.3376985, 0.3889242, 0.2222885, 0.04936324, 0.05373637, 
    0.08256884, 0.06824031, 0.003387124, 0.000143675, 0.0004490862, 
    2.30943e-07, 3.817922e-05, 0.008372841, 0.116907, 0.1334979, 0.1021679, 
    0.2544911, 0.04866105, 7.658984e-05, 0.0002418496, 0.01421122, 0.01442502,
  0.195779, 0.2012843, 0.2128918, 0.005810488, 0.00231066, 0.001882669, 
    0.05443487, 0.4313566, 0.363771, 0.2750777, 0.1516251, 0.2275442, 
    0.2341273, 0.2164084, 0.1462378, 0.1589688, 0.08910045, 0.03523981, 
    0.01395734, 0.1015765, 0.4025173, 0.2993756, 0.2244197, 0.2151609, 
    0.07409122, 0.03676455, 0.06603928, 0.1762267, 0.2259765,
  0.02571313, 0.001466722, 0.02105871, 0.0001284683, 0.0008988863, 
    0.05811001, 0.2955947, 0.1080443, 0.1845802, 0.1037915, 0.1250874, 
    0.2016102, 0.1634454, 0.1260611, 0.1643809, 0.07262982, 0.02419649, 
    0.0003363722, 1.178638e-05, 0.02178317, 0.09769652, 0.1642781, 0.1175136, 
    0.1491293, 0.113839, 0.0959965, 0.02292762, 0.03344668, 0.09540364,
  -0.000278643, 0.007335052, -1.280992e-05, 1.702528e-07, -2.018554e-08, 
    -3.441332e-07, 0.0008961465, 0.02491216, 0.03358477, 0.09771904, 
    0.06250069, 0.08337539, 0.07186376, 0.06168536, 0.1026312, 0.06155504, 
    0.07676835, 0.01812267, -4.54597e-05, -2.874414e-08, 0.1490287, 
    0.09013045, 0.1150171, 0.1508469, 0.105406, 0.06557196, 0.004732423, 
    0.04533057, -8.94811e-05,
  -7.32171e-05, 0.01893015, 0.0004415498, -5.965979e-07, -2.329603e-06, 
    3.164448e-08, 0.0008047171, 0.02038849, 0.03336634, 0.05133025, 
    0.1444806, 0.2890726, 0.2118115, 0.158334, 0.1373554, 0.1298776, 
    0.03691267, 0.04818593, 0.002745195, 0.0004091563, 0.002949607, 
    0.07631186, 0.1179093, 0.0841558, 0.1380204, 0.08866523, 0.04012673, 
    0.01135456, 0.006352791,
  0.003631037, 0.01218928, 0.0001374039, 0.005006263, 6.772145e-05, 
    0.007409104, 0, 0.001045049, -0.0002428122, 0.01162701, 0.01820865, 
    0.04310532, 0.1058781, 0.09469559, 0.05310086, 0.03586793, 0.0841722, 
    0.0230548, 0.006348117, -1.129444e-05, 0.0009048363, 0.001366872, 
    0.03382373, 0.02210381, 0.09593081, 0.08367006, 0.1190697, 0.0244062, 
    0.008563079,
  0.005955471, -0.0001232398, 0.01659709, 0.004737367, 0.001480343, 
    0.002571292, -0.0001346269, -5.276394e-06, 0.0006244323, 0, 0.001063884, 
    0.001195096, 0, 0.000461701, 4.86872e-05, 0.01917479, 0.007199819, 
    0.009046273, 0.00206119, 0.002872981, -6.08238e-05, 6.391622e-05, 
    0.00488334, 0.008329883, 0.02161482, 0.02327725, 0.007018192, 0.01357275, 
    0.006272207,
  0, 0, 0, 0, 0, 0, -2.065593e-05, 0, 0, 0, 0, 0, 0, 0, -0.0001539925, 
    0.0007769507, 0.002624897, 3.047478e-07, 0, -8.81887e-07, 0, 0, 0, 0, 0, 
    0, 0, 0.0002375295, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2.968351e-06, 
    6.23839e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0012555, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0.0001128219, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2.185013e-05, 
    0, 0, 0, 0.001492544, 0, 0, 0, 0, 0, 0, 0, 0,
  -0.000212524, 0.0007261047, 0.0004271235, 0.003491475, 0.01364786, 
    0.01806204, 0.007320741, 0.002388022, 0.0005521967, -4.293605e-08, 
    -1.610229e-08, 0, 0, 0, 0.001794725, -2.856193e-06, -6.561764e-06, 
    0.0002028327, 0.004817259, 0.02291728, 0.01364525, 0.002515226, 
    -4.923673e-05, 0, 0, 0.01058432, -2.415125e-05, 0.01072487, 0.003490653,
  0.005550643, -0.0002473691, 0.01536631, 0.04636763, 0.01745265, 0.04810005, 
    0.01798196, 0.0002308258, 3.892277e-05, -3.539882e-06, 0.0001915115, 
    0.004401715, 0.0006996469, 0.01056032, 0.02474169, 0.000586227, 
    0.01453071, 0.03787788, 0.04837025, 0.04835417, 0.03443607, 0.006312389, 
    0.007016912, 0.00560658, 0.01249316, 0.05571977, 0.1398248, 0.05286327, 
    0.04144603,
  0.0314547, 0.01563042, 0.001693787, 0.01518095, 0.006262513, 0.0007355028, 
    0, -7.218796e-12, -2.408072e-06, 2.962852e-06, 1.181647e-06, 
    0.0001833867, 7.377825e-05, 0.01267969, 0.02745987, 0.05742505, 
    0.1032669, 0.1438936, 0.2052511, 0.08319508, 0.01576865, 0.005212894, 
    0.009560726, 0.003560172, 0.03897148, 0.1236222, 0.1155006, 0.08712741, 
    0.03236922,
  6.504109e-07, -4.847057e-09, 0.004551251, 3.606462e-09, 0, 8.17973e-07, 
    2.383294e-06, 0.000187409, 6.414128e-07, 1.443346e-06, 3.694294e-07, 
    7.959815e-08, 0.0242716, 0.0003248113, 0.0520361, 0.09456342, 0.07949885, 
    0.04366774, 0.005034926, 0.001501832, 4.183709e-06, 4.516347e-06, 
    5.188113e-06, 0.02146341, 0.04576332, 0.02913424, 7.138371e-05, 
    1.329651e-06, 0.0005733626,
  3.107181e-06, -0.0001005045, 0.007043804, -1.083374e-07, 0.001433314, 
    0.008993691, 0.04978114, 0.03532213, 0.0001772587, 0.0002013065, 
    0.02529155, 0.06541547, 0.08095811, 0.09111534, 0.06720223, 0.0514086, 
    0.01440323, -1.187251e-06, 1.115947e-07, 1.018986e-06, 0.0001237734, 
    2.651102e-05, 1.187694e-05, 0.04014425, 0.08601261, 1.949084e-07, 
    2.281921e-05, 1.017279e-06, 3.914681e-07,
  0.04484333, 0.4237855, 0.3317067, 3.707069e-05, -6.557468e-06, 0.1322542, 
    0.05277207, 0.2920913, 0.2952164, 0.1902576, 0.02906302, 0.04322685, 
    0.05624986, 0.05714918, 0.001780121, 3.685134e-05, 1.105784e-05, 
    1.963917e-07, 1.353686e-05, 0.0001658563, 0.03392575, 0.04437008, 
    0.06977642, 0.1845555, 0.01479543, 1.591843e-05, 8.818254e-05, 
    0.009485572, 0.0001894673,
  0.16146, 0.1770663, 0.1587191, 0.0478235, 0.0003584392, 0.0001997155, 
    0.02820143, 0.2831612, 0.2705197, 0.1652895, 0.08456632, 0.1825651, 
    0.1940501, 0.1773217, 0.1130664, 0.1414105, 0.06132503, 0.03042285, 
    0.01121696, 0.0588362, 0.3339477, 0.2716013, 0.2020226, 0.1615073, 
    0.04431618, 0.02689998, 0.0504982, 0.142856, 0.181641,
  0.0180251, 0.001133297, 0.0109574, 7.430837e-05, 4.658639e-05, 0.03965333, 
    0.278272, 0.09829264, 0.1477356, 0.09742524, 0.1111351, 0.1717256, 
    0.124678, 0.06728816, 0.09433033, 0.05201406, 0.009290464, 4.334966e-05, 
    3.337328e-06, 0.01887358, 0.07093906, 0.1291341, 0.09179159, 0.1320087, 
    0.09877668, 0.07090716, 0.02050185, 0.01206608, 0.07827715,
  0.05298829, 0.05735752, -1.28873e-05, 6.894522e-08, -3.211121e-07, 
    -8.686669e-08, 0.0008348611, 0.03691689, 0.07788781, 0.09561247, 
    0.05491146, 0.07157657, 0.07988232, 0.03676108, 0.07417894, 0.05252945, 
    0.09604724, 0.01713099, -2.10271e-05, -1.453745e-08, 0.13918, 0.0842119, 
    0.08686908, 0.1295632, 0.09762635, 0.05787867, 0.06514171, 0.03964994, 
    0.003536727,
  0.02969535, 0.08444995, 0.01443322, 0.0001655031, 0.005754536, 
    4.309078e-05, 0.003844248, 0.04698141, 0.07384987, 0.06271491, 0.1954382, 
    0.2786908, 0.1841433, 0.1293028, 0.1313256, 0.212273, 0.1374963, 
    0.1395395, 0.03178154, 0.01701049, 0.04907688, 0.1496761, 0.1359463, 
    0.1117332, 0.1365539, 0.1222479, 0.07951911, 0.06003671, 0.06654363,
  0.03173342, 0.03114397, 0.04974955, 0.01084139, 0.0005506889, 0.01321961, 
    -0.000120301, 0.003081718, 0.0001634776, 0.02838358, 0.05142065, 
    0.05987913, 0.1037621, 0.1627682, 0.09334933, 0.1016868, 0.2020319, 
    0.1528583, 0.09329973, 0.002598813, 0.006221223, 0.03987186, 0.06017161, 
    0.06941773, 0.1816126, 0.2111601, 0.2205481, 0.1501554, 0.06088417,
  0.04034531, 0.003515583, 0.0242811, 0.01196237, 0.005728521, 0.006315696, 
    0.001891506, 0.0009258752, 0.00550517, 0, 0.009812183, 0.003725166, 
    -0.00118059, 0.004419698, 0.005893641, 0.02112687, 0.03408017, 
    0.02463562, 0.007994924, 0.007242628, 0.0002868268, 0.006280979, 
    0.006380437, 0.03035249, 0.03504318, 0.04747842, 0.03747872, 0.02210844, 
    0.03572343,
  -7.772876e-05, -9.598072e-07, 0, 0.0002598108, 0.0002646709, -3.482144e-07, 
    0.005344946, 0, 0, 0, 0, 0, 0, 0, 0.001450556, 0.0117761, 0.0231778, 
    0.02573747, 0.01995892, 0.02627414, 0.009325264, -0.0002548732, 
    1.987189e-06, -0.0002671809, -8.291662e-06, 0, 0, 0.004333836, 
    -1.053144e-06,
  0, 0, 0, 0, -2.559616e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2.375575e-08, 
    -4.47368e-05, 0.0009700392, 2.848399e-07, -4.281916e-09, -4.719884e-09, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.006984909, 0, 0, 0, 0,
  0, 0, 0, 0, -2.79164e-06, -5.574048e-06, -0.0001653288, 1.111069e-05, 
    0.0003926097, 0, 0, 0, 0, 0, 0, 0, 0.000140055, 0, 0.0006648292, 
    0.003091948, 0.00337375, 0.002013693, 0, 1.710514e-05, 2.902491e-05, 0, 
    0, 0, 0,
  0.006120497, 0.02254388, 0.003127952, 0.04443217, 0.08655572, 0.06923747, 
    0.03795301, 0.02657444, 0.005128387, 0.0004238832, -2.992275e-05, 
    -0.0004159988, 0.001854902, 0.0001470161, 0.007348649, 0.0001663783, 
    0.000420818, 0.007146083, 0.01626161, 0.04077836, 0.03068827, 0.01158597, 
    0.001683106, -5.958192e-05, 0.004041539, 0.01509295, 0.004658725, 
    0.02830583, 0.0156633,
  0.0821572, 0.06627182, 0.1082187, 0.1353223, 0.1033843, 0.09937891, 
    0.05450792, 0.03117116, 0.004380841, 0.0007759898, 0.008788151, 
    0.01816925, 0.01171844, 0.06572554, 0.05793155, 0.04491566, 0.02606161, 
    0.06096146, 0.08439592, 0.0789875, 0.09119371, 0.03263963, 0.02692216, 
    0.02108501, 0.03677014, 0.08215047, 0.1777552, 0.09839027, 0.1256494,
  0.05304899, 0.01324056, 0.03083273, 0.01203144, 0.001214866, 0.000517749, 
    0.0001148869, -3.840613e-06, -4.446949e-05, 0.0002447642, -5.408503e-06, 
    0.003368908, 0.0002176512, 0.02878058, 0.04945525, 0.08373594, 0.1243616, 
    0.1674685, 0.2214384, 0.1214272, 0.02581058, 0.02517729, 0.01357283, 
    0.005578378, 0.04521052, 0.1040125, 0.07088528, 0.04352599, 0.05596747,
  6.926513e-07, -2.044716e-05, 0.007353407, 7.855738e-07, -7.745788e-11, 
    3.455987e-07, 5.897559e-06, 0.0004757539, 1.739776e-07, 8.390308e-07, 
    3.138504e-07, -6.772619e-07, 0.01156095, 0.005977035, 0.06336536, 
    0.08091575, 0.048471, 0.04651533, 0.001800603, 1.898625e-05, 
    4.810113e-07, 1.335174e-06, 6.021622e-07, 0.01699459, 0.04325987, 
    0.01500749, 7.277801e-06, -2.086732e-07, 1.011202e-06,
  1.653804e-06, -5.469883e-05, 0.00550653, -3.148719e-07, 0.001563827, 
    0.001899227, 0.044336, 0.02039987, -5.220843e-06, 0.0006174754, 
    0.02991663, 0.0447509, 0.07634034, 0.09120772, 0.06604571, 0.0395008, 
    0.01194454, 3.764368e-07, -6.34124e-09, 2.046265e-06, 1.413438e-05, 
    1.664864e-06, 1.15405e-05, 0.03547679, 0.02362158, -4.031841e-07, 
    3.194823e-06, 3.812847e-07, 1.470695e-08,
  0.007519629, 0.3839654, 0.2367418, -9.980934e-07, 0.0003804743, 0.1265106, 
    0.04468421, 0.2431766, 0.2324222, 0.1836341, 0.02262318, 0.04101873, 
    0.05789433, 0.05131845, 0.003251283, 1.006493e-06, 4.937165e-06, 
    7.679126e-08, 3.110118e-06, 2.935715e-06, 0.0007145194, 0.01446011, 
    0.05129245, 0.1696827, 0.004476364, 1.83022e-06, 2.743839e-05, 
    0.0006956785, -3.872884e-05,
  0.1452968, 0.1775984, 0.1402108, 0.03147945, 0.0007863665, 0.0001235962, 
    0.01908278, 0.1432884, 0.2162461, 0.113305, 0.05083248, 0.1685981, 
    0.1688596, 0.1502518, 0.1193275, 0.1511043, 0.0515867, 0.02821117, 
    0.01043611, 0.04709674, 0.2784464, 0.2566211, 0.1746921, 0.1352786, 
    0.038876, 0.02280528, 0.04275943, 0.1385308, 0.1709292,
  0.02150327, 0.0007482755, 0.003785497, 5.250462e-05, 2.516912e-05, 
    0.02763034, 0.2770939, 0.08176255, 0.1404101, 0.08229797, 0.09269437, 
    0.1492788, 0.1090086, 0.05252239, 0.07954659, 0.03635963, 0.00102502, 
    1.891912e-06, 9.410824e-07, 0.01591142, 0.04993341, 0.1258877, 0.0840098, 
    0.1150387, 0.07986093, 0.05352274, 0.02793665, 0.002753596, 0.07628677,
  0.04883644, 0.02512616, -5.450352e-07, 2.332317e-07, -4.118863e-09, 
    3.694631e-08, 0.001235138, 0.108972, 0.1458862, 0.1191092, 0.04943356, 
    0.06625677, 0.07139302, 0.02584215, 0.0691496, 0.03669675, 0.06575503, 
    0.00993646, 0.0003026986, -7.651349e-07, 0.1170593, 0.0808137, 
    0.07977337, 0.1119082, 0.08684866, 0.03244987, 0.04086819, 0.02404607, 
    0.009160484,
  0.109493, 0.116786, 0.02531766, 0.001411273, 0.02494824, 0.01275106, 
    0.01060052, 0.1218321, 0.1251729, 0.1172491, 0.2237948, 0.2717805, 
    0.1717906, 0.1158787, 0.110568, 0.2405566, 0.1430975, 0.1057208, 
    0.0236574, 0.04868699, 0.1340138, 0.1344187, 0.1030095, 0.1126548, 
    0.1365498, 0.09674596, 0.07183652, 0.05848883, 0.08585039,
  0.06667004, 0.1619975, 0.1535149, 0.08532826, 0.06333537, 0.08675205, 
    0.01624576, 0.006437869, 0.009621928, 0.0441739, 0.08647832, 0.1256555, 
    0.137962, 0.190685, 0.1436604, 0.09346177, 0.2368679, 0.2418214, 
    0.1796789, 0.05122094, 0.04700966, 0.1379354, 0.1285497, 0.09428123, 
    0.1827978, 0.2058198, 0.2164999, 0.1950472, 0.1314497,
  0.1007648, 0.0369077, 0.05636443, 0.04670456, 0.02552355, 0.02389573, 
    0.08490101, 0.03263997, 0.01588801, 0.02322624, 0.03869565, 0.03510408, 
    0.02858406, 0.03108389, 0.03651362, 0.06113816, 0.0502281, 0.07712855, 
    0.03396033, 0.04015234, 0.04585412, 0.09179386, 0.03908613, 0.06777912, 
    0.07345571, 0.09441884, 0.08777432, 0.05502687, 0.09001204,
  0.00756898, 0.01021862, 0.0004474391, 0.004498954, 0.003807863, 
    -0.0002932216, 0.008349958, -0.0004665253, 0, 0, -1.389781e-10, 0, 0, 
    0.002698348, 0.01925397, 0.01994147, 0.04035382, 0.02494221, 0.03021627, 
    0.03425408, 0.03142706, 0.01627851, -3.085882e-05, 0.005570211, 
    0.04092983, -8.749276e-05, 8.080952e-06, 0.03365395, 0.01289797,
  0.001686445, -0.0001615789, 0.0005604056, 0.0002539717, -2.703648e-05, 0, 
    0, -2.724304e-05, 0.001919897, -3.743836e-05, 0, 0, 0, 0, 0, 
    0.0001564089, 0.001526601, 0.005170454, 0.01130772, 0.01194367, 
    0.0004459496, -7.01617e-05, -3.831844e-08, 0, 0, 0, -2.022726e-09, 
    -0.0006520745, 0.002490528,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -5.582838e-06, 
    -0.0002498452, 0.0005127584, 0.006662949, 0.02151997, 0.0003892461, 
    -4.353896e-06, 0, 0,
  0.004352794, 0, 0, -2.908622e-05, -7.808371e-05, -0.0001892905, 0.01024659, 
    0.01689331, 0.01250726, 0.004378003, -7.89294e-05, -2.027341e-05, 
    0.001305674, 0.007671513, 0.003440336, 0.00515745, -7.370303e-06, 
    0.0003426307, 0.008842719, 0.01551838, 0.0167994, 0.02489088, 
    0.002813788, 0.004727062, 0.0003473928, -0.000187116, -7.917527e-08, 
    0.001197308, 0.004149506,
  0.04437295, 0.05256199, 0.06555577, 0.1046025, 0.1517474, 0.1387542, 
    0.1000607, 0.08263572, 0.0302997, 0.008729478, 0.01624111, 0.07028932, 
    0.08482974, 0.03833789, 0.04435672, 0.03414779, 0.05723745, 0.07196823, 
    0.0484411, 0.1008836, 0.07798184, 0.06861364, 0.02917676, 0.002457773, 
    0.01765311, 0.05348302, 0.04843235, 0.08243094, 0.0592146,
  0.1670038, 0.08759395, 0.1256422, 0.1776876, 0.1244804, 0.09311369, 
    0.09706864, 0.07029553, 0.0546635, 0.04304499, 0.04387235, 0.06830946, 
    0.0740568, 0.1103968, 0.1070245, 0.1030234, 0.08604164, 0.09589823, 
    0.2026392, 0.1117443, 0.1318256, 0.07076079, 0.06529252, 0.05535943, 
    0.08478033, 0.1041735, 0.185898, 0.1215696, 0.1803023,
  0.0592203, 0.01088839, 0.0293907, 0.008903911, 0.00117981, 4.615748e-05, 
    0.0001002564, -0.0002108465, 0.001633536, 0.003071728, -6.923876e-05, 
    0.006962928, 0.006639921, 0.03857655, 0.07421983, 0.08309681, 0.110474, 
    0.1306459, 0.1959325, 0.1063422, 0.03360489, 0.03346195, 0.003250043, 
    0.001164301, 0.04674978, 0.09122545, 0.0504178, 0.02734526, 0.06137502,
  1.021738e-06, -3.205624e-05, 0.01281667, 6.19297e-06, -1.321917e-08, 
    0.004876672, 1.416372e-06, 4.169203e-05, 2.545768e-07, 9.087318e-07, 
    3.648017e-08, -1.121325e-07, 0.002787425, 0.02954721, 0.04945672, 
    0.08134001, 0.03253839, 0.05031991, 0.0004941507, 6.543029e-07, 
    9.720218e-09, 8.853354e-08, 1.042742e-07, 0.0154416, 0.0257, 0.00790257, 
    3.381075e-06, -1.076957e-05, 1.457706e-07,
  6.80142e-07, -3.704585e-05, 0.004544664, -1.070025e-06, 0.003598237, 
    0.0001495138, 0.03390273, 0.01251581, 6.146621e-05, 0.001028296, 
    0.024651, 0.03252478, 0.07587424, 0.1048041, 0.07263488, 0.02753184, 
    0.0110517, -1.106453e-06, -6.076538e-10, 7.623341e-06, 3.008806e-06, 
    1.328188e-06, 1.903179e-05, 0.03028994, 0.00764321, -8.034508e-10, 
    8.778078e-07, 9.647847e-08, -2.154482e-09,
  8.922828e-05, 0.3544326, 0.1618172, 0.004394645, 0.0008697346, 0.121415, 
    0.03119583, 0.1801972, 0.1650366, 0.1741786, 0.01687449, 0.03989585, 
    0.05416001, 0.04700607, 0.003420954, 4.669376e-06, 9.279735e-07, 
    -1.815847e-08, 1.908287e-06, -1.607542e-05, 5.240417e-05, 0.0004986056, 
    0.02019683, 0.1392588, 0.003664742, -3.031916e-06, 1.68304e-06, 
    2.340056e-05, -2.958301e-05,
  0.1302167, 0.1644838, 0.1100064, 0.02489359, 0.0006215021, 0.0001544459, 
    0.01109966, 0.07462925, 0.1885847, 0.08469539, 0.03296272, 0.1382789, 
    0.1330498, 0.1213482, 0.1051281, 0.1428341, 0.04863888, 0.02728384, 
    0.01216307, 0.04851434, 0.2582169, 0.2563232, 0.132835, 0.0891647, 
    0.03235311, 0.02293468, 0.04122049, 0.1229917, 0.1498977,
  0.02467402, 0.001897666, 0.001927655, 7.989743e-05, 0.0004268007, 
    0.01440809, 0.2460148, 0.07078046, 0.1113753, 0.07767992, 0.07067221, 
    0.1321961, 0.08438548, 0.03972094, 0.05935884, 0.02156097, 5.495119e-05, 
    1.47174e-06, 5.07009e-07, 0.03654095, 0.04370767, 0.1128239, 0.05883781, 
    0.09068654, 0.06425635, 0.035186, 0.03662129, 0.004406611, 0.06195192,
  0.04986061, 0.003684017, 2.955137e-07, 1.850731e-07, -3.031301e-09, 
    -3.18201e-09, 0.001503137, 0.1262938, 0.1564493, 0.1547771, 0.0471922, 
    0.06096628, 0.03772934, 0.01837681, 0.06132415, 0.02831568, 0.04063828, 
    0.007672336, 5.299905e-05, 0.0001213609, 0.08731989, 0.07688213, 
    0.07777312, 0.09765104, 0.080499, 0.02384126, 0.01487581, 0.01084427, 
    0.003629289,
  0.09217095, 0.09654217, 0.01160937, 0.004354103, 0.02018909, 0.01433068, 
    0.01869087, 0.1685341, 0.144258, 0.1281746, 0.1952289, 0.2847063, 
    0.1681185, 0.1189108, 0.09491388, 0.2727026, 0.1357157, 0.1548562, 
    0.01696879, 0.0450391, 0.1122592, 0.1132618, 0.09815412, 0.102399, 
    0.1324287, 0.08986675, 0.06358892, 0.05923165, 0.07265365,
  0.07865754, 0.1847446, 0.1533006, 0.09752891, 0.1209291, 0.1393588, 
    0.07407992, 0.02491433, 0.05243056, 0.1499371, 0.1461688, 0.1547573, 
    0.1489108, 0.2101862, 0.1859258, 0.08936717, 0.263602, 0.2384644, 
    0.1764297, 0.1251759, 0.06978551, 0.1186282, 0.1459869, 0.1380101, 
    0.1758459, 0.2203249, 0.212239, 0.1754131, 0.1523981,
  0.1785842, 0.1116786, 0.1080474, 0.07827853, 0.1046738, 0.1274136, 
    0.1334945, 0.1725447, 0.1302369, 0.08896595, 0.06277017, 0.07087589, 
    0.08593298, 0.1543414, 0.1078526, 0.138423, 0.1320042, 0.1218198, 
    0.08905508, 0.1062995, 0.0891538, 0.1889369, 0.1293627, 0.1121254, 
    0.1321984, 0.1355752, 0.1319107, 0.1127958, 0.1417204,
  0.07759313, 0.09188836, 0.05047585, 0.1205244, 0.1814469, 0.1545419, 
    0.1235698, 0.1142913, 0.05084669, 0.01022939, -2.272847e-05, 
    6.317787e-07, 0.03112485, 0.0285545, 0.07527772, 0.09381387, 0.08933777, 
    0.08521629, 0.05793643, 0.05939127, 0.0476357, 0.03330191, 0.02324012, 
    0.03659752, 0.09732071, 0.0004183001, -0.0004368837, 0.1159859, 0.08994251,
  0.07643438, 0.09712832, 0.06498238, 0.0557156, 0.04553844, 0.0441667, 
    0.05430964, 0.05502839, 0.02941821, 0.01563545, -0.0003071315, 
    -8.047418e-06, 0, -5.25384e-08, 2.614355e-05, 0.003864535, 0.007719086, 
    0.01461229, 0.03203524, 0.03327991, 0.01684444, 0.004718182, 
    -1.510452e-05, -3.142456e-05, -7.75979e-06, -8.551686e-08, -0.0008588847, 
    0.008958942, 0.0830179,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.0002575941, -0.0001521201, 0,
  8.244292e-05, -1.368634e-09, 0.001459625, 0, 0, 0, 0, 0, 0, 0, 0, 
    -1.36214e-05, 0, -0.0002532503, 0.0005876645, -0.0001187477, 
    -7.569337e-06, 0.0005612294, 0, -0.0002345146, 0.001859936, 0.01500141, 
    0.01589538, 0.0356832, 0.03641725, 0.003014192, 0.01291342, 0.005793047, 
    0.00363584,
  0.01621065, 0.01325015, 0.009164746, 0.001762977, 0.004503425, 0.004744656, 
    0.01910269, 0.01927995, 0.01754301, 0.02172567, 0.0261391, 0.03708328, 
    0.08943389, 0.08645912, 0.06409238, 0.09036602, 0.05022256, 0.05098448, 
    0.06985004, 0.04923541, 0.04461487, 0.04750696, 0.05413108, 0.05370731, 
    0.01167445, 0.01848437, 0.01811857, 0.01620262, 0.01609768,
  0.1404595, 0.1945732, 0.1399602, 0.1862548, 0.2031359, 0.178386, 0.1245392, 
    0.1163618, 0.1031017, 0.1080012, 0.1850027, 0.1607433, 0.1575132, 
    0.1179593, 0.12195, 0.129959, 0.1713773, 0.1641282, 0.116544, 0.1978455, 
    0.1429028, 0.1444495, 0.1143686, 0.02807393, 0.09579283, 0.1265555, 
    0.1031268, 0.1434926, 0.1143896,
  0.1830064, 0.07426605, 0.1228591, 0.1743293, 0.1106474, 0.08183158, 
    0.09760936, 0.08154, 0.08190662, 0.07441615, 0.05354047, 0.07507192, 
    0.111284, 0.1762907, 0.1379772, 0.1400137, 0.09261221, 0.130638, 
    0.176416, 0.1266518, 0.1300219, 0.08663389, 0.1048963, 0.07762992, 
    0.07160719, 0.1139585, 0.1877197, 0.1178174, 0.1909529,
  0.05459714, 0.002732979, 0.02149316, 0.007143259, 0.000814941, 
    3.386465e-07, -0.0001577174, -0.0003247228, 0.006020704, 0.00606382, 
    0.001143274, 0.007581932, 0.01648219, 0.04546443, 0.08647644, 0.08775508, 
    0.08504562, 0.115452, 0.190336, 0.07879324, 0.02040818, 0.01290687, 
    0.00742619, 0.0004617572, 0.04504066, 0.0715385, 0.03585004, 0.02549034, 
    0.06327885,
  8.244555e-08, 0.0002656494, 0.01565116, 3.30392e-06, -6.284069e-08, 
    0.03088222, 2.508651e-08, 4.647039e-06, 2.607263e-07, 8.966808e-07, 
    3.743366e-08, -7.840559e-08, 0.0003982145, 0.03297278, 0.04491251, 
    0.1003389, 0.01825735, 0.05228291, 0.0003087972, -1.757247e-06, 
    8.314495e-09, -1.01759e-09, 7.687567e-09, 0.01485259, 0.0177462, 
    0.004193466, 6.021911e-06, -1.725946e-05, 6.976687e-08,
  8.130264e-07, 0.001278263, 0.001692184, 4.374866e-05, 0.006482663, 
    9.261135e-05, 0.03633749, 0.009628806, 0.0003296344, 0.001014365, 
    0.0415735, 0.04730447, 0.07915378, 0.09400374, 0.06286325, 0.02079912, 
    0.01214129, -9.509512e-07, -1.151028e-10, 9.699078e-07, 8.668969e-07, 
    5.442404e-07, 6.820333e-06, 0.02532366, 0.004567268, 8.163468e-10, 
    2.202434e-07, 9.440868e-09, 3.707733e-08,
  2.960982e-05, 0.3308604, 0.1276382, 0.004688219, 0.001733068, 0.1053225, 
    0.02483333, 0.1278336, 0.1013206, 0.1852408, 0.0152672, 0.03224632, 
    0.04679271, 0.02912142, 0.003998375, 8.608507e-05, 2.419901e-06, 
    -7.230108e-05, 9.33255e-07, -4.503708e-05, 2.066331e-05, 1.249032e-05, 
    0.01976725, 0.1027835, 0.004621179, -5.523299e-06, -3.004095e-06, 
    6.727482e-06, 0.0001027874,
  0.1195713, 0.144977, 0.1007283, 0.03350395, 0.0020628, 0.0002446976, 
    0.0100987, 0.03392482, 0.1311782, 0.06927292, 0.02018187, 0.09970843, 
    0.08971174, 0.09396007, 0.07524487, 0.1355635, 0.04752563, 0.03087427, 
    0.02162312, 0.08119112, 0.2095206, 0.2233824, 0.1133011, 0.06300244, 
    0.0284627, 0.01779374, 0.04204962, 0.1164092, 0.1299341,
  0.02163659, 0.001016158, 0.0007337934, 0.0001827125, 0.000345647, 
    0.02578207, 0.2252446, 0.07034454, 0.08221637, 0.07723999, 0.06273636, 
    0.1079848, 0.07416972, 0.02725865, 0.03934196, 0.01405944, 2.1879e-05, 
    9.720195e-07, 4.202476e-07, 0.03114378, 0.04069696, 0.1113136, 
    0.03486471, 0.06266452, 0.05204769, 0.0264225, 0.05042759, 0.005934304, 
    0.04138745,
  0.05629255, 0.0009045877, -4.395543e-09, 5.611501e-07, -4.954727e-06, 
    3.655635e-08, 0.00137537, 0.1192354, 0.1603317, 0.1384244, 0.04329308, 
    0.04849989, 0.01693552, 0.01339313, 0.05979107, 0.02339469, 0.02696785, 
    0.001303592, 2.862464e-07, -0.0003084954, 0.05624734, 0.0636835, 
    0.06401791, 0.07552569, 0.0732417, 0.01973888, 0.009878812, 0.002343996, 
    0.0002046875,
  0.08372659, 0.08676704, 0.005203185, 0.0009878618, 0.01795897, 0.01164285, 
    0.03727466, 0.155909, 0.1443948, 0.1030665, 0.1626038, 0.281274, 
    0.1678591, 0.1279538, 0.07738332, 0.2525151, 0.1263546, 0.09326328, 
    0.02154527, 0.03753123, 0.06844945, 0.09216188, 0.09506085, 0.1061288, 
    0.1090073, 0.0828578, 0.05228153, 0.04931766, 0.05790665,
  0.0713489, 0.1778243, 0.1218531, 0.08990803, 0.1378455, 0.1308855, 
    0.07422689, 0.08719853, 0.104102, 0.1766649, 0.1638168, 0.1509781, 
    0.141587, 0.1994739, 0.1936497, 0.07793047, 0.2844319, 0.2267087, 
    0.1537412, 0.1724116, 0.07888865, 0.1034292, 0.148176, 0.1498551, 
    0.1695126, 0.2189882, 0.2100904, 0.1675226, 0.1434947,
  0.2268323, 0.1771106, 0.1046122, 0.1739678, 0.1831806, 0.1164882, 0.142357, 
    0.1514059, 0.1668819, 0.1698716, 0.1337842, 0.1572963, 0.1522925, 
    0.2001516, 0.2014118, 0.1624949, 0.1762423, 0.1632712, 0.1909468, 
    0.1177393, 0.1093536, 0.2358723, 0.2053809, 0.1919386, 0.1863008, 
    0.1568464, 0.1764897, 0.1435834, 0.1699783,
  0.1731318, 0.1289409, 0.1408645, 0.1591129, 0.2275261, 0.2374209, 
    0.1584163, 0.1298855, 0.1168236, 0.1506743, 0.1216562, 0.05791252, 
    0.1457512, 0.1228066, 0.181269, 0.1695896, 0.1540414, 0.1539028, 
    0.1024491, 0.09434773, 0.06645777, 0.0575452, 0.09757356, 0.09578184, 
    0.3013163, 0.00900265, 0.0006252165, 0.2405534, 0.1432007,
  0.2359238, 0.2416182, 0.1631989, 0.1643782, 0.205925, 0.1991929, 0.19584, 
    0.1646097, 0.12326, 0.09685346, 0.09918784, 0.0709975, 0.05792988, 
    0.03720869, 0.03853146, 0.04481362, 0.05863006, 0.06052231, 0.07648761, 
    0.06979404, 0.05720327, 0.05936535, 0.01787164, -0.005321569, 0.01338144, 
    0.0002701214, -0.006337801, 0.05409595, 0.2134636,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -1.273836e-06, -7.898413e-05, -1.384659e-05, 0, 0.0007139671, 
    -0.0003978056, 0,
  0.001088132, 0.0007343091, 0.001922605, 0, 0, -1.130502e-06, 0, 0, 0, 0, 0, 
    -8.651164e-05, -0.0008985366, 0.0290863, 0.0205415, 0.01469441, 
    0.01570494, 0.03878737, 0.02432441, 0.009434808, 0.02956103, 0.04994059, 
    0.03633443, 0.0540526, 0.06647019, 0.01011393, 0.02537846, 0.02296496, 
    0.01994431,
  0.03140083, 0.03022461, 0.0337887, 0.02962383, 0.03783871, 0.06189762, 
    0.05511387, 0.05274033, 0.03954377, 0.03463724, 0.09312331, 0.1290346, 
    0.1759838, 0.1968818, 0.1976639, 0.2186037, 0.2086553, 0.2129203, 
    0.1190631, 0.1295784, 0.1139706, 0.1327161, 0.1069964, 0.1178002, 
    0.07866285, 0.08319294, 0.0994657, 0.09412542, 0.06223729,
  0.1745311, 0.2340149, 0.1867585, 0.2593757, 0.1997257, 0.2129529, 
    0.1691349, 0.1597626, 0.1222144, 0.1638419, 0.228879, 0.1789383, 
    0.1756095, 0.1467202, 0.2008925, 0.1883934, 0.269045, 0.2355218, 
    0.1867297, 0.2640748, 0.1876992, 0.1738072, 0.1836369, 0.09980794, 
    0.1640404, 0.160219, 0.1342512, 0.1956406, 0.1497535,
  0.1785156, 0.06588217, 0.1173188, 0.1665338, 0.09274056, 0.08301188, 
    0.09029996, 0.07160185, 0.08721937, 0.06847364, 0.04096261, 0.08592106, 
    0.1027756, 0.1658609, 0.1635518, 0.1657492, 0.1021343, 0.1301434, 
    0.1636051, 0.1432729, 0.1445767, 0.09527171, 0.09690836, 0.09121819, 
    0.05745954, 0.1059824, 0.1752177, 0.1299662, 0.1878653,
  0.0397926, 0.0001970544, 0.01912154, 0.01653535, 0.0001552537, 
    -1.168831e-07, 0.0004491494, -2.401645e-06, 0.0004104377, 0.005228907, 
    0.01858916, 0.02686951, 0.02977557, 0.05318963, 0.07262437, 0.07262092, 
    0.07557462, 0.1056299, 0.1607572, 0.06139555, 0.02249454, 0.004637263, 
    0.003038802, 3.650737e-07, 0.0398306, 0.05132221, 0.03086003, 0.02550745, 
    0.06020246,
  -1.287904e-10, 0.0005303516, 0.01270431, 5.017436e-06, -1.057448e-07, 
    0.03199779, -1.413756e-10, 1.65656e-05, -9.763691e-07, 6.72707e-07, 
    5.056987e-08, 2.446127e-07, 0.0003116939, 0.02499851, 0.03823582, 
    0.09889045, 0.01812586, 0.04332804, 0.0003158146, -5.903531e-07, 
    8.51673e-09, 0, 4.177795e-09, 0.01393055, 0.01058249, 0.003936441, 
    1.40459e-05, -2.309934e-05, 8.110716e-08,
  9.682627e-07, 0.01857753, -4.415616e-05, 3.03688e-06, 0.00783738, 
    0.00108244, 0.0479868, 0.00724169, 0.001944058, 0.001261078, 0.04340086, 
    0.07555945, 0.1231319, 0.09239445, 0.04148389, 0.01699835, 0.01085569, 
    1.907827e-06, -2.072663e-10, 6.710694e-08, 6.380612e-07, 1.293706e-07, 
    6.072999e-07, 0.02229769, 0.003542786, -4.130456e-08, 4.362872e-08, 
    5.870823e-08, 1.43325e-07,
  3.086189e-05, 0.3126931, 0.1025762, 0.0015595, 0.002729127, 0.1049786, 
    0.02123045, 0.09992811, 0.05904272, 0.1910844, 0.01497216, 0.02722768, 
    0.04049416, 0.01868117, 0.005607827, 0.0003294993, 2.90769e-06, 
    -0.0003609874, -3.803908e-05, -0.0001570121, 1.39802e-05, 7.077911e-06, 
    0.02096911, 0.0630054, 0.004131121, 6.740282e-05, -2.192262e-05, 
    1.183616e-06, 0.0008765057,
  0.105352, 0.1243853, 0.09929667, 0.03372238, 0.001266839, 0.0004101091, 
    0.01925243, 0.01830996, 0.1093969, 0.06303877, 0.01403695, 0.07711811, 
    0.06510556, 0.08400699, 0.05856688, 0.1278795, 0.04506319, 0.0389397, 
    0.03965239, 0.1161039, 0.1970336, 0.1995053, 0.1046254, 0.0478173, 
    0.0237884, 0.01810777, 0.04647452, 0.1176086, 0.1205169,
  0.01825218, 0.0003248967, 0.0008352581, 0.0005828422, -0.0001196248, 
    0.03295984, 0.1549293, 0.0727318, 0.07713509, 0.07667296, 0.06248755, 
    0.09283188, 0.07591156, 0.02076999, 0.0246228, 0.009108104, 1.968195e-05, 
    5.181813e-07, 2.58813e-07, 0.03516343, 0.04289772, 0.1229507, 0.02408224, 
    0.04319005, 0.04275001, 0.02456844, 0.04097736, 0.002448467, 0.02695793,
  0.04501541, 0.00010882, -2.367821e-08, 2.105205e-05, -8.256912e-05, 
    1.397109e-07, 0.002614713, 0.1159983, 0.1698685, 0.1293501, 0.02670874, 
    0.04102875, 0.008371621, 0.01168892, 0.06126606, 0.01469798, 0.007086596, 
    6.890108e-05, 1.112742e-07, -8.215749e-06, 0.03624954, 0.04425017, 
    0.05162879, 0.06485709, 0.06211931, 0.01498685, 0.004935028, 
    0.0002823401, 0.0001838286,
  0.07329497, 0.09744885, 0.002813227, 0.0006482484, 0.01961153, 0.01440866, 
    0.05308104, 0.1286577, 0.1257223, 0.08959647, 0.1277234, 0.2991087, 
    0.1495327, 0.1189784, 0.08501613, 0.2407863, 0.1315385, 0.08264218, 
    0.01195421, 0.03295407, 0.0435022, 0.0805774, 0.07193665, 0.1042686, 
    0.08773591, 0.07454459, 0.05471452, 0.04544111, 0.05229941,
  0.09494635, 0.1588848, 0.1038463, 0.07980019, 0.1288817, 0.1251832, 
    0.06462777, 0.1531074, 0.128148, 0.1802269, 0.1655576, 0.145065, 
    0.1323215, 0.1822795, 0.1916468, 0.08147597, 0.2801344, 0.2362154, 
    0.1283452, 0.1669905, 0.064562, 0.09489482, 0.1553646, 0.1502883, 
    0.1587088, 0.2093449, 0.2167154, 0.1730816, 0.1353691,
  0.2265398, 0.1679593, 0.09565294, 0.1861423, 0.1944321, 0.1264954, 
    0.1704942, 0.1643908, 0.145611, 0.1922811, 0.169961, 0.2010878, 
    0.2083834, 0.2357863, 0.2538171, 0.2022719, 0.1832991, 0.2448014, 
    0.2168505, 0.122764, 0.1318335, 0.2754331, 0.1952765, 0.2248686, 
    0.2200687, 0.1827665, 0.1780764, 0.1401166, 0.2078236,
  0.1792959, 0.1336493, 0.1367046, 0.1559825, 0.2246149, 0.220747, 0.1686718, 
    0.1718772, 0.1239762, 0.1935838, 0.1933984, 0.2861784, 0.1912655, 
    0.153163, 0.1830528, 0.1869801, 0.1787496, 0.1686693, 0.148032, 
    0.1625717, 0.1486743, 0.09061512, 0.107946, 0.2397374, 0.28728, 
    0.04462345, 0.007487915, 0.2543853, 0.1742598,
  0.2164436, 0.2262177, 0.1640487, 0.1847697, 0.1954056, 0.1891074, 
    0.2168184, 0.1998473, 0.1957247, 0.2406262, 0.1861622, 0.1202528, 
    0.1361821, 0.1303764, 0.1474222, 0.167566, 0.1792014, 0.2142248, 
    0.2864307, 0.2299627, 0.1417428, 0.1148179, 0.1194222, 0.04555225, 
    0.06826707, 0.01528847, 0.04558136, 0.09566537, 0.2164414,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0009559893, 0.009289428, 
    0.01338478, 0.006847128, -0.0001567107, 0, 0, -1.029607e-05, 
    -2.37549e-05, 0.005845896, 0.02014387, 0.01549128, -0.002040306, 
    0.003887674, 0.0004156315, 0,
  0.03255113, 0.01408489, 0.002110112, 0.00015368, 0, -1.151054e-05, 
    0.002137916, 0, 0, 0, -7.931794e-06, -0.0001321345, -0.001456764, 
    0.07616261, 0.06445645, 0.1102654, 0.1486306, 0.1587438, 0.1225869, 
    0.09055531, 0.1479684, 0.144379, 0.1173922, 0.1529213, 0.1480081, 
    0.06362839, 0.08735957, 0.08167297, 0.05713629,
  0.08600756, 0.08226428, 0.1101318, 0.1349257, 0.1170842, 0.1249883, 
    0.132968, 0.13191, 0.1240577, 0.1231044, 0.1837767, 0.2173877, 0.2638418, 
    0.2826684, 0.2302327, 0.258091, 0.2203215, 0.2479028, 0.154677, 
    0.1634713, 0.1414946, 0.1662584, 0.1420278, 0.2013805, 0.129875, 
    0.1449054, 0.1725979, 0.1723801, 0.1546719,
  0.1998429, 0.2385704, 0.1964974, 0.2587271, 0.1877317, 0.2179644, 
    0.1782655, 0.1729868, 0.1541744, 0.1893644, 0.2325385, 0.1659132, 
    0.1643752, 0.1473496, 0.1872419, 0.1656623, 0.2346627, 0.2173793, 
    0.1653388, 0.255952, 0.2115837, 0.1985952, 0.2109848, 0.1446075, 
    0.1722205, 0.1635314, 0.1400156, 0.2169211, 0.1890142,
  0.1628711, 0.0471398, 0.1014014, 0.155616, 0.08891612, 0.09880986, 
    0.07865139, 0.07255448, 0.08376348, 0.05089762, 0.03288807, 0.08629031, 
    0.08362816, 0.153976, 0.1633612, 0.170631, 0.1208374, 0.1233946, 
    0.1515959, 0.1445485, 0.1535165, 0.108135, 0.1042108, 0.09258106, 
    0.05240696, 0.09068654, 0.165191, 0.1345918, 0.1849553,
  0.02517771, 0.006832821, 0.02103112, 0.03128442, 0.0001300451, 
    -1.206743e-06, 6.536466e-05, -3.910823e-06, 0.002519084, 0.002456705, 
    0.02886264, 0.0327038, 0.03726212, 0.05351573, 0.0836475, 0.07153564, 
    0.08706171, 0.09708226, 0.1509838, 0.04019548, 0.006513648, 0.0008845515, 
    0.00261068, 7.503121e-06, 0.04085176, 0.04398606, 0.03640475, 0.03224321, 
    0.05864939,
  -8.709874e-10, 0.005536149, 0.01247857, 1.356548e-05, 3.373459e-09, 
    0.02657236, -7.634258e-10, 8.44649e-05, 0.001570772, 3.701637e-07, 
    3.646786e-05, 3.729915e-07, 0.001057482, 0.03301488, 0.03374865, 
    0.1039295, 0.01842229, 0.03433499, 0.000162758, -1.775387e-08, 0, 0, 
    -6.728715e-10, 0.01315064, 0.01082281, 0.003337371, -9.293541e-06, 
    -3.079531e-05, 5.556704e-08,
  7.010624e-07, 0.002600953, 0.0005336548, 3.472627e-05, 0.006272528, 
    0.003142352, 0.08190067, 0.005582591, 0.0005887139, 0.001482489, 
    0.05496723, 0.08819896, 0.1219462, 0.09609143, 0.04596931, 0.01889108, 
    0.008927466, 3.072992e-06, -3.765745e-11, 8.747404e-08, 2.74926e-07, 
    4.106163e-08, 9.498328e-08, 0.02597135, 0.003261597, -9.975198e-09, 
    1.200435e-08, 2.088788e-07, 2.850946e-07,
  0.001288551, 0.2831298, 0.1121101, 0.0008002315, 0.004439885, 0.1014911, 
    0.01802232, 0.08673562, 0.03829002, 0.1881365, 0.01281051, 0.02391378, 
    0.03814082, 0.01245556, 0.007623957, 0.0008233875, 1.75306e-06, 
    0.00126826, -4.364881e-05, -0.0002701944, 5.372736e-06, 1.871654e-05, 
    0.02273245, 0.04557413, 0.00457358, -4.685858e-06, -0.0001725964, 
    0.0001444899, 0.023762,
  0.09773288, 0.1110727, 0.1034499, 0.03587617, 0.001686066, 0.001395943, 
    0.01955926, 0.01292055, 0.1092634, 0.06392315, 0.01244593, 0.06997038, 
    0.04873344, 0.07591532, 0.05057405, 0.1375424, 0.04220562, 0.04085184, 
    0.06947252, 0.150978, 0.1816717, 0.1907647, 0.101133, 0.0341064, 
    0.02126289, 0.02388197, 0.06289927, 0.1231535, 0.1052176,
  0.0111329, 0.0001130521, 0.002079949, 0.005020065, 0.000967481, 0.0538042, 
    0.1124859, 0.07091884, 0.08006097, 0.1019658, 0.06408799, 0.09749957, 
    0.07127766, 0.01615913, 0.0212446, 0.007257588, 3.782174e-06, 
    3.630181e-07, 1.83257e-07, 0.03476035, 0.05013414, 0.1210806, 0.02688266, 
    0.03336256, 0.03194165, 0.02631474, 0.02572925, 0.002967364, 0.01609751,
  0.03677626, 6.51103e-05, -6.649224e-09, 0.0003649908, -5.58007e-05, 
    4.580668e-07, 0.004080381, 0.1178464, 0.1857017, 0.1519774, 0.02781812, 
    0.03904164, 0.005397531, 0.01009043, 0.0607483, 0.01593835, 0.002923646, 
    1.241958e-05, 1.490243e-07, 1.801777e-06, 0.02877783, 0.04007664, 
    0.05404813, 0.06054135, 0.04800972, 0.01423852, 0.002144341, 
    9.450346e-05, 0.0004549884,
  0.05762864, 0.1008554, 0.001897165, 0.0009336254, 0.02952151, 0.01631093, 
    0.06628253, 0.08494575, 0.106849, 0.0883086, 0.1071966, 0.2716167, 
    0.1441074, 0.1161401, 0.07976461, 0.2335515, 0.1402645, 0.04091617, 
    0.01526533, 0.04469186, 0.03004481, 0.06554601, 0.06388532, 0.09845846, 
    0.07121695, 0.06465635, 0.03386308, 0.03422206, 0.05704035,
  0.1139599, 0.140574, 0.0929988, 0.07416172, 0.1070908, 0.113779, 
    0.05525174, 0.1408853, 0.1235067, 0.176456, 0.1728683, 0.1394771, 
    0.1167893, 0.1724974, 0.1760979, 0.09245095, 0.2411283, 0.1877753, 
    0.1117495, 0.1506571, 0.05611403, 0.1022895, 0.1632217, 0.1592155, 
    0.1459693, 0.1834633, 0.2026066, 0.1632164, 0.1196674,
  0.222276, 0.1591095, 0.08578467, 0.1898562, 0.1998816, 0.1371398, 
    0.1815174, 0.1560539, 0.1564923, 0.1616112, 0.149658, 0.1961209, 
    0.2102982, 0.2266909, 0.2774293, 0.1894106, 0.1832862, 0.2685518, 
    0.2156182, 0.1262224, 0.139268, 0.271683, 0.1949468, 0.2076899, 
    0.2237696, 0.2139609, 0.1950855, 0.1489942, 0.2116767,
  0.1990415, 0.1453434, 0.1342958, 0.1496907, 0.2256528, 0.1999715, 
    0.1660565, 0.1859032, 0.1202695, 0.1789489, 0.2184197, 0.3027516, 
    0.2037962, 0.1489665, 0.1765875, 0.1827321, 0.1837126, 0.1650389, 
    0.1392704, 0.1569501, 0.2281071, 0.1270196, 0.1819586, 0.2988392, 
    0.2909982, 0.09933571, 0.05501365, 0.2373412, 0.1718337,
  0.2342883, 0.2264026, 0.1437218, 0.176181, 0.1765239, 0.2008672, 0.2209391, 
    0.2029933, 0.211063, 0.2642492, 0.2421577, 0.1862845, 0.1994606, 
    0.1955737, 0.2067921, 0.2224499, 0.216176, 0.2504413, 0.2919049, 
    0.2999569, 0.214535, 0.2014034, 0.1491679, 0.1183645, 0.1176416, 
    0.05568337, 0.08772965, 0.1029366, 0.2162222,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0186984, 0.02237584, 0.02739592, 
    0.03178817, 0.009728521, -4.929684e-06, 0, -0.0002762178, 7.403832e-05, 
    0.01327787, 0.06995887, 0.07836303, 0.06330281, 0.08336211, 0.002450158, 0,
  0.05621566, 0.04271669, 0.03825869, 0.007050585, -0.0006058022, 
    0.001594678, 0.02115606, -2.37819e-05, 0, -0.0002620796, -0.0003444215, 
    -0.0007237952, 0.0399087, 0.1564193, 0.1846301, 0.2188504, 0.2002299, 
    0.1972947, 0.1734235, 0.144171, 0.1924332, 0.2198751, 0.1981903, 
    0.2512149, 0.2543611, 0.1804585, 0.2255116, 0.2128289, 0.09930044,
  0.1248484, 0.1539992, 0.161495, 0.18548, 0.1521859, 0.1370395, 0.1652842, 
    0.1796788, 0.1700308, 0.1653229, 0.2362459, 0.2563834, 0.2780423, 
    0.3346305, 0.2520688, 0.2458199, 0.2013527, 0.2233376, 0.1643698, 
    0.1697789, 0.1573278, 0.1826009, 0.1748748, 0.2091739, 0.1493018, 
    0.1697384, 0.1996614, 0.1955847, 0.1931482,
  0.1827416, 0.2331168, 0.2192074, 0.2293481, 0.1768212, 0.2277075, 
    0.1919828, 0.1813964, 0.1649918, 0.1885373, 0.2221263, 0.1587296, 
    0.1687148, 0.1319144, 0.1828976, 0.1650435, 0.1954274, 0.189199, 
    0.169038, 0.2331422, 0.2082843, 0.2008815, 0.203267, 0.1742532, 
    0.1676851, 0.1478301, 0.1415205, 0.2105684, 0.1817723,
  0.1506315, 0.04790118, 0.09245105, 0.1547906, 0.09421881, 0.1093855, 
    0.07638486, 0.0729273, 0.07187413, 0.0418519, 0.0307408, 0.09196207, 
    0.07496416, 0.1474874, 0.1648602, 0.1537031, 0.1114498, 0.1218826, 
    0.1413934, 0.1247572, 0.1436071, 0.1144573, 0.1265144, 0.1015672, 
    0.04582537, 0.08424783, 0.1520818, 0.1302688, 0.1884001,
  0.01793558, 0.04792703, 0.02919008, 0.03289016, 0.0008851046, 
    -5.865792e-06, -4.946281e-05, -6.508708e-05, 0.008953364, 0.0002415318, 
    0.03192912, 0.03189416, 0.04352977, 0.04898271, 0.08649088, 0.06668667, 
    0.07515891, 0.0935782, 0.1415527, 0.0208316, -0.0002354332, 0.0006155267, 
    0.004098723, 0.0002414039, 0.03811695, 0.0470182, 0.04444235, 0.02941484, 
    0.04380623,
  -4.830252e-07, 0.03691711, 0.02010229, 9.10711e-06, 2.157142e-05, 
    0.005188209, -2.720657e-08, 0.0001108258, 0.01242069, 3.574186e-07, 
    0.005900317, 3.054489e-05, -0.0001812375, 0.02662997, 0.02166866, 
    0.1032948, 0.01319754, 0.03576724, 8.714909e-05, -1.424688e-10, 
    -6.777505e-10, 0, 1.377164e-10, 0.01330158, 0.01466887, 0.003725583, 
    -1.724604e-05, -2.040926e-05, 3.713688e-08,
  1.330441e-06, 0.0006754529, 0.0009477608, 0.0006729201, 0.006394929, 
    0.003052183, 0.09360848, 0.01234487, 3.75694e-05, 0.002777694, 
    0.05223954, 0.07768493, 0.1329925, 0.08779202, 0.03952368, 0.02700802, 
    0.01171693, 4.194121e-06, 3.52118e-10, 1.120445e-07, 8.330478e-08, 
    3.356777e-08, 1.71587e-06, 0.01753247, 0.003203207, -2.742699e-07, 
    -4.31876e-10, 1.122336e-07, 3.302363e-07,
  0.0003174907, 0.2513346, 0.1383806, 0.001154175, 0.007295889, 0.1034207, 
    0.01836438, 0.08381839, 0.03658431, 0.1805496, 0.01191165, 0.02181282, 
    0.03428904, 0.01364423, 0.008038126, 0.000503098, 1.561853e-05, 
    -0.0003064925, -1.078022e-06, -3.112895e-05, 7.678367e-06, -6.525339e-05, 
    0.01580887, 0.04814012, 0.005084975, 0.001487688, 0.0016769, 0.005256912, 
    0.03888046,
  0.1005951, 0.1005655, 0.1218909, 0.04075311, 0.004376489, 0.002897571, 
    0.01745322, 0.01025014, 0.09538253, 0.05708433, 0.01273706, 0.0593701, 
    0.05042892, 0.06977348, 0.03263135, 0.1030732, 0.04433431, 0.04516818, 
    0.0956927, 0.1802861, 0.1771272, 0.1613935, 0.09825209, 0.02949361, 
    0.01607687, 0.03121625, 0.07290057, 0.1406193, 0.09150643,
  0.003729269, 0.0002308855, 0.003068517, 0.01363256, 0.0004988319, 
    0.04694985, 0.1063353, 0.09304176, 0.09689599, 0.08248716, 0.0718597, 
    0.1085806, 0.07870124, 0.0150065, 0.0193304, 0.006733042, 6.101913e-07, 
    2.871147e-07, 4.358707e-08, 0.03009192, 0.05560162, 0.1268734, 
    0.02061102, 0.02621885, 0.02541338, 0.02252324, 0.02552795, 0.007238248, 
    0.004218307,
  0.03062582, 1.722043e-05, -2.783605e-09, 0.001284903, 4.96315e-05, 
    2.432253e-06, 0.005995242, 0.1181146, 0.2267113, 0.1589625, 0.02700239, 
    0.04330088, 0.004188082, 0.01050161, 0.0634658, 0.008221178, 0.003869148, 
    -7.066561e-06, -2.244092e-06, 8.258058e-08, 0.02928428, 0.03474536, 
    0.04844175, 0.05584081, 0.04180484, 0.01313347, 0.001233781, 
    0.0001432211, 0.0009548774,
  0.03998243, 0.1100192, 0.002691538, 0.0008663221, 0.04058241, 0.01111101, 
    0.08471932, 0.0495788, 0.08728843, 0.07114577, 0.09238925, 0.2386966, 
    0.132826, 0.1072139, 0.08013383, 0.2165751, 0.1518045, 0.02669151, 
    0.02410375, 0.03989143, 0.02252581, 0.0656881, 0.06233599, 0.1089562, 
    0.07076022, 0.05802242, 0.03007933, 0.02545695, 0.04882599,
  0.1023048, 0.1391, 0.07479621, 0.07244176, 0.07262159, 0.111842, 
    0.05344884, 0.1415407, 0.1159399, 0.1676368, 0.1698627, 0.1378026, 
    0.1153166, 0.1782855, 0.165566, 0.09479601, 0.2060965, 0.1790558, 
    0.102678, 0.1440648, 0.07519802, 0.08737984, 0.1666157, 0.1727715, 
    0.148815, 0.1782303, 0.1930297, 0.1494105, 0.1127476,
  0.2239791, 0.1563893, 0.09056982, 0.2095859, 0.2086965, 0.1286865, 
    0.1608282, 0.1576753, 0.1377044, 0.1465981, 0.132256, 0.1858456, 
    0.2391199, 0.2186011, 0.2679935, 0.1746974, 0.1764776, 0.2571865, 
    0.2111523, 0.1386654, 0.1414496, 0.270297, 0.1826146, 0.1917763, 
    0.2335339, 0.2187484, 0.1848542, 0.1452822, 0.2156494,
  0.1949754, 0.133223, 0.1297504, 0.1558762, 0.2216658, 0.1857842, 0.1554404, 
    0.167868, 0.1024064, 0.1498868, 0.2329322, 0.3127941, 0.1924814, 
    0.140002, 0.1734704, 0.1866025, 0.1869798, 0.1544901, 0.1352877, 
    0.163027, 0.2231558, 0.1289799, 0.1644356, 0.34744, 0.2956541, 0.1928753, 
    0.1282203, 0.2129216, 0.1765098,
  0.2379533, 0.2483655, 0.1589699, 0.1825073, 0.1728231, 0.1904887, 
    0.2297182, 0.2143516, 0.2158141, 0.276591, 0.2400675, 0.2019466, 
    0.2110179, 0.2133274, 0.2129011, 0.2410421, 0.2209241, 0.251885, 
    0.2843365, 0.2934458, 0.2172515, 0.1916183, 0.1914969, 0.1372048, 
    0.1430651, 0.06938305, 0.1322705, 0.09834686, 0.2164108,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  -0.0001932691, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.607209e-06, 0.03113188, 
    0.01762464, 0.08388175, 0.141597, 0.07682228, 0.01270827, -0.0001839001, 
    0.0004596472, 0.001663108, 0.03737138, 0.1768541, 0.247742, 0.1984508, 
    0.2015998, 0.052665, 0.001845623,
  0.09259649, 0.07750648, 0.09437451, 0.1031508, 0.0004808668, -0.0005078397, 
    0.05288551, -0.001423931, -0.00104734, -0.0006396698, -0.0004727656, 
    -0.000623994, 0.09779768, 0.2693312, 0.2763922, 0.2688053, 0.2300174, 
    0.2193038, 0.2253796, 0.1932921, 0.2137737, 0.2816904, 0.2377364, 
    0.3223028, 0.339445, 0.2354551, 0.2839001, 0.2361687, 0.1618522,
  0.1930191, 0.1977347, 0.187555, 0.1751412, 0.1763943, 0.1931723, 0.2318454, 
    0.2153134, 0.2511412, 0.2272412, 0.317736, 0.3080942, 0.2967879, 
    0.3560344, 0.2481331, 0.2271405, 0.1833601, 0.2176362, 0.1645149, 
    0.1758105, 0.1632928, 0.1930552, 0.1929481, 0.218225, 0.1709972, 
    0.1719209, 0.1917537, 0.2088901, 0.1962691,
  0.1746222, 0.2211088, 0.2219157, 0.2197501, 0.156168, 0.2345378, 0.2087121, 
    0.2132953, 0.182073, 0.1861496, 0.223146, 0.1582191, 0.161651, 0.1262537, 
    0.1734519, 0.1461145, 0.1633285, 0.1868772, 0.1473005, 0.2112639, 
    0.206196, 0.2003909, 0.1883136, 0.1724888, 0.1623419, 0.1430843, 
    0.145727, 0.1986113, 0.1856014,
  0.1378476, 0.05170231, 0.08410297, 0.1512189, 0.09719548, 0.1005751, 
    0.08014077, 0.08152366, 0.06830805, 0.04947658, 0.03419271, 0.0993292, 
    0.0716927, 0.1552039, 0.1643809, 0.1375174, 0.1113345, 0.1144111, 
    0.1389788, 0.1178819, 0.1334309, 0.1016576, 0.1331214, 0.1124343, 
    0.04116326, 0.08221264, 0.1492217, 0.1220143, 0.1943901,
  0.02013496, 0.1009307, 0.0414133, 0.04291018, 3.784071e-05, 0.0001070338, 
    6.856145e-05, -1.526577e-05, 0.01158871, -0.0003634549, 0.05195168, 
    0.03226193, 0.0533781, 0.05023335, 0.08945871, 0.06403553, 0.07812408, 
    0.07757796, 0.1378689, 0.02406768, 0.00010025, 0.005192944, 0.007058829, 
    0.002135807, 0.04097206, 0.07938095, 0.05302084, 0.03471953, 0.0437543,
  -1.962654e-05, 0.04783062, 0.0184736, -6.545627e-05, 0.0002734833, 
    4.118824e-05, -9.607867e-08, 0.0003491523, 0.007826331, -1.346633e-07, 
    0.01382995, 0.001452204, -8.217611e-06, 0.02588792, 0.0146217, 
    0.09231886, 0.007007827, 0.03806167, 7.309017e-05, 1.746474e-09, 
    6.46445e-11, 7.456213e-09, 6.483166e-09, 0.006166946, 0.01753151, 
    0.004489328, -8.986884e-05, 9.372315e-05, 7.791277e-08,
  9.078274e-07, 0.00160449, 0.002219474, 0.0009719539, 0.008696624, 
    0.004040352, 0.107321, 0.02454207, 0.004851763, 0.004321068, 0.04381393, 
    0.0712898, 0.1494938, 0.0759723, 0.03786209, 0.02984167, 0.01112206, 
    1.48132e-05, 7.041304e-09, 2.759027e-07, 4.486814e-07, 1.046669e-07, 
    -1.447824e-05, 0.01089482, 0.003375409, -7.022207e-07, 1.596261e-08, 
    1.134341e-08, 4.453002e-08,
  0.0002849716, 0.2200037, 0.1666166, 0.002920405, 0.008086806, 0.08736902, 
    0.02127283, 0.08405735, 0.04773394, 0.1908281, 0.01101745, 0.02410137, 
    0.03694985, 0.01474921, 0.009109497, 0.0005753965, -1.3388e-05, 
    0.003082759, -0.0002136692, 1.705191e-05, 3.423358e-05, 0.0005347374, 
    0.01074102, 0.0500611, 0.0179992, 0.01277042, 0.007785153, 0.02031202, 
    0.02711342,
  0.1208975, 0.09730022, 0.1191958, 0.05407107, 0.02071298, 0.003399121, 
    0.01831294, 0.009395031, 0.1035511, 0.07302144, 0.01274965, 0.05361117, 
    0.05908697, 0.07814791, 0.03054637, 0.08549255, 0.06737006, 0.07881843, 
    0.1313889, 0.2023316, 0.198252, 0.1420839, 0.1061829, 0.02828209, 
    0.01122656, 0.03673425, 0.08659489, 0.1442758, 0.1110422,
  0.002181719, 0.000224626, 0.004435877, 0.009839566, 0.0002953552, 
    0.05170481, 0.118438, 0.1142072, 0.1039942, 0.07794152, 0.09193464, 
    0.1184709, 0.08658778, 0.01308269, 0.01763835, 0.007477636, 2.220038e-06, 
    4.519527e-07, 5.761556e-07, 0.02870192, 0.05885012, 0.1367936, 
    0.01934159, 0.02871395, 0.02806741, 0.02406729, 0.02481805, 0.007176918, 
    0.003896694,
  0.02702767, 6.764376e-06, -3.242753e-08, 0.003557777, 2.172487e-06, 
    2.744e-06, 0.004131822, 0.1188511, 0.2435891, 0.1618287, 0.03194169, 
    0.05984448, 0.005215028, 0.01350324, 0.06807743, 0.01044676, 0.004640475, 
    -1.601187e-05, -8.390748e-08, 1.429262e-08, 0.02532898, 0.03367953, 
    0.03999564, 0.05630493, 0.03885495, 0.0120133, 0.000992434, 6.489763e-05, 
    0.01821781,
  0.02640937, 0.1120441, 0.004399098, 0.001038743, 0.04926569, 0.006753348, 
    0.108392, 0.02994329, 0.05780808, 0.06042744, 0.07757303, 0.2067023, 
    0.1024358, 0.09167799, 0.07094035, 0.2067282, 0.1514156, 0.02426797, 
    0.02297391, 0.03907971, 0.01985278, 0.06666534, 0.06614818, 0.09954008, 
    0.06224094, 0.04666291, 0.02329734, 0.02313086, 0.05007917,
  0.1072767, 0.1236246, 0.05806587, 0.07808358, 0.0712045, 0.1203739, 
    0.0479792, 0.1369155, 0.1089022, 0.1600045, 0.1730326, 0.1360983, 
    0.1269942, 0.1636493, 0.1576793, 0.100322, 0.1720062, 0.1636922, 
    0.09940491, 0.1293686, 0.0789728, 0.06456359, 0.1811534, 0.2091782, 
    0.1507567, 0.1671469, 0.1733677, 0.1504885, 0.1211578,
  0.1988799, 0.1753696, 0.103024, 0.2011641, 0.202806, 0.125425, 0.1667423, 
    0.1531177, 0.1305815, 0.1427492, 0.1088614, 0.1797095, 0.2449315, 
    0.2110521, 0.2424981, 0.1563375, 0.1643898, 0.2582018, 0.2080684, 
    0.1457265, 0.1418004, 0.2557264, 0.1579117, 0.1904726, 0.2332184, 
    0.2495152, 0.1814504, 0.1452748, 0.2164755,
  0.2100366, 0.1210607, 0.134673, 0.1788705, 0.2056508, 0.1788835, 0.1449765, 
    0.1559133, 0.1017494, 0.1244242, 0.2194381, 0.3240569, 0.1929936, 
    0.1230741, 0.1788354, 0.1997275, 0.1847311, 0.159743, 0.1332646, 
    0.1622547, 0.2343638, 0.1367847, 0.159145, 0.3712396, 0.2921071, 
    0.2608474, 0.2199782, 0.1930858, 0.1680984,
  0.2347307, 0.2946844, 0.1584135, 0.166253, 0.1663224, 0.1843624, 0.2485068, 
    0.2243792, 0.2175722, 0.2629529, 0.2379997, 0.2114309, 0.2014056, 
    0.2044181, 0.2102268, 0.2464422, 0.2257733, 0.2513877, 0.2654928, 
    0.2833364, 0.2247903, 0.1905356, 0.1993301, 0.1477959, 0.1476597, 
    0.07139699, 0.1492638, 0.10562, 0.2147295,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0.005609978, -0.0002503169, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0001601886, 
    0.04981837, 0.1252723, 0.1786596, 0.2564222, 0.2240963, 0.06970733, 
    0.005141483, 0.002679867, 0.008471049, 0.08394138, 0.4066095, 0.3409633, 
    0.2910407, 0.2827602, 0.1653398, 0.02004628,
  0.09210042, 0.1137624, 0.1578389, 0.1976864, 0.009129276, 0.0167356, 
    0.1089693, -0.002444005, 0.006371729, -0.001019434, 0.008491925, 
    0.02643275, 0.1930095, 0.3278041, 0.3206082, 0.282805, 0.2313943, 
    0.2449362, 0.2408957, 0.2115295, 0.2159115, 0.2842766, 0.2917811, 
    0.3777226, 0.3589024, 0.2601565, 0.2800458, 0.2066398, 0.1702221,
  0.2170846, 0.2166208, 0.2075956, 0.1994408, 0.227399, 0.2730325, 0.2581166, 
    0.2318114, 0.2824144, 0.2617541, 0.3387246, 0.3218257, 0.2847776, 
    0.3378609, 0.2289626, 0.2155595, 0.1801178, 0.2195603, 0.1899001, 
    0.1749854, 0.1677236, 0.1832977, 0.2149843, 0.2095333, 0.1639281, 
    0.1469427, 0.1711556, 0.2068303, 0.2023566,
  0.1804987, 0.2187161, 0.2342312, 0.2193685, 0.1462757, 0.2385216, 
    0.2325028, 0.2135312, 0.1903518, 0.174884, 0.2129265, 0.1535285, 
    0.1431518, 0.1241271, 0.1695988, 0.1569417, 0.1467415, 0.1998345, 
    0.1640092, 0.2361966, 0.1952315, 0.1966462, 0.1811646, 0.1452677, 
    0.1587827, 0.1388708, 0.1460987, 0.182533, 0.1911448,
  0.1228434, 0.05343987, 0.08126599, 0.1372669, 0.09028103, 0.0963304, 
    0.09484945, 0.0832248, 0.08105981, 0.03834118, 0.03755886, 0.09521898, 
    0.06515391, 0.150901, 0.1642954, 0.146042, 0.1078638, 0.1009009, 
    0.1404358, 0.1134275, 0.1517928, 0.09897759, 0.134258, 0.1144176, 
    0.04255579, 0.08966551, 0.1418463, 0.1256314, 0.2043877,
  0.006534607, 0.0468374, 0.06868159, 0.04073212, 0.0009579503, 1.060874e-05, 
    7.041089e-06, 0.0002726808, 0.01260361, 0.0008333903, 0.05143288, 
    0.03556148, 0.05927424, 0.04821818, 0.08727936, 0.06091414, 0.09573873, 
    0.06193547, 0.1104062, 0.01794767, 0.001196548, 0.007314016, 0.006450934, 
    0.003858604, 0.0591227, 0.09147376, 0.05873913, 0.04777599, 0.03637968,
  0.006656339, 0.0616261, 0.03928814, -0.00014923, 0.002240115, 2.477715e-06, 
    8.796467e-06, 0.0007986964, 0.01052537, -2.006508e-05, 0.01403028, 
    0.0121221, -3.660653e-05, 0.01863964, 0.01071923, 0.04107021, 
    0.008973435, 0.04449844, 0.0001089748, 1.898485e-08, 2.377683e-09, 
    3.794327e-08, 3.423158e-08, 0.001318991, 0.02804084, 0.02373099, 
    -9.066897e-05, 5.453759e-05, -1.42361e-07,
  0.0001288363, 0.01654625, 0.02537144, 0.002650202, 0.01132067, 0.006234037, 
    0.1057924, 0.04227562, 0.001918483, 0.002641988, 0.04607492, 0.06526045, 
    0.1590268, 0.09168962, 0.05523846, 0.03450132, 0.01623805, 1.598483e-05, 
    1.100631e-07, 1.1239e-06, 2.050097e-06, 4.482609e-07, 0.01742957, 
    0.01396565, 0.005569399, 0.0003237924, 1.255769e-07, 1.978996e-07, 
    -2.225195e-06,
  0.0006298737, 0.221525, 0.2178126, 0.006885036, 0.007463691, 0.06789599, 
    0.0263669, 0.09445174, 0.0676873, 0.205368, 0.01718107, 0.02559888, 
    0.04519869, 0.01673674, 0.009618374, 0.0007956653, 0.000446771, 
    4.345518e-05, 0.005620541, 0.003061236, 7.259684e-05, 0.001839211, 
    0.01929688, 0.08208774, 0.01942895, 0.02461117, 0.02164051, 0.04316683, 
    0.05527189,
  0.1515358, 0.1182297, 0.1356333, 0.06458159, 0.03354166, 0.003226812, 
    0.02284254, 0.02246764, 0.1323779, 0.09275302, 0.02459943, 0.06085445, 
    0.08428358, 0.1125298, 0.03888997, 0.0939028, 0.08298805, 0.1030953, 
    0.1704253, 0.2295479, 0.2261347, 0.1437421, 0.1302885, 0.03954776, 
    0.01189063, 0.06753908, 0.1080785, 0.1515259, 0.1627026,
  0.01109866, 0.002077583, 0.006900019, 0.00701909, 6.668313e-06, 0.04161285, 
    0.1606648, 0.1434783, 0.1295919, 0.08556122, 0.1088542, 0.1465246, 
    0.1028268, 0.01810633, 0.01816714, 0.009086588, 0.0001382376, 
    -9.571846e-07, 8.860276e-05, 0.03559075, 0.07903792, 0.1487283, 
    0.02382856, 0.0497689, 0.03777384, 0.03314404, 0.03407455, 0.006755273, 
    0.01354236,
  0.0171252, 3.602702e-05, -1.074306e-08, 0.0009761574, -1.633096e-05, 
    -2.691949e-06, 0.007100471, 0.1168979, 0.2886184, 0.1545499, 0.03844196, 
    0.07868493, 0.01247696, 0.01668562, 0.07435846, 0.0143983, 0.008464086, 
    0.0004290248, 7.118577e-08, -6.386323e-06, 0.02956602, 0.03860595, 
    0.04215898, 0.06505472, 0.03877791, 0.01588079, 0.001851321, 
    4.571573e-05, 0.02057158,
  0.02037349, 0.1083285, 0.004370081, 0.001711305, 0.02804222, 0.0033179, 
    0.128195, 0.01943132, 0.03173742, 0.05292117, 0.07372504, 0.1879258, 
    0.08852434, 0.09931348, 0.07910249, 0.2022309, 0.1564105, 0.01879694, 
    0.02419587, 0.04163012, 0.02160712, 0.07946788, 0.06548449, 0.09311651, 
    0.06145899, 0.04242829, 0.02370125, 0.0236642, 0.05114909,
  0.1220128, 0.1300929, 0.06690317, 0.09846871, 0.05861011, 0.1171858, 
    0.04875804, 0.1445031, 0.1012068, 0.1549959, 0.1819608, 0.1344486, 
    0.1505746, 0.1506096, 0.1480244, 0.1010357, 0.1585155, 0.153744, 
    0.1024511, 0.1255051, 0.0917279, 0.05461068, 0.1670204, 0.2186961, 
    0.1677682, 0.1656637, 0.1628014, 0.1605188, 0.1124214,
  0.1822769, 0.1672217, 0.1256933, 0.2049564, 0.2027016, 0.1326703, 
    0.1821418, 0.1695487, 0.12595, 0.1459519, 0.1069246, 0.1747878, 
    0.2422337, 0.2482966, 0.2240897, 0.1628431, 0.1924592, 0.2712919, 
    0.2113993, 0.1494499, 0.1546697, 0.2410163, 0.1363731, 0.2108593, 
    0.2514739, 0.2505441, 0.182708, 0.1592898, 0.2316697,
  0.1928056, 0.1687786, 0.2125898, 0.2031268, 0.2188856, 0.1851666, 
    0.1599227, 0.163868, 0.1158917, 0.102563, 0.2241328, 0.3363956, 
    0.2116344, 0.104506, 0.1849539, 0.2033423, 0.1813703, 0.1364873, 
    0.153122, 0.2029937, 0.2768741, 0.1552159, 0.1674314, 0.4028688, 
    0.3171192, 0.2508635, 0.2520431, 0.1706029, 0.1592673,
  0.2305821, 0.2758291, 0.1441715, 0.1357474, 0.1581227, 0.1721994, 
    0.2483583, 0.2557112, 0.2230004, 0.2650136, 0.2188571, 0.2475672, 
    0.2148829, 0.2025687, 0.1936351, 0.2636327, 0.2283809, 0.2769536, 
    0.3016342, 0.3036765, 0.2371347, 0.1971571, 0.1965032, 0.1526608, 
    0.1584077, 0.07557491, 0.1765553, 0.1162792, 0.1931869,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0.0198053, -0.0006658328, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0007743601, 
    0.1040212, 0.1785383, 0.2098343, 0.3303642, 0.3803357, 0.2083119, 
    0.0468756, 0.01569324, 0.01443031, 0.1411374, 0.4277402, 0.3264049, 
    0.295381, 0.3255879, 0.2127011, 0.05479253,
  0.1068183, 0.1488088, 0.1822903, 0.2738638, 0.03005056, 0.07342856, 
    0.1168554, 0.0138848, 0.02101504, 0.01523235, 0.04815968, 0.09314139, 
    0.2606888, 0.3127004, 0.3336199, 0.2824786, 0.2341878, 0.2483574, 
    0.2603002, 0.2222094, 0.1962748, 0.2764073, 0.2921081, 0.3787252, 
    0.3509228, 0.2722236, 0.2700009, 0.190951, 0.1643065,
  0.2229205, 0.2116136, 0.2072465, 0.194821, 0.2148107, 0.2638952, 0.2640925, 
    0.2310546, 0.2919533, 0.2632712, 0.3245529, 0.3297111, 0.2744252, 
    0.3312131, 0.2301931, 0.2100819, 0.1904683, 0.2323835, 0.2019675, 
    0.1905397, 0.1757919, 0.188453, 0.211493, 0.2062858, 0.1559137, 
    0.1374955, 0.1792248, 0.2084432, 0.210417,
  0.192369, 0.2183493, 0.232483, 0.2177239, 0.148304, 0.2514353, 0.2293643, 
    0.2170507, 0.1907243, 0.1808549, 0.2088542, 0.1568134, 0.1507953, 
    0.1249175, 0.1596463, 0.1706552, 0.1377454, 0.2061643, 0.1451873, 
    0.2295306, 0.1652521, 0.1836164, 0.1911477, 0.1488516, 0.1733943, 
    0.119064, 0.1490582, 0.1848415, 0.1830282,
  0.1399421, 0.07096621, 0.08048107, 0.1180983, 0.1203548, 0.09262341, 
    0.100307, 0.09441002, 0.100122, 0.06828782, 0.0363762, 0.09050176, 
    0.06046362, 0.1423695, 0.1638054, 0.1381872, 0.1007195, 0.09067483, 
    0.1395643, 0.1127241, 0.1476191, 0.1062425, 0.1391525, 0.1180936, 
    0.04019274, 0.09688655, 0.1247154, 0.1256209, 0.2091729,
  0.009616911, 0.01882699, 0.08267803, 0.04568318, 0.0005344151, 
    3.394521e-07, 1.122515e-06, 0.0008090514, 0.01300582, 0.004162418, 
    0.02381644, 0.013883, 0.04160329, 0.04962125, 0.08139982, 0.05765456, 
    0.08719029, 0.05647578, 0.1000764, 0.01938028, 0.009530242, 0.0139554, 
    0.008106885, 0.0003874357, 0.086454, 0.08756006, 0.06716388, 0.04364276, 
    0.02642873,
  0.0005708264, 0.04577995, 0.05734449, 0.01015565, 0.003182638, 
    2.444527e-05, 0.0004929531, 0.001695793, 0.007518121, 0.00175392, 
    0.01444817, 0.0001970505, -0.0001564793, 0.01763507, 0.01631801, 
    0.0153338, 0.01098655, 0.044047, 0.0003946405, 6.454054e-08, 
    -1.604766e-07, 8.983277e-08, 9.083254e-08, 0.0006241476, 0.06899171, 
    0.05579908, -0.0001640034, 8.871199e-06, -7.092105e-05,
  0.004854818, 0.02647231, 0.06686329, 0.00108336, 0.01450124, 0.008072554, 
    0.1073266, 0.05388772, 0.002040065, 0.004885528, 0.05252334, 0.07668103, 
    0.1726636, 0.1161445, 0.07736105, 0.03655286, 0.01603367, 0.000249073, 
    2.972465e-07, 7.871907e-07, 1.422527e-06, 1.179973e-06, 0.02410002, 
    0.02089161, 0.04859502, 0.005098551, -1.101707e-05, -2.666679e-07, 
    4.92027e-06,
  0.004964636, 0.2543111, 0.2706682, 0.009656488, 0.005600689, 0.06013967, 
    0.03947891, 0.1085827, 0.09743052, 0.2463737, 0.02021273, 0.03609181, 
    0.06131574, 0.01461553, 0.007459326, 0.0007634062, 0.0009539856, 
    0.001888323, 0.0005600011, 0.001949371, 0.0004560341, 0.008243219, 
    0.03944908, 0.1319383, 0.01733719, 0.0125784, 0.02138488, 0.04843388, 
    0.05841389,
  0.1830695, 0.1362131, 0.1745832, 0.1095398, 0.02929453, 0.005103341, 
    0.02495961, 0.03428485, 0.1674272, 0.09209697, 0.03446813, 0.07000169, 
    0.09463526, 0.1211689, 0.04840351, 0.09672961, 0.08995557, 0.132818, 
    0.2034576, 0.2728717, 0.2777713, 0.1570219, 0.1663622, 0.05761937, 
    0.01305133, 0.08360817, 0.121817, 0.1855712, 0.2228939,
  0.04004848, 0.0127613, 0.02700875, 0.0007197079, -9.809402e-07, 0.02429882, 
    0.2347358, 0.1417779, 0.1901174, 0.09229968, 0.107395, 0.1554641, 
    0.09998979, 0.02546833, 0.02222241, 0.01138856, 0.000311312, 1.53603e-07, 
    0.002256461, 0.04990512, 0.09430963, 0.1730669, 0.02544756, 0.06612587, 
    0.03990293, 0.03981962, 0.03738961, 0.00957258, 0.006715202,
  0.004680577, 0.0001237082, 1.477296e-07, 0.0002462621, -1.422022e-05, 
    1.256537e-07, 0.0169179, 0.1173361, 0.317759, 0.1431042, 0.05410228, 
    0.08859444, 0.01783664, 0.01717939, 0.08440869, 0.02023252, 0.01505621, 
    0.002286287, 4.366229e-08, 3.194898e-05, 0.03538831, 0.04728505, 
    0.04668676, 0.07686731, 0.03712206, 0.02275962, 0.004026697, 
    0.0001012034, 0.002658512,
  0.02001166, 0.0817812, 0.002664643, 0.004436571, 0.02493682, 0.0009688904, 
    0.1437806, 0.0296304, 0.01885612, 0.05114074, 0.06235447, 0.1774117, 
    0.08546495, 0.1150233, 0.08598018, 0.2218471, 0.1444413, 0.01720421, 
    0.02309696, 0.04733129, 0.03401071, 0.1030251, 0.06365149, 0.09471183, 
    0.07765584, 0.04875837, 0.02932577, 0.02525837, 0.05113405,
  0.111752, 0.1313239, 0.05108858, 0.104576, 0.06140718, 0.1161534, 
    0.06247177, 0.1542922, 0.09202699, 0.1468796, 0.1862999, 0.1423693, 
    0.1417351, 0.1449462, 0.154506, 0.1010462, 0.1820743, 0.1645333, 
    0.1196564, 0.123349, 0.09140956, 0.04916963, 0.1861384, 0.2531313, 
    0.1761451, 0.1730437, 0.1682985, 0.1572075, 0.129981,
  0.167502, 0.1643115, 0.1445998, 0.2304738, 0.2036979, 0.1640193, 0.1915648, 
    0.197355, 0.1642046, 0.1514023, 0.1226395, 0.1714758, 0.2519739, 
    0.2038397, 0.2346458, 0.1962722, 0.1756232, 0.269553, 0.2032088, 
    0.1612765, 0.151247, 0.2423153, 0.1139548, 0.2166965, 0.2519546, 
    0.2569594, 0.1854103, 0.1682901, 0.2257616,
  0.2266965, 0.1392037, 0.1748659, 0.2092038, 0.2226083, 0.1909127, 
    0.1436713, 0.1990921, 0.1204364, 0.1147183, 0.2617364, 0.3470425, 
    0.2304156, 0.07814389, 0.2106727, 0.2605719, 0.179454, 0.1434396, 
    0.1733893, 0.2259771, 0.2790221, 0.1537107, 0.2038822, 0.4333624, 
    0.3315025, 0.274539, 0.2459888, 0.1428994, 0.1685406,
  0.2430798, 0.3037958, 0.1520932, 0.127903, 0.1707864, 0.1963449, 0.2210908, 
    0.193981, 0.1874723, 0.2249796, 0.1898467, 0.2381294, 0.2333036, 
    0.2144899, 0.1969815, 0.2446576, 0.2377111, 0.3363011, 0.3157205, 
    0.3523034, 0.245949, 0.2263789, 0.2080346, 0.1818749, 0.1539356, 
    0.09474195, 0.2006361, 0.1098094, 0.1892828,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0.04101567, 0.007911535, -3.335803e-05, 0, 0, 0, 0, 0, 0, 0, 0, 
    -6.895672e-05, 0.004097829, 0.1085807, 0.1615594, 0.1952975, 0.3251413, 
    0.4762108, 0.2975515, 0.1554651, 0.04727457, 0.04992796, 0.234644, 
    0.4365792, 0.3223517, 0.2886956, 0.3435734, 0.263093, 0.1016451,
  0.1230837, 0.1575885, 0.208096, 0.2705946, 0.08766499, 0.1132723, 
    0.1203815, 0.03706499, 0.03045635, 0.05915035, 0.1129605, 0.1744511, 
    0.2871938, 0.3132901, 0.3328926, 0.294424, 0.23033, 0.2295714, 0.2585745, 
    0.2236701, 0.2143966, 0.2916622, 0.2986987, 0.3733242, 0.335507, 
    0.2752874, 0.273625, 0.1935488, 0.1937956,
  0.2121679, 0.2129779, 0.2010785, 0.1952406, 0.2101979, 0.2455373, 
    0.2588196, 0.2464787, 0.2914113, 0.2683506, 0.3271485, 0.3205576, 
    0.2716875, 0.3207052, 0.240241, 0.2473964, 0.1974766, 0.2199072, 
    0.1843951, 0.1902572, 0.1608282, 0.1846936, 0.217994, 0.1863065, 
    0.1568887, 0.1356605, 0.1874633, 0.2240495, 0.1941746,
  0.2044773, 0.2139414, 0.2387855, 0.2188399, 0.1555509, 0.249117, 0.2402787, 
    0.2403031, 0.1945298, 0.1936246, 0.2175243, 0.1651445, 0.1442737, 
    0.09928794, 0.1492794, 0.1641124, 0.1505566, 0.2174841, 0.1395405, 
    0.2199795, 0.1628658, 0.1782922, 0.1973056, 0.1540943, 0.1715974, 
    0.1267371, 0.1596746, 0.2215079, 0.2073312,
  0.139585, 0.07392289, 0.08115745, 0.08657075, 0.1287856, 0.1063515, 
    0.1052999, 0.09311929, 0.0944728, 0.05440195, 0.03344529, 0.07701814, 
    0.05453215, 0.1404523, 0.1655707, 0.1349701, 0.0847922, 0.08982084, 
    0.1416249, 0.1314853, 0.1468463, 0.1062664, 0.1372368, 0.1335737, 
    0.03294422, 0.1019714, 0.1284512, 0.1323468, 0.2035547,
  0.01458981, 0.002502626, 0.07872028, 0.0302855, 0.00685708, 5.652753e-08, 
    1.212854e-05, 0.005533041, 0.01614735, 0.01013346, 0.002063518, 
    0.001617026, 0.02956375, 0.05237338, 0.07704412, 0.063682, 0.09318534, 
    0.0848612, 0.09198257, 0.02101332, 0.02353485, 0.02111537, 0.00993125, 
    -8.475806e-05, 0.07124484, 0.08563469, 0.07892016, 0.03988087, 0.03781448,
  1.038764e-05, 0.01713439, 0.05530167, 0.01313023, 0.009774829, 
    0.0004928957, 0.0007948225, 0.01009699, 0.003595087, 0.006211569, 
    0.002525919, -0.0001486079, -4.083072e-06, 0.01824482, 0.02866637, 
    0.007073569, 0.01761018, 0.04305724, 0.0007812986, 8.037656e-07, 
    1.442065e-05, 8.017161e-08, 7.706186e-08, 1.689305e-05, 0.03487622, 
    0.06807052, -5.720342e-05, -7.184422e-06, 0.0002555546,
  0.0003382926, 0.01505688, 0.1373121, 0.01507591, 0.01955128, 0.01085166, 
    0.09359442, 0.04578051, 0.00138424, 0.004256894, 0.06187119, 0.0583774, 
    0.1768923, 0.09631234, 0.08273774, 0.03834963, 0.01957839, 0.00442698, 
    -1.050462e-07, 8.354003e-07, 4.836363e-07, -9.042857e-06, 0.004922189, 
    0.02103985, 0.0635433, 0.008350319, -4.620552e-06, -6.976257e-06, 
    0.0008508106,
  0.00910346, 0.2914233, 0.285762, 0.003997425, 0.003467024, 0.06320641, 
    0.04873548, 0.1040064, 0.108814, 0.269754, 0.02303799, 0.02288364, 
    0.04956454, 0.0104387, 0.005379784, 0.0009667329, 0.006744791, 
    0.006997597, 0.000561744, -1.685566e-05, 0.004740586, 0.01379691, 
    0.06054346, 0.1363685, 0.01955943, 0.003967883, 0.03054524, 0.03587488, 
    0.03438487,
  0.1686145, 0.1553642, 0.1823131, 0.1435502, 0.02590785, 0.005067615, 
    0.0286545, 0.02556222, 0.09705741, 0.08244734, 0.01648935, 0.04993026, 
    0.06244887, 0.07489637, 0.04561517, 0.08432363, 0.08054544, 0.1459433, 
    0.2186412, 0.3009471, 0.2683811, 0.1341311, 0.1663863, 0.05745567, 
    0.01398718, 0.09070452, 0.1050669, 0.1582709, 0.2505098,
  0.01191033, 0.01035499, 0.02111218, -1.633655e-05, -3.579671e-05, 
    0.0009404725, 0.1937349, 0.1161934, 0.1997792, 0.0772867, 0.08305343, 
    0.1142698, 0.07241999, 0.01884869, 0.01945908, 0.01745964, 0.0002875245, 
    1.165718e-07, 0.003414848, 0.07060728, 0.07504462, 0.1736888, 0.0209661, 
    0.05149412, 0.04259695, 0.0369211, 0.01948656, 0.004599015, 0.009388478,
  0.0007367432, 0.00214927, 1.045103e-07, 5.838087e-06, -1.462452e-05, 
    6.492883e-08, 0.01115703, 0.1575795, 0.3476508, 0.1092763, 0.04763659, 
    0.0704161, 0.01315818, 0.01254312, 0.08349103, 0.02948003, 0.02415848, 
    0.007329513, 1.197912e-07, 0.0001123133, 0.04531777, 0.04339929, 
    0.05040973, 0.07968696, 0.02983277, 0.02456338, 0.006196853, 
    0.0005275329, 0.0009128751,
  0.02071145, 0.06107464, 0.002693369, 0.006405677, 0.02386452, 0.002017867, 
    0.1471791, 0.04431803, 0.01623348, 0.05529284, 0.06793459, 0.1668556, 
    0.07503944, 0.1212881, 0.1087514, 0.2490409, 0.1572359, 0.02362735, 
    0.02141407, 0.0420118, 0.03591105, 0.121428, 0.06514873, 0.08791195, 
    0.1044649, 0.057871, 0.02937669, 0.02913377, 0.0524246,
  0.1205106, 0.1348218, 0.05389487, 0.1198074, 0.05070014, 0.1047907, 
    0.09933325, 0.1747996, 0.09012134, 0.1451825, 0.1873453, 0.1617253, 
    0.1391083, 0.1633506, 0.1537447, 0.1141808, 0.1781267, 0.163461, 
    0.1300603, 0.1165252, 0.08379655, 0.04584024, 0.1877652, 0.2439342, 
    0.1860651, 0.1787761, 0.1811151, 0.1829584, 0.135678,
  0.147339, 0.1812294, 0.1445311, 0.2308137, 0.2146551, 0.1708624, 0.1741904, 
    0.2205664, 0.1777963, 0.1612143, 0.136632, 0.1626914, 0.2806723, 
    0.2344005, 0.2585697, 0.1748624, 0.1781844, 0.2870449, 0.2018446, 
    0.153237, 0.1514782, 0.2437257, 0.1252456, 0.2180271, 0.2648697, 
    0.2493094, 0.1847226, 0.1447162, 0.2506408,
  0.2383045, 0.1715236, 0.2069423, 0.2788766, 0.1947863, 0.1688907, 
    0.1700796, 0.195997, 0.1377279, 0.1424008, 0.2860364, 0.3215451, 
    0.2724694, 0.07339759, 0.2833817, 0.2181662, 0.1649227, 0.1626386, 
    0.1641021, 0.2115846, 0.2746212, 0.1645807, 0.2781232, 0.4608624, 
    0.4283363, 0.2780771, 0.2433456, 0.1505504, 0.1705872,
  0.2264269, 0.2786391, 0.1707991, 0.1142585, 0.157577, 0.1340359, 0.1682592, 
    0.208552, 0.1986358, 0.2397067, 0.2250613, 0.2163212, 0.2094604, 
    0.193167, 0.2083898, 0.2773102, 0.2621888, 0.3649536, 0.2913596, 
    0.3135833, 0.2529915, 0.2578996, 0.2460899, 0.2055236, 0.1734423, 
    0.0974906, 0.1991168, 0.1093424, 0.222407,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -0.0006140085, -0.0006140085, -0.0006140085, -0.0006140085, 
    -0.0006140085, -0.0006140085, -0.0006140085, 0,
  0.0587402, 0.02080031, 0.007980447, -7.705275e-05, 0, 0, 0, 0, 0, 0, 0, 
    -3.355611e-05, 0.005867464, 0.09526716, 0.1453089, 0.1858137, 0.3213037, 
    0.4907294, 0.3595784, 0.2419223, 0.1354974, 0.1387511, 0.3256739, 
    0.4574776, 0.329329, 0.2834647, 0.3595687, 0.2928575, 0.1387347,
  0.1250119, 0.161029, 0.2300327, 0.2706223, 0.1641059, 0.1322392, 0.119005, 
    0.08338922, 0.04063734, 0.1522038, 0.1562215, 0.2493568, 0.2854571, 
    0.3261677, 0.3389609, 0.3204831, 0.2478416, 0.2252771, 0.2537132, 
    0.2421527, 0.2257674, 0.3071064, 0.3168046, 0.3806976, 0.3340107, 
    0.2695908, 0.2757413, 0.2087835, 0.2057953,
  0.233788, 0.2027328, 0.194837, 0.2069649, 0.2226895, 0.2315557, 0.2649736, 
    0.2492239, 0.2913394, 0.3028927, 0.3322695, 0.3318517, 0.2856741, 
    0.3024654, 0.24117, 0.2419432, 0.2095994, 0.2215709, 0.1939352, 
    0.1877173, 0.1744502, 0.1992458, 0.2473806, 0.1767224, 0.1686895, 
    0.1592581, 0.20771, 0.2362508, 0.1906633,
  0.2088311, 0.1866422, 0.2193136, 0.2075711, 0.1746519, 0.2645933, 
    0.2626338, 0.2490129, 0.2093461, 0.2121809, 0.2192804, 0.1703931, 
    0.1329725, 0.1045904, 0.1481384, 0.1759513, 0.1845663, 0.2205437, 
    0.1598907, 0.2045065, 0.1601121, 0.179582, 0.2042268, 0.1704859, 
    0.1640922, 0.1406925, 0.1680297, 0.1811844, 0.1883042,
  0.1471079, 0.0906788, 0.09438726, 0.07941726, 0.1333566, 0.1166163, 
    0.1163383, 0.1056961, 0.09732816, 0.0658685, 0.02786607, 0.07260723, 
    0.04616156, 0.1494806, 0.1656211, 0.1309196, 0.08801226, 0.08697423, 
    0.1487397, 0.1188051, 0.1215161, 0.1065009, 0.1421608, 0.1553621, 
    0.03253783, 0.1004148, 0.1391725, 0.1425186, 0.2165176,
  0.02059992, 0.0002937597, 0.05335486, 0.01205266, 0.01611389, 1.75691e-05, 
    0.0008938058, 0.02756331, 0.02096695, 0.01422537, 3.375125e-05, 
    0.0002471028, 0.0267277, 0.05869583, 0.07348815, 0.06887992, 0.09833577, 
    0.07982365, 0.08630622, 0.02726363, 0.04117725, 0.03370073, 0.01174904, 
    9.168602e-05, 0.04776629, 0.07340699, 0.08831944, 0.04407282, 0.03962584,
  6.201553e-07, 0.001770974, 0.03544472, 0.0007882372, 0.02098805, 
    0.001518697, 0.0004505165, 0.003742649, 0.0006540635, 0.006072858, 
    2.2021e-05, 0.0002850228, 1.920725e-05, 0.04886241, 0.04549134, 
    0.01085527, 0.02989551, 0.05332256, 0.004817892, 5.775084e-05, 
    0.001079326, 2.199223e-08, 6.178509e-08, 6.749018e-06, 0.02112919, 
    0.04727641, 1.335716e-06, 4.147607e-05, 0.0005623655,
  4.392823e-06, 0.001635565, 0.09649104, 0.05028196, 0.02714824, 0.01113314, 
    0.07482478, 0.03563841, 0.003881497, 0.002074166, 0.06390597, 0.04431351, 
    0.1842551, 0.09501173, 0.08800332, 0.03804506, 0.02656498, 0.007935842, 
    0.0003842163, 2.912694e-06, 3.489191e-07, -3.101673e-07, 0.001703017, 
    0.01346757, 0.04771278, 0.001368703, 0.0001157184, 1.995417e-06, 
    5.549533e-05,
  0.005356304, 0.2373178, 0.2036132, 0.003529427, 0.002686925, 0.05526966, 
    0.0413773, 0.07790115, 0.08931752, 0.2298435, 0.02510829, 0.01828358, 
    0.03891955, 0.01131898, 0.007299302, 0.001231783, 0.0009966389, 
    0.005171416, 3.143218e-05, 9.576007e-05, 0.0007463417, 0.01210642, 
    0.07668377, 0.09160546, 0.07853904, 0.003274364, 0.005647433, 0.0273049, 
    0.01641609,
  0.1271519, 0.1161774, 0.1080406, 0.1972757, 0.03712158, 0.004648292, 
    0.04459264, 0.02577988, 0.06498706, 0.06633369, 0.01231833, 0.03959771, 
    0.0478189, 0.05054324, 0.0436487, 0.06805002, 0.07949179, 0.1524276, 
    0.2327691, 0.3180936, 0.27323, 0.1211107, 0.1466348, 0.04557937, 
    0.01378145, 0.08751552, 0.1024923, 0.1088808, 0.2048694,
  0.0009200315, 0.001747131, 0.02424657, -2.544995e-05, -1.329953e-06, 
    -0.0002536196, 0.1566571, 0.1046375, 0.1878494, 0.07692289, 0.07093669, 
    0.08941232, 0.06138205, 0.01592313, 0.01822375, 0.02784718, 0.001423745, 
    -2.746036e-08, 0.002120746, 0.06492194, 0.06327822, 0.1777301, 0.0205148, 
    0.04129808, 0.04212731, 0.03148492, 0.003435131, 0.0003009237, 0.00230006,
  5.872541e-05, 0.003220856, 3.41461e-08, 1.059661e-06, -3.150444e-07, 
    2.954863e-08, 0.009820134, 0.2179612, 0.4026799, 0.09966561, 0.03670778, 
    0.07270924, 0.01007439, 0.009339614, 0.06828667, 0.03144483, 0.03088142, 
    0.01244919, 3.077778e-07, 0.0001254204, 0.06570998, 0.04526663, 
    0.04504803, 0.06942736, 0.02211153, 0.02844206, 0.006550278, 
    0.0009295942, 0.0005072132,
  0.02959085, 0.0511785, 0.002432102, 0.01603389, 0.01783785, 0.001587529, 
    0.1373374, 0.02724391, 0.01400833, 0.07301768, 0.06977794, 0.1605223, 
    0.076153, 0.1261173, 0.1073076, 0.2677661, 0.1576725, 0.04401994, 
    0.01314064, 0.03154784, 0.0517364, 0.1347059, 0.06718103, 0.07130253, 
    0.1027381, 0.06645016, 0.03372869, 0.03609851, 0.05045394,
  0.1214534, 0.1474862, 0.06087271, 0.1240616, 0.07255767, 0.1022632, 
    0.1206831, 0.1871363, 0.09561338, 0.1480598, 0.1744221, 0.1623239, 
    0.1415219, 0.167985, 0.1395796, 0.1054077, 0.1633472, 0.1664141, 
    0.1292879, 0.1183729, 0.1012, 0.04757468, 0.2226062, 0.2442973, 
    0.1799092, 0.1678949, 0.1987845, 0.2025128, 0.1439489,
  0.1494687, 0.1848138, 0.1295155, 0.2242147, 0.2634709, 0.1681761, 
    0.1573041, 0.2324756, 0.1785985, 0.2075286, 0.140331, 0.1626662, 
    0.3143168, 0.2306866, 0.2519771, 0.1762549, 0.1790208, 0.3073692, 
    0.1909579, 0.1407466, 0.1295628, 0.247363, 0.1146404, 0.1947466, 
    0.2970098, 0.2544243, 0.2015109, 0.1767268, 0.2492499,
  0.2604291, 0.1413232, 0.2584516, 0.2664461, 0.2261519, 0.1982167, 0.168117, 
    0.1531867, 0.1282557, 0.1684431, 0.3135808, 0.3340585, 0.2354162, 
    0.08961886, 0.3058482, 0.2298748, 0.1234095, 0.1563711, 0.1719134, 
    0.2604659, 0.2667056, 0.1374137, 0.3190317, 0.4536086, 0.396341, 
    0.290571, 0.2503838, 0.1399593, 0.151591,
  0.2415016, 0.2827227, 0.2356288, 0.1182184, 0.1265038, 0.176968, 0.2045761, 
    0.1930165, 0.1665271, 0.2709765, 0.2706094, 0.2534204, 0.2605419, 
    0.258276, 0.2489748, 0.3236983, 0.2633617, 0.3252949, 0.4157144, 
    0.3517084, 0.307364, 0.2721251, 0.2926622, 0.2355062, 0.2203614, 
    0.1412023, 0.2008214, 0.1125299, 0.2170012,
  0.001833516, 0.001156008, 0.0004785001, -0.0001990077, -0.0008765154, 
    -0.001554023, -0.002231531, 0.0001304686, 0.0001304686, 0.0001304686, 
    0.0001304686, 0.0001304686, 0.0001304686, 0.0001304686, -0.00242491, 
    -0.001654084, -0.0008832574, -0.0001124309, 0.0006583956, 0.001429222, 
    0.002200048, 0.002375565, 0.002282246, 0.002188927, 0.002095608, 
    0.00200229, 0.001908971, 0.001815652, 0.002375522,
  0.07647536, 0.03489848, 0.02510806, 0.00157916, 0, -9.324479e-07, 0, 0, 0, 
    0, 0, -0.0001472514, 0.002650928, 0.08133718, 0.1347611, 0.1785739, 
    0.3194836, 0.4694613, 0.4010493, 0.2851418, 0.2264029, 0.2837436, 
    0.3356674, 0.4679502, 0.3388142, 0.2825948, 0.3537048, 0.3110055, 
    0.1754355,
  0.1194645, 0.1665313, 0.2399783, 0.2593425, 0.2266139, 0.1397555, 
    0.1195791, 0.1425375, 0.1007601, 0.2723774, 0.2722411, 0.3057319, 
    0.2573773, 0.3377521, 0.3328564, 0.3159906, 0.251451, 0.2464013, 
    0.3123328, 0.3351609, 0.2821195, 0.328741, 0.2908233, 0.3833501, 
    0.2982525, 0.2644976, 0.2763142, 0.213345, 0.2101713,
  0.2100382, 0.2164904, 0.1915359, 0.2129172, 0.2193811, 0.2072737, 
    0.2955477, 0.2829805, 0.3116067, 0.3284143, 0.3233945, 0.3402365, 
    0.2656104, 0.3052772, 0.2422157, 0.2531235, 0.2252015, 0.2439469, 
    0.2166169, 0.22339, 0.2072238, 0.2252359, 0.2518632, 0.2051163, 
    0.1647159, 0.1623776, 0.1794368, 0.2305652, 0.202709,
  0.273238, 0.2036696, 0.2452988, 0.2003014, 0.2081518, 0.2738146, 0.2754861, 
    0.2642042, 0.207036, 0.2308053, 0.2136631, 0.159924, 0.1506741, 
    0.1187799, 0.1568574, 0.182195, 0.1883599, 0.2757801, 0.2144421, 
    0.2253504, 0.1724708, 0.2115472, 0.2365697, 0.1765059, 0.1545928, 
    0.1453731, 0.2055678, 0.2540051, 0.2204777,
  0.1508853, 0.135826, 0.1039711, 0.07385278, 0.1266462, 0.131007, 0.1314936, 
    0.1280248, 0.1008748, 0.08948378, 0.02872214, 0.07185324, 0.05414193, 
    0.1562239, 0.1713548, 0.1462066, 0.1118002, 0.0853911, 0.1678423, 
    0.1157188, 0.1101999, 0.1205265, 0.1652999, 0.1769242, 0.04124972, 
    0.1082487, 0.153211, 0.1683573, 0.2234579,
  0.02478536, -9.438155e-06, 0.04182207, 0.01058897, 0.02269346, 0.001853396, 
    0.007374474, 0.02899787, 0.02950861, 0.01458375, 0.0002284542, 
    8.505618e-06, 0.03141194, 0.0702555, 0.1072817, 0.09178548, 0.1088241, 
    0.1034356, 0.09320333, 0.04178584, 0.05671261, 0.04496034, 0.01610824, 
    0.0008057898, 0.03276881, 0.06952889, 0.08953035, 0.05142376, 0.04309557,
  3.646695e-08, 0.0003008201, 0.06757394, 0.005545137, 0.04276783, 
    0.007018921, 0.003303615, 0.001306403, 3.842993e-05, 0.001289729, 
    -2.422842e-06, -3.479212e-05, 1.1377e-05, 0.05139669, 0.03016726, 
    0.007461706, 0.04418514, 0.0577635, 0.02574305, 0.01128513, 0.00143967, 
    0.0001602856, 5.764891e-08, 3.512517e-06, 0.01923965, 0.01379087, 
    0.0006943824, 0.0002142442, 0.002865122,
  1.165835e-06, -0.0004912462, 0.0449942, 0.1427341, 0.0304802, 0.01111574, 
    0.06286444, 0.03186963, 0.005579358, 0.001221807, 0.06128595, 0.0446938, 
    0.2108176, 0.097049, 0.08350445, 0.03857398, 0.03702633, 0.01368609, 
    0.007387158, 2.663921e-05, 7.640176e-07, -1.066662e-07, 0.0004772643, 
    0.01315983, 0.016814, 4.821052e-05, 0.005968009, 6.35408e-06, 1.334746e-06,
  0.001928414, 0.1943994, 0.130474, 0.01036807, 0.002742698, 0.04815048, 
    0.03249428, 0.07161468, 0.08067434, 0.2187595, 0.0233999, 0.0198013, 
    0.03272701, 0.01444753, 0.01360105, 0.00319121, 0.001139864, 
    0.0005895642, 1.082581e-05, 4.973312e-05, 1.738121e-05, 0.01285146, 
    0.093305, 0.07546187, 0.1358178, 0.001885566, 0.004751223, 0.008435127, 
    0.001365529,
  0.1042962, 0.09693925, 0.07309131, 0.2612237, 0.04172579, 0.007064523, 
    0.06951988, 0.02719011, 0.04652961, 0.05982839, 0.0127139, 0.03795064, 
    0.0419773, 0.04291828, 0.04710279, 0.05843877, 0.1058688, 0.1893725, 
    0.2526208, 0.3215852, 0.2429081, 0.1154382, 0.1406438, 0.04155741, 
    0.01395364, 0.06908228, 0.09754371, 0.09662526, 0.1707393,
  0.0001531588, 8.038354e-05, 0.02925284, -1.733157e-05, -4.016148e-07, 
    -3.837491e-05, 0.1235345, 0.1114727, 0.2321734, 0.09386296, 0.07020234, 
    0.07572134, 0.05878037, 0.01790572, 0.02224801, 0.03850217, 0.006735058, 
    -1.899427e-05, 0.0009312472, 0.08462735, 0.06207132, 0.2056344, 0.022362, 
    0.04047018, 0.04265096, 0.03256647, 0.0003493621, 8.619647e-05, 
    0.000966338,
  2.602926e-06, 0.00124912, 2.69192e-08, 4.03209e-07, -4.941842e-08, 
    5.506359e-09, 0.01761992, 0.2985283, 0.4299231, 0.1026779, 0.03335024, 
    0.07352785, 0.0100239, 0.009858779, 0.06152725, 0.03020532, 0.04141927, 
    0.01981013, 4.852982e-07, 1.503983e-05, 0.08240108, 0.07755803, 
    0.05817365, 0.07914077, 0.02260021, 0.0368103, 0.01067476, 0.001045964, 
    -0.0001315439,
  0.03542497, 0.03486475, 0.001828649, 0.02374757, 0.007603129, 0.0009397747, 
    0.126838, 0.01401128, 0.02049115, 0.09299497, 0.06807565, 0.1419085, 
    0.07824692, 0.1140614, 0.1273014, 0.2760114, 0.1814464, 0.04944073, 
    0.0117245, 0.01087341, 0.06170644, 0.1280023, 0.07059369, 0.05891525, 
    0.1034674, 0.07606493, 0.03721988, 0.04435008, 0.0609454,
  0.1284322, 0.159899, 0.08547057, 0.1744499, 0.06563474, 0.1081732, 
    0.1791676, 0.2214481, 0.0888363, 0.1485593, 0.1710051, 0.1776279, 
    0.1620098, 0.1902487, 0.1428175, 0.1272002, 0.1728563, 0.1753898, 
    0.175827, 0.1251006, 0.1024121, 0.06951205, 0.2666713, 0.2610887, 
    0.1969434, 0.1613555, 0.2003626, 0.2184679, 0.1673542,
  0.1790364, 0.174217, 0.1739199, 0.2178084, 0.275099, 0.231245, 0.1603736, 
    0.214631, 0.1628873, 0.2097183, 0.22229, 0.1977596, 0.347939, 0.2339197, 
    0.2176016, 0.2124136, 0.1893728, 0.3169803, 0.2102986, 0.1520991, 
    0.1407766, 0.2725354, 0.1119229, 0.1941313, 0.2758224, 0.2480116, 
    0.2044826, 0.1823896, 0.2563127,
  0.3287213, 0.1809971, 0.2885613, 0.2946563, 0.3279235, 0.2203107, 
    0.1597587, 0.1665642, 0.1161581, 0.21119, 0.3426311, 0.3561343, 
    0.2416705, 0.1224742, 0.3539127, 0.1826747, 0.1491568, 0.1797685, 
    0.1529745, 0.2023404, 0.2753762, 0.1809116, 0.2706555, 0.4600051, 
    0.3307786, 0.3376185, 0.2561281, 0.1295853, 0.2115568,
  0.2405384, 0.2452959, 0.2013528, 0.1790768, 0.1404622, 0.1746421, 
    0.1868562, 0.2188511, 0.1721359, 0.1936071, 0.2857971, 0.3321667, 
    0.3492135, 0.3058443, 0.2448408, 0.2927376, 0.329673, 0.3723194, 
    0.4307334, 0.4071378, 0.3241114, 0.275574, 0.3419109, 0.2710873, 
    0.236402, 0.1522152, 0.1982482, 0.1275119, 0.2732365,
  0.005529186, 0.003127942, 0.0007266969, -0.001674548, -0.004075793, 
    -0.006477037, -0.008878282, 0.0006949429, 0.0007294692, 0.0007639954, 
    0.0007985216, 0.0008330478, 0.0008675741, 0.0009021003, -0.00455424, 
    -0.002519206, -0.0004841725, 0.001550861, 0.003585895, 0.005620929, 
    0.007655963, 0.01678466, 0.01711635, 0.01744803, 0.01777972, 0.0181114, 
    0.01844308, 0.01877477, 0.007450182,
  0.1005232, 0.04536717, 0.03780172, 0.02064471, 0.002177879, 0.0001568273, 
    2.240687e-05, 0, 0, 0, 0, 0.0008722527, 0.0257108, 0.07649966, 0.1082523, 
    0.1753649, 0.3203958, 0.4656482, 0.4079669, 0.3307453, 0.2643465, 
    0.3511878, 0.3533748, 0.471619, 0.3368057, 0.2737024, 0.3638711, 
    0.3243768, 0.2199409,
  0.1151861, 0.1765355, 0.2443689, 0.271779, 0.2586676, 0.1457113, 0.1185395, 
    0.1746323, 0.2095954, 0.332473, 0.3370849, 0.3373283, 0.2654972, 
    0.3320278, 0.3231967, 0.3020106, 0.2727212, 0.2493472, 0.2821052, 
    0.2735667, 0.2509601, 0.2965024, 0.2724393, 0.3939649, 0.2906246, 
    0.2942443, 0.2832165, 0.2138755, 0.2150802,
  0.2120051, 0.2295197, 0.1953373, 0.2314692, 0.2510425, 0.2061928, 
    0.2904891, 0.2996019, 0.2908891, 0.3048035, 0.3430057, 0.3411899, 
    0.2745343, 0.2968875, 0.257347, 0.307386, 0.255047, 0.2593087, 0.2247029, 
    0.2305101, 0.2201558, 0.231218, 0.2764083, 0.2405448, 0.1700011, 
    0.1550437, 0.2206765, 0.2476677, 0.2220909,
  0.2711019, 0.2172044, 0.2331717, 0.188812, 0.2233507, 0.2733836, 0.2909996, 
    0.2807744, 0.2095127, 0.2614607, 0.2234371, 0.1649413, 0.1636327, 
    0.1454007, 0.1673947, 0.2240168, 0.2202487, 0.3171369, 0.270533, 
    0.2407273, 0.1757329, 0.2511944, 0.2422253, 0.1759522, 0.1640587, 
    0.1798452, 0.2456326, 0.2218184, 0.2021066,
  0.1810287, 0.1597624, 0.1237984, 0.08129104, 0.1270927, 0.1718986, 
    0.1534842, 0.1340266, 0.1264397, 0.1079144, 0.0552119, 0.07662986, 
    0.0630728, 0.1571974, 0.1779497, 0.1412042, 0.1236706, 0.1001433, 
    0.2032137, 0.1476832, 0.130528, 0.1320854, 0.1985454, 0.1952839, 
    0.0262208, 0.1313977, 0.1708941, 0.1938994, 0.2304471,
  0.0320908, -0.000110095, 0.02401772, 0.008613284, 0.03512571, 0.009197719, 
    0.01672961, 0.03090089, 0.04185235, 0.009847257, -1.240581e-05, 
    -7.791127e-05, 0.03288909, 0.08052668, 0.1132891, 0.1005679, 0.1134829, 
    0.1164381, 0.1095526, 0.0581337, 0.06398343, 0.07976664, 0.02815642, 
    0.0009700824, 0.02660134, 0.06981777, 0.09707059, 0.05332248, 0.0525204,
  1.356271e-08, 6.754205e-05, 0.008383289, 0.001416912, 0.05867517, 0.033001, 
    0.004233577, 0.001429052, 1.866653e-05, 0.0002583269, -8.575476e-07, 
    -6.432585e-07, 0.0001824406, 0.06998571, 0.03326912, 0.007286044, 
    0.03765712, 0.07747815, 0.05885469, 0.05392614, 0.0130949, 0.003273241, 
    1.076127e-07, 2.048126e-06, 0.006007873, 0.006615003, 0.02055701, 
    0.00135201, 0.003986807,
  1.647701e-07, -0.0004683446, 0.01913212, 0.1794364, 0.04252485, 0.0106861, 
    0.0574735, 0.04748915, 0.008979148, 0.001760994, 0.04905617, 0.04566856, 
    0.2351873, 0.09431642, 0.06983246, 0.04033105, 0.0407984, 0.02068028, 
    0.008180354, 0.001146854, 2.581437e-06, 1.071465e-07, 3.068793e-05, 
    0.01272035, 0.004327673, -9.21027e-06, 0.02104434, 0.0006496399, 
    8.62377e-07,
  0.0001052793, 0.1702121, 0.09863594, 0.03301815, 0.006082571, 0.04117366, 
    0.02694633, 0.06973396, 0.07369472, 0.2110744, 0.02171067, 0.02048333, 
    0.0301824, 0.01594152, 0.01458872, 0.007055535, 0.002889855, 
    0.0009259439, 7.409132e-05, 1.913696e-05, 1.562092e-05, 0.01029392, 
    0.08055643, 0.06466585, 0.1162968, 0.0009840024, 0.005910411, 
    5.465436e-05, 9.290364e-05,
  0.07650749, 0.08188152, 0.05606735, 0.2593557, 0.01671974, 0.0051364, 
    0.07904291, 0.02900453, 0.03795865, 0.05101476, 0.01376115, 0.03624804, 
    0.04133359, 0.04003523, 0.04481767, 0.0556262, 0.1260603, 0.186698, 
    0.2716695, 0.3169089, 0.2149885, 0.1153746, 0.1431211, 0.04304097, 
    0.01633373, 0.05345106, 0.07938009, 0.07363835, 0.152669,
  2.232362e-05, 4.1128e-06, 0.01750815, -1.336629e-05, -4.868187e-07, 
    -1.260199e-06, 0.09832024, 0.1179191, 0.2368885, 0.1039789, 0.07089383, 
    0.07304586, 0.05203622, 0.01971501, 0.02218514, 0.03739905, 0.0255324, 
    0.0005468963, 0.003137563, 0.09715462, 0.05946757, 0.2294027, 0.0209076, 
    0.03792662, 0.03842419, 0.04331903, 0.0001666848, 4.955646e-05, 
    0.0003719759,
  4.264403e-06, 0.0002524523, 7.183042e-05, 2.273125e-07, -2.307782e-08, 
    1.608537e-09, 0.005945625, 0.3165406, 0.4294893, 0.09590238, 0.03398895, 
    0.07868769, 0.01349348, 0.01306072, 0.06040238, 0.03339549, 0.05435874, 
    0.02013835, 0.000437617, -6.694996e-07, 0.06664899, 0.08583584, 
    0.05203283, 0.07452536, 0.02425893, 0.03725917, 0.019228, 0.001819669, 
    -3.071247e-05,
  0.03271645, 0.0201264, 0.003481828, 0.03083046, 0.002095358, -2.525027e-05, 
    0.1099697, 0.0098116, 0.01080811, 0.08708869, 0.07058375, 0.134164, 
    0.07722776, 0.13693, 0.1260494, 0.2837209, 0.1714579, 0.06630038, 
    0.01330169, 0.003419608, 0.05046268, 0.1227902, 0.07025225, 0.06330252, 
    0.1110068, 0.08359996, 0.03879655, 0.05321606, 0.06110597,
  0.127199, 0.1707396, 0.07576134, 0.1689656, 0.07037221, 0.1300482, 
    0.1576387, 0.2036495, 0.07730092, 0.1607858, 0.179096, 0.2036876, 
    0.1805606, 0.1906329, 0.1650139, 0.1887846, 0.195072, 0.1971885, 
    0.184556, 0.1569083, 0.1129083, 0.07642302, 0.2785999, 0.2790411, 
    0.1995703, 0.1698214, 0.2069459, 0.2313512, 0.1666382,
  0.2040172, 0.1742638, 0.2020045, 0.2748092, 0.3352232, 0.2041918, 
    0.1898999, 0.2775393, 0.150717, 0.1949362, 0.2340097, 0.2315235, 
    0.3373347, 0.2521609, 0.2742676, 0.2304952, 0.2134119, 0.3255211, 
    0.2213709, 0.1881293, 0.1720818, 0.3194876, 0.1365678, 0.2300209, 
    0.3255662, 0.2489393, 0.2291991, 0.2076753, 0.2648271,
  0.3309936, 0.1716998, 0.259591, 0.2803484, 0.3010642, 0.207457, 0.155356, 
    0.182154, 0.1170753, 0.2792285, 0.4133455, 0.4333017, 0.1901002, 
    0.1474883, 0.2931549, 0.2058492, 0.2355324, 0.2101434, 0.1561885, 
    0.1949898, 0.2068182, 0.1636546, 0.3169241, 0.4302333, 0.3669583, 
    0.3873476, 0.2593691, 0.1462138, 0.2445074,
  0.2412694, 0.2192696, 0.1533562, 0.1541149, 0.1328902, 0.1137029, 
    0.1411327, 0.1683849, 0.1423879, 0.198415, 0.3009819, 0.2806513, 
    0.2417809, 0.229215, 0.2100829, 0.2865367, 0.2989309, 0.2676682, 
    0.3713276, 0.4429687, 0.3242337, 0.2595077, 0.3142441, 0.2873918, 
    0.2613695, 0.1639883, 0.1997855, 0.1341373, 0.2720466,
  0.03075307, 0.02672863, 0.02270419, 0.01867975, 0.01465531, 0.01063087, 
    0.006606435, 0.007592264, 0.007053259, 0.006514254, 0.00597525, 
    0.005436246, 0.004897241, 0.004358237, 0.001995303, 0.006630994, 
    0.01126669, 0.01590238, 0.02053807, 0.02517376, 0.02980945, 0.03598514, 
    0.0359129, 0.03584065, 0.0357684, 0.03569615, 0.0356239, 0.03555166, 
    0.03397262,
  0.1389418, 0.06027723, 0.04431556, 0.02851085, 0.007830996, 0.0005465415, 
    9.787298e-06, -1.911436e-06, 0, 0, -0.0007519519, 0.02976606, 0.02772136, 
    0.08193622, 0.09905991, 0.1564675, 0.3447239, 0.4590985, 0.4059911, 
    0.342512, 0.3064207, 0.3878246, 0.3774493, 0.4607448, 0.3242897, 
    0.2493565, 0.3601713, 0.3190837, 0.244112,
  0.1289874, 0.1658173, 0.2494069, 0.2754923, 0.2869496, 0.1417523, 
    0.1266822, 0.1769311, 0.2721239, 0.3573496, 0.3414056, 0.3434828, 
    0.2559159, 0.3418925, 0.3375087, 0.3129952, 0.2743818, 0.2611759, 
    0.2867086, 0.2643564, 0.215721, 0.276178, 0.2910385, 0.3954065, 
    0.2943494, 0.2926241, 0.2608023, 0.1856834, 0.2023271,
  0.2521562, 0.1855132, 0.2034334, 0.2672359, 0.2923257, 0.2443373, 
    0.3280085, 0.3229318, 0.3143474, 0.3560909, 0.3765007, 0.366001, 
    0.2958362, 0.3055243, 0.2614895, 0.3392722, 0.2749325, 0.2615091, 
    0.2535357, 0.2149359, 0.2186989, 0.2449225, 0.3234287, 0.2321293, 
    0.2061728, 0.1399523, 0.2046946, 0.2266737, 0.2484037,
  0.2474904, 0.2044286, 0.2143398, 0.1971817, 0.2276836, 0.2949913, 
    0.3034806, 0.3074273, 0.2216318, 0.2584576, 0.2636236, 0.1873678, 
    0.1655806, 0.1610634, 0.2107718, 0.220898, 0.2285195, 0.2621903, 
    0.2673247, 0.2978846, 0.207243, 0.2478515, 0.2557019, 0.1712242, 
    0.1879699, 0.1909861, 0.2149599, 0.2177547, 0.2318229,
  0.1954959, 0.1681815, 0.1464512, 0.09535921, 0.1318531, 0.1988344, 
    0.1574898, 0.1787806, 0.1567592, 0.1296879, 0.08287417, 0.09675433, 
    0.06816357, 0.1927506, 0.1930585, 0.156937, 0.1519146, 0.1269842, 
    0.2074186, 0.1763072, 0.1832049, 0.1698112, 0.2038569, 0.2232794, 
    0.02613217, 0.1342467, 0.1834795, 0.2059232, 0.2535377,
  0.03461768, 0.0002482166, 0.007996898, 0.02328973, 0.02871296, 0.02943171, 
    0.01764766, 0.04448528, 0.04375869, 0.01099834, -8.904622e-05, 
    -9.134402e-05, 0.03017223, 0.094731, 0.09339295, 0.1006647, 0.1227322, 
    0.1526162, 0.08413967, 0.0658455, 0.09635753, 0.1427589, 0.05162931, 
    0.001458359, 0.02606478, 0.06364027, 0.09730942, 0.05702161, 0.06747837,
  -4.627899e-07, 2.179279e-06, 0.001379876, 0.0007333254, 0.05090511, 
    0.05191828, 0.02314581, 0.004687021, 0.01098427, 5.365543e-05, 
    -1.204369e-07, -9.181851e-09, 0.001351729, 0.1041742, 0.0476479, 
    0.01484824, 0.03039078, 0.07314532, 0.04780534, 0.06471232, 0.04296776, 
    0.00783251, 7.068776e-08, 2.411259e-06, 0.004111765, 0.001928612, 
    0.034792, 0.01504487, 0.009992298,
  7.978789e-08, -0.000173021, 0.003168482, 0.1460926, 0.04673343, 0.01405784, 
    0.05538591, 0.06982853, 0.0124321, 0.003109116, 0.04349631, 0.04785701, 
    0.2479115, 0.09023162, 0.05517622, 0.03575943, 0.03591955, 0.02400373, 
    0.009770884, 0.0122523, 5.825724e-05, 5.109147e-07, 8.996147e-06, 
    0.01200109, 0.002634341, -2.654473e-05, 0.03708266, 0.0009214146, 
    8.645841e-07,
  0.0002492362, 0.1654136, 0.07952537, 0.03263509, 0.01191049, 0.03796534, 
    0.0232556, 0.0644137, 0.06728536, 0.2084106, 0.02436076, 0.01988786, 
    0.02665181, 0.0169333, 0.01356727, 0.01615734, 0.01011394, 0.009132866, 
    0.002790533, 0.0001514901, 4.939462e-05, 0.007735413, 0.04972196, 
    0.05949114, 0.03905394, 0.00105437, 0.01155507, 0.000418045, -1.651656e-05,
  0.05694303, 0.07870446, 0.04772411, 0.2241238, 0.006793058, 0.005614719, 
    0.08029379, 0.0276266, 0.03076608, 0.04313954, 0.01426396, 0.03932777, 
    0.03632559, 0.03782116, 0.03789623, 0.05196637, 0.1338331, 0.1729033, 
    0.2824615, 0.3107769, 0.1965048, 0.1173184, 0.1474839, 0.0498366, 
    0.0185821, 0.03910546, 0.06513776, 0.0663086, 0.141027,
  -5.389967e-07, 1.019022e-06, 0.00483201, -1.53112e-05, -4.828983e-07, 
    8.193814e-06, 0.07424577, 0.1165224, 0.2434722, 0.100072, 0.07367443, 
    0.07273782, 0.0456997, 0.01941237, 0.02097692, 0.03033847, 0.06141961, 
    0.01828724, 0.009296999, 0.1201164, 0.05323125, 0.2325665, 0.0193267, 
    0.02984276, 0.03622757, 0.04184837, 0.0009291442, 3.019728e-05, 
    0.0001323053,
  2.485908e-06, 5.106231e-05, 0.0001073717, 1.51291e-07, -1.365322e-08, 
    3.884493e-10, 0.002403821, 0.2454945, 0.4342431, 0.1071688, 0.03374971, 
    0.08263223, 0.01703392, 0.02562304, 0.05903713, 0.02937358, 0.06239573, 
    0.03821415, 0.007478826, -6.042226e-06, 0.04672026, 0.07100063, 
    0.03864912, 0.06587023, 0.02811994, 0.03319521, 0.03624824, 0.004381073, 
    -9.476362e-05,
  0.02341702, 0.01760759, 0.00145399, 0.03862656, 0.00178944, -3.140541e-05, 
    0.09439593, 0.0046634, 0.006134491, 0.103848, 0.08153173, 0.1367388, 
    0.09299397, 0.1629537, 0.1574394, 0.2927031, 0.1582604, 0.08662982, 
    0.006036938, 0.00098455, 0.03275576, 0.05736083, 0.07160265, 0.06592484, 
    0.1225619, 0.08255691, 0.05347643, 0.07515145, 0.0462748,
  0.1244504, 0.1741103, 0.06000031, 0.1311942, 0.06026094, 0.1244556, 
    0.1498201, 0.2007293, 0.08081446, 0.1584947, 0.1828771, 0.2264091, 
    0.160631, 0.1868469, 0.1726782, 0.2199703, 0.2195994, 0.1810519, 
    0.1496999, 0.1616036, 0.1180666, 0.08892821, 0.2467567, 0.3275275, 
    0.1955728, 0.1867333, 0.2197979, 0.269169, 0.1633933,
  0.2177271, 0.1901635, 0.1947473, 0.2760732, 0.3028327, 0.1971757, 
    0.2136864, 0.2186167, 0.1773723, 0.2262623, 0.2243017, 0.2341603, 
    0.3038625, 0.2574506, 0.2870544, 0.2230112, 0.255989, 0.3297948, 
    0.2663962, 0.1662053, 0.1701866, 0.2994697, 0.1751465, 0.2382305, 
    0.359878, 0.2122706, 0.2552864, 0.2111647, 0.2807839,
  0.2809982, 0.2216419, 0.2771038, 0.2343986, 0.2699746, 0.2611783, 
    0.1833668, 0.2350364, 0.1517662, 0.2864436, 0.4064387, 0.4077676, 
    0.1334633, 0.192318, 0.2261245, 0.1921876, 0.1563346, 0.2112367, 
    0.1379831, 0.2216662, 0.2082816, 0.2143798, 0.359923, 0.4538781, 
    0.3309464, 0.3609003, 0.22772, 0.1820098, 0.214588,
  0.2382369, 0.2205017, 0.1236013, 0.09242239, 0.1297504, 0.1179355, 
    0.1180084, 0.1485324, 0.1256966, 0.2353938, 0.2162688, 0.1888677, 
    0.2043615, 0.2367793, 0.2163151, 0.3341617, 0.2454124, 0.2744105, 
    0.3574058, 0.391171, 0.3010404, 0.2619051, 0.2320397, 0.3454236, 
    0.282161, 0.2818694, 0.1812389, 0.1265854, 0.231156,
  0.07431089, 0.06730748, 0.06030407, 0.05330066, 0.04629725, 0.03929384, 
    0.03229044, 0.0435973, 0.04282419, 0.04205107, 0.04127796, 0.04050484, 
    0.03973172, 0.03895861, -0.0002885437, 0.01147191, 0.02323236, 
    0.03499281, 0.04675326, 0.05851372, 0.07027417, 0.1220781, 0.1180942, 
    0.1141102, 0.1101263, 0.1061424, 0.1021585, 0.09817454, 0.07991362,
  0.1732562, 0.08541671, 0.04595749, 0.03111274, 0.009095764, -0.0003444556, 
    0.003862443, -6.127153e-05, -7.111904e-06, -5.148581e-05, -0.001657828, 
    0.03313326, 0.04365393, 0.08002091, 0.1000286, 0.1496243, 0.3388016, 
    0.4627903, 0.4086493, 0.3256359, 0.3458649, 0.4054938, 0.3798548, 
    0.4638514, 0.3041305, 0.2324222, 0.3481521, 0.3000687, 0.271527,
  0.1466881, 0.1732305, 0.2413886, 0.260507, 0.2991045, 0.1403336, 0.1169346, 
    0.1952205, 0.3085006, 0.3677857, 0.3394767, 0.3133852, 0.2552348, 
    0.358905, 0.3799954, 0.3096713, 0.2618289, 0.2482179, 0.3114217, 
    0.2709908, 0.2108407, 0.2615442, 0.2945946, 0.4080103, 0.2557031, 
    0.2704881, 0.2687582, 0.1931678, 0.2112357,
  0.2543906, 0.2059079, 0.2080717, 0.3084827, 0.345741, 0.2890138, 0.3616968, 
    0.3494098, 0.3514276, 0.4646564, 0.4131786, 0.3611138, 0.3149605, 
    0.363124, 0.3030156, 0.3354198, 0.3349261, 0.3009046, 0.2806856, 
    0.2992234, 0.2608744, 0.3161592, 0.3557258, 0.2368624, 0.2195873, 
    0.1554045, 0.2514131, 0.2883708, 0.2262398,
  0.2939183, 0.2468044, 0.2512011, 0.2406513, 0.2623397, 0.3341675, 
    0.3057934, 0.3180012, 0.2671947, 0.3086397, 0.2635188, 0.2148467, 
    0.2221612, 0.2132787, 0.2437327, 0.2406601, 0.2979321, 0.3328438, 
    0.3416271, 0.3933671, 0.2683054, 0.2347552, 0.3136841, 0.2029435, 
    0.1838885, 0.1656857, 0.2285894, 0.2622769, 0.2427071,
  0.2333917, 0.2143048, 0.1832414, 0.1263702, 0.189884, 0.2508043, 0.1978209, 
    0.2398535, 0.2128705, 0.201907, 0.1004973, 0.1311408, 0.07045393, 
    0.2357156, 0.2047371, 0.2085132, 0.1726491, 0.185303, 0.2035611, 
    0.2125457, 0.2275536, 0.1950603, 0.2147501, 0.251075, 0.04341839, 
    0.1691288, 0.2303462, 0.232372, 0.2965875,
  0.06982718, 0.01528461, 0.003268119, 0.04787118, 0.03074016, 0.04597864, 
    0.0331888, 0.06657109, 0.06744877, 0.02601721, -0.0001348545, 
    -1.06029e-05, 0.01825172, 0.1148634, 0.1081305, 0.1059383, 0.1242651, 
    0.1622152, 0.08311082, 0.05894334, 0.159716, 0.1735889, 0.1056475, 
    0.000898465, 0.03016936, 0.05293081, 0.09996013, 0.08961099, 0.0833924,
  -1.411863e-05, 8.607262e-07, 0.0003336534, 0.001126461, 0.03916772, 
    0.05315551, 0.06757045, 0.03127221, 0.02195351, 0.0002048376, 
    2.009975e-08, 3.688461e-09, 0.05386658, 0.1268316, 0.07128432, 
    0.01497813, 0.02814509, 0.07738552, 0.03091303, 0.04625978, 0.08221256, 
    0.02686788, 1.118744e-05, 2.465938e-06, 0.001355976, 0.0007386891, 
    0.0547546, 0.05905259, 0.0176417,
  1.638152e-06, -5.610984e-05, 0.0005008285, 0.09670761, 0.04487142, 
    0.01967358, 0.06153359, 0.0711432, 0.01394955, 0.007191752, 0.04248311, 
    0.06816103, 0.2519761, 0.08233263, 0.04049455, 0.03160925, 0.0316078, 
    0.02072173, 0.0104494, 0.02488891, 0.006477505, 3.102792e-05, 
    1.534443e-06, 0.01255529, 0.001796226, 6.880336e-07, 0.04953949, 
    0.0110036, 1.638116e-06,
  0.0009668152, 0.1646043, 0.06456368, 0.03463247, 0.02151822, 0.03564264, 
    0.02125935, 0.05694669, 0.05957048, 0.2144113, 0.0242341, 0.01762881, 
    0.02280928, 0.01831892, 0.01510747, 0.01523424, 0.01685803, 0.01807575, 
    0.01530096, 0.00402881, 0.0001367982, 0.001910471, 0.020493, 0.05674592, 
    0.01293143, 0.002049824, 0.01700345, 0.004526397, 8.847763e-05,
  0.05122317, 0.07801046, 0.03993502, 0.1827939, 0.001856541, 0.004680024, 
    0.07068893, 0.02643862, 0.02321012, 0.03542954, 0.01469106, 0.0383081, 
    0.02928406, 0.03210848, 0.03258336, 0.04464503, 0.1258708, 0.1687814, 
    0.2787388, 0.2898288, 0.1712811, 0.1126548, 0.1498639, 0.06066702, 
    0.01960175, 0.03537303, 0.05535164, 0.05971316, 0.122237,
  -7.81846e-07, 3.665185e-07, 0.001902678, 0.000158933, -4.477739e-07, 
    -1.347894e-05, 0.06308197, 0.1088817, 0.2638234, 0.1007599, 0.06226614, 
    0.06321181, 0.03880348, 0.0195293, 0.02059871, 0.0278569, 0.05810255, 
    0.08256998, 0.003141408, 0.1561354, 0.05408909, 0.2318213, 0.01843393, 
    0.02192335, 0.034855, 0.03721653, 0.01018262, 1.429321e-05, 6.824129e-05,
  1.642692e-06, 1.315777e-05, 4.239934e-05, 1.099568e-07, -8.376738e-09, 
    5.290341e-11, 0.0004297852, 0.1964973, 0.4486237, 0.1045467, 0.03451004, 
    0.07378199, 0.02061787, 0.02190036, 0.04789451, 0.04279676, 0.0607513, 
    0.07856577, 0.01652828, -2.162464e-06, 0.03371767, 0.04481453, 
    0.04338362, 0.06067742, 0.04085915, 0.02967767, 0.0469427, 0.01302559, 
    -0.0001493083,
  0.01795151, 0.01940579, 0.00400048, 0.05604896, 0.002619343, -5.423813e-06, 
    0.07963482, 0.001607105, 0.004215862, 0.08849474, 0.08387627, 0.1282052, 
    0.1236873, 0.1667167, 0.1906794, 0.3167116, 0.1928132, 0.1383516, 
    0.01261725, 0.0001214485, 0.02658992, 0.0269152, 0.07432641, 0.1085657, 
    0.1415939, 0.1302102, 0.08949497, 0.1004276, 0.05155107,
  0.1470694, 0.1593872, 0.05868125, 0.143937, 0.07508241, 0.1021049, 
    0.1084321, 0.1941706, 0.08398169, 0.1473528, 0.1839581, 0.237919, 
    0.158993, 0.2134386, 0.1885004, 0.2154383, 0.2265206, 0.2259726, 
    0.1799877, 0.1561515, 0.130183, 0.09315621, 0.245836, 0.347319, 
    0.2096131, 0.2003604, 0.2522953, 0.29174, 0.1484606,
  0.2388815, 0.1935776, 0.1735095, 0.2905797, 0.279832, 0.19961, 0.1725309, 
    0.1851496, 0.1843573, 0.2971689, 0.2271365, 0.2810159, 0.2920443, 
    0.274476, 0.3156728, 0.2750612, 0.2563109, 0.351535, 0.2896383, 
    0.1790378, 0.1812547, 0.295948, 0.2627467, 0.2748823, 0.3844668, 
    0.184706, 0.3306986, 0.2579961, 0.3227421,
  0.3129343, 0.2110513, 0.3248868, 0.2810824, 0.3538919, 0.1815505, 
    0.1589836, 0.2236538, 0.1830431, 0.3156222, 0.4210799, 0.4195206, 
    0.1626163, 0.2249069, 0.2262324, 0.2415245, 0.1680119, 0.1826887, 
    0.1833944, 0.2670967, 0.2166854, 0.2697132, 0.3152452, 0.4547046, 
    0.2978854, 0.3534817, 0.2501428, 0.1628248, 0.2857421,
  0.2251528, 0.2192052, 0.1857569, 0.1329374, 0.1812272, 0.1559338, 
    0.1506066, 0.1507406, 0.1600844, 0.1807833, 0.2522063, 0.2169681, 
    0.2139033, 0.2808799, 0.268885, 0.3043515, 0.2749271, 0.3419413, 
    0.3899472, 0.3780125, 0.3158312, 0.3316482, 0.2168928, 0.3023241, 
    0.301083, 0.2670924, 0.1956307, 0.1407169, 0.2120166,
  0.13739, 0.1291475, 0.1209049, 0.1126623, 0.1044197, 0.09617709, 
    0.08793449, 0.08277111, 0.08440508, 0.08603905, 0.08767302, 0.08930699, 
    0.09094096, 0.09257493, 0.07846242, 0.09329171, 0.108121, 0.1229503, 
    0.1377796, 0.1526089, 0.1674381, 0.2091756, 0.200955, 0.1927343, 
    0.1845136, 0.176293, 0.1680723, 0.1598516, 0.1439841,
  0.2023837, 0.1321262, 0.05491048, 0.03349486, 0.008662321, -0.00129946, 
    0.006284385, 0.0006961452, 0.003199973, 0.007109885, 0.009927452, 
    0.05558569, 0.06251793, 0.06831723, 0.1085572, 0.1326181, 0.3116684, 
    0.478104, 0.4451499, 0.3144446, 0.3741811, 0.4093955, 0.3836781, 
    0.4467451, 0.294459, 0.2266338, 0.333922, 0.2795829, 0.2891826,
  0.1488972, 0.1708384, 0.2393283, 0.2501229, 0.2867453, 0.1399146, 
    0.1027296, 0.2124843, 0.3302119, 0.3854171, 0.3271461, 0.2936323, 
    0.2511319, 0.3302704, 0.3887299, 0.3144372, 0.2470692, 0.2373237, 
    0.2888996, 0.2754263, 0.210268, 0.274511, 0.3204896, 0.4228413, 
    0.2306338, 0.2721877, 0.3190709, 0.2181195, 0.2271617,
  0.2626636, 0.2373839, 0.2701308, 0.4207704, 0.4261359, 0.3135641, 
    0.3634737, 0.3458591, 0.3635194, 0.4828605, 0.3802526, 0.3143046, 
    0.3216594, 0.3372388, 0.3199877, 0.3561246, 0.3636583, 0.3857305, 
    0.3916565, 0.3530456, 0.3674555, 0.3476231, 0.3926513, 0.2886963, 
    0.2956287, 0.1953092, 0.3117241, 0.3276382, 0.2463285,
  0.3565422, 0.3296855, 0.3634605, 0.2943151, 0.3311492, 0.3663196, 
    0.3276026, 0.3120556, 0.2674044, 0.3120311, 0.274129, 0.2460068, 
    0.3185298, 0.3107761, 0.3263381, 0.336086, 0.2985975, 0.4325283, 
    0.4064496, 0.4066143, 0.2965398, 0.2493389, 0.3728314, 0.230648, 
    0.1855781, 0.2116403, 0.3286255, 0.3322092, 0.2971406,
  0.3241813, 0.1891334, 0.2110811, 0.1952285, 0.2702565, 0.2713623, 
    0.2614786, 0.2206423, 0.2495448, 0.2141756, 0.1211088, 0.1346246, 
    0.1119746, 0.2746186, 0.2529892, 0.2669271, 0.1748958, 0.2662031, 
    0.2948335, 0.2661768, 0.2835056, 0.2235017, 0.2181734, 0.282302, 
    0.06863407, 0.1560509, 0.2591302, 0.335646, 0.3251947,
  0.1076475, 0.03822297, 0.001386873, 0.09088421, 0.05087084, 0.08802218, 
    0.09279126, 0.08454019, 0.1655371, 0.06001174, 0.0005107262, 
    2.554104e-06, 0.01256648, 0.1780708, 0.1563617, 0.1534309, 0.1409838, 
    0.1873041, 0.1446559, 0.1639615, 0.1770005, 0.1986955, 0.1759281, 
    0.002496709, 0.03779695, 0.1176914, 0.1661339, 0.1601615, 0.1416098,
  0.000574798, 2.041468e-07, 7.973306e-05, 0.005713483, 0.042557, 0.05182599, 
    0.126399, 0.1378319, 0.06193157, 0.0003173519, 8.523886e-09, 
    1.787193e-09, 0.09657551, 0.1381199, 0.08460295, 0.0223322, 0.05010423, 
    0.08476403, 0.03503681, 0.05066842, 0.1465059, 0.3169098, 0.07831353, 
    8.261536e-07, 0.0007431727, 0.0005263531, 0.08630284, 0.1304783, 0.1030526,
  1.404247e-05, 0.0001071593, 0.0001220939, 0.05800681, 0.04674672, 
    0.02556581, 0.06535821, 0.06463712, 0.02954032, 0.02957933, 0.04196752, 
    0.07955135, 0.2297867, 0.07300439, 0.03429684, 0.03158445, 0.03101067, 
    0.02495694, 0.01546974, 0.02525871, 0.04164493, 0.01053761, 3.35018e-06, 
    0.01145961, 0.00104095, 3.097272e-09, 0.05649609, 0.08854702, 0.0001329132,
  0.01146382, 0.1720658, 0.05589397, 0.03294958, 0.02711609, 0.03716628, 
    0.02310224, 0.04905798, 0.05297385, 0.2208867, 0.02319337, 0.01788374, 
    0.02401388, 0.02233554, 0.01937986, 0.01374844, 0.01712765, 0.01683774, 
    0.02369863, 0.02700617, 0.004181264, 0.0004249213, 0.008666172, 
    0.05364805, 0.007143456, 0.004905305, 0.02083903, 0.0183539, 0.003839063,
  0.04584373, 0.06956729, 0.02777992, 0.1378981, 0.0001828627, 0.006571749, 
    0.06144964, 0.02879012, 0.020146, 0.02996642, 0.01496334, 0.03788802, 
    0.02557865, 0.0284168, 0.02965779, 0.04316589, 0.1051544, 0.1469893, 
    0.2520833, 0.2565865, 0.1461678, 0.09372325, 0.1559492, 0.05969953, 
    0.02264899, 0.031447, 0.05716297, 0.05497781, 0.1178357,
  -5.18444e-07, 1.922265e-07, 6.419271e-05, 0.0005638553, -3.802528e-07, 
    -3.740958e-05, 0.05156835, 0.09714387, 0.2633452, 0.113306, 0.06278432, 
    0.05530758, 0.0348804, 0.02185282, 0.02384376, 0.02992276, 0.05674107, 
    0.1487294, 0.02500474, 0.1748543, 0.05667802, 0.2258062, 0.02211746, 
    0.02454565, 0.0394815, 0.03854682, 0.01775677, -2.146035e-05, 3.0716e-05,
  1.136667e-06, 2.714303e-06, 3.196413e-05, 8.526924e-08, -6.009561e-09, 
    -1.560212e-11, -3.895174e-05, 0.1777948, 0.4655047, 0.122942, 0.03575813, 
    0.08595965, 0.02705235, 0.05827654, 0.06451593, 0.106751, 0.07371217, 
    0.1121674, 0.1012194, -6.869033e-06, 0.02256686, 0.03710071, 0.06957291, 
    0.05804297, 0.03802956, 0.03601857, 0.05329117, 0.07800706, 0.0012998,
  0.01515259, 0.01884665, 0.004776714, 0.08339152, 0.001000885, 
    -2.592025e-06, 0.06314831, -2.226175e-05, 0.001735528, 0.06717302, 
    0.08944507, 0.1307765, 0.1452228, 0.1810976, 0.223646, 0.3787556, 
    0.2577367, 0.1990214, 0.05157809, -8.235875e-05, 0.0163848, 0.02167817, 
    0.08696273, 0.138681, 0.182581, 0.152444, 0.1521559, 0.2057094, 0.05772036,
  0.1727493, 0.168885, 0.05728019, 0.1259896, 0.04582364, 0.07770689, 
    0.09793709, 0.1879329, 0.1027286, 0.1425102, 0.1340915, 0.2133402, 
    0.181307, 0.237434, 0.2642808, 0.2351754, 0.2401305, 0.2486455, 
    0.2047004, 0.1643645, 0.1207296, 0.08464331, 0.256885, 0.3660543, 
    0.2018899, 0.2094257, 0.3174714, 0.2834112, 0.1710171,
  0.2819978, 0.2169685, 0.239817, 0.2597709, 0.2784396, 0.2247833, 0.1614042, 
    0.1724066, 0.1891694, 0.3328036, 0.2792212, 0.3216231, 0.3176599, 
    0.4003282, 0.3768623, 0.3683471, 0.3033965, 0.3742708, 0.3148095, 
    0.1929451, 0.2262985, 0.2830875, 0.4086622, 0.3315172, 0.441129, 
    0.1671761, 0.3590569, 0.2722186, 0.3552965,
  0.3476051, 0.3009394, 0.3528638, 0.3409331, 0.4040375, 0.216343, 0.2011106, 
    0.1967962, 0.1761584, 0.4349975, 0.4097056, 0.4620698, 0.2693544, 
    0.3030103, 0.3349178, 0.2408721, 0.2316797, 0.2414467, 0.2594195, 
    0.3559497, 0.3796694, 0.3687994, 0.3832137, 0.44775, 0.3216747, 
    0.3746468, 0.2607035, 0.1737813, 0.4050836,
  0.2272309, 0.2462976, 0.2441442, 0.1804565, 0.222769, 0.2037449, 0.2118389, 
    0.2065288, 0.2712457, 0.2624949, 0.3350611, 0.3238932, 0.3294708, 
    0.3708914, 0.3904172, 0.3710391, 0.3996067, 0.4323914, 0.4613145, 
    0.483986, 0.4195098, 0.3677654, 0.2978303, 0.2773727, 0.225267, 
    0.2748976, 0.2043737, 0.1828617, 0.2312562,
  0.1638758, 0.155448, 0.1470203, 0.1385925, 0.1301648, 0.121737, 0.1133093, 
    0.1323165, 0.137756, 0.1431956, 0.1486351, 0.1540747, 0.1595142, 
    0.1649538, 0.1747637, 0.1870399, 0.1993161, 0.2115923, 0.2238684, 
    0.2361446, 0.2484208, 0.2362301, 0.2269422, 0.2176542, 0.2083662, 
    0.1990782, 0.1897902, 0.1805022, 0.170618,
  0.2326793, 0.1633229, 0.06369261, 0.03966782, 0.007511571, -0.001745113, 
    0.002980092, 0.005347523, 0.004278996, 0.008727815, 0.02275307, 
    0.08280959, 0.09385412, 0.06713123, 0.1052049, 0.1248096, 0.292928, 
    0.4867602, 0.4517043, 0.315919, 0.386428, 0.4013686, 0.3626745, 
    0.4108987, 0.3026397, 0.2235744, 0.2985362, 0.2428082, 0.2928989,
  0.1657897, 0.1524919, 0.2276944, 0.2318842, 0.2543149, 0.134455, 
    0.07628104, 0.2275018, 0.3346779, 0.3961068, 0.3283449, 0.2712892, 
    0.2327825, 0.2865151, 0.3767106, 0.3087866, 0.2513007, 0.2353504, 
    0.2716961, 0.2836015, 0.2499778, 0.2966481, 0.3334723, 0.4426018, 
    0.2148911, 0.2683932, 0.3168673, 0.2525544, 0.2581429,
  0.3062772, 0.2858591, 0.4042987, 0.4324662, 0.4045802, 0.3323407, 
    0.3753296, 0.347918, 0.3715112, 0.4468762, 0.3123349, 0.3085023, 
    0.3735193, 0.2985651, 0.2910382, 0.3448298, 0.3716519, 0.452399, 
    0.4165414, 0.4066304, 0.4205409, 0.2857496, 0.3609547, 0.3154448, 
    0.3950054, 0.2618237, 0.3695093, 0.3879559, 0.3370309,
  0.4088067, 0.3513134, 0.3904786, 0.3148902, 0.3603281, 0.3454298, 
    0.3093149, 0.2867869, 0.2520432, 0.2813716, 0.2818932, 0.23793, 
    0.2325072, 0.234094, 0.3078991, 0.316439, 0.331008, 0.4091124, 0.3958351, 
    0.4411854, 0.3137072, 0.269743, 0.3464892, 0.2380996, 0.2219249, 
    0.2650352, 0.3347467, 0.3751327, 0.4498834,
  0.2549471, 0.2113999, 0.1673733, 0.2067034, 0.2991565, 0.2646797, 0.203168, 
    0.2175677, 0.2958781, 0.2776806, 0.1353937, 0.1140963, 0.06498095, 
    0.2167153, 0.3305631, 0.2630419, 0.2191033, 0.2231781, 0.286401, 
    0.2658257, 0.2337737, 0.1715535, 0.1818748, 0.3369967, 0.08133449, 
    0.1385486, 0.2448151, 0.350602, 0.3347663,
  0.2402462, 0.06549629, 0.001666789, 0.08333573, 0.07965352, 0.1701309, 
    0.1668936, 0.1426898, 0.2004453, 0.06206641, 0.0007818926, 2.833398e-06, 
    0.01181943, 0.2427074, 0.1787805, 0.1804791, 0.1487676, 0.2479509, 
    0.1884579, 0.1246731, 0.1780373, 0.2118924, 0.1813386, 0.006562364, 
    0.0369544, 0.1194473, 0.212869, 0.2014035, 0.1377925,
  0.154377, -8.276752e-08, 4.068361e-06, 0.01173884, 0.05862113, 0.05207556, 
    0.1134878, 0.2450821, 0.2030085, 0.0002597567, 4.849593e-09, 
    1.484097e-09, 0.1033355, 0.1696794, 0.08926201, 0.0320079, 0.06690672, 
    0.09552398, 0.04903804, 0.0592514, 0.2902693, 0.4995239, 0.4592336, 
    -3.25379e-06, 0.004253324, 0.001986967, 0.09727678, 0.2588501, 0.328237,
  0.00407592, 0.00377297, 5.25379e-05, 0.03164453, 0.05894441, 0.03914395, 
    0.08088186, 0.06648228, 0.07095776, 0.0590079, 0.03939104, 0.07799046, 
    0.1943945, 0.06664231, 0.03770012, 0.03785838, 0.039281, 0.04844719, 
    0.03576902, 0.05329755, 0.1156868, 0.1213445, 0.000106424, 0.00814472, 
    0.0005613167, 6.07254e-09, 0.0719808, 0.1151381, 0.05650128,
  0.08040487, 0.1768032, 0.04824834, 0.04132451, 0.03174422, 0.04777652, 
    0.02904631, 0.04818639, 0.03736554, 0.214661, 0.03005955, 0.02728298, 
    0.03052335, 0.02795962, 0.06722488, 0.01297762, 0.01546329, 0.0133743, 
    0.02000115, 0.04409166, 0.04379128, 0.001928254, 0.0003949394, 
    0.04290821, 0.003073467, 0.008841122, 0.03872241, 0.02955981, 0.04151357,
  0.03620253, 0.0599573, 0.0184453, 0.1073407, -9.69944e-06, 0.01370122, 
    0.05503879, 0.03681378, 0.01734454, 0.03032429, 0.01975237, 0.03956924, 
    0.02981513, 0.02843011, 0.03325088, 0.04792331, 0.09218582, 0.1320604, 
    0.2190544, 0.2179568, 0.1242042, 0.08362809, 0.1494317, 0.05292007, 
    0.03902401, 0.04067571, 0.0672603, 0.05045455, 0.1007715,
  -1.430967e-07, 1.223339e-07, -1.846123e-05, 0.00039179, -2.743633e-07, 
    0.001046218, 0.03343014, 0.08870486, 0.280604, 0.1083854, 0.09145373, 
    0.05328107, 0.03486986, 0.02962056, 0.03606514, 0.0383477, 0.07187794, 
    0.146911, 0.1908986, 0.1787338, 0.05054569, 0.219087, 0.03490217, 
    0.02306124, 0.06466612, 0.06812293, 0.0425726, 9.9594e-05, 2.240634e-05,
  8.135775e-07, 6.172392e-07, 6.455924e-05, 6.971182e-08, -4.572697e-09, 
    -2.309531e-11, -0.0002074249, 0.1812234, 0.4726347, 0.09097728, 
    0.08081472, 0.08836111, 0.03440847, 0.03637258, 0.1046411, 0.0871539, 
    0.1010334, 0.1193379, 0.2965296, -8.848009e-06, 0.01167966, 0.03345157, 
    0.06897461, 0.06127387, 0.0338925, 0.05981185, 0.07563483, 0.1544109, 
    0.001043369,
  0.01043394, 0.02102758, 0.001240227, 0.1099952, 0.001457952, 5.075647e-07, 
    0.05722196, -0.0002435802, 0.0003339482, 0.04532952, 0.1021946, 
    0.1223649, 0.1982961, 0.2168994, 0.2342019, 0.3328447, 0.3226025, 
    0.2804579, 0.1060034, -2.570621e-05, 0.01146779, 0.01508374, 0.0789519, 
    0.1283314, 0.1528009, 0.160899, 0.1776096, 0.2244416, 0.07409423,
  0.1574741, 0.1892459, 0.1054093, 0.08473093, 0.0343331, 0.04905848, 
    0.08156396, 0.1861303, 0.08077233, 0.1457454, 0.1272122, 0.1878205, 
    0.2014828, 0.2392265, 0.3251772, 0.2643621, 0.2507632, 0.2945868, 
    0.3261979, 0.1694139, 0.08499553, 0.06452664, 0.2264907, 0.3599196, 
    0.2056893, 0.2008413, 0.3074515, 0.2780381, 0.169903,
  0.2946238, 0.2383115, 0.2254474, 0.2510526, 0.3121091, 0.2190577, 
    0.1562705, 0.1615171, 0.1494913, 0.2969541, 0.2748616, 0.3307357, 
    0.3379728, 0.4284784, 0.4267826, 0.4478391, 0.3598983, 0.3750978, 
    0.2499956, 0.1581782, 0.2470569, 0.3284573, 0.4432566, 0.4377921, 
    0.4019381, 0.1556942, 0.3547899, 0.2337012, 0.3689635,
  0.4581095, 0.3700868, 0.3490402, 0.4523157, 0.4653219, 0.2490733, 
    0.2698511, 0.192431, 0.1819676, 0.4020588, 0.4330642, 0.4317448, 
    0.3972999, 0.4448601, 0.4173881, 0.3334342, 0.3106656, 0.3758415, 
    0.4049458, 0.4492811, 0.3832651, 0.4046016, 0.4361414, 0.4642161, 
    0.4075064, 0.3844916, 0.2442994, 0.2308061, 0.4409229,
  0.2939896, 0.3093304, 0.2863096, 0.2648871, 0.2633431, 0.3283283, 
    0.3379484, 0.3325352, 0.3339479, 0.3593763, 0.3888218, 0.3701375, 
    0.4087505, 0.5100312, 0.4650306, 0.5436209, 0.4216835, 0.4051633, 
    0.5311138, 0.5343727, 0.4062364, 0.3568178, 0.367343, 0.2860811, 
    0.2246675, 0.3042181, 0.2124405, 0.2243173, 0.3197888,
  0.1769939, 0.1683514, 0.1597088, 0.1510663, 0.1424238, 0.1337813, 
    0.1251387, 0.1367756, 0.1443138, 0.151852, 0.1593902, 0.1669284, 
    0.1744666, 0.1820048, 0.2011254, 0.2116886, 0.2222519, 0.2328152, 
    0.2433784, 0.2539417, 0.264505, 0.2513355, 0.2418765, 0.2324176, 
    0.2229586, 0.2134997, 0.2040407, 0.1945817, 0.1839079,
  0.2709692, 0.2048606, 0.08718245, 0.04682407, 0.006832914, -0.002083171, 
    0.0008083291, 0.008532166, 0.003760719, 0.008008083, 0.03137816, 
    0.1147099, 0.1003208, 0.06301719, 0.09933925, 0.1368201, 0.2794501, 
    0.4795203, 0.4331973, 0.3102197, 0.3971698, 0.4074228, 0.3496194, 
    0.3871045, 0.3194788, 0.2568716, 0.2343201, 0.2104316, 0.2896751,
  0.206956, 0.1254877, 0.2180273, 0.1867498, 0.2267101, 0.1140011, 
    0.05249501, 0.2394705, 0.3433881, 0.4079851, 0.3596981, 0.2393182, 
    0.2014238, 0.2679214, 0.358533, 0.2994851, 0.2635975, 0.2897434, 
    0.3101231, 0.3213541, 0.3003851, 0.3169717, 0.3445542, 0.4801241, 
    0.2241509, 0.2451175, 0.3198145, 0.3200276, 0.3025771,
  0.3304856, 0.3203914, 0.4976746, 0.3546766, 0.3319938, 0.3893563, 
    0.3640315, 0.3804782, 0.3681886, 0.3502494, 0.2615631, 0.3137259, 
    0.3591446, 0.3302401, 0.2708112, 0.365585, 0.405055, 0.5088868, 
    0.5295823, 0.3926065, 0.3303169, 0.2529984, 0.3145931, 0.2728069, 
    0.3581426, 0.36849, 0.4412068, 0.4333045, 0.3805476,
  0.3815507, 0.346741, 0.3086114, 0.3476048, 0.3515756, 0.3146468, 0.3007096, 
    0.2384919, 0.224223, 0.2663761, 0.277835, 0.2524365, 0.2089132, 
    0.1529396, 0.2572274, 0.2752566, 0.2990109, 0.3841646, 0.3744034, 
    0.4037545, 0.2912012, 0.3149019, 0.3076998, 0.2472011, 0.2422039, 
    0.275508, 0.4100983, 0.4078, 0.4089667,
  0.2211805, 0.1548791, 0.1459289, 0.213236, 0.2623112, 0.2473563, 0.1910358, 
    0.2200834, 0.25269, 0.2639386, 0.1867111, 0.08042394, 0.03147722, 
    0.1918235, 0.3417184, 0.1792322, 0.1600145, 0.2126303, 0.249395, 
    0.2077446, 0.1539885, 0.1132059, 0.1536665, 0.3724274, 0.04700146, 
    0.0967976, 0.1986301, 0.2809609, 0.3175092,
  0.2100817, 0.1108808, 0.001722048, 0.1065306, 0.1346427, 0.2321327, 
    0.2676567, 0.1394482, 0.1606991, 0.05453586, 0.001254225, 1.858382e-07, 
    0.009941881, 0.1704058, 0.1685904, 0.1192787, 0.1335479, 0.2628016, 
    0.1395525, 0.09390806, 0.1618882, 0.144152, 0.276512, 0.01474188, 
    0.02832489, 0.134043, 0.2021993, 0.2091629, 0.2493885,
  0.4353931, -5.120293e-05, -2.514805e-05, 0.05984955, 0.03562203, 
    0.02326316, 0.04954963, 0.09368052, 0.225308, 0.002294203, 4.245305e-09, 
    1.192548e-09, 0.03470473, 0.1583494, 0.1222445, 0.04225844, 0.06303574, 
    0.09103943, 0.0292819, 0.02249445, 0.1365288, 0.2466199, 0.5192481, 
    -0.0001708294, 0.006054765, 0.002543918, 0.07302498, 0.1511264, 0.3037639,
  0.1272427, 0.03775164, 2.843015e-05, 0.0246781, 0.05306284, 0.04733373, 
    0.07119409, 0.0485867, 0.08135885, 0.04432585, 0.03710325, 0.05755077, 
    0.1967345, 0.07928858, 0.05135774, 0.0366613, 0.05195577, 0.0355731, 
    0.03238244, 0.02979322, 0.1076596, 0.4053147, 0.04026021, 0.003033384, 
    0.0002088945, 2.999132e-09, 0.06715357, 0.1731525, 0.5134017,
  0.1576495, 0.1653083, 0.04828524, 0.05678992, 0.0464328, 0.07275484, 
    0.03527706, 0.05187188, 0.02824134, 0.1684339, 0.05494427, 0.1088827, 
    0.07727784, 0.07094152, 0.05211741, 0.06904844, 0.0457326, 0.01585463, 
    0.02847772, 0.02639362, 0.09487272, 0.02488595, 9.745151e-05, 0.01637707, 
    0.00108219, 0.05044534, 0.06640527, 0.09064192, 0.1482647,
  0.02339356, 0.04961086, 0.01211967, 0.08896594, 3.593587e-06, 0.02550614, 
    0.05591941, 0.04173797, 0.0163607, 0.03865594, 0.01629991, 0.1096809, 
    0.04803324, 0.05893281, 0.04230573, 0.09681944, 0.1158846, 0.173228, 
    0.1955955, 0.1886847, 0.1224107, 0.09944712, 0.1374347, 0.04421819, 
    0.05090957, 0.07282992, 0.08603735, 0.06537707, 0.07503749,
  -3.69665e-08, 8.935684e-08, -5.719379e-06, 0.001072768, -1.36714e-07, 
    0.03242565, 0.0184057, 0.08106496, 0.2255426, 0.1062609, 0.08380388, 
    0.05214364, 0.05438342, 0.0367066, 0.06852809, 0.04163893, 0.01837109, 
    0.09913608, 0.3787131, 0.1814733, 0.04352421, 0.2233013, 0.0896375, 
    0.0154856, 0.05101946, 0.1244498, 0.1427134, 0.0482625, 1.425929e-05,
  6.382444e-07, -4.977726e-07, 0.0004905873, 6.014317e-08, -3.728261e-09, 
    -1.847424e-11, -0.0002585443, 0.1871978, 0.4752476, 0.0644649, 0.1189078, 
    0.06976204, 0.06156262, 0.05269416, 0.1222606, 0.07112834, 0.09588251, 
    0.1048115, 0.2521158, -0.000241792, 0.006898972, 0.04604946, 0.06680182, 
    0.06911419, 0.05546105, 0.115033, 0.1473487, 0.1979498, 0.003234633,
  0.008308296, 0.01088204, 0.0007970331, 0.1374166, -0.0001351638, 
    1.056057e-07, 0.05419903, -7.8276e-05, -2.757226e-05, 0.03540642, 
    0.1077981, 0.132671, 0.225788, 0.2352268, 0.2387818, 0.3395599, 
    0.2784823, 0.3560512, 0.2535674, -0.0002933783, 0.003077209, 0.0126455, 
    0.07724778, 0.1052136, 0.1448225, 0.132411, 0.1770377, 0.191938, 0.0640585,
  0.1512838, 0.1883568, 0.1019585, 0.1204627, 0.02405337, 0.03220119, 
    0.06479028, 0.1911477, 0.06990301, 0.1429186, 0.1086695, 0.1744246, 
    0.2011542, 0.2618784, 0.2699456, 0.2690237, 0.2579178, 0.3385993, 
    0.3526078, 0.1578384, 0.07277445, 0.05259613, 0.1879742, 0.3553158, 
    0.2115093, 0.197757, 0.3061194, 0.2512805, 0.1316994,
  0.2337158, 0.2200069, 0.1907329, 0.2434518, 0.3000402, 0.1979067, 
    0.1620542, 0.1606784, 0.155371, 0.2935757, 0.2636222, 0.3643886, 
    0.3482319, 0.3971318, 0.4594614, 0.3782218, 0.3420652, 0.3646409, 
    0.2530638, 0.1564132, 0.2036559, 0.3067963, 0.2830062, 0.3650174, 
    0.3755399, 0.1404438, 0.2983708, 0.1984126, 0.3115785,
  0.5962761, 0.3755931, 0.3463587, 0.5752741, 0.4855492, 0.2932017, 
    0.2353511, 0.1729471, 0.2009636, 0.3113578, 0.4364478, 0.4453125, 
    0.4054301, 0.5604641, 0.4361745, 0.481178, 0.3535421, 0.426515, 
    0.3794854, 0.4463367, 0.3685122, 0.3902568, 0.4451764, 0.5003735, 
    0.4625798, 0.3738841, 0.2509699, 0.2848434, 0.4794127,
  0.3720137, 0.4757876, 0.3898276, 0.3391753, 0.3352623, 0.4028652, 0.432453, 
    0.4059367, 0.3492184, 0.4446717, 0.3774858, 0.3910284, 0.4098399, 
    0.4543129, 0.4794863, 0.5456902, 0.4210495, 0.5808713, 0.6324966, 
    0.5820041, 0.5870055, 0.3651448, 0.3767307, 0.3552192, 0.189589, 
    0.2827783, 0.1822841, 0.2253862, 0.3963511,
  0.1627824, 0.1533676, 0.1439529, 0.1345382, 0.1251235, 0.1157087, 0.106294, 
    0.1304793, 0.1386651, 0.146851, 0.1550368, 0.1632227, 0.1714085, 
    0.1795943, 0.1851411, 0.1950824, 0.2050237, 0.2149651, 0.2249064, 
    0.2348477, 0.244789, 0.2656464, 0.256934, 0.2482215, 0.2395091, 
    0.2307966, 0.2220842, 0.2133718, 0.1703141,
  0.3283429, 0.2398203, 0.1058186, 0.04966273, 0.006558859, -0.002009208, 
    -0.0004150847, 0.008717002, 0.002959435, 0.006225948, 0.02042871, 
    0.1269219, 0.1159121, 0.05338767, 0.09307045, 0.1326111, 0.2784851, 
    0.4278746, 0.3613546, 0.3137907, 0.3894423, 0.4065027, 0.3405014, 
    0.3659488, 0.3256717, 0.2702493, 0.1719903, 0.165869, 0.3147298,
  0.2164862, 0.1015814, 0.208961, 0.1200723, 0.2066663, 0.07758128, 
    0.02429113, 0.2460132, 0.3400637, 0.4043109, 0.3943339, 0.2112236, 
    0.1912141, 0.2487142, 0.3648778, 0.3340838, 0.303273, 0.3419226, 
    0.382122, 0.4117605, 0.3491449, 0.3429543, 0.3433538, 0.5212136, 
    0.2225211, 0.2490063, 0.3392973, 0.3723908, 0.3538012,
  0.4004233, 0.3298449, 0.4896056, 0.25818, 0.2456775, 0.353556, 0.3715201, 
    0.3733604, 0.387462, 0.2595669, 0.2261702, 0.3026718, 0.309734, 
    0.3435777, 0.2721914, 0.3983272, 0.4166132, 0.475961, 0.4934829, 
    0.3376491, 0.2653794, 0.2217465, 0.3021848, 0.1978337, 0.2780954, 
    0.404807, 0.4809428, 0.4678794, 0.3910112,
  0.3311986, 0.285327, 0.2756368, 0.2998655, 0.3115507, 0.3102811, 0.3041313, 
    0.2166959, 0.2056553, 0.2484614, 0.2717847, 0.2443065, 0.1564154, 
    0.1187744, 0.1996092, 0.2409839, 0.2253548, 0.3456664, 0.3560572, 
    0.3556164, 0.2530479, 0.3233478, 0.2649438, 0.2220829, 0.2050528, 
    0.2789737, 0.3664537, 0.3678867, 0.3640393,
  0.1998958, 0.1021236, 0.1253385, 0.2299664, 0.2554195, 0.2426822, 
    0.2099584, 0.2078912, 0.2128205, 0.1855164, 0.1610192, 0.05439158, 
    0.01081093, 0.1564473, 0.3027465, 0.1504287, 0.1370358, 0.179855, 
    0.2347929, 0.1614289, 0.1115061, 0.1048384, 0.102511, 0.3772224, 
    0.02992706, 0.08153404, 0.201321, 0.2239038, 0.2532693,
  0.117687, 0.07989078, 0.00189848, 0.05948839, 0.1060015, 0.2001034, 
    0.11022, 0.1166396, 0.1106121, 0.02466571, 0.000947236, -7.980255e-06, 
    0.008428925, 0.1390566, 0.130803, 0.09924068, 0.1456212, 0.2526169, 
    0.1354872, 0.08279537, 0.07947821, 0.0671906, 0.1578875, 0.01224665, 
    0.02825618, 0.1855478, 0.1707938, 0.1450598, 0.1095859,
  0.3345087, -0.0002656644, -7.587568e-05, 0.0821063, -0.002603142, 
    0.003176511, 0.009119038, 0.04943436, 0.1348065, 0.0003576444, 
    3.185477e-09, 1.066363e-09, 0.04225637, 0.1504716, 0.121505, 0.08691499, 
    0.06527781, 0.07160179, 0.004380731, 0.002970425, 0.03355701, 0.07142942, 
    0.2471927, 0.01006739, 0.002231105, 0.005366822, 0.02170639, 0.04572253, 
    0.1395729,
  0.6566697, 0.1316046, -1.708616e-05, 0.03841114, 0.03211265, 0.02326031, 
    0.03993452, 0.02490153, 0.02038042, 0.03394534, 0.03341196, 0.03090183, 
    0.1650985, 0.04872176, 0.03093785, 0.01699447, 0.01793901, 0.009524745, 
    0.009029486, 0.005943655, 0.03343786, 0.2320622, 0.3229898, 0.001024594, 
    8.242355e-05, 2.157991e-09, 0.01682282, 0.06297816, 0.2961182,
  0.2227626, 0.1300855, 0.03176198, 0.08419657, 0.1084266, 0.0445328, 
    0.03990171, 0.04795908, 0.02630859, 0.1325421, 0.07368372, 0.08214068, 
    0.02108624, 0.009378982, 0.006553534, 0.02154696, 0.03534498, 0.01369765, 
    0.01977187, 0.02033466, 0.1079186, 0.2192797, 0.007893268, 0.006226044, 
    0.0004576931, 0.04816216, 0.02315443, 0.06039965, 0.2313906,
  0.02199833, 0.04455578, 0.007976329, 0.07253775, -2.23556e-05, 0.01651301, 
    0.06392604, 0.0154927, 0.007400974, 0.02347705, 0.007247198, 0.07036366, 
    0.02455568, 0.03545435, 0.04731011, 0.0625922, 0.08399506, 0.1291327, 
    0.1929165, 0.1710203, 0.0853347, 0.1022155, 0.1302323, 0.03177051, 
    0.01530876, 0.06379984, 0.07866678, 0.09712671, 0.05544246,
  -6.803482e-09, 7.147256e-08, -2.478297e-06, 0.0007631115, -8.638479e-08, 
    0.1153546, 0.007338321, 0.060241, 0.1662616, 0.06488705, 0.05799856, 
    0.03536989, 0.01843883, 0.01894801, 0.01202441, 0.009801448, 0.001952413, 
    0.02391888, 0.238748, 0.2805836, 0.1167526, 0.2272006, 0.0142755, 
    0.004303295, 0.01653854, 0.05184696, 0.2582843, 0.05193456, 6.681663e-06,
  5.12526e-07, -1.80581e-06, 0.0008902926, 2.35212e-08, -3.174571e-09, 
    -1.247455e-11, -0.0001711714, 0.1977955, 0.459596, 0.04081022, 0.109162, 
    0.07106198, 0.09725545, 0.08141997, 0.1102694, 0.02862631, 0.02697743, 
    0.05277672, 0.1990636, 0.0949804, 0.009191312, 0.04152598, 0.05136135, 
    0.08801003, 0.03993007, 0.03968807, 0.1037655, 0.2107341, 0.007722893,
  0.007764409, 0.01200942, 0.001267225, 0.1623894, -5.738917e-05, 
    1.380794e-07, 0.05464099, -3.891938e-05, -0.0001048043, 0.03084256, 
    0.1075885, 0.1408056, 0.2531608, 0.2714737, 0.2832913, 0.3575037, 
    0.319885, 0.485438, 0.3447931, -0.0001985881, 0.0007299475, 0.01421877, 
    0.06736746, 0.1011315, 0.120863, 0.09085923, 0.1110763, 0.1105808, 
    0.06600659,
  0.1405039, 0.193321, 0.07823834, 0.09310251, 0.01884537, 0.02321334, 
    0.04985013, 0.1735476, 0.06111899, 0.1276982, 0.09766195, 0.1531581, 
    0.2514925, 0.288965, 0.2153295, 0.247965, 0.3640836, 0.3874159, 
    0.3164511, 0.1527314, 0.06838347, 0.0467851, 0.1586142, 0.3642437, 
    0.2312606, 0.2313852, 0.2874381, 0.2899397, 0.2381084,
  0.227497, 0.2140478, 0.1485918, 0.2136116, 0.2610229, 0.1942424, 0.1402614, 
    0.1650417, 0.1468312, 0.2754752, 0.2949329, 0.4043514, 0.3496628, 
    0.3168833, 0.4350245, 0.2999626, 0.3363222, 0.3262349, 0.2776241, 
    0.1274263, 0.1601704, 0.2450735, 0.1842118, 0.2879336, 0.3070965, 
    0.1415158, 0.2336843, 0.202595, 0.2752084,
  0.5548936, 0.3718927, 0.3762659, 0.5050893, 0.5038002, 0.4559486, 
    0.2901371, 0.1537699, 0.198724, 0.3015185, 0.4568879, 0.3963665, 
    0.3443986, 0.3959266, 0.4110488, 0.5255138, 0.3823013, 0.3410685, 
    0.2652977, 0.2800653, 0.2773463, 0.3322983, 0.4220889, 0.5693249, 
    0.3529633, 0.3483982, 0.2634162, 0.2349583, 0.4407094,
  0.516044, 0.4611923, 0.3716557, 0.4502541, 0.6232545, 0.6009263, 0.5102425, 
    0.5125871, 0.4134673, 0.4787112, 0.4748983, 0.4159659, 0.390334, 
    0.4191258, 0.4492417, 0.457946, 0.5005398, 0.6697321, 0.674874, 
    0.6070851, 0.5257869, 0.3535691, 0.3336369, 0.4136617, 0.2053947, 
    0.2599289, 0.1779601, 0.210715, 0.4171565,
  0.1071833, 0.09966077, 0.09213826, 0.08461574, 0.07709323, 0.06957072, 
    0.0620482, 0.08131493, 0.08782962, 0.09434431, 0.100859, 0.1073737, 
    0.1138884, 0.1204031, 0.1215387, 0.1318093, 0.1420798, 0.1523503, 
    0.1626208, 0.1728913, 0.1831619, 0.220881, 0.2116183, 0.2023556, 
    0.1930929, 0.1838302, 0.1745675, 0.1653048, 0.1132013,
  0.376786, 0.2500581, 0.108879, 0.04858341, 0.008203343, -0.00156629, 
    -0.0009501062, 0.006773934, 0.001677631, 0.00621052, -0.000450193, 
    0.05015385, 0.1621375, 0.03258133, 0.1000492, 0.1529423, 0.2953073, 
    0.3803053, 0.2942122, 0.303974, 0.3887955, 0.3905901, 0.3035333, 
    0.3436016, 0.2904228, 0.2541756, 0.1394766, 0.1300714, 0.3480587,
  0.2050579, 0.08777669, 0.1977443, 0.07130629, 0.1846612, 0.05621444, 
    0.01271388, 0.2543811, 0.3138034, 0.3862553, 0.3882153, 0.2005509, 
    0.186819, 0.2334109, 0.3792098, 0.3899134, 0.3621162, 0.3613284, 
    0.4040295, 0.4288669, 0.3911832, 0.3628666, 0.3715639, 0.5458872, 
    0.1854264, 0.2666951, 0.3840308, 0.4216106, 0.3821778,
  0.4532976, 0.3607229, 0.4157429, 0.2007694, 0.1859258, 0.3331094, 
    0.3690787, 0.358353, 0.4374087, 0.2080903, 0.1921411, 0.2625461, 
    0.2789718, 0.3407941, 0.2700348, 0.3928788, 0.4160706, 0.4141642, 
    0.4272743, 0.2961442, 0.2331138, 0.1883493, 0.2653806, 0.1526884, 
    0.2418977, 0.3869914, 0.4511596, 0.4570873, 0.4376522,
  0.2893733, 0.2730506, 0.257395, 0.2641115, 0.3161264, 0.3109989, 0.2852567, 
    0.1845194, 0.18336, 0.223354, 0.2217361, 0.2103256, 0.1116881, 
    0.09168414, 0.1542136, 0.1976151, 0.1832636, 0.3091955, 0.3202629, 
    0.3197013, 0.2130879, 0.2732998, 0.2186298, 0.1926696, 0.1476842, 
    0.2532709, 0.3257191, 0.327504, 0.3456584,
  0.1435175, 0.05744475, 0.1055908, 0.2228325, 0.3114324, 0.2591526, 
    0.1887854, 0.1627165, 0.1689415, 0.1193568, 0.09568422, 0.03114657, 
    0.004639427, 0.1349951, 0.2560093, 0.1319256, 0.09981222, 0.1370311, 
    0.2064146, 0.1500284, 0.09999492, 0.09020763, 0.06350511, 0.3760928, 
    0.02727393, 0.0778136, 0.1799176, 0.1871881, 0.2070103,
  0.0401798, 0.06165554, 0.001507318, 0.03199954, 0.05773722, 0.05809092, 
    0.03067872, 0.04554814, 0.041822, 0.01139585, 0.000967415, -7.334338e-06, 
    0.004726309, 0.1074243, 0.1131227, 0.09213208, 0.1707719, 0.1925006, 
    0.1427309, 0.03856785, 0.04125284, 0.03403964, 0.04881516, 0.007194397, 
    0.02305757, 0.1727762, 0.1160919, 0.07597697, 0.04439417,
  0.1490793, -0.0002325591, -4.788854e-05, 0.01618676, -0.005013535, 
    4.429885e-05, 0.001997464, 0.01141027, 0.04211195, 0.03668114, 
    2.680132e-09, 1.004201e-09, 0.0125634, 0.1075931, 0.07660772, 0.05722876, 
    0.01853078, 0.03292903, 9.324739e-05, 8.934e-05, 0.009555503, 0.02105277, 
    0.09657203, 0.007488798, 0.0006578356, 0.0107773, 0.005761473, 0.0106791, 
    0.04439323,
  0.3338654, 0.2517762, -2.445974e-05, 0.07404733, 0.01353688, 0.006363459, 
    0.0163635, 0.008945512, 0.003271038, 0.008804336, 0.03043731, 0.01387561, 
    0.1383137, 0.02526538, 0.006695583, 0.004364282, 0.00313465, 
    0.0005970419, 0.000167793, 0.000372068, 0.008274235, 0.07453538, 
    0.271051, 0.0003822142, 6.281838e-05, 3.013844e-09, -0.001385904, 
    0.01584699, 0.1091526,
  0.1126254, 0.115701, 0.02399758, 0.06866293, 0.04734962, 0.01290448, 
    0.006967011, 0.03302392, 0.03409408, 0.09782939, 0.0232187, 0.01388738, 
    0.004936871, 0.00125424, 0.001339198, 0.002855623, 0.007874687, 
    0.005080881, 0.01035066, 0.008354266, 0.04870433, 0.4322486, 0.2625342, 
    0.005786779, 0.0001825912, 0.01039418, 0.003863716, 0.008776238, 0.1140787,
  0.01043118, 0.04032415, 0.00944911, 0.0691168, 9.462381e-05, 0.003984241, 
    0.07405902, 0.002287379, 0.001719405, 0.01151337, 0.002558161, 
    0.02332886, 0.005363793, 0.01467801, 0.01046328, 0.0264516, 0.03865182, 
    0.05469094, 0.1172363, 0.1285311, 0.04139373, 0.04654983, 0.139081, 
    0.02101775, 0.001674107, 0.009611499, 0.02342915, 0.08566321, 0.04112235,
  1.515786e-08, 6.123334e-08, -9.038921e-07, -1.898022e-05, -3.361427e-08, 
    0.1141421, 0.0124649, 0.04147357, 0.1225876, 0.03378896, 0.01363725, 
    0.01451342, 0.005175884, 0.002524293, 0.002282762, 0.001273999, 
    0.0005257457, 0.004795067, 0.08524543, 0.2394238, 0.1132519, 0.1982319, 
    0.002199973, -0.001429288, 0.008104066, 0.01606907, 0.1060211, 
    0.03919309, 3.354936e-06,
  4.4058e-07, -4.394171e-07, 0.001103656, -4.076015e-09, -2.786995e-09, 
    -6.452212e-12, -0.000107033, 0.2186494, 0.4295152, 0.02577658, 0.131733, 
    0.05879422, 0.03631099, 0.01980252, 0.03412485, 0.005002028, 0.009287518, 
    0.01140866, 0.09001593, 0.1803189, 0.006275743, 0.03666794, 0.03236854, 
    0.01907418, 0.007690797, 0.005324461, 0.03397936, 0.06945728, 0.009706294,
  0.006067213, 0.01405108, 0.0008966605, 0.1786521, -0.0006935283, 
    1.413277e-07, 0.05077956, -1.954887e-05, -0.0001143575, 0.03536437, 
    0.1131307, 0.139359, 0.2911339, 0.2251884, 0.2848199, 0.3451349, 
    0.4400224, 0.3860143, 0.2391516, -0.0001872423, 0.000227492, 0.01752603, 
    0.05743454, 0.1913331, 0.1106031, 0.06773193, 0.06388123, 0.055458, 
    0.08234094,
  0.1165296, 0.1906086, 0.07713931, 0.07228025, 0.009456499, 0.02304226, 
    0.04510289, 0.1585986, 0.04984926, 0.1249497, 0.08531275, 0.1318238, 
    0.2837071, 0.2765419, 0.191469, 0.2325971, 0.3283311, 0.3708577, 
    0.2686975, 0.14974, 0.06242053, 0.03927083, 0.1465424, 0.3546459, 
    0.231022, 0.2152899, 0.2432119, 0.2749272, 0.248442,
  0.1822082, 0.1865852, 0.1231004, 0.1895229, 0.2457983, 0.1886553, 
    0.1292096, 0.1642596, 0.1595416, 0.2697184, 0.2826131, 0.4867558, 
    0.3595545, 0.2463436, 0.323202, 0.243059, 0.3391978, 0.3091789, 
    0.2721076, 0.1045348, 0.1167016, 0.2175068, 0.146411, 0.25352, 0.2884328, 
    0.1416021, 0.1719816, 0.1889522, 0.250982,
  0.4408545, 0.285698, 0.4285069, 0.4082269, 0.518561, 0.4184025, 0.2982705, 
    0.1382513, 0.1668213, 0.2898064, 0.4608445, 0.3093411, 0.2745626, 
    0.291315, 0.3981331, 0.4614066, 0.3063945, 0.2254501, 0.1825158, 
    0.1975631, 0.2000637, 0.2729875, 0.3668205, 0.5639579, 0.2612004, 
    0.3210898, 0.2813911, 0.1683582, 0.3786636,
  0.5019649, 0.3509988, 0.3417594, 0.5301498, 0.6213882, 0.4944558, 
    0.4467674, 0.4633129, 0.3476168, 0.4485941, 0.5073003, 0.4870974, 
    0.3745873, 0.3924603, 0.4087968, 0.4763803, 0.558163, 0.6280761, 
    0.6534455, 0.5910249, 0.4519307, 0.3151381, 0.3157205, 0.4099686, 
    0.2250774, 0.227114, 0.1660449, 0.2495571, 0.321776,
  0.03902563, 0.03444779, 0.02986995, 0.02529211, 0.02071427, 0.01613643, 
    0.01155859, 0.007268183, 0.01094732, 0.01462646, 0.0183056, 0.02198473, 
    0.02566387, 0.02934301, 0.02826621, 0.03537732, 0.04248843, 0.04959954, 
    0.05671065, 0.06382176, 0.07093286, 0.09519928, 0.08898687, 0.08277447, 
    0.07656206, 0.07034966, 0.06413725, 0.05792485, 0.0426879,
  0.3743533, 0.2554266, 0.07068674, 0.04296578, 0.01176426, -0.001063608, 
    -0.0004101217, 0.002774992, 0, 4.322697e-08, 0.0003100704, 0.004178217, 
    0.09437196, 0.02069548, 0.09876377, 0.1636771, 0.3106797, 0.3473177, 
    0.2591503, 0.2829072, 0.3999667, 0.3898751, 0.2673358, 0.3015658, 
    0.2846472, 0.2715274, 0.1235612, 0.1003396, 0.3498499,
  0.2079294, 0.05854652, 0.1858455, 0.04618436, 0.1365521, 0.04734992, 
    0.007593418, 0.2484554, 0.2740844, 0.3610884, 0.3686335, 0.1889289, 
    0.1790931, 0.2110733, 0.3806112, 0.3982924, 0.3672453, 0.3684395, 
    0.3948084, 0.4132564, 0.402675, 0.3471712, 0.3731859, 0.5616183, 
    0.1612624, 0.2918908, 0.4413913, 0.4583928, 0.3857821,
  0.4607058, 0.3801884, 0.3587768, 0.1412958, 0.1441917, 0.2931004, 
    0.3582031, 0.3417588, 0.4436844, 0.1665449, 0.1538751, 0.2112226, 
    0.2574953, 0.2998883, 0.2349366, 0.3626872, 0.3778323, 0.4151976, 
    0.3463516, 0.2413986, 0.1867117, 0.1506468, 0.2197734, 0.1292185, 
    0.1904445, 0.3412109, 0.3944959, 0.4101813, 0.4422119,
  0.2531416, 0.2654851, 0.2297752, 0.2352923, 0.3207599, 0.2957677, 0.251272, 
    0.154199, 0.1518168, 0.1739017, 0.1608201, 0.1483674, 0.08006571, 
    0.08672587, 0.1192933, 0.1508294, 0.1538935, 0.2746782, 0.2837679, 
    0.2786584, 0.1851519, 0.2213029, 0.1730926, 0.1502339, 0.1137564, 
    0.2082216, 0.2745337, 0.288844, 0.2937009,
  0.08636735, 0.02758659, 0.07984145, 0.2063917, 0.3041397, 0.2359676, 
    0.1320667, 0.1037354, 0.1093704, 0.07726787, 0.06852756, 0.01176832, 
    0.001735589, 0.130704, 0.1957016, 0.09480333, 0.06300317, 0.1078541, 
    0.1730717, 0.1329678, 0.0943809, 0.06086583, 0.04213547, 0.3488035, 
    0.02629333, 0.08024866, 0.1500771, 0.1528927, 0.1811743,
  0.01563308, 0.03375869, 0.0006454607, 0.01881297, 0.03432137, 0.02150126, 
    0.01292242, 0.01691279, 0.01827264, 0.006219178, 0.0003131763, 
    -2.426943e-06, 0.002743773, 0.07550274, 0.09663888, 0.06894597, 
    0.1201096, 0.1462334, 0.1299466, 0.02233634, 0.01996366, 0.01906324, 
    0.01948651, 0.004934036, 0.01577268, 0.1272664, 0.06138196, 0.04414026, 
    0.01859309,
  0.06803046, 0.003896046, -2.304386e-05, 0.005847496, -0.00323247, 
    -4.481341e-06, 0.0008596667, 0.004069531, 0.01833054, 0.03005102, 
    2.548936e-09, 8.112008e-10, 0.003882108, 0.06423672, 0.03909357, 
    0.01861708, 0.00421316, 0.01196735, 1.21171e-05, 1.669684e-05, 
    0.004007128, 0.008630028, 0.04269059, 0.002478987, 0.000232376, 
    0.01928765, 0.0006852811, 0.004187872, 0.01561665,
  0.1526489, 0.1875226, -1.10571e-05, 0.102045, 0.004599625, 0.001174689, 
    0.005842085, 0.00200212, 0.001321584, -0.0004862093, 0.02295758, 
    0.005519901, 0.08251915, 0.005494458, 0.0007049447, 0.001092137, 
    0.0007285844, 7.716962e-05, 3.391463e-05, 0.0001439589, 0.003156315, 
    0.02666608, 0.1240693, 0.0001314461, 4.268125e-05, 2.770724e-09, 
    -0.0008321773, 0.006876248, 0.03896581,
  0.02988976, 0.1153478, 0.01849927, 0.0536918, 0.01113303, 0.00459603, 
    0.0008131607, 0.01685274, 0.05446725, 0.08868192, 0.00296735, 0.00277788, 
    0.0004451519, 0.0003480251, 0.0004487283, 0.0008863567, 0.0008676705, 
    0.0001823107, 0.0009957009, 0.0002377757, 0.008551643, 0.192164, 
    0.1519393, 0.003401942, 9.436563e-05, 0.003742176, 0.0005791213, 
    0.002195285, 0.03666733,
  0.006393651, 0.03717532, 0.005090754, 0.07293997, 0.0001093621, 
    0.0002638881, 0.07928658, 0.0001112334, -0.000182524, 0.003210509, 
    0.0002988458, 0.009790001, 0.001982248, 0.003664267, 0.002239091, 
    0.01256731, 0.01483286, 0.0358611, 0.0738427, 0.07207111, 0.02126611, 
    0.01613147, 0.1452657, 0.02101539, 0.0002419444, 0.002019048, 
    0.006739485, 0.02497184, 0.04062102,
  2.302525e-08, 5.497796e-08, -2.842321e-07, -3.244838e-05, -5.97538e-09, 
    0.03843379, 0.01412807, 0.01699277, 0.1016805, 0.01871827, 0.00492778, 
    0.004198453, 0.0004575359, 0.0002411043, 0.0006027832, 0.0002069616, 
    0.0002552751, 0.001674788, 0.03226627, 0.1430264, 0.02641182, 0.1481608, 
    0.0007244023, -0.001357579, 0.001780542, 0.005158043, 0.03935984, 
    0.02378105, 1.169822e-06,
  3.865432e-07, -8.389028e-08, 0.0008215257, -1.731301e-07, -2.512672e-09, 
    -2.552849e-12, -4.572381e-05, 0.2239306, 0.4020128, 0.01264483, 
    0.1023089, 0.0170732, 0.00652356, 0.003139872, 0.0145418, 0.001371108, 
    0.003054444, 0.003445065, 0.03509464, 0.3412298, 0.004716374, 0.03350693, 
    0.02320577, 0.006556605, 0.002117232, 0.001694628, 0.01061542, 
    0.02784757, 0.01165869,
  0.005422704, 0.006264664, 0.0007275678, 0.1921651, -0.0006707797, 
    1.259491e-07, 0.05009093, -1.067063e-05, -0.000118013, 0.03384661, 
    0.1148848, 0.1189468, 0.2616117, 0.1564682, 0.2239337, 0.3123583, 
    0.3839548, 0.2301962, 0.1217217, -0.0004194719, -0.0001072203, 
    0.01564086, 0.04816553, 0.215771, 0.07382898, 0.04445662, 0.03156888, 
    0.0251844, 0.04703708,
  0.1112779, 0.1858965, 0.06472179, 0.06642793, 0.005450625, 0.01816199, 
    0.03540243, 0.1485992, 0.04482795, 0.1169122, 0.07511751, 0.116416, 
    0.3021788, 0.2568784, 0.1554403, 0.2170979, 0.2398961, 0.2993101, 
    0.2379196, 0.1412956, 0.05198733, 0.03048917, 0.1309188, 0.3358182, 
    0.2219183, 0.2025488, 0.2164576, 0.1993369, 0.1471898,
  0.1445996, 0.1679891, 0.102869, 0.1686244, 0.2431676, 0.1660069, 0.1081128, 
    0.1471468, 0.1443687, 0.2749631, 0.2479581, 0.5148211, 0.3721544, 
    0.1924167, 0.2229656, 0.2003016, 0.3333714, 0.2919663, 0.2472277, 
    0.09344645, 0.0944268, 0.218584, 0.1346645, 0.2260523, 0.2226256, 
    0.1348556, 0.1388598, 0.1451352, 0.2295698,
  0.3747641, 0.1994705, 0.411213, 0.379921, 0.4757541, 0.3984627, 0.2798426, 
    0.122352, 0.1376154, 0.3227793, 0.4455402, 0.2891106, 0.2315361, 
    0.2172782, 0.3799407, 0.3968136, 0.2351199, 0.1635815, 0.1443317, 
    0.1383326, 0.151627, 0.2373375, 0.346527, 0.5298992, 0.1926695, 
    0.2882898, 0.2757225, 0.1394832, 0.3290235,
  0.3994712, 0.2602627, 0.2776151, 0.5238792, 0.5345031, 0.4247889, 
    0.3823933, 0.4453475, 0.4019013, 0.4220996, 0.4617663, 0.4213852, 
    0.3503832, 0.3936303, 0.3781984, 0.4615545, 0.5781999, 0.5375566, 
    0.6052253, 0.5378357, 0.3811573, 0.2947503, 0.2882873, 0.440109, 
    0.2256171, 0.191379, 0.1393496, 0.2666414, 0.2604823,
  0.0139429, 0.01239912, 0.01085534, 0.009311559, 0.007767776, 0.006223995, 
    0.004680214, 0.003103154, 0.003904388, 0.004705622, 0.005506855, 
    0.006308089, 0.007109323, 0.007910557, -0.005517403, -0.003404077, 
    -0.001290751, 0.0008225752, 0.002935901, 0.005049227, 0.007162553, 
    0.01520381, 0.01383303, 0.01246225, 0.01109148, 0.009720699, 0.008349921, 
    0.006979142, 0.01517793,
  0.3576486, 0.1941382, 0.05037564, 0.03553027, 0.01256274, -0.0003693032, 
    0.000369646, -1.183333e-05, 0, 0, 0.0001886849, 0.0002562384, 0.04003898, 
    0.01537835, 0.1273077, 0.220227, 0.4003574, 0.3127176, 0.2153338, 
    0.259621, 0.4160917, 0.3728743, 0.2116871, 0.2161072, 0.3096504, 
    0.3532621, 0.1574726, 0.06778955, 0.3315965,
  0.2335092, 0.06036537, 0.1660816, 0.02717229, 0.0925056, 0.03025878, 
    0.005354778, 0.2121627, 0.2187839, 0.2796257, 0.3153344, 0.1627791, 
    0.1716361, 0.1766937, 0.4053934, 0.3624079, 0.3319769, 0.348407, 
    0.3643908, 0.3698371, 0.3868639, 0.3184499, 0.3328719, 0.5472578, 
    0.1464648, 0.3396728, 0.478958, 0.4494811, 0.3991836,
  0.4051651, 0.3686641, 0.2859069, 0.1011413, 0.1037275, 0.2234954, 
    0.3105081, 0.289959, 0.3555326, 0.1215709, 0.1136464, 0.164046, 
    0.2175711, 0.2347166, 0.1868396, 0.3140136, 0.3372697, 0.3619724, 
    0.2612751, 0.1862101, 0.1471916, 0.1207511, 0.1646986, 0.1038258, 
    0.1484154, 0.2739754, 0.3481253, 0.3591714, 0.3997738,
  0.2151961, 0.2230945, 0.18926, 0.1907298, 0.2808014, 0.2471411, 0.214833, 
    0.1222119, 0.1163738, 0.1312736, 0.1134681, 0.10571, 0.05218265, 
    0.06413941, 0.1034041, 0.1075186, 0.1053567, 0.2354083, 0.2004799, 
    0.1934711, 0.150383, 0.1674422, 0.1234485, 0.1140532, 0.09008657, 
    0.1550007, 0.1960395, 0.2415234, 0.2357297,
  0.05473449, 0.01208654, 0.05466366, 0.1659021, 0.2384114, 0.1720271, 
    0.08314568, 0.04842003, 0.05807048, 0.04962969, 0.0357185, 0.004516731, 
    0.0008125997, 0.1035312, 0.1404628, 0.06560028, 0.03404408, 0.0791771, 
    0.1276117, 0.09834651, 0.07546798, 0.03808068, 0.02708143, 0.3119815, 
    0.02592773, 0.07504171, 0.1209194, 0.1154051, 0.1479628,
  0.008462261, 0.01999993, 0.001660665, 0.008130322, 0.01563449, 0.01244605, 
    0.008151026, 0.009807062, 0.01005756, 0.003604457, 0.0002115794, 
    -1.023838e-06, 0.002350944, 0.06110956, 0.06499438, 0.05072258, 
    0.05115118, 0.1132645, 0.09072519, 0.0108735, 0.01066199, 0.00931114, 
    0.01145849, 0.003870622, 0.02003362, 0.07600799, 0.03551513, 0.02165359, 
    0.01025892,
  0.03737497, 0.01127854, -1.0078e-05, 0.003259304, -0.002452424, 
    -3.860705e-06, 0.0004759339, 0.002306079, 0.0104272, 0.01352051, 
    2.241585e-09, 8.049694e-10, 0.001885224, 0.03412242, 0.01627923, 
    0.005129841, 0.001728842, 0.002732452, 2.323838e-06, 7.731696e-06, 
    0.002171017, 0.004677684, 0.02357549, 0.0007218699, 0.0001014108, 
    0.02750301, 0.0003378379, 0.002231671, 0.007371108,
  0.07930963, 0.09054422, -3.28854e-06, 0.07781829, 0.001076845, 
    0.0002285007, 0.00170157, 0.0003643224, 0.0007372515, -0.002938048, 
    0.01576157, 0.001987767, 0.03955892, 0.001453565, 5.785219e-05, 
    0.0003351354, 0.0002689375, 3.722776e-05, 1.226889e-05, 7.517132e-05, 
    0.001632362, 0.01321394, 0.06634095, 4.976116e-05, 2.258371e-05, 
    2.573917e-09, -0.0003239097, 0.003941364, 0.01870758,
  0.0141279, 0.1209385, 0.01567256, 0.03679582, 0.002214077, 0.001528232, 
    0.0001906054, 0.008610872, 0.04840546, 0.09508356, 0.0009831309, 
    0.001170237, 0.0001198134, 0.0001731093, 0.0002368339, 0.0004422221, 
    0.0003825508, 4.291575e-05, 0.0003254822, 7.115714e-05, 0.003511856, 
    0.07465459, 0.0835043, 0.001778637, 3.15574e-05, 0.001934311, 
    0.0002739039, 0.001057664, 0.01558763,
  0.006588286, 0.02924228, 0.003293254, 0.0704538, 3.799808e-05, 
    0.0001179761, 0.05178648, 3.136122e-05, -0.0007786829, 0.001018448, 
    5.630827e-05, 0.006184647, 0.0006476337, 0.001069786, 0.0008392367, 
    0.006670709, 0.006177826, 0.02729012, 0.04676232, 0.03538409, 
    0.008203685, 0.004489123, 0.131013, 0.02254349, 0.0001243957, 
    0.0008345933, 0.003491104, 0.00815436, 0.03555949,
  2.28332e-08, 5.118512e-08, 1.68293e-09, -2.174529e-05, 1.067561e-09, 
    0.0227705, 0.009893697, 0.005379069, 0.0865983, 0.006455512, 0.001102657, 
    0.001386247, 7.495435e-05, 4.516183e-05, 0.0002576026, 0.0001000849, 
    0.0001537017, 0.000817752, 0.01595824, 0.09246057, 0.008442727, 
    0.1147387, 0.0004093087, -0.000956991, 0.0003335119, 0.002426735, 
    0.0183421, 0.006546583, 4.872019e-07,
  3.451158e-07, -2.560724e-09, 0.002394087, -5.66037e-07, -2.327857e-09, 
    -4.621688e-13, -2.840734e-05, 0.2158701, 0.3730426, 0.005193538, 
    0.04210884, 0.00586454, 0.002219813, 0.001354451, 0.008367853, 
    0.0007098577, 0.001120662, 0.001614867, 0.01780895, 0.2906144, 
    0.003587104, 0.02263919, 0.01687476, 0.003455265, 0.001073573, 
    0.0009173107, 0.004861163, 0.01549279, 0.01126202,
  0.006150763, 0.00289611, 0.001102707, 0.198507, -0.0005856216, 
    1.131096e-07, 0.04851818, -6.651163e-06, -0.0001094785, 0.02413129, 
    0.109568, 0.101432, 0.2178756, 0.09894124, 0.1792909, 0.2992654, 
    0.2521363, 0.1394574, 0.05967029, -0.000695179, 0.0009613843, 0.02196738, 
    0.0379617, 0.1656706, 0.04305058, 0.0188438, 0.01752149, 0.01151026, 
    0.0408175,
  0.08348903, 0.1674329, 0.04623181, 0.04267226, 0.002846289, 0.00974731, 
    0.02331669, 0.1356548, 0.0448195, 0.1057959, 0.07002884, 0.1134216, 
    0.3186502, 0.2211625, 0.1148704, 0.1626873, 0.1948453, 0.234399, 
    0.2135725, 0.1295465, 0.04070124, 0.02340386, 0.105689, 0.2956748, 
    0.2009241, 0.1793791, 0.1796061, 0.1461329, 0.07160599,
  0.09377108, 0.1473263, 0.08036285, 0.1413986, 0.2277474, 0.1451168, 
    0.0890256, 0.1279083, 0.125756, 0.24607, 0.2167537, 0.4749074, 0.3549899, 
    0.1546055, 0.166162, 0.1615388, 0.3200022, 0.261358, 0.2150889, 
    0.08718788, 0.07311445, 0.1993553, 0.1104517, 0.1906336, 0.176829, 
    0.1109891, 0.1089643, 0.1120644, 0.1931513,
  0.2969346, 0.1452786, 0.3685127, 0.3186673, 0.4152998, 0.4085528, 
    0.2547143, 0.1157845, 0.1058951, 0.3026055, 0.4019043, 0.274993, 
    0.2063554, 0.1497229, 0.356308, 0.3458415, 0.1913816, 0.1241279, 
    0.1202439, 0.1156097, 0.1219298, 0.230461, 0.3176731, 0.4882957, 
    0.1503403, 0.242992, 0.2778396, 0.1236891, 0.2806125,
  0.3275327, 0.1873821, 0.2290134, 0.4606558, 0.4505898, 0.3779551, 0.3851, 
    0.4310238, 0.3516751, 0.4109846, 0.4096284, 0.3323447, 0.3045441, 
    0.3651707, 0.3458505, 0.4196856, 0.5214607, 0.4717741, 0.5056869, 
    0.4788397, 0.338834, 0.2843435, 0.266714, 0.4411269, 0.2138896, 
    0.1895387, 0.1119184, 0.2761692, 0.2236894,
  0.003736889, 0.002856296, 0.001975704, 0.001095111, 0.000214518, 
    -0.0006660748, -0.001546668, 0.002776114, 0.00317247, 0.003568826, 
    0.003965182, 0.004361539, 0.004757895, 0.005154251, 0.003606171, 
    0.003667156, 0.00372814, 0.003789125, 0.00385011, 0.003911094, 
    0.003972079, 0.001109662, 0.001532914, 0.001956166, 0.002379418, 
    0.00280267, 0.003225921, 0.003649173, 0.004441363,
  0.3155184, 0.1105515, 0.04750528, 0.02455648, -0.0002711116, -0.0001335762, 
    -9.562079e-05, -5.199884e-06, 0, 0, -2.557833e-05, 0.0001830383, 
    0.007240409, 0.007845214, 0.1240581, 0.2940464, 0.3630969, 0.2378851, 
    0.1864622, 0.220329, 0.4030984, 0.3606331, 0.1600921, 0.1537883, 
    0.2858936, 0.4627224, 0.1481314, 0.03535135, 0.3339429,
  0.2219373, 0.05515671, 0.1384101, 0.01797376, 0.07224756, 0.01505441, 
    0.001866735, 0.08195688, 0.1010874, 0.201274, 0.2549312, 0.1280451, 
    0.1608997, 0.1432764, 0.4002452, 0.3204313, 0.2798788, 0.2888318, 
    0.3121083, 0.3082992, 0.331701, 0.285779, 0.2845663, 0.5052727, 
    0.1259156, 0.3461349, 0.4580262, 0.4035431, 0.3584214,
  0.3450655, 0.3119288, 0.2396354, 0.07974333, 0.07739447, 0.1752901, 
    0.2511943, 0.2434592, 0.2907659, 0.08827892, 0.08740055, 0.1259451, 
    0.1728206, 0.1786191, 0.1336281, 0.2353894, 0.2659449, 0.2959935, 
    0.1997336, 0.1443391, 0.1148003, 0.08499257, 0.1122621, 0.07646077, 
    0.1033087, 0.2166335, 0.3007387, 0.3116063, 0.3367729,
  0.1685411, 0.1807451, 0.1498007, 0.1496282, 0.2450138, 0.2054263, 
    0.1707754, 0.09461921, 0.08840878, 0.0938559, 0.07654964, 0.06207943, 
    0.0274704, 0.03867181, 0.07602347, 0.07013851, 0.06908454, 0.16825, 
    0.1322168, 0.1272038, 0.1011192, 0.1111142, 0.07325611, 0.08838344, 
    0.06652845, 0.1094039, 0.1357317, 0.188714, 0.1801424,
  0.03191224, 0.006042657, 0.03748558, 0.1161262, 0.1668864, 0.108804, 
    0.04613664, 0.02425577, 0.0279887, 0.02376086, 0.02056759, 0.002079335, 
    0.0004960737, 0.0654689, 0.09780758, 0.04161268, 0.01738193, 0.05131432, 
    0.08910346, 0.05608888, 0.046062, 0.01963093, 0.01508298, 0.2815142, 
    0.02312379, 0.05796743, 0.08290649, 0.07631639, 0.09557495,
  0.005781463, 0.01105056, 0.001835457, 0.004005357, 0.007966259, 0.0089436, 
    0.005938165, 0.00696254, 0.006742452, 0.002286891, 0.0001315075, 
    -5.424579e-07, 0.002012022, 0.04147471, 0.03680277, 0.03459184, 
    0.02149666, 0.07853905, 0.0493287, 0.005378548, 0.005824877, 0.005062636, 
    0.00810209, 0.002572728, 0.01892258, 0.044826, 0.01849332, 0.008786707, 
    0.006335865,
  0.02527937, 0.01594723, -4.92394e-06, 0.002160524, -0.001880817, 
    -2.348894e-06, 0.0003097514, 0.001552007, 0.00692662, 0.007341718, 
    2.156514e-09, 8.007304e-10, 0.001199628, 0.01910496, 0.007072756, 
    0.00263416, 0.001077937, 0.0008357398, 8.442703e-07, 4.763386e-06, 
    0.001388082, 0.003000727, 0.01551879, 0.0003328445, 5.616006e-05, 
    0.02643785, 0.0002656406, 0.001418542, 0.004349464,
  0.04973468, 0.03987334, -5.220455e-07, 0.04544014, 0.0002808806, 
    8.99684e-05, 0.0005970046, 0.000119617, 0.0004886647, -0.002061228, 
    0.01134388, 0.0008583934, 0.01740916, 0.000505114, 2.166639e-05, 
    0.0001128034, 0.0001402249, 2.421712e-05, 5.652124e-06, 4.794133e-05, 
    0.001032398, 0.008177642, 0.04216978, 6.378777e-06, 1.648742e-05, 
    2.569395e-09, -5.645613e-05, 0.002637556, 0.01136944,
  0.008644702, 0.1012491, 0.0141192, 0.02421293, 0.001081644, 0.0006176094, 
    9.519233e-05, 0.003969621, 0.03941641, 0.0936022, 0.000543837, 
    0.0007016383, 7.154057e-05, 0.0001179885, 0.0001494245, 0.0002726256, 
    0.0002208498, 2.302189e-05, 0.0001993401, 3.793473e-05, 0.002041586, 
    0.03895691, 0.05567389, 0.00271354, 1.650724e-05, 0.001217873, 
    0.0001668192, 0.0006371709, 0.009275289,
  0.006845125, 0.01967198, 0.001503213, 0.06066836, 6.531409e-06, 
    7.124562e-05, 0.02620265, 1.621668e-05, -0.0006692375, 0.0003535394, 
    3.145547e-05, 0.003465908, 0.0002347837, 0.0003752642, 0.0004040185, 
    0.003274376, 0.002767465, 0.01548596, 0.0228376, 0.01540196, 0.003012788, 
    0.001396079, 0.1070477, 0.02014594, 7.761258e-05, 0.0005269127, 
    0.001820052, 0.003099947, 0.02822481,
  2.151836e-08, 4.862098e-08, 1.895887e-07, -9.751497e-06, 1.233702e-09, 
    0.01036678, 0.004320151, 0.001870996, 0.07136505, 0.001809423, 
    0.0004767904, 0.0006371168, 2.643258e-05, 2.103723e-05, 0.0001619691, 
    6.292171e-05, 0.0001058859, 0.0004874459, 0.0098465, 0.0545815, 
    0.004322196, 0.08874526, 0.0002803142, -0.00075345, 0.0001163883, 
    0.001470503, 0.0107721, 0.003864022, 4.767388e-07,
  3.102085e-07, 9.110777e-09, 0.001815239, -1.566804e-06, -2.184201e-09, 
    -1.59794e-12, -2.127846e-05, 0.2019789, 0.3359544, 0.0020438, 0.0186787, 
    0.0022268, 0.001268886, 0.0008035175, 0.004170883, 0.0004751298, 
    0.0006281328, 0.0009744129, 0.01119232, 0.2453265, 0.002816004, 
    0.01422054, 0.0124575, 0.001751922, 0.0006782208, 0.0006027832, 
    0.00294697, 0.01032967, 0.01009599,
  0.003236781, 0.001319799, 0.002217887, 0.1864209, -0.0004826154, 
    1.043647e-07, 0.04692253, -5.996547e-06, -9.412594e-05, 0.01542872, 
    0.09941863, 0.07131217, 0.1648524, 0.05902606, 0.1414181, 0.2417962, 
    0.1822184, 0.08267833, 0.02712678, -0.0007796437, 0.001077523, 0.0206972, 
    0.02835197, 0.1157084, 0.0262452, 0.008779295, 0.009036114, 0.005849188, 
    0.03116481,
  0.06537853, 0.1461382, 0.0337928, 0.0210534, 0.001438831, 0.005910226, 
    0.01424527, 0.1221339, 0.03819445, 0.09531938, 0.06112992, 0.09919222, 
    0.285264, 0.1612043, 0.07387621, 0.1103601, 0.1408245, 0.1704185, 
    0.1674169, 0.11641, 0.0311359, 0.01833726, 0.07590474, 0.2491471, 
    0.1729893, 0.1544274, 0.1350389, 0.09975893, 0.03994841,
  0.05706474, 0.1233246, 0.06428637, 0.1092787, 0.2040037, 0.1246349, 
    0.085255, 0.1184696, 0.1126516, 0.2122347, 0.188727, 0.4305404, 
    0.3237029, 0.1240236, 0.1101531, 0.1129556, 0.2852738, 0.2283037, 
    0.171789, 0.08352036, 0.05415738, 0.1713167, 0.1085615, 0.1576535, 
    0.1355905, 0.08537903, 0.07030265, 0.07158214, 0.1339284,
  0.2026295, 0.09383702, 0.3213419, 0.2413969, 0.3807599, 0.3810441, 
    0.2198802, 0.09167758, 0.08663023, 0.2818621, 0.3604425, 0.2467697, 
    0.1770662, 0.1135985, 0.3282428, 0.283469, 0.1602551, 0.09793293, 
    0.1077427, 0.08437998, 0.1060288, 0.223979, 0.2536725, 0.4320511, 
    0.1194392, 0.1951574, 0.3162378, 0.1116937, 0.2201346,
  0.2738764, 0.1479804, 0.1859513, 0.3896585, 0.3698917, 0.324673, 0.3612355, 
    0.360703, 0.2968535, 0.3421609, 0.3342979, 0.2628648, 0.2511535, 
    0.3127277, 0.2984854, 0.3811968, 0.4211059, 0.3776793, 0.3742726, 
    0.3917092, 0.2767253, 0.2702001, 0.2536348, 0.4402015, 0.1991628, 
    0.1669793, 0.09957137, 0.281178, 0.1886972,
  0.003819135, 0.003142179, 0.002465224, 0.001788269, 0.001111314, 
    0.000434359, -0.0002425961, 0.003241599, 0.003495853, 0.003750108, 
    0.004004363, 0.004258618, 0.004512873, 0.004767127, 0.004509426, 
    0.004523278, 0.00453713, 0.004550982, 0.004564834, 0.004578686, 
    0.004592538, 0.0007925794, 0.001201428, 0.001610276, 0.002019124, 
    0.002427973, 0.002836821, 0.003245669, 0.004360699,
  0.1553686, 0.08050427, 0.0407288, -0.0002639237, 0.0001251885, 
    -9.101311e-05, -2.250747e-05, -7.461053e-06, 0, 0, -3.346679e-05, 
    6.804585e-05, 0.002530398, 0.006888913, 0.1412957, 0.1931391, 0.2423929, 
    0.2056163, 0.1573303, 0.2379702, 0.3692866, 0.3259633, 0.140346, 
    0.1125768, 0.2581019, 0.51518, 0.1553565, 0.02319781, 0.2447443,
  0.2135884, 0.05397429, 0.1148087, 0.01349876, 0.04032787, 0.001896541, 
    0.001024347, 0.05244254, 0.06106132, 0.1571665, 0.2333026, 0.1262256, 
    0.1505608, 0.1277974, 0.387876, 0.2898442, 0.2431999, 0.2561851, 
    0.2662772, 0.2739618, 0.2901891, 0.2456549, 0.2504569, 0.480491, 
    0.1148431, 0.3012463, 0.3970309, 0.3661534, 0.3055148,
  0.2934735, 0.2697783, 0.2088771, 0.06764031, 0.06338418, 0.1587075, 
    0.2135084, 0.2116599, 0.2497585, 0.06714898, 0.0712823, 0.1037504, 
    0.1429775, 0.1447857, 0.102822, 0.1831512, 0.2139286, 0.2473008, 
    0.1640072, 0.1184225, 0.09429681, 0.06155035, 0.0821843, 0.06101586, 
    0.0754097, 0.1852608, 0.2697184, 0.2722197, 0.2942137,
  0.1379347, 0.1457973, 0.1257117, 0.1269654, 0.2172241, 0.1769031, 0.144235, 
    0.07675672, 0.07078373, 0.07042611, 0.05412274, 0.04113529, 0.0172563, 
    0.0260619, 0.05613623, 0.04650661, 0.04893037, 0.1165627, 0.09326405, 
    0.08916218, 0.06703526, 0.0782723, 0.04970111, 0.07454968, 0.04604862, 
    0.08065914, 0.09908826, 0.1540549, 0.1454641,
  0.01932624, 0.003920194, 0.02414923, 0.08189567, 0.1162445, 0.06915977, 
    0.02835916, 0.01446872, 0.01641707, 0.01303746, 0.01357195, 0.001356811, 
    0.0003891802, 0.04323959, 0.06731949, 0.02730411, 0.01044665, 0.03536182, 
    0.0641173, 0.03330531, 0.02786696, 0.01111843, 0.008934745, 0.2559241, 
    0.02059643, 0.04292997, 0.05333056, 0.05001746, 0.059235,
  0.004452038, 0.006125439, 0.001311856, 0.002643352, 0.005459478, 
    0.007104287, 0.004724242, 0.005478043, 0.00514482, 0.001637894, 
    7.780913e-05, -3.390098e-07, 0.003811689, 0.02151093, 0.02118501, 
    0.02100698, 0.01108867, 0.05537861, 0.0263437, 0.003396653, 0.004060823, 
    0.003109048, 0.006376928, 0.001964048, 0.01973752, 0.02717119, 
    0.01019718, 0.004955941, 0.004502774,
  0.01926525, 0.01247335, -2.801335e-06, 0.001612136, -0.001294757, 
    -1.511662e-06, 0.0002296251, 0.001179808, 0.005194379, 0.005007437, 
    1.794815e-09, 6.22939e-10, 0.0008806245, 0.01132278, 0.00385965, 
    0.001794819, 0.000781216, 0.00044078, 6.144894e-07, 3.460611e-06, 
    0.001009355, 0.002197167, 0.01159041, 0.0002162656, 3.399159e-05, 
    0.02156162, 0.0002050973, 0.001038009, 0.003033266,
  0.03570634, 0.02450622, 1.292388e-06, 0.02925684, 0.0001416247, 
    5.251772e-05, 0.0003254984, 6.687815e-05, 0.0003665082, -0.001122638, 
    0.008660459, 0.0004038264, 0.008730619, 0.0002840869, 2.197237e-05, 
    6.175796e-05, 9.427936e-05, 1.820059e-05, 3.963124e-06, 3.52854e-05, 
    0.0007530965, 0.005862866, 0.03081483, 0.0001165083, 7.303317e-07, 
    1.78611e-09, -1.415476e-05, 0.001983327, 0.008069658,
  0.006209671, 0.08666948, 0.007437394, 0.01689755, 0.0007411733, 
    0.0003747001, 6.265928e-05, 0.001726707, 0.02800334, 0.08501744, 
    0.0003670935, 0.0005032273, 5.736344e-05, 8.744924e-05, 0.0001078363, 
    0.0001948946, 0.0001523907, 1.449389e-05, 0.0001429314, 2.383716e-05, 
    0.001435986, 0.0263686, 0.04194942, 0.002560446, 0.0004331195, 
    0.0008791141, 0.0001188145, 0.0004467886, 0.00657043,
  0.005206272, 0.01269704, 0.0006488048, 0.04596044, 3.681729e-06, 
    5.087613e-05, 0.01056637, 1.148805e-05, -0.0005451152, 0.000173386, 
    2.56054e-05, 0.00162377, 0.0001200596, 0.0002249864, 0.0002584191, 
    0.001629793, 0.001188907, 0.007299223, 0.01008093, 0.006523796, 
    0.001340549, 0.0006337736, 0.09982968, 0.02542086, 5.598547e-05, 
    0.0003855105, 0.001012956, 0.001521382, 0.02460389,
  2.091317e-08, 4.693804e-08, 3.787417e-07, -5.253439e-06, -2.722159e-09, 
    0.007018875, 0.002231013, 0.000790251, 0.05933426, 0.0002969424, 
    0.000331182, 0.0003967551, 1.577923e-05, 1.401493e-05, 0.0001176137, 
    4.538108e-05, 8.093928e-05, 0.0003372546, 0.007055872, 0.03242201, 
    0.002808335, 0.07347889, 0.0002101385, -0.0007445678, 6.891258e-05, 
    0.001043041, 0.007497014, 0.002756617, 4.71636e-07,
  2.76725e-07, -1.41823e-09, 0.0009565597, -1.192653e-06, -2.069974e-09, 
    5.025899e-13, 1.379696e-05, 0.1913283, 0.3157946, 0.0006451642, 
    0.008035798, 0.001256278, 0.0008929985, 0.0005673224, 0.002400775, 
    0.0003582924, 0.0004435229, 0.0006810466, 0.008084643, 0.2151629, 
    0.002136626, 0.009186903, 0.00953103, 0.001035229, 0.000496267, 
    0.000448122, 0.002077378, 0.007725562, 0.008608704,
  0.003537771, 0.0004948738, 0.00194768, 0.1643892, -0.0004157931, 
    9.736086e-08, 0.03980559, -5.958437e-06, -7.999223e-05, 0.009457372, 
    0.09212705, 0.04442267, 0.1193417, 0.0332902, 0.09902311, 0.1961842, 
    0.1210087, 0.05348473, 0.01590272, -0.0006816112, 0.001029054, 
    0.01923574, 0.02302472, 0.0876166, 0.01538, 0.004716441, 0.00503685, 
    0.003475408, 0.02568825,
  0.05509068, 0.1329514, 0.02712157, 0.01397068, 0.0008903274, 0.00382111, 
    0.01004193, 0.110069, 0.03200189, 0.08740754, 0.05124319, 0.09236155, 
    0.2267124, 0.1104851, 0.0489149, 0.0783808, 0.1013773, 0.1265672, 
    0.1225096, 0.1046525, 0.02466727, 0.01459681, 0.05744834, 0.2137086, 
    0.1528896, 0.1366321, 0.09895774, 0.06976143, 0.02348821,
  0.03127541, 0.1090543, 0.05611869, 0.08466429, 0.1816419, 0.1145236, 
    0.09385228, 0.1118407, 0.1093246, 0.1853277, 0.1666375, 0.3948859, 
    0.2885139, 0.09763764, 0.07251853, 0.07856914, 0.2531888, 0.2078321, 
    0.1463688, 0.08651069, 0.04179794, 0.1547283, 0.0802228, 0.1324429, 
    0.09909874, 0.06868625, 0.04524011, 0.04390335, 0.08667119,
  0.1425009, 0.06479212, 0.2821758, 0.1792904, 0.3039806, 0.3670667, 
    0.2019491, 0.07213214, 0.07864101, 0.2481142, 0.3280602, 0.2112177, 
    0.1467987, 0.09394217, 0.2923476, 0.2363642, 0.1386977, 0.07898208, 
    0.1000953, 0.06768727, 0.08985867, 0.2158392, 0.209711, 0.3877951, 
    0.1041354, 0.1584189, 0.3371793, 0.1004131, 0.149319,
  0.2320642, 0.126463, 0.1644245, 0.3221795, 0.3031285, 0.2836593, 0.3107771, 
    0.3041341, 0.2432539, 0.2875484, 0.2778439, 0.2132147, 0.2242019, 
    0.253729, 0.238665, 0.306133, 0.3475943, 0.3126805, 0.2919859, 0.3088323, 
    0.2228272, 0.244165, 0.223107, 0.4284109, 0.1948333, 0.1376496, 
    0.1018691, 0.2721912, 0.1605067,
  0.003320626, 0.002881413, 0.0024422, 0.002002987, 0.001563774, 0.001124562, 
    0.0006853486, 0.002813518, 0.002984601, 0.003155684, 0.003326768, 
    0.003497851, 0.003668934, 0.003840018, 0.003009143, 0.003090714, 
    0.003172285, 0.003253856, 0.003335427, 0.003416998, 0.003498569, 
    0.002061245, 0.002247803, 0.002434362, 0.00262092, 0.002807479, 
    0.002994037, 0.003180596, 0.003671996,
  0.1088076, 0.06422083, 0.0333178, 0.0002694232, 0.0001337228, 
    -6.779541e-05, -7.778181e-06, 0, 0, 0, 0, 4.570744e-05, 0.002271257, 
    0.007510916, 0.1465315, 0.1443805, 0.1869206, 0.2067975, 0.1461458, 
    0.2309783, 0.3462894, 0.3476567, 0.1326597, 0.109943, 0.2296435, 
    0.4849829, 0.1806402, 0.01967364, 0.1545289,
  0.2187068, 0.06199373, 0.1192345, 0.01405487, 0.03119725, 0.001935636, 
    0.0008166452, 0.05080759, 0.04252151, 0.1412032, 0.2234609, 0.1213923, 
    0.1484918, 0.1198968, 0.3695937, 0.279541, 0.2299487, 0.2420967, 
    0.2437592, 0.2616797, 0.2699751, 0.2292188, 0.2321997, 0.4594262, 
    0.1145559, 0.2688296, 0.3646346, 0.3324635, 0.2738591,
  0.2651681, 0.2565277, 0.1957878, 0.06235538, 0.05700532, 0.1550545, 
    0.1999467, 0.192549, 0.2336275, 0.05753819, 0.06290932, 0.09159563, 
    0.1292365, 0.1247614, 0.08710536, 0.156083, 0.1892149, 0.209489, 
    0.1441044, 0.1033905, 0.08295741, 0.05060146, 0.06684031, 0.05104585, 
    0.0654726, 0.1738234, 0.2521498, 0.2618544, 0.2629887,
  0.1196772, 0.1237653, 0.1071916, 0.1101366, 0.1908886, 0.1460116, 
    0.1229368, 0.06743973, 0.06254821, 0.05840267, 0.04319919, 0.0328713, 
    0.01337161, 0.01969066, 0.04397645, 0.03400395, 0.03875128, 0.09032985, 
    0.07427839, 0.07142764, 0.05081134, 0.06009049, 0.0384374, 0.08507214, 
    0.03750523, 0.06714066, 0.08334164, 0.1314708, 0.1242915,
  0.01398892, 0.003134116, 0.01674322, 0.06332438, 0.08723795, 0.04814954, 
    0.02032713, 0.01084372, 0.01177469, 0.008944328, 0.01052482, 0.001111812, 
    0.0003366728, 0.03342858, 0.0524445, 0.01993284, 0.007788775, 0.02757322, 
    0.04896837, 0.02402189, 0.01893965, 0.007698941, 0.00597404, 0.2560371, 
    0.01913097, 0.03530036, 0.03726174, 0.03628533, 0.03914427,
  0.003786181, 0.004602996, 0.001161776, 0.002127242, 0.004064945, 
    0.00610732, 0.004077869, 0.004688052, 0.004335911, 0.001326204, 
    5.042654e-05, -2.504564e-07, 0.0104638, 0.01214025, 0.01469577, 
    0.0127401, 0.006981164, 0.03826591, 0.01683871, 0.002612008, 0.003354277, 
    0.002365843, 0.005503102, 0.001761406, 0.01799162, 0.01744792, 
    0.006241574, 0.003682114, 0.003697502,
  0.01627467, 0.01034669, -1.830922e-06, 0.001340753, -0.001154056, 
    -1.109241e-06, 0.0001952691, 0.001015686, 0.004373522, 0.003923961, 
    2.606243e-09, 8.108241e-10, 0.0007279897, 0.006656304, 0.002329252, 
    0.00141139, 0.0006415147, 0.0003245189, 5.889449e-07, 2.943088e-06, 
    0.000835003, 0.001833102, 0.009751328, 0.0001720311, 2.124262e-05, 
    0.0276056, 0.0001747898, 0.0008670269, 0.00244002,
  0.02894951, 0.01826295, 5.430545e-05, 0.02422391, 9.924651e-05, 
    3.976524e-05, 0.0002438431, 5.041673e-05, 0.0003110589, -0.0008627353, 
    0.006974521, 0.0002398136, 0.005780548, 0.0002133597, 1.997421e-05, 
    4.496423e-05, 7.52503e-05, 1.533391e-05, 3.272691e-06, 2.954437e-05, 
    0.0006305439, 0.004810985, 0.02526773, 0.001905992, -6.557784e-05, 
    3.494385e-09, -3.34952e-06, 0.001668095, 0.006578744,
  0.005024767, 0.141858, 0.01181095, 0.0157199, 0.0005778833, 0.0002856049, 
    4.788283e-05, 0.001070972, 0.03008652, 0.1002269, 0.000292354, 
    0.0004054788, 4.841165e-05, 7.104927e-05, 8.889342e-05, 0.0001584697, 
    0.000123446, 1.159545e-05, 0.0001169946, 1.908238e-05, 0.001086529, 
    0.02070277, 0.03490636, 0.01269109, 0.01000013, 0.0007150445, 
    9.806909e-05, 0.0003611401, 0.005259892,
  0.02401781, 0.01177665, 0.0004746697, 0.03774611, 2.367236e-06, 
    4.194554e-05, 0.007082628, 9.527664e-06, -0.002675497, 0.0001141469, 
    2.276867e-05, 0.001037136, 8.011462e-05, 0.0001774975, 0.0001964989, 
    0.001055171, 0.0007418109, 0.004205625, 0.005866924, 0.003669359, 
    0.0008791086, 0.0004403481, 0.1809745, 0.0336783, 4.658565e-05, 
    0.0003153807, 0.0007200966, 0.001117809, 0.05544249,
  2.061497e-08, 4.601446e-08, 3.704901e-07, -3.48562e-06, -4.597066e-09, 
    0.005420384, 0.002241872, 0.0004636892, 0.08762575, -0.0005657641, 
    0.0002706963, 0.0002899315, 1.227177e-05, 1.127768e-05, 9.682441e-05, 
    3.672204e-05, 6.897024e-05, 0.0002677308, 0.005737025, 0.02048004, 
    0.002200407, 0.06850349, 0.0001747107, -0.001401252, 5.268484e-05, 
    0.0008470214, 0.006012137, 0.002239605, 4.747498e-07,
  2.643216e-07, -1.009343e-07, 0.0003638579, -8.551532e-07, -1.993659e-09, 
    -8.423672e-13, 0.0009863127, 0.2003131, 0.3193026, 0.0003554288, 
    0.005455408, 0.0009252085, 0.000684209, 0.0004573705, 0.001824945, 
    0.0003025235, 0.000362527, 0.0005451186, 0.006613772, 0.1951818, 
    0.003535163, 0.01609218, 0.01811511, 0.0007695077, 0.0004081772, 
    0.0003697446, 0.001566297, 0.006444085, 0.00724651,
  0.005201503, 9.139995e-05, 0.001852798, 0.1496998, -0.0003978137, 
    1.388032e-07, 0.03556325, -6.279655e-06, -7.313363e-05, 0.005553214, 
    0.1040227, 0.02246264, 0.09644511, 0.02165798, 0.0673503, 0.1450304, 
    0.08046195, 0.03405457, 0.01205792, -0.0006412414, 0.0009901352, 
    0.0175861, 0.03166685, 0.06300797, 0.009608836, 0.00315331, 0.003583136, 
    0.002492334, 0.02322591,
  0.04810804, 0.1392524, 0.02964419, 0.0137056, 0.0007092635, 0.002786851, 
    0.008365285, 0.1102908, 0.03495772, 0.09374462, 0.07906664, 0.1156687, 
    0.1885257, 0.08242727, 0.03539357, 0.06206406, 0.07216369, 0.09656575, 
    0.08306634, 0.09949249, 0.02219866, 0.01381304, 0.06243599, 0.2327989, 
    0.1482402, 0.1162484, 0.07721621, 0.04939017, 0.01620917,
  0.0193737, 0.1176959, 0.06454857, 0.07251874, 0.2048796, 0.1336188, 
    0.1294816, 0.1507027, 0.1428714, 0.2039389, 0.1726635, 0.4003625, 
    0.2789664, 0.09985127, 0.05666051, 0.05757917, 0.2682154, 0.1971971, 
    0.1553149, 0.09548647, 0.03979564, 0.1732617, 0.06102396, 0.1316631, 
    0.07901314, 0.06137848, 0.03194381, 0.02978408, 0.06098969,
  0.1048398, 0.04720428, 0.2867671, 0.1345722, 0.2389545, 0.3395731, 
    0.2085911, 0.07579644, 0.08560295, 0.2417577, 0.3300693, 0.2182861, 
    0.1381454, 0.08115135, 0.251444, 0.2095014, 0.1282192, 0.06852756, 
    0.09413262, 0.05744017, 0.07482473, 0.1982665, 0.1935615, 0.3577109, 
    0.08508095, 0.1369215, 0.3803146, 0.08859442, 0.1114508,
  0.204938, 0.1102418, 0.1504271, 0.2742644, 0.2667171, 0.2511892, 0.2675401, 
    0.2717261, 0.2061752, 0.2592616, 0.2371298, 0.1834888, 0.1958585, 
    0.2137551, 0.1998409, 0.2496639, 0.3016909, 0.2708806, 0.2476508, 
    0.2668933, 0.1907983, 0.2317434, 0.216931, 0.3968654, 0.1845884, 
    0.1239521, 0.1240149, 0.2633601, 0.1487926,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6.154653e-05, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2.230827e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, -8.124457e-06, 0, 0, 0, 0, 0, -6.048856e-06, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.473911e-05, 0, 
    -4.159544e-06, 0, -7.22978e-06, 0, 0, 0.001278043, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -3.775271e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -3.746029e-05, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0.002037907, 0, 0, 0, -4.805837e-11, 0, -3.249783e-05, 0, 0, 0, 0, 0, 
    -3.021615e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2.899475e-05, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, -1.68484e-05, 0, 0, -3.862627e-05, -5.324242e-06, 
    -3.945397e-05, 0.0005304427, 0.0003213612, -9.10747e-06, 0, 0, 
    0.0007594192, 0, -2.570566e-05, 0, 0.0009071177, 0, 0, 0.003324798, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -5.905418e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -6.16363e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, -8.164448e-06, -9.222302e-05, 0, 0, 0, 0, 0, 0, 0.002850032, 
    0.0004145993, 0, 0, 0, 0, 0, 0, 0, 0, -3.281154e-06, 0, 0, 0, 0, 0,
  0, 0.003485011, 0.0004134018, 0, 0, 7.396915e-06, 0, -9.210917e-05, 0, 0, 
    0, 0, -1.470585e-05, -7.522603e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -4.790024e-05, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, -0.0001934672, -1.626908e-05, 0.0002041936, 
    -8.050026e-05, -5.324242e-06, 0.0006348848, 0.002867679, 0.0009811906, 
    -2.845141e-05, 0.0003236224, 0.0001292403, 0.005234789, 0.00130743, 
    -4.513313e-05, 0.000205271, 0.004460293, -4.364609e-06, 0, 0.006271483, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2.285427e-06, 2.323892e-05, -4.880111e-05, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0009548934, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.237933e-05, 0.0001382474, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -4.257934e-05, -3.926973e-05, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -3.58668e-05, 0, 
    -9.548405e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, -0.000113998, -0.0001706786, 0, 0, 0, 0, 0, -5.15609e-05, 
    0.002780244, 0.0004354316, 0, 0, 0, 0, 0, 0, 0, 0, 0.0005932897, 0, 0, 0, 
    0, 0,
  0, 0.01002971, 0.001664266, 0, 0, 6.87446e-05, 0, -6.193431e-05, 
    -5.170505e-05, 0, 0, 0.0004441048, 1.476801e-06, 0.002098887, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, -4.875969e-05, 0, 0, 0, 0, 0,
  0, 0, 0, -4.733762e-06, 0, 0, 0.0003653515, -7.829882e-05, 0.002984954, 
    -0.0003136916, -6.193804e-05, 0.00296518, 0.01055276, 0.004036393, 
    0.001501552, 0.002707099, 0.001730951, 0.01144197, 0.003315308, 
    0.0009236381, 0.0006626823, 0.008623817, -8.377289e-05, -1.513061e-05, 
    0.009140997, -7.446614e-06, -4.477482e-05, 0, 0,
  0, 0, 0, 0, 0, 3.463354e-05, 0, 0, -4.053793e-06, 0, -8.71263e-06, 
    0.009462229, 0.0001458888, 0, 0, 0, 0, -3.483986e-05, 0, 0, 8.93318e-06, 
    0, 0, 0, 0, 0.003073286, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0001221773, 0.0001541064, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0.0008987286, -1.153022e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.0008223205, 0.0005174491, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.00161295, 0, 0.002619454, 
    -8.733144e-06, 0, 0, 0, 0, 0, 0, 1.319225e-05, 0, 0, 0,
  0, 0, 0, 0, 7.001641e-06, -0.0002179434, -0.0003626918, 0, 0, 0, 0, 
    -1.511857e-05, -0.000115819, 0.004648985, 0.0004502205, -0.0001070642, 
    -4.6193e-05, 0, 0, 0, 0, 0, 0, 0.002714153, 0.001607177, 0, 0, 0, 0,
  -1.466606e-05, 0.02170042, 0.004930328, 0, 0, 0.002380342, 0, 2.832318e-05, 
    -0.0001160036, -5.875896e-06, 0, 0.0004504337, 6.921834e-05, 0.003720431, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, -9.541083e-05, 0, 0, 0, -7.539543e-07, 0,
  0, 0, 0, -7.235114e-05, 0, 0, 0.002614645, -0.0001911795, 0.004731748, 
    0.001613482, -0.0001395924, 0.006626505, 0.02589686, 0.01284367, 
    0.004752196, 0.005168595, 0.002994629, 0.02283999, 0.01271249, 
    0.002013281, 0.0007777871, 0.01510597, -0.0002040116, 0.0001043803, 
    0.01113865, -9.575576e-06, 0.0001777333, 0, 0.0008380768,
  0, 0, 0, 0, 0, -5.377397e-05, 0, -1.136579e-05, -1.688352e-05, 0, 
    4.279487e-06, 0.02060095, 1.097489e-06, 0, 0, 0, 0, 0.0001277738, 0, 0, 
    -2.195077e-06, 0, 0, 0, 0, 0.005810348, -1.719154e-05, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.002014353, 0.001698202, -0.0002171198, 
    0.0002811451, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5.361647e-06, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2.050048e-07, -8.007573e-05, 
    0.0002938849, 0, -2.749047e-05, 0, -3.07239e-05, 0, 0, 0, 0, 0, 0, 
    -7.079433e-06, -2.060131e-06, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -3.546825e-05, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, -2.199679e-06, 0.0005697064, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, -1.92331e-07, 0, 0, 0, 0, 0, -7.346438e-07, 0, 0, 0,
  0, 0, 0, 0.002086059, -2.151592e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -1.137266e-05, 0, 0.0005502679, 0, 0, 0, 0, 0, 0.001613034, 0.009255762, 
    -7.977227e-05, 0, 0,
  0, 0, 0, 0, -9.07396e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.002535058, 
    -5.599033e-06, 0.009054874, -0.0001135785, 0, 0, 0, 0, 0, 0, 0.000923129, 
    0, 0, 0,
  0, 0, -3.03104e-06, 0, 0.0002061646, 0.0008643484, -0.0006286228, 0, 0, 0, 
    0, -3.887605e-05, 0.001419847, 0.01091112, 0.001879948, -0.0002262013, 
    0.0007708458, 0, 0, 0, 0, 0, 0, 0.00348147, 0.003175766, 0, 0, 0, 0,
  -1.023825e-05, 0.03901584, 0.007523295, 0, 0, 0.008115639, -1.655378e-05, 
    0.0003466931, 6.642511e-05, -7.734417e-05, 0, 0.001054631, 0.000765299, 
    0.005482585, 0, 0, -7.07513e-05, 0, 0, 0, 0, 0, 0, -0.0001005474, 0, 0, 
    1.264087e-05, -3.015817e-06, 0,
  0, 0, 0, 0.001060588, 0, 0, 0.01248701, -0.000332502, 0.01316785, 
    0.008674879, -2.086291e-05, 0.01202101, 0.0527008, 0.02442395, 
    0.01276899, 0.00736049, 0.007120233, 0.04429347, 0.02600222, 0.003604661, 
    0.001870811, 0.02054843, -0.0001113665, 0.001064699, 0.01382474, 
    -0.0001026354, 0.0006018525, 6.350077e-05, 0.004012785,
  0, 0, 0, 0, 0, 2.17432e-05, 0, -2.007388e-05, -4.461769e-05, 0, 
    0.000671945, 0.04025114, 0.001429707, 0, 0, 0, 0, 0.0001436479, 0, 0, 
    0.001019017, 0, 0, 0.0003210425, 0, 0.008555872, 0.000200173, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.004737178, 0.009894996, 0.001115953, 
    0.005714893, 0.000489917, -9.199701e-06, 0, 0, 0, 0, 0, -2.388851e-06, 0, 
    0, 0.0001846026, 6.966882e-05, 0, 0, 0,
  0.0002117478, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.00690899, -2.793508e-05, 
    0.004268022, 0.0003827955, 0.0002362297, 0.001459308, 0.0002579224, 0, 0, 
    0, 0.0008457053, 1.386227e-05, -1.601597e-05, -1.234525e-05, 
    -2.345549e-05, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001620328, 1.996909e-05, 
    0, 0, 0, 0, 0, 0, -5.944255e-06, -1.620665e-05, -1.641839e-05, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -8.283734e-08, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, -8.417326e-06, -9.483421e-05, 0.003013554, 0, 0, 0, 0, 0, 
    -7.770896e-06, 0, 0, 0, 0, 0, 0, 0, -1.932181e-05, 0, 0, 0, 0, 0, 
    -4.342528e-05, 0.0005838685, -1.370676e-05, 0,
  0, 0, 0, 0.005964808, 0.001146854, -9.813507e-05, 0, 0, 0, 0, 0, 
    9.148133e-08, 0, -6.688224e-05, 0, 0, -7.529155e-05, 9.379969e-05, 
    0.00424098, 0, 0, 0, 0, 0, 0.005959458, 0.02317924, 0.00698821, 
    -3.592245e-05, 0,
  0, 0, 0, 0, 0.0005245007, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.16945e-06, 
    0.00578032, 0.002565152, 0.01672463, 0.0009269739, -2.131626e-10, 0, 0, 
    0, 0, 6.753168e-05, 0.002150024, 0, 0, 0,
  0, 0, 0.0001729791, 0, 0.0002104842, 0.007530023, 0.00089591, 
    -2.713417e-09, 0, 0, -1.17255e-05, 0.0009087505, 0.008564995, 0.0289155, 
    0.004091152, 7.777872e-05, 0.005259351, -4.674541e-07, 0, 0, 0, 0, 0, 
    0.01254683, 0.003647172, -1.73789e-05, 0, 0, 0,
  -2.222054e-05, 0.0535721, 0.009296576, 0, 0, 0.01273187, -1.997011e-05, 
    0.005597047, 0.002854858, -0.0003477282, 1.6702e-06, 0.004457449, 
    0.003180751, 0.01477889, 6.126216e-05, 0, 1.41665e-05, 1.690321e-05, 0, 
    0, 0, 0, 0, 0.0006158881, 1.247173e-05, 0, 0.0002808356, -9.473518e-06, 0,
  -2.922517e-06, -6.987437e-05, 0, 0.003564832, 0, -2.799214e-05, 0.02262449, 
    0.001194254, 0.02272264, 0.02262762, 0.002350844, 0.03107737, 0.08468135, 
    0.04377565, 0.02465922, 0.01418589, 0.01154306, 0.07044664, 0.03933512, 
    0.004706346, 0.0101724, 0.02801808, 0.00134183, 0.002861159, 0.01522644, 
    0.0005850727, 0.001923547, 0.0005648978, 0.006854399,
  0, 0, 0, 0, 0, 0.0005612855, 0, 0.0002734376, 0.0003246772, -9.776336e-06, 
    0.005797841, 0.06234131, 0.00451015, 3.162252e-06, -3.517175e-05, 0, 
    0.0004886505, 0.001887342, -7.102082e-05, -1.447528e-06, 0.003840614, 0, 
    0, 0.001269351, -1.106857e-05, 0.0140011, 0.006463624, 0, 0,
  0, 0, 0, 0, -3.281094e-06, 0, 0, 0, 0, -1.951687e-06, 0.008171594, 
    0.01924532, 0.007580761, 0.007162415, 0.003827887, -0.0001507932, 0, 
    -1.955179e-06, 0.001689198, 0.001089921, 0, -3.471797e-05, 0, 
    7.021369e-05, 0.004367831, 0.001803382, 0, 0, 0,
  0.002932993, -2.125861e-05, 0, 0, 0, 0, 0, 0, 0, 0, -2.220659e-07, 
    0.01662751, 0.003262526, 0.0118318, 0.009447232, 0.005534354, 
    0.008717801, 0.002070515, -4.234319e-06, 0, 0, 0.007612242, 0.002016948, 
    -7.690994e-05, 0.0003263234, 4.638613e-05, 3.308472e-06, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.004522455, 1.131958e-05, 
    -3.442536e-05, 0, 0, 0, 0, 0, 0.0001649018, 0.002814214, 0.001026422, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001533309, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.0002713795, 0.00022405, 0, 0,
  0.000468781, 0, 0, 0.001177552, 0.004417126, 0.00965946, -6.753759e-05, 0, 
    0, 0, 0, 0.0009620117, 8.644633e-07, 0, -0.0001149707, 0.0008108442, 
    -8.457001e-05, 0, -1.930583e-05, 0.002366903, 0, -0.0001117906, 0, 0, 
    0.0007610258, 0.003075541, 0.00279487, 0.0002069432, 0,
  0, -8.676979e-06, 0, 0.01735349, 0.008713471, -0.0002777867, 0, 0, 0, 0, 0, 
    1.091543e-05, 0.0001482691, 0.002607029, -3.041329e-05, -0.0002869304, 
    0.0004811305, 0.003446381, 0.006529305, 0.008456564, -0.0001358793, 0, 0, 
    0, 0.008864949, 0.04487341, 0.02177853, 0.002423359, -7.46001e-05,
  -2.065315e-08, 0, -8.181607e-08, 0, 0.002049988, -1.207767e-05, 0, 0, 0, 0, 
    0, -4.038598e-06, 0, 8.344582e-05, 0.01414967, 0.01521016, 0.01321562, 
    0.02728179, 0.01023018, 2.374379e-06, 3.246809e-07, 0, 0, -1.945958e-07, 
    0.001442324, 0.004655788, 0.0001682155, 0.0002669793, 0,
  -7.808379e-11, -7.634983e-06, 0.001874851, 1.730244e-06, 0.001957393, 
    0.02761164, 0.006427294, -3.692296e-06, -8.14341e-05, 0, 0.0004753706, 
    0.01137991, 0.02003518, 0.05733931, 0.01550451, 0.002950328, 0.01248125, 
    -1.900691e-06, 1.465055e-06, 0, 0, 0, 4.357912e-06, 0.03877023, 
    0.02348846, -8.628765e-06, 9.205347e-13, 3.760673e-05, 0,
  0.002318193, 0.0818291, 0.01780833, 1.190218e-06, 0, 0.01751716, 
    -6.658394e-05, 0.01796366, 0.02188402, 0.0008889588, 8.823394e-05, 
    0.03201738, 0.02078764, 0.03635707, 0.002617325, -4.514715e-07, 
    0.0009277871, 4.194567e-05, -2.265389e-09, 0.0007886316, 0, 1.138436e-09, 
    1.501623e-06, 0.02776584, 0.0003903206, 0, 0.0005438441, 0.0002137605, 0,
  0.0005448502, -0.0001122829, -2.291691e-05, 0.005756396, -5.896568e-06, 
    -4.654878e-05, 0.03749493, 0.01335108, 0.04127442, 0.05701391, 
    0.01850343, 0.09147985, 0.152297, 0.08883747, 0.07177011, 0.0397744, 
    0.0255538, 0.1209549, 0.05641986, 0.008883711, 0.023582, 0.04716664, 
    0.01737471, 0.009455622, 0.02008289, 0.005849622, 0.009520432, 
    0.00452943, 0.01471451,
  0, 0, 0, 2.3632e-08, 0, 0.002382667, 0.0008695854, 0.0002978086, 
    0.001939991, 0.001133015, 0.01490649, 0.08691359, 0.01597263, 
    0.0003250625, 7.830313e-05, 7.33987e-07, 0.0008937166, 0.01499063, 
    0.0007047275, -1.397774e-05, 0.007754121, -1.146729e-05, 0.0009832721, 
    0.001317032, 0.000165608, 0.01915116, 0.0231182, 0, -5.601354e-07,
  0, 0, 0, 0, -4.600456e-05, 0, 0, 0, 0, -0.000107439, 0.008086122, 
    0.03658487, 0.02375228, 0.01558038, 0.009474615, 0.002693438, 
    -1.130155e-05, -0.0001152142, 0.00433208, 0.006731394, -1.901041e-07, 
    -1.769022e-06, -0.0001285136, 0.001282097, 0.009687481, 0.004871356, 0, 
    0, 0,
  0.003608176, 0.000413155, 0, 0, 0, 0, 0, 0, 0, 0, -1.641613e-05, 
    0.02903231, 0.02071198, 0.02643006, 0.02725625, 0.02024204, 0.01216145, 
    0.003068692, -1.687286e-05, 0, 0, 0.01088612, 0.004052694, -4.27958e-05, 
    0.01102805, 0.001182183, 4.30764e-05, -1.473008e-05, 0,
  0, 0.000810867, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.867921e-06, -1.383207e-07, 
    -8.902604e-13, 0, 0.0001235237, 0.01477786, 0.003305629, 0.004441083, 0, 
    0, 0, 0, 0, 0.003772656, 0.01416999, 0.01264662, -5.116748e-05, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -6.252631e-06, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.0001470491,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0.0008526851, -4.749107e-05, 0.0002978597, 0, 0, 0, 0, 0, 
    0.002936447, 0, 0.0001810187, 5.823267e-05, 0, 0, 0.0003224351, 0, 0, 0, 
    0, 0, 0.002883485, 0.002779997, -8.709419e-05, 0,
  0.004229086, 0.0001653862, 0, 0.00716128, 0.01409125, 0.01883201, 
    0.0002633811, -4.975328e-05, 0, 0, 0, 0.004649748, 0.005723955, 
    0.0006955823, -0.0001491748, 0.003520981, 0.003155772, 0, 0.0008247188, 
    0.007022276, 0.001972493, 0.003004222, 0, 0, 0.004523881, 0.01542853, 
    0.009787302, 0.002420261, -2.422195e-08,
  -5.38092e-05, 0.005134628, 0, 0.02773975, 0.02144231, 0.002120439, 
    4.362387e-07, 0, 0, 0, 5.23304e-07, 3.897628e-05, 0.001452881, 
    0.004942125, 0.002179525, 0.01114151, 0.006090404, 0.01854129, 
    0.02045785, 0.02833313, 0.00371752, 0.00088633, 9.296527e-05, 
    0.0004155585, 0.0135489, 0.06256652, 0.03865841, 0.005537109, 0.0005380196,
  -1.931157e-07, -1.721718e-05, -2.835294e-07, 0, 0.005318536, 0.00180216, 
    -0.0001140851, -1.126143e-10, 0, 1.543766e-07, 2.853121e-08, 
    -0.000155014, 0.002920186, 0.001973383, 0.02256355, 0.03113489, 
    0.03448763, 0.06050353, 0.02384619, 0.00156279, 1.94038e-05, 
    -4.728641e-07, 0, 0.0002525652, 0.01477966, 0.01547122, 0.001898159, 
    0.0005702184, 6.047503e-05,
  1.255703e-06, 0.002346347, 0.002855306, 9.141023e-05, 0.002205358, 
    0.05267908, 0.02295782, 0.001475144, 0.00150851, 6.551792e-07, 
    0.004096564, 0.1330968, 0.1039139, 0.1518062, 0.1039847, 0.03752224, 
    0.01646708, -7.387129e-06, 0.0006222485, 8.614242e-05, 0, -9.41257e-08, 
    9.295915e-05, 0.1609183, 0.1510586, 0.004442388, 7.42129e-05, 
    0.0007638832, 7.623017e-09,
  0.002461913, 0.1504253, 0.06293833, 6.055135e-06, 3.931107e-05, 0.02844626, 
    0.002100163, 0.04073982, 0.1010374, 0.03039359, 0.03184727, 0.1938418, 
    0.1336404, 0.1252456, 0.03807405, 1.967908e-05, 0.002898792, 0.004493547, 
    -1.271001e-06, 0.006441772, -2.820305e-08, 3.971982e-07, 0.00381452, 
    0.1604219, 0.05540748, 2.292379e-05, 0.002552508, 0.003763855, 
    -4.661158e-08,
  0.0008758551, 0.001291924, 0.0001378319, 0.01029154, 1.629209e-05, 
    0.0001874461, 0.09536348, 0.07805668, 0.1551988, 0.1630865, 0.2094325, 
    0.3234368, 0.3433725, 0.2772901, 0.3138451, 0.1959184, 0.07226276, 
    0.2164101, 0.08864605, 0.02756639, 0.08868938, 0.1806125, 0.07481921, 
    0.05336254, 0.0262778, 0.02540853, 0.03127903, 0.02439095, 0.02379796,
  -6.357859e-06, -2.238591e-06, 0, 1.206346e-05, 2.313577e-05, 0.007264148, 
    0.007484268, 0.009802457, 0.0204885, 0.01127328, 0.0661208, 0.1429856, 
    0.09847981, 0.02448676, 0.01587882, 4.268368e-05, 0.004547739, 
    0.03458574, 0.002860447, 0.004982135, 0.05048816, 0.0004712623, 
    0.0105383, 0.01512404, 0.004343113, 0.02487275, 0.03759639, 5.389753e-05, 
    0.0006726195,
  0, 4.267582e-05, -1.266669e-08, 0, 0.0007745749, -1.179792e-05, 
    0.000286234, 0, 1.836357e-05, 0.009955749, 0.009651572, 0.1226694, 
    0.08595995, 0.0662319, 0.04077854, 0.0231505, 0.002626625, 0.005575079, 
    0.006824708, 0.01610188, -0.0003097131, 0.002369112, 0.0006245562, 
    0.0096337, 0.0176799, 0.0123723, 0, -4.235485e-07, -1.522897e-08,
  0.008502824, 0.002410972, 0, 0, -3.96583e-07, 0, 0, 0, 0.001117547, 
    -8.224234e-06, 1.881723e-05, 0.05743628, 0.04513356, 0.06048872, 
    0.05585103, 0.05702426, 0.02661494, 0.011865, 0.0003522589, -3.78256e-06, 
    0, 0.01487123, 0.007976858, 0.003725587, 0.03514434, 0.005686954, 
    0.0006571321, 0.0005391015, 0,
  -0.0001250436, 0.006517426, 0, 0.0006733249, 0, 0, -6.678056e-06, 
    -2.191134e-05, 0, 0, 0, 0.002011491, -5.176498e-05, -0.0004175072, 
    -6.058219e-05, 0.0009399068, 0.03879155, 0.01678846, 0.01262068, 
    0.001779242, 0, -2.127269e-05, 0, 0.0002798422, 0.01268291, 0.0424176, 
    0.03902155, 0.00774631, 0.0004306951,
  0, -1.629526e-06, -2.020738e-05, -2.971199e-07, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, -6.856222e-05, 0.002237587, 0, -2.550745e-05, 0, 0, 0, 0, 0, 
    -5.28491e-05, 0.002033807, 2.627006e-05, 0.004181318,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2.373168e-05, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, -8.127922e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.000795333, 
    -4.804352e-06, -1.200804e-05, 0, 0, 0, 0, 0, 0, 0, -6.057048e-05, 0,
  0, -2.893036e-05, 0, 0, -4.817276e-06, 0.003706376, 0.0006307059, 
    0.003357474, 0.002925615, 0.00157219, 0, 0, 0, 0.00589588, 0, 
    0.0005815882, 0.002364642, -3.25667e-06, 0, 0.004637642, -0.0001759585, 
    -1.809721e-05, -4.745926e-06, -2.7072e-05, 0, 0.007156576, 0.006085088, 
    0.00155117, 0.001769453,
  0.007227246, 0.008101043, -6.656576e-06, 0.01608799, 0.01946511, 0.0345266, 
    0.004840577, 0.003257046, -3.261319e-05, 2.998858e-06, 6.607141e-06, 
    0.006160913, 0.009668539, 0.005757808, 0.007304405, 0.008897091, 
    0.02150267, -1.962604e-05, 0.008334426, 0.02975969, 0.008195847, 
    0.007598162, 0.002229878, 0, 0.0127663, 0.02279166, 0.01840604, 
    0.006604852, 6.584277e-05,
  0.007690849, 0.0257948, 1.429942e-05, 0.03750616, 0.03700092, 0.003143454, 
    0.001546957, 0.0005776675, -2.550642e-07, -1.416161e-06, 0.003788394, 
    0.002709551, 0.003796239, 0.01536, 0.005952184, 0.05067482, 0.03449533, 
    0.03944916, 0.04777927, 0.04954788, 0.0148644, 0.001617744, 0.001787334, 
    0.01237649, 0.01622377, 0.1084595, 0.1327584, 0.02424241, 0.01264149,
  0.001090842, 0.01803783, -2.040001e-05, 0.005288909, 0.02474215, 0.0489381, 
    0.001036274, 0.00641484, 3.813496e-05, 7.941765e-07, 3.538068e-08, 
    0.01327586, 0.002698792, 0.00757942, 0.04226121, 0.06530717, 0.1009753, 
    0.1575678, 0.1056462, 0.04263894, 0.005282363, -2.912972e-05, 
    6.961871e-07, 0.006673899, 0.1143146, 0.1542938, 0.08776989, 0.02815145, 
    0.03167351,
  -6.60945e-07, 0.02742456, 0.03752741, 0.009256982, 0.03108388, 0.1042023, 
    0.07555123, 0.02276989, 0.0003673148, 0.0001411967, 0.01340215, 
    0.1651161, 0.09079289, 0.1290398, 0.119077, 0.08238672, 0.04978929, 
    0.001407497, 0.001762925, 5.066571e-05, 2.528663e-06, -2.830844e-07, 
    0.007280028, 0.4117788, 0.3276178, 0.0560516, 0.009058029, 0.006611784, 
    1.080636e-05,
  0.02782741, 0.4236027, 0.4617591, 0.001085752, 0.001405828, 0.06065343, 
    0.02766468, 0.08247162, 0.3814572, 0.2136742, 0.04635586, 0.1708949, 
    0.1090152, 0.1005699, 0.02181438, 8.322915e-06, 0.001461211, 0.01058052, 
    0.0002991931, 0.01652474, 8.582738e-07, 0.0001009176, 0.05917021, 
    0.3223016, 0.1002506, -0.0001872682, 0.01732626, 0.03235278, 1.135234e-05,
  0.09693069, 0.03603126, 0.02027971, 0.01737429, -0.0002360055, 0.001638163, 
    0.1949173, 0.1155525, 0.1421779, 0.153901, 0.1741362, 0.2756733, 
    0.3052783, 0.2178029, 0.3061426, 0.2096094, 0.0987168, 0.229668, 
    0.1636052, 0.03940717, 0.1045801, 0.1661924, 0.2453499, 0.2130278, 
    0.08636944, 0.1216356, 0.2113858, 0.181463, 0.1250327,
  0.02132734, 0.0005808569, -3.088277e-07, 0.03931636, 0.001508389, 
    0.02778614, 0.1046293, 0.01225851, 0.06611724, 0.00367159, 0.04244088, 
    0.1162828, 0.06850621, 0.01686865, 0.0243066, 0.06198048, 0.03929891, 
    0.1149625, 0.03030269, 0.03685702, 0.1285082, 0.02393663, 0.08293466, 
    0.0774167, 0.1333542, 0.09086684, 0.1223432, 0.08194117, 0.08018584,
  -4.39364e-05, 0.0004226215, -7.727382e-05, 6.21118e-05, 0.0019762, 
    -5.928838e-05, 0.0009189793, 0, -5.590013e-06, 0.01171873, 0.008818273, 
    0.1232511, 0.09715598, 0.06636781, 0.05479868, 0.1508081, 0.09009838, 
    0.07417782, 0.009196036, 0.02628302, 0.001367895, 0.05929639, 
    0.009627185, 0.1453826, 0.2072016, 0.08987822, -8.964436e-05, 
    0.0004981254, -1.541613e-06,
  0.01884119, 0.01117302, 6.848543e-05, 0, 0.0001039133, 0, -3.036667e-05, 0, 
    0.00146531, -3.257086e-05, 0.004392687, 0.09505755, 0.1049228, 0.1086014, 
    0.09829614, 0.1129205, 0.1087605, 0.04247093, 0.006089588, 9.40038e-05, 
    5.872241e-07, 0.02079781, 0.01345483, 0.009412672, 0.1509153, 0.02461775, 
    0.008125768, 0.01071884, 0.002200697,
  0.002333881, 0.01133558, -5.776052e-05, 0.00142004, 0, -1.261707e-10, 
    0.001894505, -0.0001150928, -1.669159e-05, 0, 0, 0.004216847, 0.01254745, 
    0.02134423, 0.002478523, 0.02109393, 0.06940535, 0.0667676, 0.0220476, 
    0.008752389, -3.162377e-05, 0.002641008, 0, 0.005098197, 0.02088063, 
    0.08799847, 0.07790595, 0.02762744, 0.009691602,
  3.750041e-06, -3.477437e-05, -1.624052e-05, -4.321315e-05, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, -6.088441e-06, 0.0006999261, 0.01907823, 0.001128063, 
    -0.0001705549, 0, 9.564106e-10, -7.906859e-11, 0, -4.651871e-05, 
    0.006889272, 0.01218781, 0.005943584, 0.006365536,
  -2.568306e-06, 0, 0, -3.103535e-05, -8.820713e-06, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.0002653598, -2.980185e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -0.0001000629,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0.0001126778, 0, 0, 0, 0, -3.203877e-05, 0.001303329, 0, -1.409163e-08, 0, 
    0, 0, 0, -1.156194e-05, -1.839784e-05, 0, 0.0005929187, 0.004073989, 
    -2.66675e-05, -7.992642e-05, 0, 0, 0, 0, 0, 0, -1.288625e-05, 
    0.001302916, 1.424058e-06,
  -8.600312e-05, 0.002879662, -2.50422e-10, 0.002432615, 0.001111046, 
    0.01049223, 0.009400349, 0.02336172, 0.01616231, 0.005197256, 
    0.004812911, -2.066462e-07, -2.078682e-07, 0.01592059, -2.964191e-06, 
    0.004008732, 0.01412573, 0.001899787, 8.61977e-05, 0.007534239, 
    0.001196792, 0.0005098435, 0.00270242, 0.003285266, 0.001010628, 
    0.0146189, 0.02254861, 0.020966, 0.01573912,
  0.01198843, 0.02787684, 0.01382851, 0.02783288, 0.0341581, 0.09388094, 
    0.01885338, 0.009858187, 0.009394729, 0.001522066, 0.002105055, 
    0.01114924, 0.01288763, 0.01348811, 0.02597441, 0.01738661, 0.04564488, 
    0.02278238, 0.02715891, 0.05331931, 0.01166047, 0.02599419, 0.003567394, 
    0.0004898785, 0.03064491, 0.06053086, 0.05920389, 0.02360861, 0.0111242,
  0.1442795, 0.12014, 0.0006925526, 0.1013228, 0.1027721, 0.05596712, 
    0.01451363, 0.01156093, 0.006372031, 0.0009471236, 0.01463893, 
    0.01428469, 0.01139756, 0.06746738, 0.02727902, 0.04903131, 0.05837103, 
    0.08010654, 0.1731202, 0.1789124, 0.1336486, 0.08314828, 0.04760943, 
    0.07740074, 0.03530291, 0.1154416, 0.1696469, 0.09145054, 0.06675019,
  0.00297471, 0.02486623, 0.04943646, 0.01302795, 0.0263453, 0.04088845, 
    0.003610602, 0.002435229, 1.450757e-05, 1.591274e-07, -7.767e-07, 
    0.01565776, 0.0005580705, 0.01355802, 0.06127937, 0.06297143, 0.121814, 
    0.1465265, 0.09546885, 0.06067665, 0.01887801, 0.0004730199, 
    1.875325e-07, 0.000215068, 0.07430492, 0.2205099, 0.07153489, 0.03869397, 
    0.02971913,
  -5.772644e-08, 0.01751463, 0.01581275, 0.004293337, 0.02891347, 0.08192154, 
    0.0472018, 0.01535471, 0.0003657402, 4.460059e-05, 0.01046728, 0.1345461, 
    0.08911414, 0.1127847, 0.08743765, 0.05794965, 0.0369058, 0.001042527, 
    0.001483273, 3.508811e-06, 6.210323e-07, -4.085778e-08, 0.001066656, 
    0.322265, 0.2837463, 0.05758401, 0.001253578, 0.0002229159, 5.157467e-06,
  0.007272589, 0.4039142, 0.3970867, 6.621162e-05, 0.0004589287, 0.04846312, 
    0.009657832, 0.0595758, 0.2998291, 0.1612985, 0.01726002, 0.1327861, 
    0.08514794, 0.08683908, 0.01163148, 8.749301e-06, 8.844979e-05, 
    0.005242162, 0.003674072, 0.006437737, 1.094441e-08, 1.974173e-05, 
    0.005884397, 0.2904998, 0.06583309, -4.18296e-05, 0.01382572, 0.01533048, 
    -5.199982e-06,
  0.054948, 0.008462191, 0.007121268, 0.06612445, -0.0001302074, 
    0.0001141467, 0.1338235, 0.08165587, 0.1333092, 0.1320014, 0.1376875, 
    0.2478198, 0.2709397, 0.1825243, 0.2495406, 0.1561266, 0.07585776, 
    0.1970091, 0.1333534, 0.03079511, 0.06588928, 0.1229969, 0.1944833, 
    0.1723161, 0.05641809, 0.09683571, 0.1623949, 0.1215471, 0.1033025,
  0.07274907, 0.007075236, 0.0009245132, 0.04590921, 0.004721183, 0.01638859, 
    0.1015632, 0.008840165, 0.06345708, 0.002709366, 0.03176167, 0.1165812, 
    0.06491967, 0.008353089, 0.01376702, 0.04242786, 0.02090819, 0.09953129, 
    0.02994878, 0.0258578, 0.1022247, 0.01197846, 0.067147, 0.0456001, 
    0.07781042, 0.07303642, 0.1104598, 0.08209716, 0.1354722,
  0.04643588, 0.05223541, 0.03665446, 0.0180293, 0.0233507, 0.02051983, 
    0.04240057, -2.704292e-09, -0.0004190379, 0.02932711, 0.006645971, 
    0.1057332, 0.1006774, 0.05603663, 0.05141873, 0.1413561, 0.1435985, 
    0.1199548, 0.06974535, 0.05353956, 0.03795728, 0.09019666, 0.04535659, 
    0.1801313, 0.1855819, 0.1145856, 0.03031624, 0.03396842, 0.01667448,
  0.04983805, 0.02542237, 0.02328041, -6.120213e-07, 0.002039386, 
    -1.285606e-06, 0.0008342382, 1.151749e-06, 0.01509318, 0.009450105, 
    0.0395234, 0.146874, 0.1668991, 0.159127, 0.1654966, 0.1816496, 
    0.1542364, 0.1825782, 0.06428349, 0.01260587, 0.0007896189, 0.02866524, 
    0.02949915, 0.04415355, 0.2027774, 0.1828251, 0.08961881, 0.04185426, 
    0.01369082,
  0.0263685, 0.03173088, 0.002930152, 0.003394079, 3.366574e-05, 
    0.0002447917, 0.004140487, 0.001708196, -4.939558e-05, 0, 0, 0.007027445, 
    0.007036131, 0.02241368, 0.01762306, 0.05611641, 0.1156381, 0.2230077, 
    0.07834657, 0.01375617, 0.0001350778, 0.005654135, 4.472047e-05, 
    0.01808425, 0.03146385, 0.1689228, 0.1619342, 0.08442163, 0.05430273,
  -2.195516e-05, 0.00195909, 0.008888017, 0.001602339, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, -0.0001886728, 0.01111894, 0.005691266, 0.07732888, 0.005783006, 
    0.0005588108, 0.002652896, 0.001250315, -7.18022e-08, 0, 0.001045732, 
    0.01386775, 0.01617171, 0.01351274, 0.007792898,
  0.003461816, 3.348381e-05, -5.893687e-05, 1.657661e-05, 0.0009637137, 
    -2.629235e-07, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0.0001425791, 0.004453013, 
    0.003909148, 0.003635485, -7.781184e-08, -7.166162e-06, 0, 0, 0, 0, 0, 0, 
    0.003199061,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.948631e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 6.944002e-05, 0, 0, 0,
  0.004819674, -4.94686e-05, 1.043529e-07, 1.637895e-06, 0, -0.0001634817, 
    0.00201298, 0.001916671, 0.00231098, 0.001452328, 0.0003085662, 
    0.002407486, 0, 0.0006570228, -5.836031e-05, -2.523685e-05, 0.006004216, 
    0.01130627, -8.956092e-05, 0.002577939, 0.0004071954, -4.44865e-05, 
    -7.70363e-05, 0, 0, 0, -5.822828e-05, 0.006984119, 0.01114218,
  0.03323768, 0.01933958, 0.01159393, 0.01427195, 0.01705297, 0.03388786, 
    0.05583064, 0.1068946, 0.07353968, 0.06482574, 0.02329493, -0.000203181, 
    0.004980431, 0.0317204, 0.01144006, 0.01090625, 0.03517194, 0.03489733, 
    0.03787866, 0.03889379, 0.009485046, 0.003376927, 0.01133459, 
    0.007664854, 0.003283121, 0.03376466, 0.08379944, 0.09911854, 0.04028513,
  0.0432969, 0.08454116, 0.09446225, 0.1094077, 0.1136143, 0.1651951, 
    0.1045442, 0.1241961, 0.07791213, 0.03128974, 0.02269509, 0.0410797, 
    0.03827015, 0.0465018, 0.04992843, 0.09238747, 0.07481126, 0.07848331, 
    0.1424062, 0.1128011, 0.09394797, 0.1121375, 0.05310669, 0.004950103, 
    0.07827707, 0.1003874, 0.08572628, 0.08368652, 0.03509214,
  0.170658, 0.07986108, 0.1073592, 0.07926821, 0.1040608, 0.05459855, 
    0.008364167, 0.01829118, 0.0190979, 0.006908237, 0.02787296, 0.03290664, 
    0.04925733, 0.1069672, 0.09902486, 0.08628297, 0.1111801, 0.1351784, 
    0.1955808, 0.1940581, 0.1500663, 0.0905179, 0.04874921, 0.04476603, 
    0.03801729, 0.09154043, 0.1548257, 0.1025215, 0.1295253,
  -8.820771e-05, 0.01253457, 0.04517744, 0.004834575, 0.01758031, 0.03240276, 
    -0.0008382612, 0.0006105812, -3.573707e-05, 1.972495e-07, -7.333203e-06, 
    0.01413224, 0.003437875, 0.02793504, 0.07899339, 0.1041078, 0.1317638, 
    0.12551, 0.06135117, 0.05180541, 0.008444253, -0.0001192002, 
    -8.055096e-08, 0.001606129, 0.05627091, 0.2113786, 0.04999089, 
    0.04256932, 0.03449589,
  -8.790285e-06, 0.01176013, 0.008453167, 0.00516537, 0.02747558, 0.0693986, 
    0.0336715, 0.01144229, 0.0002476092, 2.353752e-05, 0.01198892, 0.1074062, 
    0.0945331, 0.1056365, 0.07872812, 0.04564852, 0.03481192, 0.0008806337, 
    0.0005985305, 4.513411e-07, 2.156938e-07, -1.05814e-08, 2.938791e-05, 
    0.2601617, 0.2678149, 0.05758723, -0.0002191489, 2.045415e-06, 
    1.758762e-06,
  0.005011471, 0.3777144, 0.314098, 6.880157e-05, 0.0001205454, 0.04782583, 
    0.009229674, 0.06568663, 0.2570243, 0.1222121, 0.006266338, 0.1074543, 
    0.07863835, 0.0709248, 0.01078377, 3.912064e-06, 3.566104e-05, 
    0.0001410584, 6.808584e-05, 8.774643e-05, -7.794813e-09, 1.810523e-06, 
    0.001788152, 0.2577117, 0.04818101, 1.784157e-06, 0.01544708, 0.01620954, 
    -3.451971e-06,
  0.03940233, 0.003795958, 0.008426346, 0.05558887, -0.0001064542, 
    0.0007381511, 0.1207599, 0.07707606, 0.1285921, 0.1220458, 0.1052688, 
    0.2294669, 0.2436668, 0.1736249, 0.223092, 0.1224677, 0.0730896, 
    0.1855972, 0.1277557, 0.02809732, 0.05835875, 0.1076326, 0.1554, 
    0.1583979, 0.05129338, 0.08769264, 0.1241391, 0.09394153, 0.09182382,
  0.06891813, 0.007846132, -1.650096e-05, 0.05134358, 0.002575402, 
    0.01628389, 0.0952277, 0.006825252, 0.05791708, 0.001639761, 0.02649649, 
    0.1136119, 0.06611898, 0.008818309, 0.01081628, 0.04075762, 0.01664775, 
    0.0719488, 0.01911506, 0.02249156, 0.09075829, 0.01239563, 0.05814304, 
    0.03554769, 0.04890291, 0.05470988, 0.09092672, 0.05872404, 0.1054805,
  0.06353232, 0.06309404, 0.03522011, 0.02729819, 0.06085268, 0.0486719, 
    0.04422026, 0.0001127601, 0.0003060634, 0.050922, 0.009649179, 0.1048447, 
    0.1080131, 0.03851078, 0.04752323, 0.1210722, 0.09844281, 0.1074039, 
    0.05395793, 0.04724709, 0.06492557, 0.08074901, 0.04100748, 0.1579441, 
    0.1482915, 0.09210669, 0.01428792, 0.02099003, 0.04753463,
  0.1300811, 0.1213195, 0.07490213, 0.006354052, 0.03276289, 0.03606579, 
    0.003042254, 0.0002926448, 0.03324479, 0.06610058, 0.07733172, 0.1646449, 
    0.1952149, 0.1991205, 0.1907533, 0.1965352, 0.1895814, 0.252429, 
    0.06134152, 0.03548545, 0.002883083, 0.09038944, 0.08706465, 0.07868944, 
    0.1980634, 0.1561416, 0.08519567, 0.05378215, 0.0884219,
  0.0935254, 0.07179455, 0.04753358, 0.0680422, 0.0336526, 0.001506387, 
    0.009269623, 0.005145157, 0.0001026183, 0, 0.01248957, 0.0218324, 
    0.02344078, 0.04823169, 0.02347649, 0.1355633, 0.1690466, 0.3442525, 
    0.1253007, 0.03177927, 0.04493567, 0.05189927, 0.009056651, 0.03690003, 
    0.09742257, 0.2220709, 0.2069363, 0.1617547, 0.1059932,
  0.01998912, 0.0299809, 0.03759331, 0.01710192, 0.001225572, -2.147618e-05, 
    3.509319e-05, 0.001051317, 0, 0, 0, 0, -0.0004503627, 0, -2.907186e-05, 
    0.05130258, 0.03266778, 0.1936368, 0.06314599, 0.03065761, 0.03702148, 
    0.03190562, -1.554338e-06, 0, 0.01076935, 0.02700559, 0.0263088, 
    0.03389438, 0.02226966,
  0.01014336, 0.004301839, 0.003114497, 0.003988693, 0.001694662, 
    1.211793e-05, 0, -3.908605e-05, 0, 0, 0, 0, 0, 0, 0, -2.051654e-06, 
    0.007068919, 0.02757545, 0.0409168, 0.05552804, 0.03369017, 0.0008872714, 
    0, 0, 0.00212303, -2.802814e-06, 1.979713e-09, 0.0007982557, 0.007032488,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0.0009702836, 0, 0, 0, 0, 0, 0, 0, 0, 0, -3.418508e-06, -3.897262e-05, 0, 
    0, -8.374931e-06, 0, 0, 0, 0, 0, 0.0001637469, 0, 0, 0, 0.0001753191, 
    0.0001544585, 0, 1.997094e-05, 0.0008896661,
  0.07879104, 0.02802825, 0.01582905, 0.0002128605, -2.649917e-05, 
    0.001713003, 0.004967208, 0.01554808, 0.02100443, 0.02094062, 0.03175529, 
    0.02521291, 0.01764113, 0.01680403, 0.02515888, 0.002077352, 0.01232537, 
    0.03472816, 0.05957786, 0.07151663, 0.03331776, 0.02369933, 0.007470416, 
    -4.200122e-06, 0.006463772, 0.01341877, 0.01460532, 0.07200135, 0.0898724,
  0.05225783, 0.04736837, 0.07220235, 0.08548858, 0.09684516, 0.09732813, 
    0.1185143, 0.1882848, 0.1685832, 0.1007201, 0.06353268, 0.07307624, 
    0.06361654, 0.1092855, 0.06603733, 0.1174446, 0.1657611, 0.1165472, 
    0.1085097, 0.1161937, 0.04774794, 0.04034501, 0.04487748, 0.01684668, 
    0.01839979, 0.145746, 0.2153941, 0.1436432, 0.0942561,
  0.1268834, 0.1119025, 0.1054334, 0.1241215, 0.1105418, 0.1370815, 
    0.1078469, 0.1286001, 0.07384349, 0.03487264, 0.06835742, 0.07125488, 
    0.08936793, 0.1253446, 0.09190989, 0.1100407, 0.1457812, 0.1686313, 
    0.1704693, 0.1221727, 0.08454727, 0.1437922, 0.1055372, 0.03098302, 
    0.156615, 0.1256878, 0.1433406, 0.09785195, 0.06993268,
  0.14018, 0.06171982, 0.08081555, 0.06547764, 0.07751659, 0.04665484, 
    0.01132261, 0.01745012, 0.01636882, 0.01548904, 0.01238155, 0.04662403, 
    0.0671555, 0.1048624, 0.095149, 0.07728042, 0.1176938, 0.129481, 
    0.1744422, 0.1618956, 0.1374748, 0.06495659, 0.04346355, 0.01951304, 
    0.0314203, 0.07612251, 0.1319875, 0.08153107, 0.1418479,
  0.0001313937, 0.001691034, 0.03167742, 0.0007936795, 0.01547268, 
    0.02817864, -0.0001482785, -1.333066e-05, 0.001537522, 9.817276e-07, 
    -1.740256e-05, 0.01487098, 0.01421439, 0.01699476, 0.08725165, 
    0.09496769, 0.1276753, 0.1098759, 0.04836682, 0.05043266, 0.00383398, 
    0.001656726, -7.832958e-09, 0.00121984, 0.04148769, 0.1985514, 
    0.04449729, 0.04533179, 0.04525688,
  0.002415237, 0.009301614, 0.00554796, 0.002914724, 0.04090775, 0.06142474, 
    0.04119939, 0.007724488, 0.001219461, 2.546704e-05, 0.01829173, 
    0.09450592, 0.09833719, 0.112962, 0.06764515, 0.03725249, 0.02828904, 
    0.000911736, 0.001940157, 1.014177e-07, 9.349522e-09, 7.24136e-09, 
    9.79939e-06, 0.1834147, 0.2215343, 0.06378889, 0.0002174786, 
    3.982648e-08, 2.732243e-07,
  0.01485632, 0.3351238, 0.2114692, 0.0001232595, 9.214641e-05, 0.04813721, 
    0.01326537, 0.07285099, 0.2009061, 0.08179045, 0.007417543, 0.08189578, 
    0.06305891, 0.05477477, 0.008599176, 3.023975e-06, -1.485502e-06, 
    -0.0001003759, 9.102346e-06, -3.489682e-06, -4.592257e-09, 3.074215e-07, 
    0.0001419263, 0.200331, 0.03087485, 1.630953e-06, 0.02608491, 0.02767078, 
    -1.682395e-05,
  0.03338264, 0.003136446, 0.00948979, 0.04621346, -3.728069e-05, 
    0.001749449, 0.1091238, 0.06408951, 0.1079954, 0.1117963, 0.09072831, 
    0.2115013, 0.2090217, 0.1495344, 0.1737954, 0.09164672, 0.07817873, 
    0.2181588, 0.1155339, 0.02196715, 0.04451513, 0.0888358, 0.1161411, 
    0.1138376, 0.04868948, 0.08111927, 0.08237464, 0.05917036, 0.0827137,
  0.05606981, 0.006449059, 8.944395e-06, 0.04992353, 0.0014282, 0.01542369, 
    0.07879683, 0.005428925, 0.04534606, 0.00150367, 0.02734321, 0.1044596, 
    0.05583347, 0.009321918, 0.008863742, 0.03389751, 0.01342761, 0.02942235, 
    0.0185915, 0.02022406, 0.07666402, 0.01670194, 0.04433311, 0.02879115, 
    0.03344303, 0.05018928, 0.0674019, 0.0388637, 0.05916143,
  0.06064368, 0.04739077, 0.04701116, 0.0401292, 0.04947359, 0.03743308, 
    0.03033081, 0.0009784477, 0.01049027, 0.08417846, 0.010259, 0.1046576, 
    0.08826087, 0.03693224, 0.0311071, 0.1111431, 0.07377149, 0.07483263, 
    0.03679135, 0.04489576, 0.06302468, 0.05985652, 0.03907157, 0.1438873, 
    0.1258399, 0.07043618, 0.006039096, 0.01083333, 0.0250538,
  0.200512, 0.1455692, 0.07647753, 0.03594272, 0.109006, 0.09265514, 
    0.008057779, 0.06443663, 0.1096857, 0.1019464, 0.1066498, 0.1542286, 
    0.2047555, 0.2113865, 0.2111529, 0.1855604, 0.2078932, 0.2357123, 
    0.04712974, 0.04915344, 0.04687594, 0.09862919, 0.1410717, 0.09482846, 
    0.1896758, 0.1413829, 0.06818277, 0.05170056, 0.1116739,
  0.1443023, 0.1756753, 0.06792141, 0.08458062, 0.1227894, 0.09303654, 
    0.03799962, 0.01004435, 0.000849396, 2.941382e-09, 0.02703083, 
    0.03334847, 0.05015621, 0.07733241, 0.105419, 0.1778112, 0.1866549, 
    0.3502144, 0.1324541, 0.07295451, 0.07604495, 0.1492649, 0.08439726, 
    0.1144191, 0.1463708, 0.1936739, 0.1871031, 0.1427434, 0.1199405,
  0.07511081, 0.1151468, 0.1616979, 0.1636166, 0.07638544, 0.02882802, 
    0.04634701, 0.01176373, -1.076377e-05, 0, -1.668421e-09, 0, 0.003479881, 
    -4.787765e-06, 0.02573431, 0.113242, 0.07742464, 0.2729509, 0.1729214, 
    0.05895167, 0.06359947, 0.05608002, 0.01758434, 0.001024893, 0.04968136, 
    0.09898891, 0.1025169, 0.07750934, 0.06934606,
  0.04314004, 0.0864993, 0.03921156, 0.07359743, 0.04531528, 0.01067675, 
    0.0101258, 0.0002068315, 0, 0, 0, 0, 0, 0, 0, 0.008487873, 0.06439367, 
    0.09533471, 0.1212202, 0.1011422, 0.07641496, 0.03478659, 0.004917292, 
    -9.035629e-05, 0.005158446, 0.0001378985, -4.464146e-06, 0.02266543, 
    0.015353,
  -1.956008e-05, 0, -8.830906e-05, -1.697385e-05, 5.528163e-05, 
    -3.171595e-05, 1.271041e-06, 0, 0, 0, 0, 0, 0, 5.697395e-06, 
    -0.0001314437, 0.009701145, 0.01828459, 0.01248615, 0.009519844, 
    0.003808597, -9.32827e-05, 0, 0, 0, 0, 0, 0, -5.000555e-05, 1.16149e-05,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -1.250689e-06, 0.0001673163, 0, 0,
  0.06353374, 0.02393301, 0, 0, 0, 0, 0, 0, 0, 0, -3.418508e-06, 9.71811e-05, 
    0, -7.379648e-06, 0.002394269, -0.0007382133, 0.01024314, 0.005860687, 
    3.161594e-05, -3.006474e-05, 0.002029029, 0.01660007, 0.01036467, 
    -0.0003371493, 0.002633864, 0.0004514472, 0.0004154742, 0.02942537, 
    0.03561658,
  0.1561843, 0.1279249, 0.08645015, 0.03484046, 0.0225933, 0.02976494, 
    0.04380775, 0.05765748, 0.09503865, 0.1222147, 0.1003143, 0.08644541, 
    0.07235454, 0.06291691, 0.06808119, 0.04986924, 0.08369001, 0.2382498, 
    0.1800426, 0.1522131, 0.08420708, 0.06040798, 0.01579485, 0.05416798, 
    0.05305514, 0.0329976, 0.08791483, 0.1557216, 0.1730919,
  0.09247393, 0.09582456, 0.1013025, 0.124512, 0.1615966, 0.147976, 0.158471, 
    0.1914136, 0.2027721, 0.1136678, 0.1047586, 0.08317263, 0.09366512, 
    0.1135757, 0.1043647, 0.1804004, 0.1864113, 0.1532652, 0.1526784, 
    0.1762771, 0.1430254, 0.1180632, 0.1284663, 0.03605618, 0.0782279, 
    0.2510778, 0.2806595, 0.1526267, 0.1281582,
  0.1228324, 0.116753, 0.1056638, 0.1232817, 0.1079852, 0.1103543, 
    0.09864383, 0.1103481, 0.06522643, 0.03802672, 0.08160944, 0.0741037, 
    0.1070225, 0.1385873, 0.1146496, 0.104992, 0.1316974, 0.1485729, 
    0.1461703, 0.1085038, 0.0762298, 0.133483, 0.11617, 0.04453935, 
    0.1446111, 0.1138013, 0.1307189, 0.07916896, 0.06980284,
  0.1135685, 0.05282732, 0.04598068, 0.06595583, 0.06342957, 0.04651661, 
    0.008132763, 0.003857618, 0.005110033, 0.0009782737, 0.0001549186, 
    0.05124836, 0.07427108, 0.09956317, 0.05714221, 0.07479377, 0.1161002, 
    0.1260005, 0.1606196, 0.1274452, 0.1104374, 0.04704769, 0.02316985, 
    0.005676877, 0.03786888, 0.07379272, 0.1056891, 0.05507679, 0.1428732,
  0.003034428, -0.000353204, 0.01358667, 0.0001490961, 0.01110427, 
    0.02088611, -7.695962e-06, 2.62106e-07, 0.00442762, 0.000102948, 
    0.000682337, 0.01237866, 0.02200506, 0.0008025628, 0.06665218, 
    0.09211228, 0.122376, 0.08998037, 0.03873735, 0.03291148, 0.003319792, 
    0.0002215596, -2.489151e-09, 0.0007889949, 0.02873422, 0.1541436, 
    0.06033529, 0.04640417, 0.03380036,
  0.005580705, 0.009879513, 0.003878205, 0.004398639, 0.04019822, 0.06117307, 
    0.05805631, 0.001646033, 0.002082732, 0.0002473411, 0.02470588, 
    0.07600304, 0.08524153, 0.1067448, 0.04775378, 0.02653646, 0.02345469, 
    0.001557186, 0.0002883865, 4.327465e-08, 5.227012e-09, 7.933286e-10, 
    1.900418e-05, 0.1161485, 0.1651317, 0.0609878, 1.325749e-05, 
    1.402675e-07, 5.153318e-08,
  0.03085258, 0.3054682, 0.1384455, 7.75466e-05, 8.604572e-05, 0.0499327, 
    0.01055309, 0.07922034, 0.1509212, 0.07477067, 0.008925192, 0.05111049, 
    0.0409957, 0.04429924, 0.00567764, 8.841515e-07, -5.668875e-05, 
    0.0002211478, 4.51835e-07, -4.851896e-08, -9.905876e-10, 1.619449e-06, 
    0.0001052261, 0.1373213, 0.02007473, 2.623417e-05, 0.02678139, 
    0.01869711, -5.347889e-06,
  0.03171886, 0.005184165, 0.01149892, 0.04146799, 9.039284e-05, 0.002427968, 
    0.08107913, 0.04988754, 0.0969248, 0.1001199, 0.06423818, 0.186497, 
    0.1798747, 0.1499809, 0.1486758, 0.06518184, 0.08876189, 0.226235, 
    0.09796299, 0.02123732, 0.0336062, 0.07797959, 0.1050818, 0.06680865, 
    0.04984028, 0.07173967, 0.06040769, 0.03700441, 0.06734103,
  0.03578896, 0.002139953, -3.742236e-05, 0.03760323, 0.0005535462, 0.017193, 
    0.05043342, 0.008517916, 0.02934739, 0.001957431, 0.0269692, 0.1043333, 
    0.05021752, 0.006875375, 0.01080952, 0.02391368, 0.01519221, 0.0240946, 
    0.02616495, 0.02702855, 0.0626936, 0.0177432, 0.02536662, 0.01832137, 
    0.01854482, 0.04262308, 0.05506321, 0.02838024, 0.03710504,
  0.04691216, 0.03514475, 0.03720538, 0.02215054, 0.03815179, 0.02870839, 
    0.02185777, 0.001539272, 0.03975688, 0.07881764, 0.01194162, 0.08869093, 
    0.09004857, 0.03280963, 0.03632896, 0.09731245, 0.04446756, 0.0618519, 
    0.02209156, 0.03568185, 0.05490365, 0.04480619, 0.04606863, 0.1246678, 
    0.1037004, 0.07194802, 0.004000802, 0.007359501, 0.01380865,
  0.1828379, 0.1463865, 0.06047031, 0.04652539, 0.0874596, 0.07067599, 
    0.01817847, 0.1057028, 0.1492884, 0.1330561, 0.101571, 0.1368095, 
    0.1948939, 0.2081416, 0.2266684, 0.1816902, 0.1788543, 0.2157226, 
    0.03924046, 0.04863289, 0.08145858, 0.09840428, 0.1431688, 0.09095356, 
    0.1685541, 0.1375141, 0.07406955, 0.03890497, 0.104386,
  0.1510392, 0.1772628, 0.07354455, 0.0657314, 0.126212, 0.1167271, 
    0.1521969, 0.01312903, 0.007131487, 0.01784866, 0.1515148, 0.08127146, 
    0.09265395, 0.08545467, 0.1639875, 0.2415946, 0.1849544, 0.3326584, 
    0.1404167, 0.09739936, 0.08743499, 0.1704097, 0.1751656, 0.2030324, 
    0.1569219, 0.1628263, 0.1747505, 0.1638123, 0.1308412,
  0.1586093, 0.2481216, 0.1949701, 0.2064425, 0.1798682, 0.147026, 0.1653971, 
    0.05806973, 0.01489452, -0.0001169714, 0.02821842, -0.0005776915, 
    0.00289091, 0.02261222, 0.05634919, 0.1982542, 0.1714859, 0.3186604, 
    0.1919854, 0.07006348, 0.1090913, 0.07622662, 0.0717543, 0.06699491, 
    0.1306865, 0.1830088, 0.1479686, 0.1107003, 0.1373697,
  0.1755245, 0.203145, 0.2030386, 0.2170086, 0.1914781, 0.06684983, 
    0.02971191, 0.01461512, -0.0001414125, 0, 0.008515801, 0.004251572, 
    0.009950335, 0.004777827, 0.0008029504, 0.08457518, 0.1400468, 0.1218041, 
    0.1504307, 0.1568121, 0.1083616, 0.05099303, 0.04281148, -0.0004631804, 
    0.03799295, 0.004178385, 0.002149111, 0.1584529, 0.1283917,
  0.008006669, 0.009025078, 0.007742705, 0.001658105, 0.004271837, 
    0.006668825, 0.00615063, 0.002914533, 0.0001362301, 0, 0, -3.602694e-05, 
    0.0007587543, 0.01312804, 0.03688987, 0.04154146, 0.02232854, 0.01643128, 
    0.01309975, 0.01462344, 0.003982798, -0.0001577434, 0, -1.575015e-05, 
    -6.137484e-06, -1.389422e-05, 0, 0.0005328847, 0.002355988,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    4.373517e-05, -0.001033565, 0.03598047, 0.02568573, 0,
  0.1223514, 0.04712442, 0.01011255, 0.0006380793, -3.697379e-05, 
    -2.025425e-05, -0.0004066465, -3.810067e-05, -0.000118136, 0, 
    0.000226181, 0.0002381161, -0.00108934, 0.008972338, 0.01383896, 
    0.02114358, 0.03619846, 0.02721771, 0.01855948, 0.02067329, 0.02133183, 
    0.04139683, 0.04095863, 0.02543119, 0.0342601, 0.07340024, 0.09023687, 
    0.07181858, 0.1082628,
  0.2338834, 0.1881254, 0.1677793, 0.09098093, 0.08039209, 0.0765681, 
    0.1163617, 0.1394196, 0.1639568, 0.1642675, 0.1336232, 0.1510766, 
    0.1355885, 0.1232717, 0.09884937, 0.06977896, 0.1243599, 0.2936273, 
    0.235868, 0.217139, 0.1742585, 0.1406059, 0.1250629, 0.1893016, 
    0.1889694, 0.18777, 0.1911806, 0.2408613, 0.2613593,
  0.09097651, 0.08116375, 0.1217355, 0.1481647, 0.170866, 0.1589448, 
    0.1836238, 0.1959088, 0.2229639, 0.1249074, 0.1379106, 0.1116152, 
    0.1196911, 0.1480386, 0.1233609, 0.155939, 0.1600611, 0.1555434, 
    0.1690017, 0.1904564, 0.1657215, 0.1427956, 0.1664786, 0.08379615, 
    0.1140603, 0.2479407, 0.2649589, 0.146597, 0.1058772,
  0.107005, 0.1149706, 0.08892567, 0.1207474, 0.111494, 0.09916054, 
    0.1002253, 0.09613679, 0.05932018, 0.03577414, 0.05259769, 0.07112226, 
    0.1032538, 0.1429482, 0.1208727, 0.1020508, 0.1101641, 0.1401613, 
    0.135598, 0.08800116, 0.0713703, 0.1300395, 0.126461, 0.05994502, 
    0.1311678, 0.1053701, 0.1263977, 0.06519496, 0.0601736,
  0.08244328, 0.03091047, 0.06073391, 0.07128824, 0.05544247, 0.06414217, 
    0.01127041, -5.159445e-05, 4.980206e-05, -2.26286e-05, 0.001386769, 
    0.05934287, 0.0740178, 0.09256298, 0.06196715, 0.07820381, 0.1294118, 
    0.1241552, 0.1464049, 0.1041495, 0.09823193, 0.02391102, 0.01000059, 
    0.001070963, 0.04298927, 0.07300216, 0.09774432, 0.04192494, 0.1110094,
  0.001336297, -0.0002030537, 0.00406792, 0.0001084504, 0.01347957, 
    0.01788064, -2.536565e-05, 2.315984e-08, 0.001131527, 0.01382828, 
    0.00079114, 0.01106429, 0.04059142, -0.0008378258, 0.0518495, 0.08701251, 
    0.1194824, 0.07681729, 0.04906931, 0.03964543, 0.001270336, 0.0003666664, 
    5.814283e-10, 3.769594e-05, 0.02549334, 0.137551, 0.07055366, 0.04158899, 
    0.01308509,
  0.01228121, 0.005966699, 0.00932974, 0.003589444, 0.04942262, 0.06754303, 
    0.07620639, 0.0007617549, 0.003662078, 0.001030637, 0.02842461, 
    0.06813992, 0.09534083, 0.106402, 0.04534281, 0.01736465, 0.02455586, 
    0.000881409, 4.979169e-06, 3.225599e-08, 4.082301e-09, 0, 4.970042e-06, 
    0.08354373, 0.1127421, 0.05908559, 1.747019e-06, 4.720416e-07, 
    -3.089339e-07,
  0.03325825, 0.2778928, 0.09667919, 0.000309228, 0.001881707, 0.05096665, 
    0.007717255, 0.09716417, 0.1076211, 0.08629048, 0.00898447, 0.04193648, 
    0.02322759, 0.032747, 0.003950168, -1.80039e-06, -0.0001839215, 
    -0.0001157443, -1.155196e-05, 1.005243e-06, 2.738013e-09, 8.706168e-07, 
    0.002724601, 0.1020145, 0.01363668, 6.418203e-05, 0.022662, 0.03113988, 
    2.000608e-05,
  0.02269315, 0.01402263, 0.01202823, 0.04033354, 0.0001203346, 0.003437008, 
    0.07998285, 0.03613956, 0.07523777, 0.08712582, 0.05113776, 0.1473045, 
    0.159429, 0.1511189, 0.1301121, 0.05138446, 0.09253778, 0.2198372, 
    0.0947948, 0.0242805, 0.06029698, 0.06758134, 0.0923636, 0.03772808, 
    0.04406878, 0.05979662, 0.06256687, 0.02105435, 0.04588338,
  0.01353129, 0.0001877988, 1.08202e-05, 0.02479565, 0.0003677116, 0.0174308, 
    0.02453723, 0.003982448, 0.01459455, 0.001317641, 0.0293257, 0.1035622, 
    0.05111149, 0.005291441, 0.01112661, 0.01442379, 0.01996934, 0.01766637, 
    0.03001919, 0.03374479, 0.05510827, 0.01819824, 0.01445039, 0.01907744, 
    0.01233617, 0.03589759, 0.04088325, 0.02358762, 0.02769471,
  0.02559061, 0.03013958, 0.03600147, 0.02176579, 0.03234125, 0.02024241, 
    0.01789435, 0.003065549, 0.08451699, 0.07544919, 0.02059451, 0.08808073, 
    0.09256108, 0.02920565, 0.02437043, 0.0773571, 0.03156263, 0.04557375, 
    0.01634637, 0.02995755, 0.04691934, 0.03525383, 0.04913751, 0.102426, 
    0.08055432, 0.05979027, 0.003149794, 0.003475433, 0.009230991,
  0.1811244, 0.1682303, 0.04990474, 0.03820937, 0.07126939, 0.05573256, 
    0.05365205, 0.1075227, 0.1426139, 0.1184187, 0.0995467, 0.1191743, 
    0.1868532, 0.1841941, 0.2223903, 0.1855011, 0.1672926, 0.2035723, 
    0.03291461, 0.04297232, 0.09267386, 0.09426067, 0.1315798, 0.07982013, 
    0.1629024, 0.1122108, 0.07527743, 0.02810648, 0.1169544,
  0.1709168, 0.1971614, 0.06024136, 0.05635052, 0.1220726, 0.1033796, 
    0.1873956, 0.06827354, 0.04163897, 0.1169095, 0.2332309, 0.1464621, 
    0.1147663, 0.1260496, 0.1664569, 0.2737805, 0.1967952, 0.3307373, 
    0.1118587, 0.1003504, 0.08939511, 0.1796721, 0.1956569, 0.2165602, 
    0.1581527, 0.147754, 0.1710455, 0.1648345, 0.1511773,
  0.2080915, 0.2466742, 0.1751521, 0.1763884, 0.2243097, 0.1589994, 
    0.2159294, 0.17055, 0.06102363, 0.02734568, 0.0391577, 0.06396287, 
    0.01461608, 0.06584828, 0.09980212, 0.2922455, 0.2390588, 0.3518705, 
    0.2177365, 0.09662689, 0.1312073, 0.07688436, 0.1218528, 0.1025581, 
    0.2540922, 0.2430336, 0.2101851, 0.2397708, 0.2154774,
  0.2452923, 0.2014731, 0.2359373, 0.2346393, 0.2509518, 0.1623898, 
    0.1685091, 0.05017594, 0.005759988, 0.01039604, 0.02184008, 0.03833346, 
    0.06016435, 0.006814146, 0.01649629, 0.1891643, 0.220727, 0.1651879, 
    0.1737718, 0.1871109, 0.1517727, 0.09005862, 0.06763688, 0.02070022, 
    0.1745264, 0.0150679, 0.004135749, 0.223479, 0.207124,
  0.08018532, 0.09011235, 0.1063806, 0.1120896, 0.08309749, 0.02882805, 
    0.03788756, 0.02598342, 0.001174701, 0.006474266, 0.02135899, 0.04800432, 
    0.08478766, 0.1364774, 0.1644213, 0.1560087, 0.07669447, 0.06106672, 
    0.04357281, 0.01323161, 0.0131989, 0.05823822, 0.007099607, -0.004840795, 
    0.001368158, 0.0005676339, -0.003320933, 0.03740597, 0.129012,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  -0.0002600058, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3.862797e-06, 
    -2.941477e-05, 0, 1.900451e-08, 0, 0, 0, 0, 0, 0, 0.02524723, 0.03188253, 
    0.0340972, 0.08929046, 0.07047957, 0.006908427,
  0.2259685, 0.1108621, 0.04661576, 0.02152749, -0.0003773262, 0.0001225096, 
    0.0252098, -5.000743e-05, 3.876296e-05, -0.0004397384, 0.00309068, 
    0.003243922, 0.004747651, 0.03912864, 0.03391152, 0.07443532, 0.08609481, 
    0.06986587, 0.05105301, 0.04472946, 0.03227055, 0.0695051, 0.08269319, 
    0.07714002, 0.1605188, 0.192604, 0.213164, 0.2013229, 0.2377642,
  0.2552706, 0.1974581, 0.1783304, 0.1294609, 0.1370996, 0.1641748, 
    0.2022534, 0.2105183, 0.216462, 0.2137594, 0.1804899, 0.1708327, 
    0.2083355, 0.1887395, 0.115974, 0.1158027, 0.1333532, 0.3037711, 
    0.2525103, 0.2281203, 0.2093265, 0.2041194, 0.1796768, 0.236763, 
    0.2287195, 0.2126365, 0.2177778, 0.2461106, 0.2934343,
  0.09344848, 0.06790499, 0.1036523, 0.1656406, 0.1924451, 0.173756, 
    0.1677773, 0.2034394, 0.2171207, 0.137258, 0.1507216, 0.133699, 
    0.1166966, 0.1603203, 0.1110878, 0.1249789, 0.1554528, 0.1571825, 
    0.1472779, 0.1746594, 0.1501732, 0.1334746, 0.1568015, 0.1023087, 
    0.1154602, 0.2271682, 0.2311305, 0.149243, 0.08199634,
  0.09543779, 0.1030081, 0.07881729, 0.1075274, 0.1115928, 0.08983988, 
    0.09339935, 0.09952608, 0.06006378, 0.03041694, 0.04069503, 0.07469926, 
    0.1017836, 0.1254084, 0.1238424, 0.1150709, 0.08379859, 0.1240055, 
    0.1234016, 0.06487194, 0.07649565, 0.1184791, 0.09934101, 0.06899862, 
    0.1276526, 0.1091463, 0.1217681, 0.06988499, 0.0707845,
  0.07584538, 0.02633808, 0.08276553, 0.0767741, 0.06226635, 0.05392933, 
    0.0006091786, 0.0001128667, -9.379965e-06, 4.151648e-07, 0.01203074, 
    0.07081155, 0.0698057, 0.08627851, 0.06141888, 0.07967628, 0.1295715, 
    0.1127492, 0.1299357, 0.08093493, 0.1018749, 0.01698306, 0.001446049, 
    0.0001134147, 0.0457736, 0.07043456, 0.09898359, 0.03310381, 0.1229507,
  -2.565118e-05, 0.001025958, 0.005104928, 5.738394e-05, 0.01406861, 
    0.008110788, 5.335601e-07, 2.026695e-08, 0.004544896, 0.01242165, 
    0.0008401184, 0.005079276, 0.04281908, 4.296496e-05, 0.03651722, 
    0.08536038, 0.09858873, 0.06436718, 0.05012794, 0.03922087, 3.333111e-05, 
    3.921553e-06, 4.393023e-09, -9.69645e-05, 0.01737596, 0.1283252, 
    0.05318883, 0.0376178, 0.002953199,
  0.01024706, 0.006417965, 0.00476737, 0.0021599, 0.04393224, 0.07625466, 
    0.101579, 0.001123188, 0.004869006, 0.001735529, 0.03115663, 0.06182238, 
    0.08433533, 0.1238737, 0.0552437, 0.01341341, 0.02542634, 0.0009014224, 
    0.0008274269, 4.081572e-08, -2.572093e-10, 0, 2.045568e-06, 0.05810691, 
    0.07319433, 0.02261552, 3.918962e-06, 2.215536e-07, 2.355233e-05,
  0.03712481, 0.271827, 0.0813691, 0.002964445, 0.01238284, 0.05222254, 
    0.01003991, 0.1147674, 0.09162619, 0.07264644, 0.01302715, 0.02154885, 
    0.01803854, 0.02345176, 0.00302697, 2.295068e-05, 0.0008427492, 
    0.000108467, -1.691237e-05, 5.056889e-07, 1.151467e-07, 4.846324e-07, 
    -5.197895e-05, 0.08403199, 0.009816726, 2.140418e-05, 0.01414817, 
    0.04894614, 0.0007738433,
  0.0165837, 0.02083238, 0.01134553, 0.06578024, 0.001494088, 0.003436285, 
    0.07211777, 0.02552076, 0.07958823, 0.07087705, 0.05580924, 0.1228903, 
    0.1490433, 0.1507028, 0.1223275, 0.05669513, 0.09241801, 0.2299288, 
    0.09932311, 0.04868013, 0.07030176, 0.05960526, 0.0803744, 0.02097317, 
    0.04091524, 0.06137995, 0.05916636, 0.01330138, 0.03093874,
  0.004647234, 2.437776e-05, -8.792042e-05, 0.009548403, 0.0001503163, 
    0.01757429, 0.01349866, 0.004990789, 0.005194872, 0.005790676, 
    0.03587859, 0.09480884, 0.05216428, 0.006264569, 0.01451169, 0.008934643, 
    0.02545314, 0.01139521, 0.02961176, 0.03661771, 0.04705719, 0.02237047, 
    0.009590775, 0.01689728, 0.008965716, 0.03183217, 0.02424188, 0.02410175, 
    0.008164376,
  0.01460383, 0.02595088, 0.03644557, 0.02601229, 0.03390952, 0.01461497, 
    0.01696377, 0.007614092, 0.1122987, 0.07134453, 0.01998813, 0.06754096, 
    0.1005681, 0.04048957, 0.02921905, 0.07844321, 0.02345166, 0.05014515, 
    0.01729717, 0.02904248, 0.01839734, 0.03471006, 0.04537934, 0.08006407, 
    0.07227076, 0.05143044, 0.002436297, 0.001169512, 0.007839127,
  0.1626744, 0.1721922, 0.04293945, 0.02356694, 0.06739123, 0.05030818, 
    0.07744269, 0.1021092, 0.1371169, 0.1071148, 0.08720864, 0.09173905, 
    0.1848875, 0.181114, 0.2027132, 0.1854694, 0.1582108, 0.193421, 
    0.02288767, 0.0407385, 0.06928374, 0.08988485, 0.1290807, 0.08133478, 
    0.1593538, 0.09758458, 0.04228723, 0.01945283, 0.1332744,
  0.1714694, 0.1974475, 0.05729107, 0.05133061, 0.09916855, 0.09053767, 
    0.1936043, 0.1747059, 0.1181947, 0.1777287, 0.2599722, 0.1591378, 
    0.1187655, 0.1264532, 0.1706355, 0.2675196, 0.1887785, 0.2945721, 
    0.09813456, 0.09514841, 0.1119878, 0.1842205, 0.2120986, 0.2320316, 
    0.1779817, 0.1529451, 0.1802, 0.1569251, 0.1645732,
  0.240652, 0.2277031, 0.1411209, 0.1572774, 0.2307293, 0.1451219, 0.1950765, 
    0.252279, 0.1275615, 0.1045762, 0.1061971, 0.1159304, 0.1544756, 
    0.1730079, 0.1247004, 0.3040084, 0.288679, 0.3471559, 0.2566642, 
    0.111342, 0.1473925, 0.1482042, 0.1492144, 0.25156, 0.3317352, 0.2765087, 
    0.2377555, 0.2312093, 0.2581907,
  0.2515466, 0.1993886, 0.2492114, 0.243993, 0.2565412, 0.2080131, 0.277263, 
    0.1876031, 0.06339519, 0.03509669, 0.02148725, 0.1420914, 0.1143152, 
    0.02675537, 0.06057843, 0.2307708, 0.306103, 0.2061005, 0.204267, 
    0.2197457, 0.1790592, 0.1042594, 0.1374562, 0.07015911, 0.2351043, 
    0.04259851, 0.01229405, 0.2585516, 0.1853083,
  0.1875323, 0.1902606, 0.1772446, 0.1975018, 0.2077555, 0.1700664, 
    0.09196276, 0.04862218, 0.02430641, 0.06885735, 0.1386243, 0.2392695, 
    0.2848497, 0.2527499, 0.2195164, 0.1682937, 0.0905481, 0.07139537, 
    0.08517608, 0.0428069, 0.03190029, 0.09567691, 0.1224426, 0.03963868, 
    0.08950444, 0.01526275, 0.00131329, 0.1146317, 0.2402297,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  -0.00105901, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.002018493, 0.009831729, 
    0.006581591, 0.0002105939, -9.161779e-05, -1.008231e-12, 0, 0, 0, 
    0.001832002, 0.09578917, 0.1153807, 0.1126553, 0.1539999, 0.1141486, 
    0.03097654,
  0.3269029, 0.166958, 0.1004471, 0.07668895, -0.0007316504, 0.002427216, 
    0.05959895, 0.0001954403, 0.00389508, -0.0026224, 0.009179311, 0.010342, 
    0.009453758, 0.08683407, 0.09963597, 0.136494, 0.1788177, 0.1263314, 
    0.1217173, 0.1174321, 0.0721553, 0.1019255, 0.1123584, 0.1489295, 
    0.210992, 0.2676493, 0.271259, 0.252346, 0.3119009,
  0.2418174, 0.202824, 0.2084968, 0.1604189, 0.1736242, 0.2062328, 0.2320022, 
    0.2291424, 0.2140842, 0.2328405, 0.2173178, 0.2012139, 0.2348522, 
    0.2115172, 0.158248, 0.1917377, 0.1235226, 0.3008753, 0.2630578, 
    0.241494, 0.2546544, 0.241254, 0.2767464, 0.3069256, 0.2770993, 
    0.2208549, 0.2359489, 0.2376232, 0.2502035,
  0.09264588, 0.06900609, 0.08973976, 0.1503024, 0.2046107, 0.1808134, 
    0.1505731, 0.2038231, 0.2007636, 0.1356878, 0.1463487, 0.1220137, 
    0.1146045, 0.1664668, 0.09861646, 0.1159005, 0.1378796, 0.1413349, 
    0.1341225, 0.1710313, 0.1552766, 0.1336542, 0.1720131, 0.1075548, 
    0.1000382, 0.2171562, 0.2233512, 0.1415972, 0.08066282,
  0.08639742, 0.1021867, 0.06427651, 0.09343087, 0.1101912, 0.08978166, 
    0.09086461, 0.1071851, 0.05593526, 0.0160921, 0.03951413, 0.08024821, 
    0.09415858, 0.1125958, 0.13075, 0.1181033, 0.07964133, 0.104582, 
    0.1142147, 0.05123942, 0.09438872, 0.1136614, 0.1158797, 0.08214148, 
    0.1237257, 0.1248072, 0.1026778, 0.06584885, 0.07176946,
  0.06014534, 0.02637376, 0.08378998, 0.08750467, 0.06404339, 0.04832219, 
    -9.728091e-06, 0.001060622, -3.128664e-05, 2.104406e-07, 0.02541532, 
    0.09454697, 0.06351452, 0.07891219, 0.05526262, 0.07218429, 0.1219197, 
    0.1083584, 0.1173888, 0.05684245, 0.0933133, 0.01437396, 3.3039e-05, 
    -1.067467e-05, 0.04920549, 0.08296472, 0.1076166, 0.03500611, 0.1641583,
  0.001111876, 0.02733912, 0.01002484, 2.316013e-05, 0.01605218, 0.001323104, 
    4.665598e-09, -1.156513e-06, 0.001308765, 0.00635324, 0.00498852, 
    0.0120417, 0.04299029, 0.001893926, 0.02331478, 0.0669289, 0.08451515, 
    0.05791855, 0.05883738, 0.04273792, 0.00015313, 1.804164e-07, 
    3.215996e-09, -7.824436e-05, 0.01705682, 0.1266367, 0.05223551, 
    0.01069578, 0.001520028,
  0.003903583, 0.03369104, 0.005032727, 0.002082335, 0.03335103, 0.07416636, 
    0.1198906, 0.001576699, 0.005432476, 0.002586307, 0.03129029, 0.06161161, 
    0.09232963, 0.1366406, 0.0651923, 0.009783543, 0.02543897, 0.00161101, 
    0.0003364184, -4.469743e-09, 1.469368e-10, -4.254091e-12, 1.375009e-06, 
    0.04961623, 0.05127923, 0.004953647, 5.055757e-06, 1.454747e-07, 
    -1.883651e-06,
  0.04726302, 0.2619175, 0.08290739, 0.008617451, 0.01391151, 0.02628531, 
    0.009915277, 0.1283857, 0.07665671, 0.04724666, 0.02925275, 0.0122116, 
    0.01747003, 0.02137618, 0.003815154, 0.000628928, 0.004346486, 
    0.0001076107, -2.821247e-05, 1.04249e-06, 1.77602e-07, 1.164145e-07, 
    0.0008336871, 0.06108272, 0.005747904, 0.0002660638, 0.008716348, 
    0.06767793, 0.004024752,
  0.01118204, 0.01930049, 0.009522732, 0.08699156, 0.001056408, 0.00288306, 
    0.0625043, 0.01715886, 0.07961816, 0.0479883, 0.05673321, 0.1080724, 
    0.1376176, 0.15862, 0.1092444, 0.06496447, 0.08239661, 0.2095593, 
    0.1148169, 0.05461015, 0.09711003, 0.06213245, 0.09030961, 0.01594588, 
    0.04350218, 0.07309501, 0.07690665, 0.01032971, 0.0273386,
  0.001826589, 2.574933e-06, -7.575017e-08, 0.00861309, 9.093208e-05, 
    0.01682106, 0.008147436, 0.0052294, 0.002870767, 0.001290588, 0.04004573, 
    0.09782849, 0.05721755, 0.0138784, 0.02452185, 0.007101862, 0.03020611, 
    0.008131287, 0.02570574, 0.03140224, 0.03304375, 0.02703168, 0.007398659, 
    0.0138567, 0.007498721, 0.03116923, 0.0222655, 0.02631559, 0.003180931,
  0.01205362, 0.03511795, 0.03655021, 0.029872, 0.03636963, 0.008674596, 
    0.01723031, 0.04549636, 0.1248601, 0.06690996, 0.02934288, 0.0646445, 
    0.1031379, 0.02572996, 0.02273989, 0.082814, 0.01702976, 0.04931671, 
    0.02046538, 0.02569194, 0.01310127, 0.03271763, 0.05409999, 0.0674114, 
    0.06933245, 0.04609773, 0.001716684, 0.0008218519, 0.009417263,
  0.1442587, 0.1636377, 0.03907334, 0.01822213, 0.0641885, 0.04739276, 
    0.07561797, 0.08980106, 0.124865, 0.1122095, 0.07044882, 0.0588378, 
    0.1531947, 0.1704671, 0.1923629, 0.1825609, 0.1554161, 0.1827063, 
    0.01649129, 0.03939993, 0.05156036, 0.09348793, 0.1423989, 0.07811227, 
    0.1709515, 0.07392794, 0.0248611, 0.0199785, 0.124839,
  0.1649836, 0.1755261, 0.05712126, 0.04825692, 0.09038317, 0.06561507, 
    0.1837085, 0.2438714, 0.1793105, 0.1998481, 0.2425817, 0.1661746, 
    0.128834, 0.1459937, 0.1855875, 0.3005691, 0.2251556, 0.273494, 
    0.08988757, 0.08491222, 0.111429, 0.1772781, 0.2404829, 0.2479024, 
    0.19779, 0.1568678, 0.1828132, 0.1583443, 0.1512322,
  0.2399873, 0.2127413, 0.1359122, 0.1643452, 0.2181528, 0.1414057, 
    0.2060066, 0.2670955, 0.2342865, 0.1660708, 0.1706434, 0.2104719, 
    0.2485527, 0.1710918, 0.1380126, 0.3357177, 0.2923352, 0.3304856, 
    0.259738, 0.1067402, 0.1570252, 0.1877752, 0.2310755, 0.328728, 
    0.3494942, 0.3031851, 0.2177441, 0.25211, 0.2446804,
  0.2334988, 0.2018531, 0.2727737, 0.2528237, 0.2568502, 0.2133851, 
    0.2970237, 0.2474255, 0.1656243, 0.1206007, 0.05035959, 0.2225177, 
    0.1315188, 0.04235153, 0.07638399, 0.1957455, 0.3126991, 0.214777, 
    0.2070555, 0.2263539, 0.2079316, 0.1136822, 0.1762164, 0.1553124, 
    0.2794297, 0.06695139, 0.06836691, 0.2264228, 0.1821452,
  0.196612, 0.2137786, 0.2024709, 0.2280224, 0.2288056, 0.173057, 0.1464873, 
    0.1267847, 0.1127207, 0.1489364, 0.221495, 0.3097859, 0.3273859, 
    0.2797236, 0.2575242, 0.2275141, 0.1519991, 0.1163056, 0.113466, 
    0.05376057, 0.03336473, 0.1227196, 0.1876805, 0.1017857, 0.2027149, 
    0.07345422, 0.07536488, 0.1480335, 0.2658094,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0.02500182, -6.618957e-06, -2.141559e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.02531112, 0.04296383, 0.008222874, 0.03606141, 0.02554318, 
    0.0004905778, 0, 0, -6.181902e-05, 0.01735619, 0.1948265, 0.1775157, 
    0.2322323, 0.2956519, 0.1510964, 0.04488265,
  0.3529555, 0.1846898, 0.1345829, 0.136168, 0.002632708, 0.01590183, 
    0.1353498, 0.002181873, 0.004772749, 0.009645475, 0.01738394, 0.02185904, 
    0.06766596, 0.2372827, 0.1944392, 0.2724472, 0.2606556, 0.2487577, 
    0.2569475, 0.2259808, 0.1478534, 0.1743874, 0.1665547, 0.1907865, 
    0.2462801, 0.2779644, 0.2861262, 0.2547404, 0.3434406,
  0.2396355, 0.205517, 0.2244674, 0.178511, 0.2361029, 0.2337419, 0.2512346, 
    0.2537163, 0.2242304, 0.239052, 0.2523852, 0.2197587, 0.2342036, 
    0.2398112, 0.2031523, 0.2154096, 0.1324415, 0.2862454, 0.2639798, 
    0.2587782, 0.2440583, 0.2442377, 0.3222598, 0.3256291, 0.2648722, 
    0.2186693, 0.2395925, 0.2295444, 0.2516661,
  0.08441783, 0.0693936, 0.08097373, 0.1383843, 0.196004, 0.1704133, 
    0.1343541, 0.1966869, 0.1843816, 0.1342743, 0.1266149, 0.1014012, 
    0.1028696, 0.1634404, 0.09144316, 0.1077763, 0.1204065, 0.1355358, 
    0.1202169, 0.1746322, 0.1511097, 0.1312128, 0.1640036, 0.1188053, 
    0.09450497, 0.2191351, 0.2030647, 0.1300021, 0.07465962,
  0.07203399, 0.1089013, 0.05131976, 0.08019827, 0.1085411, 0.09917486, 
    0.08411279, 0.1103302, 0.05568823, 0.0166741, 0.04070877, 0.08614168, 
    0.0933347, 0.1206953, 0.1240221, 0.1144595, 0.07728361, 0.1045895, 
    0.09717382, 0.04156104, 0.108042, 0.1089702, 0.1135161, 0.1070207, 
    0.1060941, 0.1247806, 0.09111032, 0.0594501, 0.05472051,
  0.05003101, 0.03006331, 0.08868909, 0.09500921, 0.0606328, 0.04516371, 
    0.0006627659, 0.001572006, 0.0004164717, 1.161445e-07, 0.03621119, 
    0.08233981, 0.06963704, 0.06942467, 0.04654934, 0.05459413, 0.1041577, 
    0.09934714, 0.121354, 0.06299197, 0.06941584, 0.03091646, -1.017835e-05, 
    -3.268807e-06, 0.06140361, 0.08634574, 0.1114277, 0.03261141, 0.1976832,
  0.007646383, 0.05851043, 0.02267867, 3.254719e-05, 0.02040421, 
    0.0003058536, 1.330191e-07, -5.652654e-05, 0.0007590879, 0.006783954, 
    0.01466146, 0.03162364, 0.03995882, 0.0007270625, 0.01494887, 0.05961863, 
    0.06469955, 0.06026668, 0.06559218, 0.04996792, 3.056798e-06, 
    8.908849e-09, 2.328136e-08, -5.367063e-05, 0.02220866, 0.1272542, 
    0.05824251, 0.005946075, 0.007550809,
  0.003112973, 0.04692029, 0.01704353, 0.003422207, 0.02995475, 0.08856942, 
    0.1383472, 0.002527063, 0.008699033, 0.002403252, 0.03198206, 0.07307752, 
    0.09974483, 0.1334272, 0.0713641, 0.007022677, 0.02548519, 0.01111902, 
    0.0001129311, 5.612528e-09, 2.044356e-08, 7.414448e-09, 0.0008270904, 
    0.07373177, 0.04756105, 0.006221453, 4.002183e-06, 1.375779e-07, 
    -4.237279e-06,
  0.07352212, 0.2693551, 0.1104132, 0.006258613, 0.01210084, 0.01389423, 
    0.01064279, 0.1344287, 0.06881233, 0.02279573, 0.02242921, 0.00751197, 
    0.01831296, 0.02054577, 0.002752831, 0.0008438291, 0.00459125, 
    0.002559626, 5.241359e-05, -2.27512e-05, 6.176785e-07, -2.440791e-06, 
    0.007859993, 0.06039074, 0.005356893, 0.0001448845, 0.01046974, 
    0.06537783, 0.003263144,
  0.009262744, 0.0173095, 0.01112903, 0.09909464, 0.000485094, 0.003914819, 
    0.07721224, 0.01626217, 0.0874458, 0.04537214, 0.07213707, 0.1166174, 
    0.1382973, 0.1664239, 0.1084753, 0.06643819, 0.09413915, 0.1922709, 
    0.1230392, 0.0738492, 0.1211788, 0.06748659, 0.0839105, 0.01597038, 
    0.04505452, 0.07294069, 0.0854996, 0.01020083, 0.01898682,
  7.964842e-05, -3.879651e-06, 0.0005184577, 0.01368953, 5.318128e-05, 
    0.0196567, 0.005552032, 0.004281058, 0.002165749, 0.001414166, 
    0.04409348, 0.1121867, 0.07524221, 0.01265272, 0.02825039, 0.005530849, 
    0.01838588, 0.008415272, 0.02100214, 0.05456415, 0.02734692, 0.03560168, 
    0.00618, 0.02076529, 0.008707504, 0.03151783, 0.03562615, 0.02528783, 
    0.00109932,
  0.01561095, 0.04227525, 0.04290075, 0.03589477, 0.04204316, 0.005788571, 
    0.01590085, 0.05371606, 0.1360772, 0.06715681, 0.04916623, 0.1052225, 
    0.08568319, 0.02042377, 0.02597177, 0.09318683, 0.01304133, 0.05136917, 
    0.0236838, 0.02187381, 0.02137859, 0.02862301, 0.06517236, 0.06485835, 
    0.07682076, 0.03169808, 0.0004850282, 0.0006800771, 0.01203782,
  0.155522, 0.1303706, 0.03677774, 0.01769163, 0.05447055, 0.03778171, 
    0.07495675, 0.07984257, 0.1074314, 0.1179732, 0.05843022, 0.03774796, 
    0.1359648, 0.1625386, 0.1952205, 0.1808547, 0.1494065, 0.1711685, 
    0.0133588, 0.0355263, 0.05308562, 0.100827, 0.1310837, 0.07702459, 
    0.1645345, 0.06774551, 0.03112799, 0.01459162, 0.110091,
  0.1650025, 0.1565429, 0.0551344, 0.04735017, 0.06638163, 0.06045619, 
    0.1837388, 0.256597, 0.1928833, 0.1764964, 0.2265004, 0.1684807, 
    0.1319834, 0.164105, 0.1707713, 0.2971171, 0.2142904, 0.2539625, 
    0.07769347, 0.08369139, 0.09899371, 0.1694527, 0.2607397, 0.2873717, 
    0.1722448, 0.1495387, 0.172401, 0.1476219, 0.137986,
  0.237923, 0.2275701, 0.1419093, 0.1596889, 0.1957459, 0.146651, 0.201039, 
    0.2704029, 0.2680154, 0.2269412, 0.2259317, 0.2495508, 0.2906069, 
    0.1675092, 0.1492067, 0.3294649, 0.276361, 0.3231286, 0.258723, 
    0.1097196, 0.1514275, 0.2069973, 0.2266252, 0.3150539, 0.3608856, 
    0.314738, 0.2359273, 0.2437424, 0.2697296,
  0.2149129, 0.2055889, 0.2841034, 0.2292762, 0.2504768, 0.2197667, 
    0.3320134, 0.240447, 0.2840504, 0.2058966, 0.1682903, 0.2664557, 
    0.1043883, 0.0429771, 0.06259234, 0.1761458, 0.3127441, 0.2236601, 
    0.2072217, 0.2293689, 0.2416357, 0.1450577, 0.2414145, 0.234115, 
    0.2770413, 0.155939, 0.2021691, 0.2187202, 0.1620295,
  0.188693, 0.1995675, 0.2049417, 0.2326211, 0.237142, 0.2014658, 0.1572279, 
    0.1521576, 0.1474549, 0.1600685, 0.2163726, 0.290913, 0.280561, 
    0.2412186, 0.2408111, 0.205752, 0.1518233, 0.0899168, 0.09899339, 
    0.1037503, 0.09325836, 0.1803236, 0.2136963, 0.1045361, 0.2131185, 
    0.1113704, 0.1141525, 0.1377937, 0.2848412,
  0.000794057, 0.0004321011, 7.014522e-05, -0.0002918107, -0.0006537666, 
    -0.001015722, -0.001377678, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -0.00177872, -0.001416764, -0.001054808, -0.0006928525, -0.0003308966, 
    3.105929e-05, 0.0003930152, 0.001083622,
  0.02761946, 0.04008167, 0.00136964, 0, 0, 0, 0, 0, 0, 0, 0, 0.0005149216, 
    0.001498018, 0.07492375, 0.04465102, 0.02747609, 0.07361402, 0.08656841, 
    0.04257539, -0.0001154285, -0.0004991622, -0.0006045466, 0.04713182, 
    0.2288737, 0.1836426, 0.2322351, 0.3018312, 0.2425956, 0.07718557,
  0.3526894, 0.1798543, 0.158917, 0.2095964, 0.009888049, 0.04244858, 
    0.1944559, 0.01606549, 0.006831249, 0.04979165, 0.04625062, 0.04472161, 
    0.156907, 0.3005276, 0.2438322, 0.2794189, 0.2723829, 0.2738881, 
    0.2519001, 0.2330205, 0.1613321, 0.1833811, 0.1863762, 0.2333976, 
    0.2646981, 0.2620671, 0.2806203, 0.243215, 0.336787,
  0.2174589, 0.205011, 0.211194, 0.1958418, 0.2805728, 0.2443297, 0.2571866, 
    0.2605401, 0.2200902, 0.2467394, 0.3005285, 0.2467577, 0.2476331, 
    0.2447077, 0.2268541, 0.2247542, 0.1468758, 0.2697589, 0.259563, 
    0.2595558, 0.230831, 0.2322495, 0.320118, 0.3092927, 0.2698632, 
    0.2224655, 0.2359037, 0.2262965, 0.2022392,
  0.09081902, 0.08283918, 0.06747436, 0.1306683, 0.1739117, 0.1512523, 
    0.1293879, 0.1898019, 0.186, 0.1375763, 0.1256995, 0.1232284, 0.1080909, 
    0.1623125, 0.09332012, 0.1075404, 0.1202301, 0.1358654, 0.1328073, 
    0.1795382, 0.1588135, 0.1336624, 0.144191, 0.1245938, 0.08982126, 
    0.2179274, 0.2022814, 0.1188274, 0.05428776,
  0.06110963, 0.1110278, 0.04632967, 0.0718158, 0.1072551, 0.09715301, 
    0.08881439, 0.12311, 0.05472616, 0.02128866, 0.03770972, 0.101738, 
    0.097218, 0.1404867, 0.1250626, 0.1100596, 0.0742972, 0.08544647, 
    0.0947013, 0.05137794, 0.1113665, 0.1095553, 0.1118084, 0.1282363, 
    0.09250192, 0.1523044, 0.09627325, 0.0579078, 0.05623638,
  0.03053913, 0.01202781, 0.08679374, 0.09736198, 0.06203412, 0.0433949, 
    0.001960592, 0.003449955, 0.007744851, -1.34968e-07, 0.02268867, 
    0.06152725, 0.06963667, 0.06122844, 0.04554775, 0.04576061, 0.0833306, 
    0.09094365, 0.1156648, 0.06009032, 0.0725332, 0.05081467, -5.653265e-06, 
    -8.697953e-07, 0.07567611, 0.09511264, 0.1225733, 0.03221549, 0.1980529,
  0.005883462, 0.0282773, 0.0594512, 0.008626492, 0.03137952, 0.000916275, 
    2.510282e-06, -8.659538e-05, -7.016076e-05, 0.003163453, 0.06125836, 
    0.0662636, 0.03726438, 0.0001584249, 0.01032147, 0.06005453, 0.0519118, 
    0.0599947, 0.06335626, 0.05082623, 1.374763e-07, 1.443452e-07, 
    5.13077e-07, -2.65946e-05, 0.03360067, 0.1433474, 0.06332958, 
    0.009210132, 0.01193442,
  0.007466639, 0.06466177, 0.05970209, 0.004237937, 0.02993059, 0.1096726, 
    0.166674, 0.005210401, 0.01237271, 0.003475327, 0.0314523, 0.1026653, 
    0.1237158, 0.1635449, 0.08260377, 0.009929155, 0.0296834, 0.01756959, 
    0.0004671834, 4.559359e-07, 8.964255e-08, 1.520497e-07, 0.00726922, 
    0.09469263, 0.05862598, 0.03351359, 1.639921e-05, 1.633189e-06, 
    -0.0001868794,
  0.06070418, 0.2806258, 0.1599634, 0.006536455, 0.004115471, 0.009559457, 
    0.01485653, 0.1510245, 0.084594, 0.02429125, 0.01941359, 0.008683067, 
    0.03377485, 0.03009914, 0.00282335, 0.0005989897, 0.003309165, 
    0.002662621, 2.781335e-05, 0.0009278631, 2.657866e-06, 0.001242271, 
    0.007747116, 0.07383725, 0.00544881, 0.0008601205, 0.00916366, 
    0.04095722, 0.008499364,
  0.01174672, 0.01946035, 0.0193078, 0.1225999, 0.0003878805, 0.004319044, 
    0.0865786, 0.02541987, 0.09222201, 0.05523863, 0.1085136, 0.1539351, 
    0.152434, 0.1907453, 0.1353705, 0.08669398, 0.1100595, 0.2000768, 
    0.1393723, 0.105276, 0.1427716, 0.07459328, 0.09563431, 0.02314273, 
    0.04921067, 0.08573133, 0.0906534, 0.01623365, 0.01849817,
  0.0006518125, -1.810014e-05, 7.538374e-05, 0.01710041, 5.476553e-05, 
    0.02131301, 0.005870346, 0.004974167, 0.00808942, 0.003373109, 
    0.05138555, 0.135986, 0.08603497, 0.01468412, 0.03861357, 0.006644703, 
    0.01177174, 0.009020785, 0.01169624, 0.04814899, 0.03104245, 0.0516993, 
    0.007396783, 0.03320061, 0.01159366, 0.03641199, 0.0625882, 0.02548489, 
    0.003797722,
  0.01709815, 0.01813739, 0.03589265, 0.03833174, 0.0362967, 0.005876209, 
    0.02239304, 0.06795387, 0.1399068, 0.07494371, 0.06343524, 0.1514157, 
    0.08239641, 0.01846221, 0.02366045, 0.1109611, 0.01609896, 0.0608773, 
    0.01751084, 0.01945129, 0.03318327, 0.02836348, 0.08418505, 0.07310934, 
    0.08748363, 0.02375423, 0.0001471136, 0.001611976, 0.01608019,
  0.1548897, 0.1057881, 0.02918212, 0.01759353, 0.04485229, 0.03425301, 
    0.07814484, 0.07458636, 0.09308489, 0.1197361, 0.04463329, 0.02902662, 
    0.1164137, 0.1509431, 0.1955559, 0.1685818, 0.1540862, 0.1653812, 
    0.01559269, 0.02541293, 0.05266861, 0.1052355, 0.1219866, 0.06298426, 
    0.1576921, 0.06255288, 0.03144621, 0.01695074, 0.1072542,
  0.1625656, 0.1544669, 0.05458293, 0.04598156, 0.05914845, 0.07042481, 
    0.1706761, 0.265569, 0.2108416, 0.1618616, 0.2158198, 0.1691427, 
    0.1327781, 0.1659086, 0.1471198, 0.3384864, 0.2308906, 0.2447439, 
    0.08204433, 0.08288498, 0.09308752, 0.1703263, 0.2669841, 0.3454542, 
    0.1868198, 0.1499327, 0.1708915, 0.1418728, 0.1569157,
  0.2483864, 0.2612615, 0.1392264, 0.1482776, 0.1881799, 0.1631399, 
    0.2037299, 0.2673734, 0.2920462, 0.3212841, 0.2693087, 0.2609681, 
    0.2809566, 0.1476961, 0.173504, 0.3617159, 0.3033286, 0.3483475, 
    0.2579552, 0.1207839, 0.1561279, 0.2164179, 0.2451066, 0.2984093, 
    0.3508039, 0.3353961, 0.2341817, 0.2497634, 0.2453332,
  0.2213687, 0.193061, 0.2613391, 0.2378069, 0.2709322, 0.2195329, 0.3413912, 
    0.2783726, 0.3203548, 0.2065508, 0.1669092, 0.2519538, 0.06878425, 
    0.03900056, 0.04516227, 0.1652822, 0.2982623, 0.2333107, 0.2313164, 
    0.2397752, 0.2490838, 0.2361128, 0.2515046, 0.2524947, 0.2634243, 
    0.202252, 0.3186287, 0.2654513, 0.1724066,
  0.1538554, 0.1882906, 0.2143628, 0.2248313, 0.231305, 0.2179872, 0.1717262, 
    0.1658118, 0.1537413, 0.1549492, 0.1855281, 0.2331579, 0.2045374, 
    0.1688026, 0.1698144, 0.1326429, 0.1046323, 0.05423542, 0.07455081, 
    0.1093386, 0.11542, 0.2466859, 0.2279087, 0.1113786, 0.1832552, 
    0.1399902, 0.1430109, 0.1342938, 0.2715013,
  0.02086262, 0.01861147, 0.01636031, 0.01410916, 0.01185801, 0.009606857, 
    0.007355704, 0.01039827, 0.009474524, 0.008550775, 0.007627026, 
    0.006703277, 0.005779528, 0.004855779, -0.0007775004, -0.0001200121, 
    0.0005374762, 0.001194965, 0.001852453, 0.002509941, 0.003167429, 
    0.005874358, 0.008391771, 0.01090918, 0.0134266, 0.01594401, 0.01846143, 
    0.02097884, 0.02266354,
  0.06077183, 0.0501748, 0.04094445, 0.01330039, -0.0002163705, 0, 0, 0, 0, 
    0, 0.002631771, 0.04709768, 0.002008721, 0.1096057, 0.05402214, 
    0.03911665, 0.09509344, 0.1247465, 0.1324572, 0.05267803, -0.0006494079, 
    0.006214836, 0.09371983, 0.2343724, 0.1781559, 0.2310999, 0.3165978, 
    0.3311682, 0.1234493,
  0.3572952, 0.1822678, 0.1609335, 0.2295346, 0.04145732, 0.09443258, 
    0.2159328, 0.05361039, 0.05600931, 0.07347772, 0.1243719, 0.05070863, 
    0.2356559, 0.2978918, 0.2706795, 0.274625, 0.2792429, 0.2935703, 
    0.2827059, 0.2265109, 0.1801232, 0.1928619, 0.2129841, 0.2419756, 
    0.2854057, 0.2572238, 0.2826747, 0.2579398, 0.3629061,
  0.2047112, 0.1910809, 0.224075, 0.2033648, 0.2776314, 0.2337904, 0.2572717, 
    0.2728604, 0.2314865, 0.2556569, 0.3165686, 0.2490812, 0.2482982, 
    0.2430834, 0.2327922, 0.2540958, 0.1558649, 0.2789133, 0.2735609, 
    0.2775301, 0.2203534, 0.2394007, 0.3193186, 0.3206839, 0.2592595, 
    0.2255005, 0.2182855, 0.2320751, 0.1897958,
  0.08782694, 0.06830267, 0.06593493, 0.1258148, 0.1798149, 0.1554841, 
    0.1316046, 0.1788568, 0.1791046, 0.1360641, 0.113448, 0.09835365, 
    0.0908033, 0.1649836, 0.1084561, 0.1161557, 0.1407292, 0.128922, 
    0.116744, 0.194562, 0.1668918, 0.1595854, 0.165537, 0.1315553, 
    0.07978304, 0.1780471, 0.1865505, 0.1123337, 0.04739652,
  0.06009735, 0.1137704, 0.04345293, 0.07111938, 0.1057328, 0.1009647, 
    0.09251915, 0.1188141, 0.04602297, 0.01605574, 0.04605967, 0.1149936, 
    0.1015009, 0.1277613, 0.1345919, 0.1201055, 0.08172487, 0.06626601, 
    0.1033072, 0.04922483, 0.1231765, 0.1089603, 0.1007356, 0.1494371, 
    0.08520172, 0.1447537, 0.1076374, 0.04682611, 0.05969012,
  0.009346246, 0.0006686652, 0.07909138, 0.1039116, 0.06326839, 0.05128035, 
    0.00399141, 0.004866756, 0.01510003, 2.844075e-06, 0.006867934, 
    0.04923628, 0.06546684, 0.05671567, 0.05684018, 0.05390596, 0.06860895, 
    0.08585942, 0.1190569, 0.06876908, 0.08613136, 0.05195397, 1.027057e-05, 
    7.756432e-08, 0.09334878, 0.1051731, 0.1084416, 0.03071397, 0.1402104,
  0.009161284, 0.01274014, 0.08277175, 0.01250875, 0.03159732, 0.003241892, 
    1.639362e-05, -0.0001240442, 0.0001584946, 0.0008685459, 0.06291284, 
    0.07698051, 0.03129881, 7.763604e-05, 0.0109372, 0.07256382, 0.03795793, 
    0.0563565, 0.0727227, 0.05346301, -6.268732e-07, 2.180349e-07, 
    4.965437e-07, -1.921792e-06, 0.05850916, 0.1663212, 0.05350371, 
    0.02001071, 0.005006666,
  0.01178323, 0.06251119, 0.1653974, 0.006772026, 0.03047, 0.1249437, 
    0.2021171, 0.01171021, 0.01554374, 0.003377629, 0.0368605, 0.12155, 
    0.1319802, 0.1800103, 0.09046747, 0.01368606, 0.03298146, 0.02289712, 
    0.0002723938, 1.12461e-06, 6.520298e-08, 5.287571e-07, 0.005544203, 
    0.1169734, 0.07414363, 0.118882, 4.587711e-05, 3.096805e-05, -8.02045e-05,
  0.07314108, 0.3223689, 0.2009143, 0.006514828, 0.001909834, 0.009641754, 
    0.02182306, 0.159903, 0.1015113, 0.06017108, 0.01810788, 0.01129631, 
    0.04194744, 0.03111742, 0.003395553, 0.0004779418, 0.001891177, 
    0.01827166, -0.0004455975, 0.002367347, 0.02073015, 0.0149243, 
    0.05193923, 0.09922153, 0.008890782, 0.0009869159, 0.008688967, 
    0.03059545, 0.009247858,
  0.01688599, 0.0270482, 0.02795335, 0.1352251, 0.0003846488, 0.003800401, 
    0.09958632, 0.03758894, 0.1077311, 0.07936325, 0.1219483, 0.1573929, 
    0.1643381, 0.1891796, 0.1705924, 0.0971004, 0.1337224, 0.2267497, 
    0.1482518, 0.1137244, 0.1650019, 0.08843058, 0.1058332, 0.02783551, 
    0.05111883, 0.09907345, 0.08961864, 0.04753925, 0.02275711,
  0.008586143, -1.064141e-06, -0.0001030659, 0.01288301, 0.001518697, 
    0.02844751, 0.009655586, 0.005779416, 0.01038045, 0.007562777, 
    0.05119018, 0.1399023, 0.0905047, 0.01787321, 0.05221312, 0.01072545, 
    0.01328804, 0.0113535, 0.005818008, 0.07112786, 0.04219748, 0.06688609, 
    0.009120153, 0.04276194, 0.01215177, 0.03979944, 0.04230148, 0.04207093, 
    0.0009923676,
  0.01191147, 0.004556985, 0.03323742, 0.02925869, 0.0351425, 0.006665682, 
    0.0256543, 0.07389016, 0.144986, 0.07609206, 0.06798945, 0.1754876, 
    0.07570906, 0.01808016, 0.02049084, 0.1196982, 0.02276549, 0.07174229, 
    0.02087383, 0.01914153, 0.05418867, 0.04583159, 0.07724686, 0.08239536, 
    0.1188456, 0.02312942, 0.000353126, 0.004450877, 0.02141044,
  0.1508704, 0.09159687, 0.03063757, 0.02675897, 0.05354373, 0.02256511, 
    0.08211172, 0.0754711, 0.07384338, 0.1142736, 0.0382239, 0.01544882, 
    0.1091161, 0.1552491, 0.1951198, 0.1670877, 0.1541346, 0.1690236, 
    0.01565412, 0.01799768, 0.05098937, 0.1085331, 0.1286207, 0.06174216, 
    0.1579456, 0.09178498, 0.02973194, 0.02430892, 0.1066355,
  0.1760309, 0.1611721, 0.0600947, 0.04780789, 0.04888118, 0.07799939, 
    0.1848465, 0.2799008, 0.2059947, 0.1509705, 0.2106954, 0.174426, 
    0.1308089, 0.1849407, 0.1515903, 0.3224031, 0.2191291, 0.2324787, 
    0.07400414, 0.07865051, 0.09546705, 0.1879085, 0.2596647, 0.3594061, 
    0.1843583, 0.1440819, 0.1826109, 0.1422047, 0.1650653,
  0.2324737, 0.248024, 0.1396399, 0.126479, 0.1862034, 0.1471999, 0.2136018, 
    0.2553746, 0.286437, 0.3621215, 0.2755804, 0.2466247, 0.3043041, 
    0.1349854, 0.1615925, 0.363169, 0.3058965, 0.3444906, 0.2495031, 
    0.1376477, 0.180077, 0.2118024, 0.2565275, 0.3525611, 0.3977709, 
    0.3520835, 0.2430335, 0.270946, 0.297284,
  0.2744348, 0.1930588, 0.2582973, 0.2184221, 0.2903801, 0.2580844, 
    0.2965563, 0.3237065, 0.3159427, 0.1870161, 0.1645043, 0.2113628, 
    0.05618054, 0.02844702, 0.03645394, 0.1463981, 0.3384114, 0.2402563, 
    0.2453885, 0.2590074, 0.2693886, 0.2409961, 0.2736567, 0.2437271, 
    0.2492816, 0.2498503, 0.4002802, 0.2744169, 0.2078843,
  0.1238159, 0.1795181, 0.2194607, 0.1983255, 0.2293098, 0.2360063, 
    0.2083025, 0.1753932, 0.1288562, 0.1296453, 0.1506387, 0.178468, 
    0.1378414, 0.1259405, 0.1268826, 0.09743582, 0.07309794, 0.03166313, 
    0.05865576, 0.1192329, 0.1797798, 0.3023337, 0.2259166, 0.1086123, 
    0.1479069, 0.1331182, 0.1359458, 0.1160513, 0.2536112,
  0.05324561, 0.05175487, 0.05026412, 0.04877337, 0.04728262, 0.04579188, 
    0.04430113, 0.03961232, 0.03708759, 0.03456287, 0.03203814, 0.02951342, 
    0.0269887, 0.02446397, 0.02294404, 0.02463192, 0.0263198, 0.02800767, 
    0.02969555, 0.03138342, 0.0330713, 0.03454504, 0.03687264, 0.03920023, 
    0.04152783, 0.04385542, 0.04618302, 0.04851061, 0.05443821,
  0.09489982, 0.05906706, 0.04875644, 0.04403935, 0.02211795, 0.003767038, 0, 
    0, 0, 0.0006281925, 0.05260986, 0.05489861, 0.01447343, 0.1125931, 
    0.05369511, 0.04351455, 0.08582023, 0.1462739, 0.1790246, 0.1171134, 
    0.0774845, 0.0371461, 0.1619688, 0.252954, 0.1873938, 0.2172042, 
    0.3062699, 0.3365201, 0.1967438,
  0.3596921, 0.1912575, 0.1743017, 0.2279046, 0.1099112, 0.1528421, 
    0.2188397, 0.1355631, 0.1016506, 0.08009731, 0.158197, 0.08168036, 
    0.3058955, 0.3260557, 0.2530781, 0.2611852, 0.2852683, 0.3101826, 
    0.2955582, 0.2335931, 0.1816933, 0.2015897, 0.2317893, 0.2568805, 
    0.2770294, 0.2507036, 0.2558077, 0.2569337, 0.3612663,
  0.1775066, 0.1929166, 0.2181276, 0.2313098, 0.2884464, 0.2483898, 
    0.2659631, 0.2795462, 0.2598572, 0.2597401, 0.3151655, 0.2602979, 
    0.2543969, 0.2544345, 0.2369483, 0.2395927, 0.1579045, 0.2701888, 
    0.2829094, 0.2841776, 0.2213916, 0.2198451, 0.3255069, 0.2985335, 
    0.2379228, 0.2279936, 0.2036341, 0.2463703, 0.1666947,
  0.08918282, 0.06971398, 0.08344489, 0.1165599, 0.1736318, 0.1719529, 
    0.1375513, 0.1826105, 0.1709916, 0.1353587, 0.1470977, 0.1404292, 
    0.1051589, 0.1639192, 0.1038028, 0.1127469, 0.1452242, 0.1313345, 
    0.1165705, 0.1689241, 0.175242, 0.1829222, 0.1695139, 0.139815, 
    0.08326947, 0.1713683, 0.1705403, 0.1065223, 0.05840412,
  0.07802424, 0.114032, 0.04533769, 0.07230221, 0.0980019, 0.09524348, 
    0.09713513, 0.1200098, 0.04567196, 0.02030146, 0.06244627, 0.1126292, 
    0.102879, 0.1308696, 0.1382407, 0.1296203, 0.07489789, 0.07206076, 
    0.0946788, 0.06042631, 0.1184768, 0.1119515, 0.09777521, 0.1708872, 
    0.07866651, 0.1189103, 0.1124701, 0.05753489, 0.05455654,
  0.004610364, -4.828469e-05, 0.05691933, 0.1221882, 0.057071, 0.06552896, 
    0.005620448, 0.009351613, 0.02183737, 1.613978e-05, 0.004132103, 
    0.02981722, 0.05633896, 0.05131362, 0.06060569, 0.0517459, 0.07179498, 
    0.09132443, 0.1178687, 0.06344259, 0.09476043, 0.06214447, 0.0003409111, 
    6.171593e-07, 0.1013539, 0.1028835, 0.1108954, 0.03304007, 0.1185826,
  0.0001884082, 0.004312788, 0.03740655, 0.01424234, 0.02951043, 0.001185228, 
    8.038943e-05, -0.0001465126, 0.000498795, 0.000206898, 0.04234337, 
    0.05523749, 0.01317316, -0.001133349, 0.008387849, 0.07215443, 
    0.04018505, 0.04905755, 0.08447342, 0.05176021, 3.05026e-05, 
    1.983587e-07, 2.999114e-07, -5.276708e-06, 0.07302939, 0.1897281, 
    0.05393681, 0.00709041, 4.761158e-05,
  0.007500618, 0.05101715, 0.2047014, 0.01467161, 0.0302432, 0.1350525, 
    0.2008666, 0.01508692, 0.01982881, 0.002443918, 0.03430124, 0.06041514, 
    0.1059057, 0.1382108, 0.07057556, 0.01791747, 0.04498043, 0.01427854, 
    0.0002487825, 6.216918e-07, 2.599121e-08, 2.120116e-07, 0.0004977575, 
    0.1223874, 0.06973785, 0.2872838, 0.0003798914, 5.65423e-05, -3.037827e-05,
  0.0590958, 0.3899044, 0.191876, 0.008309368, 0.00163492, 0.01437912, 
    0.03054831, 0.1390559, 0.1147826, 0.07324437, 0.0156898, 0.00775714, 
    0.02965747, 0.02022606, 0.00276576, 0.0008644164, 4.087276e-05, 
    0.0150606, 0.007925934, 0.000384061, 0.001622339, 0.001050722, 
    0.05092279, 0.09880958, 0.03721784, 0.0002679759, 0.01107178, 0.02713684, 
    0.00554449,
  0.01235627, 0.03047947, 0.02485148, 0.145467, 0.001721433, 0.005057977, 
    0.1100128, 0.02788807, 0.1017803, 0.06275106, 0.1042201, 0.1204039, 
    0.1152383, 0.1563729, 0.1403109, 0.09842722, 0.1390616, 0.2185282, 
    0.1330861, 0.1265972, 0.168372, 0.07654212, 0.1184119, 0.02886452, 
    0.04702258, 0.09810682, 0.08705094, 0.04229725, 0.02353981,
  0.001516391, 5.457293e-07, -1.841592e-07, 0.01201134, 0.003066135, 
    0.0278351, 0.01151503, 0.006733361, 0.01987857, 0.01088968, 0.05782371, 
    0.1161787, 0.09171112, 0.02219586, 0.06079722, 0.01994825, 0.01433919, 
    0.02190711, 0.005910566, 0.05313031, 0.03829403, 0.08736189, 0.007562293, 
    0.04710478, 0.01484583, 0.04795336, 0.03263976, 0.1006844, 0.000165317,
  0.002491342, 0.004961313, 0.03064337, 0.0409269, 0.03057232, 0.00773908, 
    0.0382263, 0.0601853, 0.1647091, 0.06423523, 0.06087889, 0.1558801, 
    0.07433415, 0.02323911, 0.0220241, 0.1137927, 0.03931634, 0.07940722, 
    0.02358481, 0.0195576, 0.06196893, 0.05918923, 0.07342903, 0.08272602, 
    0.1387578, 0.02475397, 0.002958811, 0.006640965, 0.02993627,
  0.1333528, 0.09323584, 0.02682787, 0.04113925, 0.05380827, 0.01889386, 
    0.08396558, 0.08103147, 0.04747889, 0.1129877, 0.03637414, 0.008364124, 
    0.1116645, 0.1593257, 0.1914762, 0.1594988, 0.1512676, 0.191574, 
    0.01556492, 0.01809804, 0.0498954, 0.09030735, 0.1387817, 0.06190199, 
    0.1632427, 0.07495282, 0.03076578, 0.02804442, 0.1104578,
  0.1552864, 0.1449679, 0.07536182, 0.04875908, 0.04507671, 0.08116988, 
    0.1824666, 0.2990385, 0.1965166, 0.1453554, 0.2070417, 0.1862973, 
    0.1205274, 0.1864313, 0.1729899, 0.3394483, 0.2217062, 0.2371109, 
    0.06528639, 0.08469649, 0.08953345, 0.191675, 0.2911464, 0.3602361, 
    0.1835849, 0.1321795, 0.1703587, 0.1487917, 0.157987,
  0.2503554, 0.2299112, 0.1426123, 0.1300019, 0.2121672, 0.1425122, 
    0.2354984, 0.2368504, 0.3106614, 0.403553, 0.2657507, 0.2634306, 
    0.2896573, 0.1388084, 0.1469055, 0.3626493, 0.3208058, 0.349151, 
    0.2391028, 0.152671, 0.1798661, 0.2088078, 0.2517764, 0.3137598, 
    0.3487707, 0.3650973, 0.2301217, 0.2941632, 0.2500094,
  0.2588335, 0.2191966, 0.2441107, 0.2206305, 0.2478756, 0.2945825, 
    0.2726097, 0.3383731, 0.3070553, 0.1522547, 0.1623304, 0.1873175, 
    0.05056299, 0.04618929, 0.03868343, 0.1479732, 0.3470121, 0.2608631, 
    0.2370937, 0.2541459, 0.2767437, 0.2366892, 0.2734404, 0.2534281, 
    0.3033281, 0.2573591, 0.4354373, 0.2971801, 0.2165401,
  0.1114678, 0.1900897, 0.2267494, 0.1762122, 0.2284134, 0.2293001, 
    0.2402266, 0.1884741, 0.1186745, 0.109477, 0.1380704, 0.1494528, 
    0.09516045, 0.09610356, 0.09590869, 0.07971621, 0.05764133, 0.03271046, 
    0.07843918, 0.1707303, 0.2570195, 0.3455639, 0.2272005, 0.09200585, 
    0.1214718, 0.0901167, 0.1250433, 0.09035243, 0.2341114,
  0.06050764, 0.05912954, 0.05775145, 0.05637335, 0.05499526, 0.05361717, 
    0.05223907, 0.05362068, 0.05161499, 0.0496093, 0.0476036, 0.04559791, 
    0.04359222, 0.04158653, 0.03905246, 0.04067983, 0.0423072, 0.04393457, 
    0.04556194, 0.04718931, 0.04881667, 0.04713921, 0.04889563, 0.05065205, 
    0.05240846, 0.05416488, 0.0559213, 0.05767772, 0.06161011,
  0.1610091, 0.06941463, 0.0526447, 0.05229181, 0.02608456, 0.007193772, 
    9.44417e-05, 0.003173848, 0.00397575, 0.05212599, 0.07840967, 0.06002715, 
    0.0212042, 0.09488881, 0.0446897, 0.04398168, 0.0870089, 0.1472979, 
    0.202226, 0.1401693, 0.1099492, 0.1556444, 0.2090165, 0.26742, 0.2266883, 
    0.2411538, 0.3381155, 0.3214833, 0.2485244,
  0.372654, 0.2180136, 0.1800667, 0.2366283, 0.1797593, 0.2100876, 0.242537, 
    0.2337438, 0.1321367, 0.08431645, 0.1718503, 0.1226297, 0.3003684, 
    0.3466601, 0.2948352, 0.243176, 0.3036635, 0.3482781, 0.2770934, 
    0.2241637, 0.1985969, 0.2236631, 0.2664047, 0.2483398, 0.3009408, 
    0.2634811, 0.2716844, 0.2721579, 0.3658091,
  0.2169834, 0.1925371, 0.2568064, 0.2609513, 0.3185559, 0.253677, 0.2742097, 
    0.3238832, 0.3091362, 0.2801336, 0.338736, 0.2983067, 0.2743118, 
    0.2656586, 0.2436891, 0.2314933, 0.1625599, 0.2428979, 0.2535882, 
    0.2657871, 0.2374263, 0.2499174, 0.3554833, 0.2757404, 0.2150734, 
    0.1943068, 0.217816, 0.2351394, 0.1790245,
  0.09235505, 0.08676101, 0.09660213, 0.1426454, 0.1861163, 0.1605657, 
    0.1487042, 0.1658991, 0.1655695, 0.1443334, 0.1697073, 0.1292202, 
    0.1172975, 0.1598702, 0.1027354, 0.1066216, 0.1566371, 0.1171018, 
    0.1261715, 0.1706025, 0.1793264, 0.1737902, 0.1725551, 0.1429608, 
    0.08299799, 0.1683863, 0.1836326, 0.1206671, 0.07597091,
  0.08828682, 0.1218328, 0.05704239, 0.0707632, 0.1029802, 0.1030536, 
    0.09804136, 0.120725, 0.04742542, 0.03567941, 0.06831234, 0.111013, 
    0.09358744, 0.1399515, 0.1486286, 0.1560958, 0.08207233, 0.06842025, 
    0.09457492, 0.06978491, 0.1160525, 0.1278591, 0.1089642, 0.1901079, 
    0.07941412, 0.1101508, 0.1185671, 0.08785086, 0.05961024,
  0.003864591, -7.034351e-05, 0.03119648, 0.1357588, 0.05426436, 0.07533034, 
    0.01427105, 0.009856758, 0.022451, 3.73843e-05, 0.001511238, 0.01523856, 
    0.04712448, 0.05597037, 0.05599342, 0.04715012, 0.0757929, 0.09663917, 
    0.1374742, 0.0462526, 0.1155279, 0.08079961, 0.0003812283, 1.0833e-06, 
    0.09314565, 0.09582274, 0.1331987, 0.03725989, 0.1319848,
  1.13974e-05, 0.0001968378, 0.005019861, 0.02011087, 0.03368216, 
    0.007311258, 5.27186e-05, 0.0002908415, 2.878413e-05, 4.540458e-05, 
    0.008673977, 0.03369001, 0.001201446, -0.0006736793, -0.001228975, 
    0.06659851, 0.0289779, 0.04663645, 0.09175906, 0.05363451, 0.001198371, 
    1.503663e-07, 1.073493e-07, -9.817259e-06, 0.0635056, 0.2001305, 
    0.02053513, 0.0004757142, 5.60567e-06,
  0.0008759474, 0.02760054, 0.1341711, 0.03202019, 0.0333643, 0.1406336, 
    0.1898047, 0.02119477, 0.02653451, 0.001937099, 0.0324666, 0.0293604, 
    0.08720472, 0.1093191, 0.05455432, 0.02386702, 0.04936835, 0.01285301, 
    0.0008931539, -4.334739e-07, 1.360672e-08, 8.982489e-08, 1.997337e-05, 
    0.08569457, 0.03520843, 0.2034028, 0.0001033339, 3.109779e-07, 
    3.259766e-06,
  0.04620941, 0.3240361, 0.1209174, 0.01156476, 0.002056852, 0.01275906, 
    0.0347022, 0.1112552, 0.1082302, 0.0662, 0.0140538, 0.005942034, 
    0.02518566, 0.0192078, 0.003304094, 0.001360168, 0.0003754485, 
    0.0009494825, 0.003140388, 2.91236e-05, 0.0001956327, 0.01197451, 
    0.04710654, 0.05221405, 0.178837, 4.572193e-06, 0.02128768, 0.01293643, 
    0.002435318,
  0.004942507, 0.01951162, 0.009945526, 0.174894, 0.01200415, 0.009883945, 
    0.1148807, 0.0279313, 0.0849511, 0.05275898, 0.1083648, 0.09364952, 
    0.07304884, 0.1287314, 0.1207747, 0.08907718, 0.1392743, 0.2052028, 
    0.1346734, 0.1547159, 0.1676724, 0.07621706, 0.1236357, 0.02616611, 
    0.03396813, 0.0826514, 0.07987698, 0.021462, 0.01174056,
  5.585459e-05, 2.571378e-07, 7.994183e-08, 0.003241422, 0.000666324, 
    0.02165508, 0.008436332, 0.00958339, 0.0179757, 0.01494397, 0.06137351, 
    0.1049049, 0.07851332, 0.02680431, 0.06554986, 0.02706174, 0.01159774, 
    0.03908154, 0.00351679, 0.04049473, 0.02503848, 0.09472895, 0.009140532, 
    0.04164345, 0.01686569, 0.05278482, 0.009432838, 0.04628446, 0.0001096774,
  0.0001687629, 0.0127524, 0.02775365, 0.04508962, 0.02278719, 0.01026156, 
    0.02556925, 0.04143044, 0.2081615, 0.04303902, 0.06454155, 0.1352726, 
    0.07415883, 0.04060714, 0.03053644, 0.1110618, 0.0508846, 0.08873005, 
    0.02884216, 0.02233598, 0.06349243, 0.04646678, 0.04803428, 0.0767502, 
    0.1135876, 0.02509089, 0.0055227, 0.0108562, 0.03579577,
  0.1211615, 0.09845992, 0.02483614, 0.05543552, 0.06565958, 0.003151489, 
    0.09495027, 0.08166771, 0.02879757, 0.1157192, 0.03923127, 0.01016388, 
    0.1131613, 0.1626579, 0.1853789, 0.1634245, 0.1489169, 0.218216, 
    0.02313761, 0.01631536, 0.06131342, 0.09578912, 0.1261886, 0.05685303, 
    0.1702852, 0.07534291, 0.03216898, 0.03841392, 0.113305,
  0.1747559, 0.1553477, 0.04951573, 0.06233355, 0.05365459, 0.06746532, 
    0.1841983, 0.3429308, 0.1892843, 0.1428841, 0.1930179, 0.1960271, 
    0.1266391, 0.18882, 0.1752079, 0.3421787, 0.2395267, 0.234719, 
    0.06824889, 0.09860563, 0.08599125, 0.1939265, 0.2856455, 0.3658686, 
    0.1796477, 0.1327957, 0.1606661, 0.1555456, 0.1629451,
  0.2297852, 0.2258552, 0.1551605, 0.1466833, 0.1906044, 0.2040757, 
    0.2120463, 0.2361307, 0.3648379, 0.4050236, 0.3344041, 0.2917171, 
    0.2520511, 0.1465828, 0.1594083, 0.3947202, 0.3473851, 0.3431723, 
    0.2561718, 0.1410291, 0.1709691, 0.2266518, 0.2663879, 0.3331241, 
    0.374888, 0.3387478, 0.2245002, 0.2696634, 0.2831329,
  0.3179001, 0.2317808, 0.2589788, 0.2137969, 0.273975, 0.2936206, 0.249437, 
    0.3568249, 0.3007739, 0.1541902, 0.1592699, 0.1740746, 0.04285114, 
    0.09480425, 0.04534556, 0.140829, 0.351432, 0.258826, 0.2333519, 
    0.3127722, 0.2809074, 0.242699, 0.2652825, 0.257217, 0.2985041, 0.270148, 
    0.4208117, 0.2804593, 0.260038,
  0.1298002, 0.2139867, 0.2362804, 0.2064445, 0.2616715, 0.3036139, 
    0.2911625, 0.2401886, 0.1170794, 0.09385916, 0.1396845, 0.1256689, 
    0.08572262, 0.09164283, 0.08532131, 0.07370041, 0.06314813, 0.09731517, 
    0.1830755, 0.2932557, 0.3572158, 0.3689145, 0.2499154, 0.1160471, 
    0.1342899, 0.04432977, 0.1004041, 0.07867205, 0.1929312,
  0.1016514, 0.09597941, 0.09030747, 0.08463552, 0.07896357, 0.07329163, 
    0.06761968, 0.06691708, 0.06508902, 0.06326095, 0.06143289, 0.05960483, 
    0.05777676, 0.0559487, 0.05416377, 0.05815041, 0.06213705, 0.06612369, 
    0.07011033, 0.07409697, 0.07808361, 0.07330251, 0.07681588, 0.08032925, 
    0.08384261, 0.08735598, 0.09086934, 0.09438272, 0.1061889,
  0.2190153, 0.1294457, 0.08029786, 0.05605403, 0.02538587, 0.005678529, 
    0.0004595012, 0.008569361, 0.01256393, 0.07553229, 0.07948762, 
    0.06203558, 0.04183932, 0.07414501, 0.04748517, 0.04617357, 0.08805796, 
    0.1389326, 0.21123, 0.143446, 0.1341234, 0.2383387, 0.2204992, 0.2396822, 
    0.2226119, 0.2773412, 0.3428358, 0.3150208, 0.2836214,
  0.3823265, 0.1870195, 0.1914833, 0.2560827, 0.2517114, 0.2442124, 
    0.2766558, 0.2801161, 0.1386029, 0.1120938, 0.1918592, 0.1204363, 
    0.3031025, 0.3149493, 0.2873525, 0.2364704, 0.278014, 0.3060246, 
    0.2451794, 0.2686244, 0.2200837, 0.197043, 0.2510365, 0.2762868, 
    0.3337601, 0.2703323, 0.2720353, 0.2630835, 0.364261,
  0.214818, 0.2074599, 0.3065498, 0.293448, 0.3499178, 0.2651714, 0.309431, 
    0.3423664, 0.3304687, 0.3295383, 0.3612657, 0.3320201, 0.2762083, 
    0.2860331, 0.2793367, 0.2466473, 0.1794441, 0.229207, 0.2654505, 
    0.294104, 0.2567797, 0.2695435, 0.3193418, 0.2694023, 0.2218077, 
    0.2009764, 0.1906278, 0.2533879, 0.2331508,
  0.09135092, 0.09583125, 0.1045221, 0.1397264, 0.1824114, 0.1637786, 
    0.142532, 0.1748284, 0.1731982, 0.1344662, 0.1758331, 0.1625126, 
    0.1095569, 0.1602854, 0.1100736, 0.1146331, 0.1756113, 0.1377459, 
    0.1497503, 0.1933349, 0.1997766, 0.1675673, 0.1785518, 0.1511236, 
    0.1095716, 0.176371, 0.207633, 0.1134044, 0.08460694,
  0.1273597, 0.1336587, 0.06871882, 0.08961141, 0.1071605, 0.1146438, 
    0.1079785, 0.1239333, 0.06708536, 0.06418789, 0.09206141, 0.1031, 
    0.09582248, 0.1480992, 0.1695807, 0.1715574, 0.1025622, 0.07941208, 
    0.1403836, 0.08021498, 0.1370993, 0.1337542, 0.1264613, 0.1969893, 
    0.0796185, 0.1029087, 0.1439191, 0.1214284, 0.06697545,
  0.005350749, -4.41674e-05, 0.01694882, 0.1220436, 0.05883361, 0.1010042, 
    0.03671163, 0.009614594, 0.0358132, 4.62054e-05, 0.0005069905, 
    0.003869762, 0.04811959, 0.04943385, 0.0534622, 0.05227027, 0.1154972, 
    0.09454829, 0.1413723, 0.03865581, 0.1181657, 0.09087134, 0.0005559579, 
    1.295825e-06, 0.05980467, 0.09895515, 0.1546017, 0.05144455, 0.1497897,
  1.575278e-06, 4.835253e-05, 0.0006045289, 0.01485928, 0.04326186, 
    0.01503211, 0.003107728, 0.002176569, 0.00049843, 7.715007e-06, 
    0.001654249, 0.008845349, 0.000758359, -0.0001654365, -0.001726615, 
    0.06588797, 0.01821232, 0.03941627, 0.106267, 0.06167362, 0.003146129, 
    -3.403974e-07, 4.584291e-08, -7.44154e-06, 0.06447957, 0.2038058, 
    0.01244403, 0.0007975944, 2.858585e-06,
  2.306387e-05, 0.01470156, 0.05657515, 0.05704438, 0.03622133, 0.150097, 
    0.1890865, 0.02823221, 0.02479628, 0.002463351, 0.03074952, 0.01879221, 
    0.09617809, 0.1019258, 0.04531096, 0.02767221, 0.04933091, 0.01995069, 
    0.002031796, 1.250771e-05, 1.255208e-08, 2.744735e-08, 6.835273e-06, 
    0.09400754, 0.02496498, 0.09855936, 0.0001981199, 1.528057e-07, 
    1.873731e-06,
  0.05019939, 0.2854304, 0.07617902, 0.01778529, 0.004328447, 0.0118617, 
    0.03054417, 0.09687752, 0.1155244, 0.05008943, 0.01201958, 0.006522653, 
    0.02278735, 0.02392784, 0.004538942, 0.001167338, 0.006057713, 
    4.123326e-05, 0.0002288551, -3.52207e-06, 0.002288855, 0.02980589, 
    0.03476113, 0.04242748, 0.2173672, 0.0001325772, 0.02950208, 0.01014903, 
    0.0007218617,
  0.002720826, 0.007879286, 0.006950859, 0.2243319, 0.009452193, 0.01390403, 
    0.1372243, 0.03389142, 0.07902282, 0.04926326, 0.1164871, 0.08163819, 
    0.06280974, 0.1055586, 0.1136633, 0.09000991, 0.1393929, 0.1884885, 
    0.1419844, 0.1631783, 0.1760135, 0.08057568, 0.1373813, 0.02500048, 
    0.0246806, 0.06447149, 0.07300124, 0.01323752, 0.00585523,
  9.849928e-06, 8.939709e-08, 4.175383e-08, 0.001666351, 0.001078933, 
    0.02021928, 0.00646849, 0.01092975, 0.02951844, 0.01981601, 0.06836921, 
    0.1040819, 0.07425225, 0.03100249, 0.06779122, 0.04046573, 0.01749929, 
    0.05431, 0.009936447, 0.04016775, 0.02291124, 0.1285991, 0.01434812, 
    0.04395755, 0.02363233, 0.05980565, 0.01509809, 0.004561972, 5.17504e-05,
  -0.0002104395, 0.01938729, 0.02471854, 0.01916961, 0.01660071, 0.006739302, 
    0.0164003, 0.03343624, 0.2316123, 0.03273018, 0.07401866, 0.1256857, 
    0.07679491, 0.05464507, 0.03386791, 0.1112065, 0.06404318, 0.08274347, 
    0.03783263, 0.02451365, 0.06454718, 0.04064767, 0.04130864, 0.0638596, 
    0.1030639, 0.02709856, 0.01483029, 0.01234623, 0.05001433,
  0.1096025, 0.09403735, 0.02389845, 0.06238398, 0.05485686, 0.001672847, 
    0.09763388, 0.0729304, 0.01665376, 0.1167075, 0.03357814, 0.01336144, 
    0.1090266, 0.1707443, 0.1869441, 0.1898293, 0.1485827, 0.2340491, 
    0.02130179, 0.02599255, 0.08621421, 0.06969545, 0.1370924, 0.05273355, 
    0.1457488, 0.07106094, 0.03966665, 0.0521216, 0.1325795,
  0.1937212, 0.1467137, 0.05212176, 0.0590144, 0.04113348, 0.09087817, 
    0.2061044, 0.3531487, 0.1853921, 0.1191482, 0.1902222, 0.195584, 
    0.1882271, 0.2093807, 0.2136319, 0.3324922, 0.233229, 0.2369298, 
    0.07601074, 0.09152495, 0.07091869, 0.1855243, 0.3078004, 0.3779712, 
    0.1856969, 0.1374569, 0.1456305, 0.1704809, 0.1733821,
  0.2544364, 0.2337358, 0.1663826, 0.2135732, 0.1733769, 0.2014875, 
    0.2392054, 0.2904575, 0.37234, 0.413277, 0.3717654, 0.3077084, 0.2322434, 
    0.1449439, 0.2175696, 0.440578, 0.3653364, 0.3513629, 0.2602637, 
    0.1223226, 0.1716894, 0.1972519, 0.296111, 0.3095818, 0.4154197, 
    0.3251585, 0.2081838, 0.2954383, 0.2985695,
  0.3280682, 0.1936668, 0.2790784, 0.2165978, 0.295797, 0.2889369, 0.3030196, 
    0.4089164, 0.2982329, 0.1608874, 0.1621887, 0.1574762, 0.0387019, 
    0.04020789, 0.1021976, 0.1742894, 0.3395164, 0.2994311, 0.2678051, 
    0.4396632, 0.2907397, 0.2819023, 0.3464135, 0.2660054, 0.267548, 
    0.2917739, 0.3995269, 0.3098374, 0.2665044,
  0.1506769, 0.2157809, 0.2427096, 0.2383303, 0.2610755, 0.2459421, 
    0.2810974, 0.2591414, 0.1116215, 0.08194976, 0.1541339, 0.1159556, 
    0.08661973, 0.1001429, 0.09002167, 0.102868, 0.1283168, 0.2061469, 
    0.2527595, 0.2886327, 0.390117, 0.4337982, 0.3085476, 0.151798, 0.154557, 
    0.03140078, 0.08283774, 0.08840705, 0.1579153,
  0.1688053, 0.1615343, 0.1542633, 0.1469924, 0.1397214, 0.1324505, 
    0.1251795, 0.1177738, 0.1153459, 0.112918, 0.11049, 0.1080621, 0.1056341, 
    0.1032062, 0.09565765, 0.10434, 0.1130224, 0.1217048, 0.1303872, 
    0.1390696, 0.147752, 0.1822352, 0.1832517, 0.1842682, 0.1852847, 
    0.1863012, 0.1873178, 0.1883343, 0.174622,
  0.3086219, 0.1982387, 0.1308968, 0.05543637, 0.02440127, 0.003769189, 
    0.0008351377, 0.007934916, 0.03912521, 0.08373778, 0.0774003, 0.08968129, 
    0.0689217, 0.0559053, 0.0317586, 0.05011027, 0.08359471, 0.1291853, 
    0.2055065, 0.1395393, 0.1564824, 0.279589, 0.2482627, 0.2165275, 
    0.1874782, 0.2336979, 0.3579573, 0.3217088, 0.2917323,
  0.3762021, 0.1650719, 0.1833169, 0.2557912, 0.270786, 0.2435973, 0.3178859, 
    0.2700647, 0.1474518, 0.135517, 0.2250526, 0.1285765, 0.3130031, 
    0.284005, 0.2709335, 0.2380093, 0.2549139, 0.3268456, 0.2355586, 
    0.2412812, 0.2013821, 0.1972515, 0.2056596, 0.2627626, 0.3234366, 
    0.2528758, 0.2981766, 0.281687, 0.3756447,
  0.2081743, 0.2079075, 0.264419, 0.304103, 0.3442042, 0.2695917, 0.2765544, 
    0.3133759, 0.3300025, 0.3063443, 0.3730874, 0.3174243, 0.2794652, 
    0.3394487, 0.2977596, 0.2622615, 0.1933661, 0.2327154, 0.2852609, 
    0.3380404, 0.2901327, 0.2854142, 0.3504298, 0.3127439, 0.2521814, 
    0.2265845, 0.2230425, 0.2629181, 0.2096342,
  0.1089714, 0.08789726, 0.09743178, 0.1587608, 0.2156611, 0.2185439, 
    0.1790054, 0.1958431, 0.1682461, 0.1306964, 0.2251306, 0.1862358, 
    0.1367819, 0.1861229, 0.1243175, 0.1257739, 0.2667243, 0.1541945, 
    0.165599, 0.2337111, 0.2403938, 0.2024312, 0.1884847, 0.1718931, 
    0.1185445, 0.1685762, 0.222606, 0.1392707, 0.09834598,
  0.1325375, 0.145042, 0.08744094, 0.1120726, 0.1213899, 0.1379877, 
    0.1240511, 0.1225112, 0.09170719, 0.06490459, 0.08686273, 0.1186384, 
    0.09923726, 0.1634831, 0.2173189, 0.2135583, 0.1183096, 0.07816151, 
    0.1584315, 0.0918531, 0.1425578, 0.1400087, 0.1428496, 0.2076767, 
    0.08398015, 0.09591798, 0.1532979, 0.1561783, 0.07726138,
  0.0161063, -1.098462e-05, 0.008568793, 0.09155603, 0.05164063, 0.1401453, 
    0.0465883, 0.01582806, 0.03702985, 0.001114289, 9.393422e-05, 
    0.0006774964, 0.03353005, 0.05242127, 0.05113581, 0.05568844, 0.1362297, 
    0.1028697, 0.1337325, 0.04377337, 0.123975, 0.09511528, 0.001182028, 
    1.529798e-06, 0.02973908, 0.09551339, 0.1774797, 0.05196287, 0.1589983,
  6.711102e-07, -8.800741e-06, 0.0001070517, 0.01259345, 0.05538111, 
    0.026555, 0.01549144, 0.005752246, 0.004387658, 1.460421e-06, 
    0.0008393431, 0.00205556, 0.0004724073, 0.0003423745, -0.0001387809, 
    0.06659925, 0.01561673, 0.05217215, 0.1323904, 0.07320584, 0.009559873, 
    3.650619e-05, 2.388941e-08, -5.369828e-06, 0.06104586, 0.1547856, 
    0.02959841, 0.007107012, 3.743761e-05,
  1.526544e-06, 0.01188505, 0.01648122, 0.06392206, 0.03882914, 0.1709, 
    0.1932198, 0.0345003, 0.01945907, 0.003818448, 0.02941144, 0.01380055, 
    0.1147732, 0.09582486, 0.04217802, 0.03286242, 0.05527826, 0.03509883, 
    0.01039365, 0.001575445, 3.406133e-08, 1.872123e-08, 2.090889e-06, 
    0.1108228, 0.0161516, 0.04129436, 0.0002005068, 1.410438e-07, 2.359573e-07,
  0.05472899, 0.2710337, 0.05477654, 0.02653201, 0.009506865, 0.01447583, 
    0.02675652, 0.0825268, 0.1296355, 0.03902322, 0.01196592, 0.008112019, 
    0.02293184, 0.02393048, 0.008325635, 0.001602888, 0.006568863, 
    0.0006728302, 0.001026961, -2.12445e-06, 0.009897867, 0.009315418, 
    0.03034842, 0.04046384, 0.1131445, 0.000265558, 0.03991967, 0.01413028, 
    0.001626251,
  0.001717796, 0.002627186, 0.00724255, 0.205813, 0.004961305, 0.01799834, 
    0.143274, 0.03911049, 0.08872563, 0.05091386, 0.1326673, 0.07718774, 
    0.05482049, 0.08867505, 0.1003752, 0.08359122, 0.1299745, 0.1742496, 
    0.1492593, 0.174732, 0.1749992, 0.09371424, 0.1393893, 0.02769801, 
    0.02067154, 0.05378988, 0.06397244, 0.009253521, 0.002795005,
  4.133111e-06, 2.223279e-08, 2.165015e-08, 0.001006776, 0.000538628, 
    0.01794142, 0.005829909, 0.01442081, 0.0440609, 0.02477984, 0.07994878, 
    0.1028849, 0.07064237, 0.04447744, 0.06908643, 0.03628988, 0.03547281, 
    0.06051972, 0.003473953, 0.04262434, 0.01810946, 0.164684, 0.01911453, 
    0.04239794, 0.02546054, 0.05974934, 0.02827623, 0.0002420929, 1.548798e-05,
  -0.0001953986, 0.01267411, 0.02408824, 0.00634462, 0.01539062, 
    0.0009689365, 0.0126081, 0.02651319, 0.237785, 0.0345731, 0.0911813, 
    0.1183602, 0.07805479, 0.06796821, 0.03876584, 0.1178021, 0.07036526, 
    0.06576251, 0.03939131, 0.02122767, 0.06566112, 0.04764612, 0.02558078, 
    0.0733795, 0.08777446, 0.04200264, 0.03795674, 0.02155268, 0.04998066,
  0.09894089, 0.07886153, 0.02775525, 0.06269174, 0.048473, 0.004006366, 
    0.09883591, 0.06309031, 0.0115912, 0.1186423, 0.03083865, 0.01774868, 
    0.1106771, 0.1663655, 0.2042866, 0.2211555, 0.1529848, 0.2417995, 
    0.01971332, 0.01025522, 0.1151507, 0.04851322, 0.1434917, 0.06557459, 
    0.1366545, 0.06658172, 0.03543411, 0.07541322, 0.153321,
  0.2150206, 0.1578222, 0.05383332, 0.07980305, 0.05862261, 0.09446702, 
    0.2234761, 0.3504743, 0.1927598, 0.1029642, 0.1830864, 0.2074398, 
    0.2485747, 0.214104, 0.2508593, 0.3507623, 0.2503193, 0.2326302, 
    0.07892514, 0.0842889, 0.07014956, 0.1932067, 0.3324223, 0.4064561, 
    0.1938254, 0.1344663, 0.1304179, 0.2028623, 0.1858655,
  0.2596887, 0.2646725, 0.225039, 0.2147359, 0.1977593, 0.1898888, 0.2396869, 
    0.3273396, 0.3103426, 0.4186448, 0.3347175, 0.3119266, 0.2340883, 
    0.1264011, 0.2547686, 0.4729911, 0.3827205, 0.3763426, 0.2484797, 
    0.1137689, 0.1579305, 0.1488639, 0.3157718, 0.3148916, 0.3870021, 
    0.3160606, 0.2429362, 0.3255359, 0.3374773,
  0.3544769, 0.1858588, 0.2643088, 0.2442393, 0.3123955, 0.2836538, 
    0.3312578, 0.4099329, 0.3031082, 0.1329721, 0.1972244, 0.1349176, 
    0.04235013, 0.02309182, 0.1337257, 0.286725, 0.3505736, 0.2929609, 
    0.2632392, 0.36711, 0.2945449, 0.3246114, 0.2811622, 0.3288248, 
    0.2985879, 0.3016701, 0.3968316, 0.395114, 0.3294179,
  0.1646106, 0.2166565, 0.3695715, 0.3286605, 0.3842089, 0.300442, 0.317841, 
    0.2762535, 0.1601869, 0.06962105, 0.1815436, 0.1848599, 0.1165245, 
    0.09502155, 0.1159293, 0.07923021, 0.1257928, 0.1136355, 0.1623414, 
    0.204965, 0.2998519, 0.3642794, 0.3145549, 0.2357653, 0.1897551, 
    0.04306829, 0.04166709, 0.07379557, 0.1328716,
  0.2082218, 0.2005184, 0.192815, 0.1851116, 0.1774082, 0.1697049, 0.1620015, 
    0.1882103, 0.1876331, 0.1870559, 0.1864787, 0.1859015, 0.1853243, 
    0.1847471, 0.179067, 0.1857568, 0.1924467, 0.1991365, 0.2058263, 
    0.2125161, 0.2192059, 0.2045221, 0.2061129, 0.2077037, 0.2092944, 
    0.2108852, 0.212476, 0.2140668, 0.2143845,
  0.3383916, 0.255904, 0.1913064, 0.08247125, 0.02573728, 0.002834402, 
    -0.0003533246, 0.00965366, 0.05335754, 0.08355346, 0.09461291, 0.117906, 
    0.09072563, 0.03693517, 0.02343938, 0.03324118, 0.06520753, 0.1001731, 
    0.1886927, 0.1397438, 0.1644544, 0.3004429, 0.2795977, 0.2088707, 
    0.1886473, 0.2420827, 0.3737142, 0.3307593, 0.3082209,
  0.4015771, 0.1569712, 0.1836218, 0.2504888, 0.2653235, 0.2217384, 
    0.3402561, 0.2789069, 0.1689783, 0.1492416, 0.2108301, 0.1383665, 
    0.3197787, 0.2596634, 0.2232562, 0.2406688, 0.2470824, 0.341184, 
    0.2379187, 0.2412408, 0.2055573, 0.1958681, 0.2096067, 0.2517879, 
    0.3122607, 0.247877, 0.2681839, 0.303588, 0.4125538,
  0.2157138, 0.2490268, 0.3120904, 0.322574, 0.3648522, 0.2602575, 0.2595973, 
    0.291439, 0.3124475, 0.3000341, 0.4064483, 0.2929821, 0.281912, 
    0.3498214, 0.2627477, 0.2532109, 0.1823513, 0.2178234, 0.2886808, 
    0.3619096, 0.2907056, 0.3087295, 0.3602873, 0.3141506, 0.2403133, 
    0.1878236, 0.1761514, 0.2516356, 0.2137951,
  0.1080746, 0.1206318, 0.08889765, 0.1947622, 0.260545, 0.2235712, 
    0.1872234, 0.2139362, 0.2008268, 0.1768347, 0.2725855, 0.2196216, 
    0.188876, 0.2150384, 0.1364954, 0.1463524, 0.279274, 0.1601796, 
    0.1990966, 0.248096, 0.2543905, 0.2276011, 0.2136839, 0.1866499, 
    0.09181763, 0.1583514, 0.2067748, 0.1368388, 0.1394424,
  0.1609195, 0.1884238, 0.1166661, 0.1457386, 0.1580022, 0.166344, 0.1428609, 
    0.1331703, 0.09474743, 0.07068422, 0.1200781, 0.1698116, 0.1192617, 
    0.1764403, 0.270434, 0.2581317, 0.1419194, 0.07282282, 0.152736, 
    0.09788846, 0.1327071, 0.1795007, 0.1789497, 0.2211638, 0.07121956, 
    0.1039217, 0.151007, 0.179767, 0.0924018,
  0.03215461, -4.654882e-06, 0.004865719, 0.06542107, 0.03936126, 0.1480872, 
    0.0744076, 0.04089818, 0.03471336, 0.003351427, -5.421572e-05, 
    4.123251e-05, 0.02357358, 0.06953417, 0.05768784, 0.05840131, 0.1168718, 
    0.1134043, 0.154848, 0.06749601, 0.1318497, 0.104765, 0.002854966, 
    8.227021e-07, 0.01361876, 0.09574135, 0.1564573, 0.06177183, 0.1720887,
  8.696292e-07, -3.327497e-05, 1.958606e-05, 0.01409941, 0.07175714, 
    0.0511457, 0.04402227, 0.0247393, 0.01373858, 6.254627e-07, 0.0002164486, 
    0.0004362083, 0.001886705, 0.00498503, 0.001442774, 0.07143661, 
    0.02717078, 0.06206963, 0.1314428, 0.08638708, 0.03721086, 0.005117007, 
    3.160772e-07, -6.731824e-06, 0.05515706, 0.1355603, 0.05419658, 
    0.01861468, 0.003108157,
  4.910624e-07, 0.008866296, 0.005165979, 0.05275758, 0.05561331, 0.182578, 
    0.1839388, 0.04376237, 0.01655454, 0.005817073, 0.03077301, 0.01038825, 
    0.129711, 0.07901403, 0.03814595, 0.03464236, 0.04803911, 0.03530496, 
    0.0152397, 0.01417728, -2.46885e-06, 5.272276e-08, 2.475925e-06, 
    0.1065251, 0.01280772, 0.009316357, 0.006060668, 1.713991e-06, 
    3.664953e-07,
  0.05529222, 0.247771, 0.04557675, 0.03633379, 0.01328154, 0.01521741, 
    0.02104589, 0.0583109, 0.1196233, 0.03637397, 0.01584752, 0.01167471, 
    0.02087335, 0.0242844, 0.01289482, 0.005804826, 0.006119606, 0.001347945, 
    0.00222735, 1.717244e-05, 0.006218141, 0.004054411, 0.03357581, 
    0.04208612, 0.04808457, 0.0004667569, 0.03908011, 0.02137827, 0.001899132,
  0.001167184, 0.001267454, 0.003596071, 0.1706383, 0.008927825, 0.0185517, 
    0.1442493, 0.03363826, 0.08897054, 0.04479171, 0.1224863, 0.06337705, 
    0.05077028, 0.07604364, 0.08227568, 0.07124697, 0.1166419, 0.1514149, 
    0.1492207, 0.1571647, 0.1587608, 0.09351598, 0.1626608, 0.03800059, 
    0.01865458, 0.0467666, 0.05289763, 0.007211343, 0.001040014,
  1.948962e-06, 5.743313e-09, 6.036836e-09, 0.000947885, 0.0001089786, 
    0.01211721, 0.006261287, 0.01789151, 0.0475832, 0.03193856, 0.1000619, 
    0.09931653, 0.06361379, 0.04247496, 0.0624919, 0.02929627, 0.03927451, 
    0.06269597, 0.005344437, 0.04842705, 0.010243, 0.1926156, 0.02043297, 
    0.03892992, 0.022927, 0.05328034, 0.0386335, 2.120659e-06, 5.167993e-06,
  -4.597094e-05, 0.01622816, 0.02900205, 0.0004604072, 0.01029663, 
    -8.165396e-05, 0.006352849, 0.01803336, 0.2217914, 0.05281157, 0.1052704, 
    0.1486163, 0.08048355, 0.08593522, 0.04617839, 0.1288705, 0.07996739, 
    0.06200286, 0.02991951, 0.019742, 0.03088853, 0.05385488, 0.01899591, 
    0.08187639, 0.06878893, 0.04083056, 0.08165473, 0.04771901, 0.03289895,
  0.08505544, 0.06959732, 0.04141783, 0.04555067, 0.02195877, 0.0003062013, 
    0.09694897, 0.05266733, 0.01393675, 0.1285902, 0.03342117, 0.02880226, 
    0.1150625, 0.1759389, 0.2232495, 0.2255731, 0.1654211, 0.2576045, 
    0.01755028, 0.003337331, 0.149283, 0.0487234, 0.1414874, 0.09800891, 
    0.1281034, 0.05849627, 0.03586158, 0.1013622, 0.1712893,
  0.2177951, 0.1383878, 0.06737408, 0.07844356, 0.06075608, 0.06671351, 
    0.2539699, 0.3467239, 0.2025501, 0.09767608, 0.148874, 0.1960176, 
    0.241724, 0.2472239, 0.2745989, 0.3905263, 0.2588569, 0.2399331, 
    0.07206421, 0.09253244, 0.09642255, 0.188644, 0.3039054, 0.4542092, 
    0.2089728, 0.1347118, 0.1465915, 0.2477069, 0.2033305,
  0.2535224, 0.2561907, 0.1963878, 0.1642172, 0.2409403, 0.1702031, 
    0.2130646, 0.3433858, 0.2926783, 0.371085, 0.3712879, 0.3265183, 
    0.2191949, 0.1121961, 0.2704347, 0.4270817, 0.430835, 0.4024944, 
    0.2594519, 0.1202247, 0.1526275, 0.1511672, 0.3364619, 0.2999302, 
    0.376355, 0.3137952, 0.3075538, 0.3655195, 0.3517298,
  0.3621118, 0.2153492, 0.2319813, 0.2964354, 0.3085606, 0.2915199, 0.32542, 
    0.3759261, 0.3394965, 0.1858377, 0.2060235, 0.1111675, 0.06992459, 
    0.1479179, 0.1631845, 0.2627909, 0.328379, 0.2789871, 0.2971736, 
    0.3610757, 0.2754899, 0.3005059, 0.2683163, 0.3678006, 0.2619883, 
    0.3005472, 0.3900822, 0.4308878, 0.377463,
  0.1500609, 0.1911584, 0.3697571, 0.2936229, 0.3517722, 0.2768181, 
    0.2957703, 0.2363238, 0.1853734, 0.1141842, 0.1663518, 0.1233967, 
    0.1012495, 0.05940288, 0.09192303, 0.07179474, 0.1067582, 0.1401309, 
    0.1886405, 0.2747124, 0.3186925, 0.3631544, 0.3173133, 0.2332931, 
    0.1610222, 0.05713561, 0.02032449, 0.09196717, 0.1524071,
  0.2529767, 0.2434386, 0.2339004, 0.2243623, 0.2148241, 0.2052859, 
    0.1957478, 0.2129044, 0.2120874, 0.2112704, 0.2104533, 0.2096363, 
    0.2088193, 0.2080023, 0.2005827, 0.2092043, 0.2178258, 0.2264474, 
    0.2350689, 0.2436905, 0.252312, 0.2694502, 0.2711838, 0.2729174, 
    0.2746511, 0.2763847, 0.2781184, 0.2798521, 0.2606073,
  0.3649154, 0.3365712, 0.2381644, 0.1316631, 0.03900337, 0.004330896, 
    0.002410913, 0.01077964, 0.06032556, 0.0983333, 0.1281752, 0.1576566, 
    0.1168854, 0.03050733, 0.01899848, 0.04084083, 0.05720359, 0.08832102, 
    0.1618839, 0.1318914, 0.1755532, 0.3118649, 0.3029815, 0.2182861, 
    0.1945314, 0.2573647, 0.3780268, 0.3318202, 0.3335651,
  0.4122979, 0.1563845, 0.1910799, 0.233906, 0.2614537, 0.2125378, 0.3279772, 
    0.2904122, 0.1660555, 0.1582436, 0.1962922, 0.133132, 0.3199352, 
    0.2434688, 0.2261678, 0.2387602, 0.2396151, 0.3385684, 0.2666317, 
    0.2813958, 0.2624413, 0.2945359, 0.222724, 0.2477723, 0.3075363, 
    0.2353094, 0.2800523, 0.3593473, 0.4242217,
  0.2117366, 0.2246341, 0.320345, 0.3391126, 0.3832757, 0.2789916, 0.3050546, 
    0.3521585, 0.3518604, 0.3973439, 0.4342017, 0.3031739, 0.2610471, 
    0.3452353, 0.264793, 0.2371282, 0.1780808, 0.2574586, 0.3605977, 
    0.4218572, 0.3376541, 0.3448283, 0.3766055, 0.2932609, 0.2485558, 
    0.2161365, 0.1580764, 0.2554784, 0.1980679,
  0.1353705, 0.1399851, 0.1638709, 0.2751944, 0.3255439, 0.2601182, 
    0.2331864, 0.3069341, 0.2730128, 0.2150998, 0.3497871, 0.2534857, 
    0.235849, 0.221588, 0.1561651, 0.1996651, 0.2940643, 0.2009409, 
    0.2418789, 0.2628581, 0.2538435, 0.2287414, 0.2500083, 0.1926915, 
    0.07252508, 0.1845419, 0.2470696, 0.1593717, 0.2004565,
  0.2393075, 0.2078701, 0.1595328, 0.2035492, 0.2312663, 0.2271003, 
    0.2067392, 0.2047476, 0.133103, 0.1288921, 0.1824998, 0.2066884, 
    0.1172738, 0.2095083, 0.2973744, 0.2733451, 0.1748511, 0.08762929, 
    0.1879605, 0.1473612, 0.1663334, 0.2418771, 0.2456693, 0.2666044, 
    0.05934352, 0.1291434, 0.1601318, 0.1831575, 0.1191897,
  0.05407296, 0.0001487633, 0.008698117, 0.0634568, 0.04985743, 0.1745021, 
    0.1049283, 0.09395132, 0.0450964, 0.008709828, -0.0003483029, 
    1.52596e-05, 0.0194754, 0.07636311, 0.08175112, 0.07971203, 0.116523, 
    0.1186674, 0.1478725, 0.1280275, 0.1515161, 0.09493239, 0.01920653, 
    -2.211959e-06, 0.006408135, 0.1042834, 0.1499545, 0.07513601, 0.1744381,
  6.434337e-07, -1.221213e-05, 4.262061e-06, 0.01352781, 0.08133964, 
    0.057083, 0.05904191, 0.05797872, 0.03709115, -1.373803e-07, 
    4.287156e-05, 0.000144055, 0.006045475, 0.006039212, 0.00370262, 
    0.09827641, 0.03381142, 0.06031356, 0.1158755, 0.05961376, 0.05400319, 
    0.03291842, -1.123076e-06, -4.013787e-06, 0.04072682, 0.1273931, 
    0.07169721, 0.04027848, 0.01089988,
  3.975036e-06, 0.00177599, 0.00128139, 0.04536841, 0.06413873, 0.1813862, 
    0.1552089, 0.04484394, 0.01629027, 0.00720288, 0.02729212, 0.0110796, 
    0.1265516, 0.0647223, 0.03404035, 0.03233696, 0.03826406, 0.02875795, 
    0.02069164, 0.02540189, 0.001378549, 7.578046e-07, 1.074353e-06, 
    0.09953789, 0.01439892, 0.0008923489, 0.02858251, 0.0004816819, 
    2.006158e-06,
  0.06100874, 0.2142738, 0.04133868, 0.02562251, 0.01261801, 0.01729446, 
    0.01781701, 0.04281844, 0.1119322, 0.05093438, 0.01964758, 0.01390456, 
    0.0206142, 0.02391306, 0.01815334, 0.008224603, 0.01056621, 0.005603486, 
    0.008910489, 0.001641294, 0.002294174, 0.02457441, 0.03430547, 
    0.04491186, 0.02030355, 0.001229635, 0.03438033, 0.03724805, 0.004850172,
  0.001018645, 0.0009310311, 0.002260494, 0.1302081, 0.001579776, 0.02196058, 
    0.1411829, 0.02769546, 0.07592545, 0.04056863, 0.09596705, 0.04818361, 
    0.04125256, 0.06433117, 0.06842439, 0.05416051, 0.1011621, 0.1351537, 
    0.1388282, 0.1261049, 0.1388091, 0.084052, 0.1720631, 0.05002847, 
    0.01927818, 0.04272244, 0.04395196, 0.00804839, 0.0008867774,
  1.165648e-06, 3.015904e-09, 2.433855e-09, 0.0009012591, 3.753074e-05, 
    0.009317542, 0.007673536, 0.01799069, 0.0578496, 0.05164361, 0.1219574, 
    0.09738558, 0.05500356, 0.04256969, 0.05867316, 0.03112582, 0.03860598, 
    0.08222478, 0.01215975, 0.04386737, 0.006677242, 0.2103889, 0.02230219, 
    0.03663174, 0.02183009, 0.04616204, 0.03925623, 3.693287e-05, 2.5321e-06,
  -8.972101e-06, 0.02991821, 0.01137221, 6.409849e-05, 0.006762727, 
    -1.050005e-05, 0.005200801, 0.01256403, 0.231602, 0.07603349, 0.1327949, 
    0.176271, 0.09802269, 0.09462846, 0.07097704, 0.1610863, 0.1119725, 
    0.07365399, 0.03470495, 0.01662208, 0.01578278, 0.05705689, 0.01640435, 
    0.1037741, 0.05710474, 0.03854604, 0.1004776, 0.09359797, 0.0241291,
  0.07408721, 0.06276433, 0.03264727, 0.06068361, 0.01556335, -0.0002043879, 
    0.09394229, 0.03838608, 0.01426602, 0.1329006, 0.03963239, 0.03486794, 
    0.1354178, 0.1964369, 0.3229118, 0.2523555, 0.1761727, 0.2711391, 
    0.03004579, 0.002662427, 0.1093595, 0.04838808, 0.1553028, 0.09296277, 
    0.1363679, 0.05983891, 0.07717978, 0.1711044, 0.1590117,
  0.2250772, 0.1250737, 0.1044977, 0.05543462, 0.04604303, 0.09570238, 
    0.2497852, 0.3736781, 0.1959405, 0.07822435, 0.1245837, 0.2284248, 
    0.2457457, 0.286275, 0.3291024, 0.4046909, 0.2917394, 0.246219, 
    0.06216394, 0.08586217, 0.1373332, 0.1933259, 0.3246096, 0.4837034, 
    0.2129129, 0.1458626, 0.2321537, 0.2937846, 0.2120803,
  0.2867139, 0.2707257, 0.1853186, 0.1970117, 0.2395675, 0.1658421, 
    0.2225056, 0.4131998, 0.3325837, 0.3843001, 0.3647367, 0.3890155, 
    0.1782434, 0.1119147, 0.3807188, 0.445551, 0.4715201, 0.419865, 
    0.2852521, 0.1391252, 0.1440371, 0.218022, 0.4092606, 0.3508549, 
    0.4137081, 0.3064716, 0.3604023, 0.4046699, 0.3775508,
  0.4582432, 0.2902009, 0.2619062, 0.3386461, 0.347199, 0.3775786, 0.3611386, 
    0.4084714, 0.3189833, 0.2609013, 0.2233256, 0.1656286, 0.1322137, 
    0.1609569, 0.1879275, 0.246648, 0.33063, 0.2724213, 0.2916527, 0.3854245, 
    0.3329635, 0.3304577, 0.3214689, 0.3642296, 0.3300159, 0.2944497, 
    0.3609751, 0.4352212, 0.4500891,
  0.1381226, 0.2496979, 0.3079139, 0.2885074, 0.2917874, 0.2657991, 
    0.2596158, 0.2125111, 0.1975239, 0.2168619, 0.2303597, 0.1464148, 
    0.1180028, 0.06095801, 0.07390147, 0.1059359, 0.1643836, 0.1814163, 
    0.194456, 0.2579936, 0.3271325, 0.3502489, 0.3437807, 0.2508132, 
    0.1557455, 0.03916002, 0.0200682, 0.0737716, 0.2667561,
  0.3260913, 0.3162608, 0.3064305, 0.2966, 0.2867696, 0.2769392, 0.2671088, 
    0.2581458, 0.2548876, 0.2516295, 0.2483713, 0.2451131, 0.241855, 
    0.2385968, 0.2294556, 0.240081, 0.2507063, 0.2613316, 0.2719569, 
    0.2825822, 0.2932075, 0.3279814, 0.3304446, 0.3329079, 0.3353711, 
    0.3378344, 0.3402977, 0.342761, 0.3339556,
  0.3782505, 0.393324, 0.2701946, 0.1474197, 0.05458491, 0.008130983, 
    -0.001199107, 0.009671147, 0.05968565, 0.1065477, 0.1684947, 0.1748487, 
    0.1600793, 0.0134354, 0.01835049, 0.04104267, 0.0521567, 0.08920401, 
    0.1447345, 0.1301306, 0.1731942, 0.3220439, 0.3159826, 0.2687931, 
    0.2254415, 0.2661063, 0.3389843, 0.3190637, 0.3604994,
  0.4168794, 0.1481296, 0.202252, 0.2219808, 0.2454407, 0.215819, 0.2783287, 
    0.2924885, 0.1484499, 0.175723, 0.1801259, 0.1380345, 0.3137432, 
    0.2256556, 0.2523969, 0.220771, 0.3232354, 0.362581, 0.2689471, 
    0.2668324, 0.2614863, 0.2857797, 0.2224524, 0.2738506, 0.256303, 
    0.2435894, 0.3069662, 0.3653855, 0.4660079,
  0.2462331, 0.2669625, 0.3206054, 0.4188882, 0.4009955, 0.3099014, 
    0.3631021, 0.4106098, 0.4218012, 0.5177323, 0.4047038, 0.346335, 
    0.2863517, 0.337245, 0.2379809, 0.2836551, 0.2732529, 0.3633282, 
    0.3984231, 0.4150003, 0.3264111, 0.2870816, 0.350267, 0.3152242, 
    0.308045, 0.2538116, 0.2012422, 0.3036845, 0.2720781,
  0.2300528, 0.2084938, 0.253935, 0.3165095, 0.3344945, 0.2479533, 0.2995684, 
    0.336286, 0.3252207, 0.3285587, 0.4369644, 0.315474, 0.2636273, 
    0.2498072, 0.1607746, 0.2665895, 0.3046045, 0.2320058, 0.3018951, 
    0.3013418, 0.2680591, 0.249961, 0.2836632, 0.2000525, 0.06243422, 
    0.2145296, 0.2780635, 0.1957629, 0.2713118,
  0.2843421, 0.2449254, 0.197221, 0.2246833, 0.2579968, 0.2526013, 0.3252765, 
    0.2862944, 0.2296712, 0.2279672, 0.3046996, 0.2003198, 0.1407437, 
    0.2751507, 0.314083, 0.2589104, 0.2166133, 0.135518, 0.2297313, 
    0.2239682, 0.2422687, 0.2736702, 0.2450478, 0.2927415, 0.05899695, 
    0.1364366, 0.1586947, 0.1716511, 0.2149556,
  0.09273162, 0.0006571798, 0.009779352, 0.09208052, 0.07398897, 0.2151653, 
    0.1485579, 0.1576578, 0.1391081, 0.05227994, 0.0007396886, -1.910433e-05, 
    0.01575179, 0.1115587, 0.1323485, 0.1063706, 0.1128449, 0.1442173, 
    0.1531374, 0.1321598, 0.176744, 0.09992669, 0.09327548, -3.756642e-06, 
    0.008164612, 0.2162059, 0.1732753, 0.1515153, 0.2173448,
  -8.510862e-05, -4.648419e-06, -3.97979e-06, 0.03316343, 0.08443766, 
    0.07648253, 0.06941348, 0.1128544, 0.1335034, -0.0001113596, 
    7.314183e-06, 4.985292e-05, 0.0180699, 0.008315994, 0.009179235, 
    0.1046818, 0.03594136, 0.06724291, 0.1024318, 0.05145115, 0.1512948, 
    0.09396653, 0.001755824, -2.378399e-06, 0.02241605, 0.1228876, 0.1037098, 
    0.05819456, 0.01656149,
  5.913906e-05, -0.0003851358, 0.0003933268, 0.03943135, 0.06456145, 
    0.1585336, 0.1303795, 0.0437646, 0.01765274, 0.01132175, 0.02380605, 
    0.01418369, 0.1106322, 0.05017313, 0.03825949, 0.03350526, 0.03548935, 
    0.02934233, 0.02705353, 0.04074313, 0.01360724, 0.0005792095, 
    2.048393e-06, 0.08773833, 0.0165258, 0.00014594, 0.07293474, 0.01316309, 
    9.286566e-05,
  0.0628125, 0.195549, 0.04395215, 0.01902414, 0.01846774, 0.02296169, 
    0.01788936, 0.03366458, 0.1078142, 0.116354, 0.02820745, 0.01490098, 
    0.0210947, 0.03999297, 0.02573878, 0.009220075, 0.006926769, 0.01607716, 
    0.02740689, 0.01703078, 0.002487951, 0.005730566, 0.02179662, 0.0493695, 
    0.006202174, 0.007312228, 0.03952284, 0.04827359, 0.01447727,
  0.0007036129, 0.0005446949, 0.00104803, 0.08945986, 0.0008529944, 
    0.02670309, 0.1195892, 0.02941184, 0.0894214, 0.06625547, 0.06970386, 
    0.03802291, 0.03316744, 0.05360458, 0.05549037, 0.04565555, 0.08678712, 
    0.1269226, 0.1201021, 0.1061886, 0.1216285, 0.07164133, 0.1637168, 
    0.05396863, 0.02273478, 0.04332145, 0.03836202, 0.01264436, 0.0004629993,
  7.796126e-07, 1.996298e-09, 6.906002e-10, 0.0008362429, 1.431713e-05, 
    0.007856486, 0.008939207, 0.01931904, 0.0739886, 0.1141064, 0.1506091, 
    0.08567034, 0.0519001, 0.06096174, 0.06705325, 0.03108286, 0.04638275, 
    0.07938562, 0.0596036, 0.04716129, 0.007420867, 0.212659, 0.05852757, 
    0.0394109, 0.02793122, 0.05500406, 0.04974139, 0.0007144029, 1.471896e-06,
  -2.161403e-05, 0.02055252, 0.002102857, 2.412057e-05, 0.005064733, 
    4.833956e-07, 0.003489282, 0.01091748, 0.2507077, 0.07597584, 0.2707202, 
    0.2416263, 0.1010773, 0.1258263, 0.132031, 0.2568807, 0.1402635, 
    0.09635761, 0.08338089, 0.008437752, 0.01933818, 0.05635529, 0.02853481, 
    0.1425386, 0.04364595, 0.03595543, 0.09938542, 0.1526142, 0.03359443,
  0.07414108, 0.06774552, 0.04455879, 0.08090492, 0.03239276, -6.315133e-05, 
    0.095136, 0.02920403, 0.011915, 0.1100782, 0.06833982, 0.07372924, 
    0.2024706, 0.2363538, 0.3159599, 0.233898, 0.2087356, 0.2890171, 
    0.05222616, 0.003251349, 0.07633128, 0.04744599, 0.2068364, 0.1169818, 
    0.1901081, 0.1063418, 0.1680641, 0.2043557, 0.1587959,
  0.2260225, 0.1147165, 0.107958, 0.04723546, 0.05112818, 0.1996125, 
    0.2385142, 0.3954699, 0.1933837, 0.09770895, 0.1077634, 0.2385646, 
    0.293493, 0.3159483, 0.3556557, 0.4158524, 0.3114718, 0.2415614, 
    0.07363196, 0.08599152, 0.1199243, 0.2003438, 0.3467546, 0.5036428, 
    0.2074203, 0.2020022, 0.2972588, 0.252081, 0.2240116,
  0.32833, 0.2889013, 0.2401769, 0.2366002, 0.2360303, 0.1847118, 0.3471091, 
    0.4546723, 0.3634111, 0.4533292, 0.4065592, 0.4011078, 0.1728362, 
    0.1547723, 0.6513368, 0.5580739, 0.4879041, 0.4353092, 0.2822129, 
    0.145575, 0.1364299, 0.2297415, 0.3891251, 0.4065316, 0.4208529, 
    0.3318072, 0.369336, 0.4440589, 0.3705946,
  0.4881812, 0.3988849, 0.2922838, 0.371318, 0.4437523, 0.4795338, 0.3240779, 
    0.3951387, 0.3247415, 0.3237502, 0.1902719, 0.209462, 0.1148987, 
    0.1768149, 0.2509968, 0.2768358, 0.3782575, 0.3154937, 0.3343978, 
    0.4031308, 0.3157185, 0.4318042, 0.3577324, 0.4129347, 0.4362677, 
    0.3217871, 0.3415711, 0.3955775, 0.4391036,
  0.3420935, 0.3822417, 0.3625019, 0.3055596, 0.3345734, 0.3087475, 
    0.3180491, 0.2205553, 0.1327606, 0.1779936, 0.2653055, 0.1355187, 
    0.1180583, 0.06533537, 0.1065709, 0.1260606, 0.1782749, 0.1938162, 
    0.2182722, 0.3099415, 0.3022018, 0.3278868, 0.3342919, 0.2580306, 
    0.1923962, 0.05778005, 0.0184197, 0.08777241, 0.2615362,
  0.3594762, 0.3494927, 0.3395092, 0.3295258, 0.3195423, 0.3095588, 
    0.2995753, 0.3116824, 0.3079818, 0.3042811, 0.3005804, 0.2968797, 
    0.293179, 0.2894784, 0.2780112, 0.2890692, 0.3001272, 0.3111852, 
    0.3222432, 0.3333012, 0.3443592, 0.3619564, 0.3645826, 0.3672087, 
    0.3698349, 0.3724611, 0.3750873, 0.3777135, 0.367463,
  0.4146209, 0.4263366, 0.2882084, 0.1771272, 0.05923052, 0.00704297, 
    -0.003844347, 0.01207937, 0.068519, 0.1112246, 0.1915173, 0.1745727, 
    0.1713842, -0.001003598, 0.01752944, 0.02559105, 0.06272041, 0.07915971, 
    0.1409024, 0.143105, 0.1846111, 0.3237299, 0.3143751, 0.3057588, 
    0.3230667, 0.2831978, 0.3151431, 0.2905389, 0.3841317,
  0.457078, 0.1397691, 0.2007286, 0.1643631, 0.2113578, 0.2161387, 0.2132246, 
    0.2737116, 0.1310412, 0.1805045, 0.1792327, 0.1449793, 0.3018139, 
    0.1980472, 0.2564466, 0.2475097, 0.3267309, 0.3744506, 0.2766797, 
    0.3131946, 0.2860423, 0.2869046, 0.2409534, 0.2846862, 0.2257176, 
    0.2924168, 0.3330215, 0.3571973, 0.51013,
  0.3617055, 0.3664619, 0.3825527, 0.5219246, 0.424703, 0.3351289, 0.377938, 
    0.4320344, 0.4265482, 0.5068298, 0.3684216, 0.3544168, 0.3012088, 
    0.2918414, 0.2515849, 0.3070839, 0.3266016, 0.403163, 0.4090333, 
    0.393323, 0.2750543, 0.2235599, 0.365896, 0.3524036, 0.3480076, 
    0.2598837, 0.306188, 0.3769191, 0.3515481,
  0.2868038, 0.3249452, 0.2883184, 0.2981412, 0.3457671, 0.3081197, 
    0.3172885, 0.3315311, 0.3571207, 0.3388981, 0.3783354, 0.257457, 
    0.2413396, 0.2318617, 0.1998525, 0.2587206, 0.3223505, 0.3321744, 
    0.3072851, 0.3583898, 0.3019806, 0.2866365, 0.2736403, 0.2114318, 
    0.04813721, 0.1847878, 0.299686, 0.2688819, 0.3173814,
  0.3683022, 0.271532, 0.1502302, 0.2032393, 0.2446698, 0.2181013, 0.3251219, 
    0.2895007, 0.4024628, 0.2584522, 0.2319792, 0.1953384, 0.1533014, 
    0.2450764, 0.3007059, 0.2892036, 0.2118957, 0.1766098, 0.3011096, 
    0.2643396, 0.377083, 0.2768562, 0.2737348, 0.3123615, 0.0551956, 
    0.1325992, 0.1839297, 0.1626052, 0.2722358,
  0.1678924, 0.03271521, 0.01109765, 0.1136334, 0.1329403, 0.2797032, 
    0.204528, 0.2857082, 0.2374358, 0.08286674, 0.000434401, -2.854316e-06, 
    0.01265208, 0.1163793, 0.1292509, 0.1563705, 0.1887142, 0.1523176, 
    0.1360634, 0.1048791, 0.2278604, 0.1862383, 0.1591206, 6.14451e-05, 
    0.01165276, 0.2571581, 0.1505478, 0.1048304, 0.2034334,
  0.005991833, -2.125812e-06, -5.959471e-07, 0.02238348, 0.07895432, 
    0.08977121, 0.0868686, 0.1640331, 0.2169399, 0.02959906, 1.478466e-06, 
    1.317935e-05, 0.0323676, 0.02784847, 0.04297975, 0.1310469, 0.07043395, 
    0.07615083, 0.09653894, 0.08089924, 0.1738791, 0.2699814, 0.129577, 
    -1.808614e-06, 0.01598448, 0.1258623, 0.1059994, 0.126405, 0.05385855,
  0.004251065, 0.002453091, 0.0001428082, 0.03351297, 0.07161865, 0.1379507, 
    0.1213587, 0.06326784, 0.03212357, 0.04298884, 0.02408723, 0.02129805, 
    0.1140898, 0.04580266, 0.0404548, 0.05430064, 0.05150295, 0.05408129, 
    0.04824809, 0.06991562, 0.05593874, 0.03831435, 0.0003164402, 0.0743325, 
    0.01298158, 4.598304e-05, 0.1141884, 0.08678157, 0.009231663,
  0.07424875, 0.1835541, 0.03171862, 0.01513646, 0.03273679, 0.03076238, 
    0.02220472, 0.03441725, 0.08632617, 0.1464489, 0.04901275, 0.01741194, 
    0.02936579, 0.07164032, 0.1059994, 0.02964106, 0.009328689, 0.02339977, 
    0.03565707, 0.03561259, 0.03217255, 0.002021041, 0.005242554, 0.03084184, 
    0.003090258, 0.02612055, 0.05479001, 0.05906287, 0.03494465,
  0.0002877146, 0.0003098668, 0.0004059478, 0.06633785, 0.001393782, 
    0.04113995, 0.09085932, 0.03983222, 0.09354994, 0.07888781, 0.05183231, 
    0.03645472, 0.03503294, 0.05103002, 0.04483653, 0.04367556, 0.07776371, 
    0.1122937, 0.107266, 0.08675166, 0.1093413, 0.06233703, 0.1473658, 
    0.05598271, 0.03918463, 0.06140506, 0.04254284, 0.03615692, 5.636172e-05,
  5.177559e-07, 1.779119e-09, 4.604852e-10, 0.001355353, 2.693976e-06, 
    0.01732257, 0.007350798, 0.02300086, 0.0591222, 0.1451157, 0.1413791, 
    0.07304774, 0.06053447, 0.05204565, 0.07445004, 0.05290769, 0.05697124, 
    0.1309794, 0.08501918, 0.05098235, 0.01785215, 0.2519649, 0.07407123, 
    0.04863708, 0.04282998, 0.05917921, 0.07295361, 0.07248621, 8.787987e-07,
  -1.143293e-05, 0.006033475, 4.546683e-05, 1.061031e-05, 0.003496914, 
    6.928398e-07, 0.003006001, 0.01056407, 0.2591651, 0.04650778, 0.2842572, 
    0.2919859, 0.09776122, 0.131301, 0.2141228, 0.2205497, 0.1008376, 
    0.1283481, 0.1886448, 0.02833329, 0.0294224, 0.0727779, 0.06402752, 
    0.1469889, 0.04203051, 0.03953356, 0.08161234, 0.124224, 0.0427474,
  0.08198201, 0.04486507, 0.04506202, 0.09607743, 0.0152903, -6.27104e-07, 
    0.09814067, 0.02253685, 0.006818925, 0.09971566, 0.07137834, 0.07349118, 
    0.3080356, 0.2557787, 0.2278298, 0.187711, 0.2091197, 0.2929912, 
    0.0859234, 0.003963793, 0.04786376, 0.04910007, 0.1943583, 0.1044908, 
    0.2365903, 0.1457238, 0.2518618, 0.2539398, 0.1661119,
  0.2279349, 0.1298905, 0.1018593, 0.03416475, 0.08473598, 0.2025432, 
    0.2296762, 0.3848449, 0.2085978, 0.1067553, 0.09813952, 0.2179673, 
    0.2970972, 0.2805594, 0.3194109, 0.4021209, 0.3222015, 0.2660244, 
    0.09916326, 0.08682935, 0.1008782, 0.2223933, 0.3742557, 0.4713113, 
    0.2140604, 0.2378097, 0.3161647, 0.2032251, 0.1875551,
  0.3313991, 0.3153302, 0.3231592, 0.2911, 0.2937188, 0.2621479, 0.4793821, 
    0.4796742, 0.4453596, 0.5291926, 0.4189061, 0.3770899, 0.194182, 
    0.2618515, 0.5472881, 0.5490267, 0.4739889, 0.432485, 0.3070601, 
    0.1557488, 0.136484, 0.3434444, 0.3404583, 0.3885148, 0.4489334, 
    0.3244066, 0.3796648, 0.3926674, 0.3367269,
  0.4588217, 0.4405117, 0.3418474, 0.3991132, 0.4537722, 0.4437079, 
    0.3515822, 0.4696849, 0.3332796, 0.368894, 0.1867361, 0.2538708, 
    0.238827, 0.284381, 0.2916464, 0.4061089, 0.440251, 0.341651, 0.4382419, 
    0.4661019, 0.4210912, 0.4838293, 0.4096293, 0.4551011, 0.3618217, 
    0.3389635, 0.3064588, 0.354569, 0.4895184,
  0.4109537, 0.3582513, 0.3648921, 0.3657659, 0.4258032, 0.379029, 0.3679057, 
    0.2153481, 0.1326661, 0.2002007, 0.2513468, 0.1737182, 0.1641984, 
    0.117151, 0.1877598, 0.2014728, 0.2185636, 0.1832002, 0.2401592, 
    0.3359228, 0.3575948, 0.3354003, 0.4001751, 0.3632674, 0.2046788, 
    0.07373761, 0.02818353, 0.1355001, 0.2933975,
  0.3837712, 0.3730008, 0.3622304, 0.3514601, 0.3406897, 0.3299194, 0.319149, 
    0.3323781, 0.3289218, 0.3254656, 0.3220094, 0.3185531, 0.3150969, 
    0.3116406, 0.3065228, 0.3184053, 0.3302879, 0.3421704, 0.354053, 
    0.3659356, 0.3778181, 0.3885207, 0.3908647, 0.3932087, 0.3955528, 
    0.3978968, 0.4002408, 0.4025849, 0.3923874,
  0.4284412, 0.454033, 0.3079066, 0.2150985, 0.05896048, 0.01240956, 
    -0.00495091, 0.01275158, 0.0796438, 0.1057273, 0.1971084, 0.1888813, 
    0.1670415, -0.009439518, 0.01881762, 0.009515346, 0.05175849, 0.09103184, 
    0.1542049, 0.1540558, 0.2112757, 0.318365, 0.334943, 0.308842, 0.3102846, 
    0.3235135, 0.2591517, 0.2442285, 0.3974684,
  0.4630944, 0.1204476, 0.1843111, 0.1138166, 0.1807155, 0.2010882, 
    0.1350101, 0.2503929, 0.1249154, 0.1828862, 0.1847961, 0.1363241, 
    0.2726837, 0.1804961, 0.2604487, 0.2698956, 0.311865, 0.390594, 
    0.3107112, 0.3575106, 0.3003349, 0.3304343, 0.261749, 0.2977345, 
    0.1958125, 0.3280759, 0.3849286, 0.3847244, 0.5845945,
  0.445187, 0.4765649, 0.4763439, 0.5240441, 0.3733319, 0.3317989, 0.3702078, 
    0.4151335, 0.464298, 0.4642504, 0.3640779, 0.3069616, 0.3256235, 
    0.302354, 0.231925, 0.2789932, 0.3965829, 0.3660135, 0.4203026, 
    0.3762975, 0.2413142, 0.2186375, 0.3221693, 0.3661157, 0.3244488, 
    0.3148162, 0.413369, 0.4624991, 0.3929798,
  0.4600626, 0.3631949, 0.3240443, 0.266275, 0.3002196, 0.3055094, 0.3219574, 
    0.3200263, 0.3455529, 0.3460648, 0.3355872, 0.2998586, 0.1930053, 
    0.197568, 0.178397, 0.2153729, 0.3511149, 0.3018791, 0.3529805, 
    0.4026531, 0.3926128, 0.342422, 0.2523076, 0.2424543, 0.05354112, 
    0.1962841, 0.3661989, 0.3486224, 0.3926118,
  0.3544832, 0.2192749, 0.1765007, 0.1529067, 0.1959664, 0.1559416, 0.209782, 
    0.2516424, 0.3090102, 0.2831674, 0.1887007, 0.132646, 0.08288644, 
    0.178532, 0.3118463, 0.283437, 0.2000969, 0.204153, 0.3012086, 0.3781405, 
    0.2922243, 0.2663816, 0.2532696, 0.3337538, 0.0538233, 0.1164382, 
    0.1705806, 0.1534094, 0.2156718,
  0.1828699, 0.06939071, 0.00967025, 0.1292098, 0.1361956, 0.3033053, 
    0.1977846, 0.304763, 0.3827639, 0.05571637, 0.0009559173, -4.06962e-06, 
    0.01120813, 0.1022411, 0.1299709, 0.1369765, 0.1744183, 0.1939547, 
    0.1147572, 0.05538091, 0.2439616, 0.2079147, 0.2444945, 0.001869523, 
    0.01424914, 0.247995, 0.1565097, 0.05211718, 0.1601056,
  0.2173045, 4.265112e-06, -3.478756e-07, 0.047577, 0.1329392, 0.08045318, 
    0.0723981, 0.1088608, 0.1093755, 0.01745165, 4.572028e-07, 2.062103e-06, 
    0.09778935, 0.1393017, 0.1016012, 0.2191901, 0.05229557, 0.09042329, 
    0.0825867, 0.06619346, 0.1333095, 0.3355437, 0.519371, 5.731289e-06, 
    0.01496772, 0.1286263, 0.1097593, 0.1593684, 0.151912,
  0.03363908, 0.02479151, 6.394798e-05, 0.03181649, 0.08243922, 0.1336526, 
    0.1274391, 0.06671031, 0.1237126, 0.1783394, 0.02127347, 0.04179593, 
    0.1228857, 0.05209907, 0.06694147, 0.05707507, 0.1101441, 0.0804039, 
    0.09602684, 0.08293682, 0.3152198, 0.474651, 0.008282424, 0.04861136, 
    0.005377565, 1.784541e-05, 0.1889424, 0.3019119, 0.2190136,
  0.08119402, 0.1588674, 0.01480333, 0.0265707, 0.04911572, 0.06819811, 
    0.04681371, 0.08383488, 0.08077944, 0.07730268, 0.1028009, 0.09047164, 
    0.1207302, 0.03775731, 0.1171151, 0.08318101, 0.03216152, 0.04513567, 
    0.03938625, 0.08004741, 0.1196289, 0.02022219, 0.001239641, 0.01516589, 
    0.001972762, 0.1110861, 0.1020893, 0.09690307, 0.07959814,
  0.0001140732, 0.0001566823, 0.0001867183, 0.04907022, 0.008983234, 
    0.1315416, 0.08319481, 0.06230163, 0.05945384, 0.06542418, 0.04644642, 
    0.04373771, 0.05607232, 0.05741541, 0.04840353, 0.04950751, 0.1036962, 
    0.1169262, 0.1120669, 0.1309396, 0.1348258, 0.05850818, 0.1414623, 
    0.05382201, 0.06800223, 0.07290584, 0.06230429, 0.100921, -0.0002010379,
  3.967907e-07, 2.07621e-09, 4.869827e-10, 0.001862437, 1.767113e-07, 
    0.03313478, 0.003596692, 0.07355016, 0.05642553, 0.1341395, 0.1320736, 
    0.06260704, 0.05644509, 0.05296824, 0.07372514, 0.0830351, 0.06592327, 
    0.1075443, 0.1375183, 0.1893485, 0.01342216, 0.2616878, 0.06242308, 
    0.03423582, 0.05841209, 0.04459275, 0.05756495, 0.08576218, 6.32997e-07,
  -9.521094e-06, 0.001134946, 0.005960591, 4.064843e-06, 0.003798858, 
    2.850536e-07, 0.002208557, 0.009416142, 0.2556402, 0.02649497, 0.2034509, 
    0.2645365, 0.109102, 0.1377564, 0.1604287, 0.1385699, 0.07643317, 
    0.1480709, 0.3144357, 0.05059667, 0.0365138, 0.05314225, 0.07607585, 
    0.1336112, 0.05330038, 0.116679, 0.05444306, 0.07755256, 0.05729063,
  0.08881283, 0.0457799, 0.05036306, 0.1027631, 0.005087386, 4.232146e-06, 
    0.09847691, 0.01989687, 0.005830542, 0.08642723, 0.09285882, 0.05791832, 
    0.2617543, 0.2390637, 0.1906332, 0.1579243, 0.1674292, 0.3408857, 
    0.1186872, 0.004059158, 0.04362027, 0.04189541, 0.1653519, 0.08338474, 
    0.2495063, 0.1550067, 0.1692863, 0.1638823, 0.1551348,
  0.2057357, 0.1072939, 0.1502931, 0.04046734, 0.1428334, 0.1546938, 
    0.2470027, 0.4081486, 0.2088448, 0.1149596, 0.1221797, 0.1924779, 
    0.3083129, 0.2019956, 0.2548456, 0.3673176, 0.3454149, 0.3012776, 
    0.1651936, 0.08788184, 0.09766393, 0.2455512, 0.409624, 0.4912859, 
    0.2456905, 0.286711, 0.2692158, 0.1614983, 0.1344417,
  0.2546664, 0.3678982, 0.4124509, 0.3342897, 0.350206, 0.3702667, 0.5875816, 
    0.5211202, 0.5108498, 0.5650619, 0.4264564, 0.4395037, 0.2762116, 
    0.2779572, 0.3832482, 0.561614, 0.5193245, 0.4432191, 0.3219247, 
    0.2012022, 0.2124576, 0.3417892, 0.2367159, 0.3477897, 0.4047371, 
    0.2890043, 0.3121737, 0.3025109, 0.2997691,
  0.4275901, 0.3401141, 0.3528514, 0.4384787, 0.4788532, 0.4222037, 
    0.3723982, 0.45011, 0.3731194, 0.4104656, 0.2142497, 0.296876, 0.3385759, 
    0.2590331, 0.3747559, 0.5949885, 0.4346627, 0.311215, 0.426225, 0.389448, 
    0.4122185, 0.4913332, 0.3885109, 0.4810258, 0.2486318, 0.3209895, 
    0.3049425, 0.3138334, 0.5050658,
  0.3620496, 0.4627792, 0.3789185, 0.3588871, 0.4538528, 0.4196868, 
    0.3611569, 0.2849084, 0.1774686, 0.2415849, 0.3066956, 0.3508763, 
    0.3102384, 0.2050606, 0.2417493, 0.2208364, 0.2279089, 0.1320083, 
    0.2565489, 0.3683505, 0.3991112, 0.3281186, 0.3938429, 0.429397, 
    0.2575932, 0.1227164, 0.05180588, 0.2885518, 0.2980332,
  0.4011571, 0.3904168, 0.3796764, 0.3689361, 0.3581957, 0.3474553, 0.336715, 
    0.3304439, 0.3269424, 0.3234409, 0.3199395, 0.316438, 0.3129365, 
    0.3094351, 0.3059961, 0.3187625, 0.331529, 0.3442954, 0.3570619, 
    0.3698284, 0.3825948, 0.4095429, 0.4110183, 0.4124936, 0.413969, 
    0.4154443, 0.4169197, 0.4183951, 0.4097494,
  0.4379379, 0.4876425, 0.3332256, 0.2243068, 0.05525269, 0.01333514, 
    -0.005354541, 0.002617481, 0.06676145, 0.09342811, 0.1810123, 0.210725, 
    0.1718688, -0.01330459, 0.020348, 0.007666067, 0.05507647, 0.1276235, 
    0.1769833, 0.1967713, 0.2526553, 0.3084067, 0.3512322, 0.310327, 
    0.3344935, 0.3604784, 0.1921514, 0.1905759, 0.396949,
  0.4961445, 0.1026705, 0.1615391, 0.07300662, 0.1390645, 0.18424, 
    0.07128848, 0.2008493, 0.1384276, 0.1735115, 0.1818585, 0.1200408, 
    0.233419, 0.1544796, 0.2873972, 0.2983835, 0.3365327, 0.4448873, 
    0.3421892, 0.3589651, 0.3345755, 0.383714, 0.2550424, 0.3158825, 
    0.1718254, 0.379248, 0.4591102, 0.4380554, 0.5796486,
  0.5017018, 0.5117695, 0.5337996, 0.412827, 0.293701, 0.321398, 0.3680078, 
    0.4309689, 0.4784703, 0.3916059, 0.3307101, 0.260083, 0.3201582, 
    0.2683843, 0.1951321, 0.2553948, 0.3425373, 0.3598971, 0.426628, 
    0.3700473, 0.2358655, 0.2000457, 0.2840694, 0.3343823, 0.3024572, 
    0.3401085, 0.4367858, 0.5231026, 0.4613922,
  0.4682131, 0.3530695, 0.3679743, 0.2767177, 0.2526189, 0.2850045, 
    0.2891706, 0.3068145, 0.3334741, 0.3293668, 0.3524442, 0.2112354, 
    0.1264268, 0.1524941, 0.1536352, 0.206284, 0.3621465, 0.2941947, 
    0.4290781, 0.4509788, 0.3967818, 0.3467174, 0.2565017, 0.2419437, 
    0.05947336, 0.2657719, 0.4127762, 0.388299, 0.4736834,
  0.3156771, 0.1583096, 0.1208655, 0.1234735, 0.1544506, 0.1237799, 
    0.1630009, 0.2091623, 0.2027471, 0.236128, 0.1406518, 0.07160152, 
    0.0366749, 0.1743937, 0.2891487, 0.2852083, 0.2288326, 0.2052364, 
    0.2923099, 0.2805457, 0.3162882, 0.3126364, 0.1993761, 0.3557257, 
    0.0608667, 0.1489201, 0.1627852, 0.1170154, 0.2136648,
  0.1338822, 0.1146926, 0.008519578, 0.08092968, 0.1099199, 0.2433275, 
    0.1421195, 0.1650685, 0.277081, 0.01675441, 0.002704366, -1.469821e-05, 
    0.01251046, 0.05115436, 0.1019149, 0.1028785, 0.1554276, 0.1291065, 
    0.1171667, 0.02840507, 0.1676351, 0.1222051, 0.2238234, 0.00143743, 
    0.01552056, 0.2130839, 0.1335876, 0.02836959, 0.1383907,
  0.2016791, 7.4957e-05, -4.309083e-06, 0.03995418, 0.07771175, 0.03660843, 
    0.02120747, 0.03184533, 0.04407504, 0.003913014, 2.915743e-08, 
    8.333897e-06, 0.1555177, 0.08278148, 0.1327521, 0.1654729, 0.03160069, 
    0.04529612, 0.05773523, 0.03027843, 0.04637946, 0.1178029, 0.285669, 
    0.000729791, 0.01095829, 0.1245805, 0.055101, 0.05827567, 0.1380273,
  0.3544381, 0.0756693, 4.484754e-05, 0.04908657, 0.05394664, 0.08786007, 
    0.0894682, 0.01808464, 0.04944599, 0.1685504, 0.02342405, 0.0525564, 
    0.124043, 0.05155827, 0.0261416, 0.02955194, 0.03939911, 0.0223598, 
    0.03224627, 0.01849159, 0.1061975, 0.3088199, 0.475548, 0.03604427, 
    0.001417803, 1.578191e-05, 0.08506917, 0.1924789, 0.5303298,
  0.1079587, 0.1335134, 0.01022173, 0.04612935, 0.2128738, 0.05013064, 
    0.1442731, 0.06669339, 0.09475476, 0.02812857, 0.02445377, 0.1354893, 
    0.02220381, 0.00825009, 0.02044151, 0.08279106, 0.06141896, 0.03527666, 
    0.02527705, 0.06742477, 0.2181115, 0.2930567, 0.01932328, 0.005926296, 
    0.0007389951, 0.06903729, 0.0403181, 0.1150848, 0.1661726,
  3.859271e-05, 4.113483e-05, 9.78892e-05, 0.03602798, 0.02588518, 0.107672, 
    0.07841772, 0.02337349, 0.02624083, 0.0284388, 0.02257521, 0.02945128, 
    0.03962418, 0.04819051, 0.03838296, 0.03843566, 0.0643079, 0.08448181, 
    0.09345706, 0.1031142, 0.1192423, 0.08420821, 0.175357, 0.05229165, 
    0.02749376, 0.03423491, 0.05861167, 0.09651701, -0.0001675856,
  3.423662e-07, 2.631811e-09, 5.016796e-10, 0.0009031215, 2.122459e-06, 
    0.05576509, 0.001602791, 0.01969106, 0.02897597, 0.04116276, 0.07766083, 
    0.04478443, 0.02574755, 0.05244208, 0.03898688, 0.0459227, 0.02534393, 
    0.05283721, 0.1424995, 0.2362201, 0.02298818, 0.1801975, 0.01522072, 
    0.01629106, 0.00755652, 0.01740519, 0.01650642, 0.0601814, 5.235266e-07,
  -1.212327e-05, 0.0005227277, 0.0001813789, 2.252949e-06, 0.004882471, 
    1.167176e-07, 0.001683019, 0.009658335, 0.2392256, 0.01824217, 0.157442, 
    0.2367612, 0.08557327, 0.09921139, 0.08973524, 0.1097053, 0.04252083, 
    0.05824284, 0.1907963, 0.3011151, 0.0395873, 0.02974423, 0.03049695, 
    0.09864035, 0.08116611, 0.04158294, 0.03588992, 0.01719406, 0.06678733,
  0.08441326, 0.02979512, 0.04280436, 0.1077949, 0.001896204, 5.925121e-06, 
    0.09744091, 0.01437362, 0.004419518, 0.07386527, 0.1043141, 0.05040517, 
    0.2293563, 0.1889898, 0.175043, 0.131896, 0.1835856, 0.3614219, 
    0.2060775, 0.002364264, 0.04634612, 0.03726607, 0.1350073, 0.0718947, 
    0.2424052, 0.1357005, 0.1358382, 0.1019301, 0.1303827,
  0.1723759, 0.112425, 0.1852483, 0.05731955, 0.1331086, 0.09986205, 
    0.2449784, 0.3805055, 0.1983867, 0.09761158, 0.1575033, 0.2009416, 
    0.2725576, 0.134185, 0.2058925, 0.3382827, 0.3367289, 0.340533, 
    0.2296813, 0.09578592, 0.08856279, 0.1971695, 0.4240596, 0.4963729, 
    0.2335404, 0.3082671, 0.2264675, 0.1668068, 0.09764914,
  0.2228051, 0.4500422, 0.4244465, 0.3492347, 0.452472, 0.419199, 0.562004, 
    0.5078937, 0.5124549, 0.5003172, 0.4440577, 0.49573, 0.2783806, 
    0.1919352, 0.2487103, 0.5504742, 0.5726612, 0.4461408, 0.3634676, 
    0.2368666, 0.2282689, 0.2889206, 0.1701545, 0.347998, 0.3316482, 
    0.2581606, 0.23113, 0.2570071, 0.239437,
  0.3678586, 0.2563212, 0.3577372, 0.4362176, 0.4376544, 0.370481, 0.4714663, 
    0.4955721, 0.3623634, 0.4641039, 0.2311114, 0.2695084, 0.2798791, 
    0.2426487, 0.4548632, 0.5632554, 0.4724383, 0.2741537, 0.3391547, 
    0.2903713, 0.4348978, 0.5186504, 0.3780279, 0.4486567, 0.187225, 
    0.2978378, 0.3010466, 0.2732091, 0.4423014,
  0.4732055, 0.3797149, 0.4692169, 0.3738399, 0.4633228, 0.4161883, 
    0.3420325, 0.3446869, 0.2454105, 0.3316188, 0.4015019, 0.4838901, 
    0.4234051, 0.3222441, 0.3938825, 0.2717249, 0.2085907, 0.1623472, 
    0.2764181, 0.4086443, 0.4770487, 0.3273473, 0.3445909, 0.5662926, 
    0.2647136, 0.1521201, 0.07533377, 0.3029371, 0.3174112,
  0.3687391, 0.3569036, 0.3450682, 0.3332327, 0.3213972, 0.3095617, 
    0.2977262, 0.2970791, 0.2953565, 0.2936339, 0.2919113, 0.2901886, 
    0.288466, 0.2867434, 0.282182, 0.2952637, 0.3083454, 0.3214271, 
    0.3345089, 0.3475906, 0.3606723, 0.4106136, 0.41109, 0.4115664, 
    0.4120428, 0.4125192, 0.4129955, 0.4134719, 0.3782075,
  0.4419533, 0.502968, 0.3452932, 0.2212962, 0.05127155, 0.01335246, 
    -0.006394508, 0.003034604, 0.05670925, 0.09514991, 0.1390611, 0.1906914, 
    0.1949645, -0.01253211, 0.02570612, 0.02154694, 0.07583605, 0.1848233, 
    0.1987423, 0.1932791, 0.311396, 0.3146628, 0.3231878, 0.3120788, 
    0.2918105, 0.408477, 0.1518375, 0.1584128, 0.3822562,
  0.4931909, 0.09097613, 0.1319014, 0.04031795, 0.09239172, 0.1705225, 
    0.03404727, 0.1509879, 0.1386691, 0.160996, 0.172469, 0.1119673, 
    0.1724578, 0.1330788, 0.2997026, 0.3529975, 0.350062, 0.4636285, 
    0.3820677, 0.3555126, 0.3431656, 0.3590108, 0.2562813, 0.3834167, 
    0.1566209, 0.4305081, 0.5145504, 0.5022886, 0.5902165,
  0.5187011, 0.4870507, 0.5605155, 0.3193162, 0.2106089, 0.2562987, 
    0.3491558, 0.4054252, 0.4629293, 0.3322387, 0.2959277, 0.246157, 
    0.2740662, 0.2353748, 0.1663513, 0.2252602, 0.3306015, 0.3485515, 
    0.4276926, 0.3756288, 0.2404287, 0.1697063, 0.2418337, 0.2953829, 
    0.2827545, 0.3708946, 0.4693073, 0.5231357, 0.5368572,
  0.4147698, 0.3046414, 0.3432089, 0.2247581, 0.2262696, 0.2537316, 0.247569, 
    0.2771378, 0.3088971, 0.2894458, 0.2752218, 0.1294156, 0.09086986, 
    0.09842005, 0.1112199, 0.2251904, 0.3626098, 0.3787942, 0.4193061, 
    0.4217847, 0.3653789, 0.2988685, 0.2106761, 0.1924597, 0.04812489, 
    0.2604046, 0.4985103, 0.3596995, 0.4774581,
  0.2541967, 0.122358, 0.07617686, 0.09966661, 0.1255098, 0.1094333, 
    0.1595745, 0.2131904, 0.1697304, 0.1673099, 0.07992928, 0.04552461, 
    0.01686772, 0.1481611, 0.2598273, 0.2434135, 0.2395989, 0.169998, 
    0.2593627, 0.1746647, 0.2397248, 0.2760136, 0.1671507, 0.3530773, 
    0.0604182, 0.1115802, 0.1884918, 0.1051876, 0.2373418,
  0.1090785, 0.06297213, 0.00442367, 0.06961109, 0.1011282, 0.1957226, 
    0.08623012, 0.06323784, 0.1091872, 0.00654958, 0.005186773, 
    -8.125546e-06, 0.01513531, 0.03765168, 0.07926023, 0.09546313, 0.110767, 
    0.07399157, 0.1387839, 0.01964454, 0.09991282, 0.0457317, 0.09906701, 
    0.002171306, 0.01940304, 0.1979377, 0.1150244, 0.01909465, 0.1180405,
  0.1457663, -0.003665989, -1.77914e-06, 0.02069408, 0.03053638, 0.01644941, 
    0.004633128, 0.009990077, 0.01390127, 0.001671465, 1.050345e-08, 
    -2.607092e-07, 0.0553023, 0.03157058, 0.04100935, 0.09636526, 0.0114168, 
    0.02004644, 0.04422173, 0.01419957, 0.01347693, 0.04475679, 0.1040617, 
    0.026914, 0.005632579, 0.1291342, 0.02375526, 0.02128947, 0.1826952,
  0.512699, 0.2053315, 2.419434e-05, 0.0833275, 0.02207211, 0.03396154, 
    0.0536914, 0.003872739, 0.01115532, 0.03104051, 0.01208018, 0.02657562, 
    0.07833013, 0.02688796, 0.01011489, 0.006173043, 0.005446211, 
    0.003801362, 0.002746724, 0.002520329, 0.03057964, 0.1102124, 0.4212978, 
    0.02227421, 0.0006085417, 1.087808e-05, 0.02043115, 0.05536119, 0.2286514,
  0.1364456, 0.1146838, 0.008375099, 0.04717505, 0.1418705, 0.005966718, 
    0.01817991, 0.02357832, 0.08906966, 0.007896442, 0.005176165, 0.02236613, 
    0.007413236, 0.002170218, 0.005917887, 0.01383843, 0.01794109, 
    0.01690929, 0.004908396, 0.01542579, 0.1012828, 0.5715203, 0.2578862, 
    0.002612358, 0.000282516, 0.02097144, 0.007259195, 0.02095359, 0.2011509,
  1.893265e-05, 2.80283e-05, 9.140209e-05, 0.02794621, 0.04084614, 
    0.01218645, 0.05566216, 0.007838507, 0.01489827, 0.004978664, 
    0.007584536, 0.0108684, 0.02068995, 0.02403802, 0.02643529, 0.02242154, 
    0.03468169, 0.07517716, 0.05385314, 0.05596796, 0.08677719, 0.05561855, 
    0.2710536, 0.03163273, 0.00833069, 0.01837071, 0.01859293, 0.0187696, 
    -0.0001639213,
  3.214287e-07, 3.093326e-09, 5.369879e-10, 0.0002206242, 3.635717e-06, 
    0.01356285, 0.006207392, 0.003538014, 0.01843004, 0.01008512, 0.0450232, 
    0.03540749, 0.005971448, 0.01328306, 0.01429921, 0.009891806, 
    0.004358368, 0.03819354, 0.06563906, 0.1650002, 0.07647558, 0.1366532, 
    0.002120987, 0.002643348, 0.0009909597, 0.005481259, 0.004050389, 
    0.02927036, 4.60711e-07,
  -1.34338e-05, 0.0004588293, 1.59679e-05, 1.676469e-06, 0.001736287, 
    7.554528e-08, 0.001262013, 0.005643739, 0.2124443, 0.01800432, 0.1159298, 
    0.2058658, 0.06107633, 0.07340092, 0.05264043, 0.06530306, 0.01727893, 
    0.02406072, 0.08430471, 0.3025029, 0.03496508, 0.01727579, 0.01421149, 
    0.05619637, 0.04685836, 0.00996457, 0.006641938, 0.003445982, 0.0764247,
  0.06044205, 0.0155255, 0.03025673, 0.09494511, -0.0002585256, 3.962812e-06, 
    0.08708284, 0.01024977, 0.002828737, 0.0672719, 0.1000115, 0.0297451, 
    0.1811705, 0.1595082, 0.143354, 0.111519, 0.1987977, 0.389883, 0.4652945, 
    0.0003139784, 0.04357747, 0.02937701, 0.1196491, 0.06059264, 0.2203256, 
    0.1193523, 0.09217304, 0.07513481, 0.09406406,
  0.130279, 0.119494, 0.1563088, 0.06030194, 0.09965602, 0.08963615, 
    0.2209447, 0.3382098, 0.1663773, 0.09336004, 0.1618354, 0.2335874, 
    0.2279054, 0.09485158, 0.1594094, 0.3097217, 0.2910945, 0.4087386, 
    0.3239917, 0.1201735, 0.08160648, 0.1496805, 0.3752493, 0.5167453, 
    0.2204024, 0.2684461, 0.1982409, 0.1348683, 0.07680754,
  0.1871134, 0.5453229, 0.4487002, 0.3812311, 0.5544403, 0.4342655, 
    0.5044224, 0.4880956, 0.4697851, 0.4343133, 0.4066494, 0.5566297, 
    0.2894199, 0.1357876, 0.1613068, 0.5079533, 0.6245975, 0.4264641, 
    0.4239499, 0.2781139, 0.2873174, 0.2466642, 0.1187524, 0.3616424, 
    0.2691352, 0.228372, 0.1691129, 0.2019416, 0.2096089,
  0.3020937, 0.1970429, 0.39248, 0.397191, 0.4128465, 0.3154859, 0.5262301, 
    0.5800613, 0.3428121, 0.4835581, 0.2705797, 0.3247803, 0.2140126, 
    0.2591623, 0.4130277, 0.4999444, 0.5221508, 0.2986518, 0.2712528, 
    0.2280259, 0.4469479, 0.5368671, 0.3735945, 0.4203551, 0.12705, 
    0.2657523, 0.3376901, 0.2070636, 0.3884433,
  0.4458711, 0.3223206, 0.4645796, 0.3576745, 0.4865402, 0.3672934, 
    0.3427358, 0.362883, 0.3867911, 0.4704109, 0.5031629, 0.4772614, 
    0.5066708, 0.4458327, 0.4930153, 0.400587, 0.3827448, 0.3371817, 
    0.4717416, 0.5617194, 0.5170814, 0.3111561, 0.3119049, 0.6222464, 
    0.2307646, 0.2048974, 0.07227916, 0.298639, 0.3680839,
  0.3176644, 0.307829, 0.2979935, 0.2881581, 0.2783226, 0.2684872, 0.2586517, 
    0.2122488, 0.2127047, 0.2131605, 0.2136164, 0.2140723, 0.2145281, 
    0.214984, 0.2187635, 0.2282443, 0.237725, 0.2472058, 0.2566866, 
    0.2661674, 0.2756482, 0.3185237, 0.3184226, 0.3183214, 0.3182202, 
    0.318119, 0.3180178, 0.3179166, 0.3255328,
  0.422233, 0.4866165, 0.3236612, 0.2017286, 0.0533503, 0.009776613, 
    -0.005108756, 0.006055201, 0.03585017, 0.06384519, 0.08432591, 0.1042749, 
    0.2373538, -0.008515546, 0.04352887, 0.04308631, 0.1312361, 0.2164659, 
    0.1936801, 0.1803326, 0.3194492, 0.3126574, 0.2920103, 0.2685625, 
    0.2469226, 0.4451488, 0.1223205, 0.1287345, 0.3453165,
  0.4669122, 0.07980765, 0.1151464, 0.01870627, 0.05492458, 0.1381796, 
    0.01531256, 0.09472045, 0.120872, 0.1412736, 0.148165, 0.09956892, 
    0.1161371, 0.09992841, 0.2949974, 0.3629529, 0.3558673, 0.4345193, 
    0.3625433, 0.3455211, 0.3300619, 0.348706, 0.2521071, 0.3999777, 
    0.161632, 0.4525117, 0.509997, 0.4910749, 0.5550396,
  0.4908776, 0.448508, 0.5182695, 0.2352116, 0.1474304, 0.2320146, 0.2889876, 
    0.3695264, 0.416174, 0.2904668, 0.2588224, 0.2237737, 0.2241112, 
    0.2195845, 0.1279917, 0.2043506, 0.3121765, 0.3421637, 0.4067375, 
    0.3484944, 0.2109314, 0.1361675, 0.2062034, 0.2409675, 0.2706289, 
    0.4065346, 0.4645884, 0.5100975, 0.5337751,
  0.3542493, 0.2698013, 0.2616516, 0.1539374, 0.1852533, 0.1972122, 
    0.2051692, 0.228435, 0.2727667, 0.2356867, 0.1992597, 0.08657648, 
    0.05706197, 0.06852791, 0.08239746, 0.2058255, 0.3207579, 0.3452578, 
    0.3670657, 0.3664609, 0.3013524, 0.2132034, 0.1539076, 0.1448019, 
    0.03290029, 0.2331578, 0.5245925, 0.35392, 0.46772,
  0.1880944, 0.09638884, 0.04307881, 0.08088212, 0.1051637, 0.0866602, 
    0.1453358, 0.1664405, 0.1474217, 0.119759, 0.05003601, 0.02842254, 
    0.01040442, 0.1086107, 0.2336147, 0.1838409, 0.187813, 0.1537476, 
    0.2170594, 0.1529108, 0.1684068, 0.2242572, 0.1356511, 0.3427378, 
    0.05966081, 0.09615067, 0.1808818, 0.09885381, 0.2060634,
  0.06808885, 0.03207226, 0.001869636, 0.05079028, 0.06374007, 0.1563319, 
    0.05211329, 0.02803674, 0.04787856, 0.003528521, 0.00265912, 
    -1.864558e-06, 0.01492215, 0.03180308, 0.05757897, 0.0771651, 0.07840354, 
    0.0464217, 0.1214723, 0.01027024, 0.05863903, 0.0135106, 0.04372505, 
    0.0007150202, 0.02481875, 0.1423786, 0.08196148, 0.01447447, 0.1025905,
  0.05898117, 0.007765987, -5.700479e-07, 0.006288357, 0.01124188, 
    0.008426056, 0.001374171, 0.00336205, 0.005824671, 0.0009407232, 
    1.589701e-08, -5.290589e-07, 0.02190886, 0.01006025, 0.01206229, 
    0.05174258, 0.00209719, 0.01113099, 0.02009843, 0.01310418, 0.005101156, 
    0.01741066, 0.04564751, 0.01677295, 0.003503075, 0.1161673, 0.01174545, 
    0.00961529, 0.09578894,
  0.2304241, 0.09583212, 9.607101e-06, 0.1155406, 0.005121364, 0.007190798, 
    0.02456864, 0.0007367511, 0.003242366, 0.01004398, 0.004567724, 
    0.004216939, 0.03733721, 0.006743196, 0.005016001, 0.0004663864, 
    0.0009847158, 0.0009805274, 0.0006558824, 0.000993156, 0.01161351, 
    0.04139627, 0.1583548, 0.01602709, 0.0004481673, 2.320669e-06, 
    0.00512493, 0.01919841, 0.08977224,
  0.03374876, 0.1235105, 0.006944756, 0.03120963, 0.02735189, 0.0009017069, 
    0.005425033, 0.01046907, 0.07031322, 0.003835203, 0.001277208, 
    0.005587649, 0.001847102, 0.0005947467, 0.001795148, 0.005049064, 
    0.002436619, 0.003318101, 0.0002993599, 0.00308041, 0.02178002, 
    0.2217942, 0.1694423, 0.001854236, 0.0001956515, 0.006596077, 
    0.001454916, 0.002696267, 0.05438004,
  1.65139e-05, 2.818469e-05, 6.29936e-05, 0.01599967, 0.03514025, 
    0.003127126, 0.04634216, 0.0009995963, 0.007546286, 0.0006338227, 
    0.001191283, 0.003395492, 0.008964668, 0.01044549, 0.01290115, 
    0.005229636, 0.009526696, 0.04339281, 0.03941269, 0.01683552, 0.04077837, 
    0.0175045, 0.2631142, 0.01483302, 0.003617847, 0.003503252, 0.004872094, 
    0.003606812, -0.0001802788,
  3.029366e-07, 3.303112e-09, 5.80882e-10, -3.920342e-05, 1.617896e-06, 
    0.003227064, 0.007171091, 0.001008565, 0.01092244, 0.003685851, 
    0.02222161, 0.01056719, 0.0008263471, 0.002748501, 0.003970732, 
    0.002139501, 0.0009430745, 0.01117558, 0.02157259, 0.08415186, 
    0.01473454, 0.1072209, 0.0006379969, -0.0008400539, 0.0002816484, 
    0.001078971, 0.001434066, 0.007750235, 4.280249e-07,
  -2.094304e-05, 2.966969e-05, -2.287176e-05, 1.406447e-06, 0.0004077366, 
    6.704872e-08, 0.0008989014, 0.003603613, 0.1859577, 0.01989814, 
    0.07747938, 0.1408337, 0.03728522, 0.02984624, 0.02189457, 0.04609839, 
    0.007324733, 0.01277843, 0.03973502, 0.225659, 0.02858683, 0.0138121, 
    0.01038097, 0.0213339, 0.02434678, 0.003981688, 0.001128635, 0.001073907, 
    0.07317824,
  0.04894012, 0.00732678, 0.02066713, 0.0907087, -0.001266728, 1.9552e-06, 
    0.07059006, 0.006653429, 0.001814176, 0.0580344, 0.09617451, 0.01772914, 
    0.1418121, 0.1385061, 0.1123494, 0.08841456, 0.1808905, 0.3323011, 
    0.3375421, 0.00135495, 0.04041015, 0.02330335, 0.1187156, 0.05402049, 
    0.1789702, 0.1052979, 0.05548613, 0.05159538, 0.07202418,
  0.09244727, 0.1556971, 0.1622568, 0.1265649, 0.08979266, 0.07832267, 
    0.1764107, 0.2871163, 0.1279199, 0.09082054, 0.1655703, 0.2620376, 
    0.1854408, 0.05936433, 0.121254, 0.2882462, 0.2377859, 0.3971016, 
    0.3916941, 0.1416951, 0.0693121, 0.1098716, 0.3064429, 0.5117496, 
    0.1914597, 0.2146591, 0.1778275, 0.1018161, 0.06050482,
  0.1439909, 0.5620277, 0.4008927, 0.4110936, 0.58039, 0.3942644, 0.4288454, 
    0.4902914, 0.4076455, 0.3743381, 0.3543484, 0.5572488, 0.2907425, 
    0.1221648, 0.1091173, 0.4485219, 0.6478743, 0.4046048, 0.4067494, 
    0.2733743, 0.259895, 0.1874986, 0.09318814, 0.381217, 0.2113606, 
    0.1956189, 0.1163229, 0.1553174, 0.1790616,
  0.2612858, 0.1544652, 0.3917586, 0.3481296, 0.3836988, 0.2721657, 0.577482, 
    0.6023906, 0.3292715, 0.5126985, 0.3252585, 0.3154621, 0.2355002, 
    0.2233808, 0.3787042, 0.4379407, 0.5734391, 0.3299545, 0.2229544, 
    0.1902992, 0.3973699, 0.5201549, 0.3934427, 0.4350571, 0.09529673, 
    0.2094208, 0.3735697, 0.1429891, 0.3470527,
  0.3960688, 0.2551997, 0.3863824, 0.3411411, 0.389217, 0.3552572, 0.373395, 
    0.3957369, 0.4739106, 0.5682777, 0.5943586, 0.5232859, 0.5136658, 
    0.4729515, 0.5078768, 0.5394704, 0.5759344, 0.6414928, 0.6816387, 
    0.6905626, 0.5653968, 0.3064269, 0.2949937, 0.6020629, 0.2030613, 
    0.2260658, 0.05756183, 0.3254219, 0.4518593,
  0.2415785, 0.2322704, 0.2229622, 0.2136541, 0.2043459, 0.1950378, 
    0.1857296, 0.1573247, 0.1593292, 0.1613338, 0.1633383, 0.1653429, 
    0.1673474, 0.169352, 0.1819609, 0.1890661, 0.1961713, 0.2032765, 
    0.2103816, 0.2174868, 0.224592, 0.2496219, 0.2498203, 0.2500187, 
    0.2502171, 0.2504156, 0.250614, 0.2508124, 0.2490251,
  0.3670374, 0.4349916, 0.2706092, 0.1777086, 0.0587694, 0.002015429, 
    -0.001513353, 0.009392481, 0.03089148, 0.04127084, 0.06783509, 
    0.07461668, 0.1946911, -0.003636626, 0.06448599, 0.2063838, 0.265135, 
    0.2500308, 0.1905358, 0.1889943, 0.3268748, 0.3267424, 0.2468797, 
    0.2158811, 0.2771341, 0.4896464, 0.1202201, 0.1068302, 0.3101336,
  0.4483697, 0.07225443, 0.09784575, 0.01419885, 0.03223802, 0.104692, 
    0.007699213, 0.05727031, 0.09919143, 0.1147117, 0.1169153, 0.09484456, 
    0.08282038, 0.0866776, 0.2741874, 0.339586, 0.3394513, 0.3962393, 
    0.3288692, 0.3259272, 0.2942671, 0.3794539, 0.2550367, 0.3579538, 
    0.1504823, 0.4321795, 0.4514183, 0.4535568, 0.517407,
  0.4462974, 0.3796625, 0.4169348, 0.1633319, 0.09522523, 0.1603434, 
    0.2386068, 0.3110862, 0.3458228, 0.2368751, 0.2192548, 0.1712491, 
    0.1891579, 0.1838551, 0.09011851, 0.1674889, 0.2395269, 0.3329077, 
    0.3634958, 0.2958074, 0.1719389, 0.1107312, 0.1704928, 0.1897963, 
    0.2631232, 0.3819176, 0.434517, 0.4602929, 0.4669515,
  0.3143908, 0.2404651, 0.1869293, 0.108051, 0.1369961, 0.1429683, 0.1558297, 
    0.1812805, 0.2208367, 0.1691598, 0.1380311, 0.05292534, 0.03072283, 
    0.04969559, 0.05785089, 0.1599299, 0.2671852, 0.2509514, 0.2878932, 
    0.2971539, 0.2252168, 0.1319485, 0.09744254, 0.1096067, 0.01956576, 
    0.205365, 0.4642463, 0.3323246, 0.454789,
  0.1273991, 0.0702565, 0.02279001, 0.06331521, 0.07887229, 0.06213869, 
    0.1104111, 0.1082386, 0.1296353, 0.08212858, 0.03172302, 0.01478213, 
    0.008585016, 0.0699994, 0.1929322, 0.1445548, 0.1480285, 0.1110126, 
    0.1631208, 0.1256615, 0.1174241, 0.1723536, 0.1027477, 0.3188817, 
    0.05718733, 0.08307479, 0.1459369, 0.08013079, 0.1564499,
  0.03546108, 0.01673029, 0.0006919007, 0.02978923, 0.0388835, 0.1059333, 
    0.03009155, 0.01463514, 0.02698377, 0.00226876, 0.001135794, 
    -2.069741e-07, 0.01324672, 0.02374706, 0.03160537, 0.04103729, 
    0.05462705, 0.03089621, 0.1101142, 0.006503329, 0.02912431, 0.005187488, 
    0.02148698, 0.0002462929, 0.02368125, 0.08981489, 0.06320423, 
    0.009416196, 0.07196698,
  0.02757891, 0.003592575, -2.243444e-07, 0.002457513, 0.001895668, 
    0.0035057, 0.0007735569, 0.001693566, 0.003368472, 0.0006226902, 
    1.470136e-08, -1.992875e-07, 0.008383151, 0.003958362, 0.005243564, 
    0.01965133, 0.0004959517, 0.005281306, 0.008488565, 0.007363019, 
    0.002660478, 0.008751464, 0.02610712, 0.008800058, 0.003299634, 
    0.1023052, 0.00413252, 0.003493462, 0.04471533,
  0.1105679, 0.031155, 5.662167e-06, 0.1061028, 0.001054625, 0.00143399, 
    0.008501126, 0.0002146395, 0.001739829, 0.005423687, 0.001476904, 
    0.00107907, 0.01412698, 0.002403834, 0.002347655, 1.583782e-05, 
    0.0001147762, 0.0005106403, 0.00034222, 0.0005449522, 0.006227451, 
    0.02094655, 0.07837852, 0.01145921, 0.0001894417, 2.59284e-07, 
    0.002483749, 0.009433866, 0.04156594,
  0.01272394, 0.1193518, 0.01352167, 0.0191037, 0.01150138, 0.0003689234, 
    0.002720105, 0.005940972, 0.05671922, 0.00610156, 0.0006352687, 
    0.002363221, 0.0007350366, 0.0002461973, 0.0008676922, 0.002624372, 
    0.0009529347, 0.0005538422, 0.0001138807, 0.001349437, 0.008162991, 
    0.1011649, 0.09641343, 0.001235425, 0.000101923, 0.003020108, 
    0.0004528686, 0.001074434, 0.02241882,
  9.566319e-06, 1.573296e-05, 2.849835e-05, 0.02110265, 0.02404552, 
    0.001530901, 0.03194289, 0.000310198, 0.002773885, 0.0002543556, 
    0.0001176742, 0.001027195, 0.003500936, 0.004066691, 0.005181202, 
    0.00128212, 0.002517336, 0.02280099, 0.02588734, 0.005137098, 0.0130265, 
    0.004822503, 0.2133584, 0.01250743, 0.001849815, 0.0009210407, 0.0020869, 
    0.001496814, -0.0003465707,
  2.858527e-07, 3.292161e-09, 5.998726e-10, -2.903973e-05, -3.565141e-07, 
    0.001349877, 0.006716126, 0.0005662544, 0.01033124, 0.00192085, 
    0.009074482, 0.002745463, 0.0001853562, 0.0009067348, 0.0009316905, 
    0.001067147, 0.0003500074, 0.004147834, 0.008512255, 0.05595232, 
    0.005575842, 0.0879577, 0.0003630787, -0.0008735982, 0.0001445667, 
    0.0002048476, 0.0006715285, 0.003975617, 4.12195e-07,
  -1.345383e-05, -1.625516e-05, -1.648887e-05, 1.282072e-06, -0.0003091044, 
    6.339317e-08, 0.0005236187, 0.003107129, 0.1640778, 0.01013649, 
    0.05282569, 0.09428664, 0.02106967, 0.01505672, 0.01045839, 0.03657856, 
    0.002320525, 0.008136029, 0.01809707, 0.1639053, 0.02582054, 0.01051084, 
    0.009318009, 0.02510891, 0.009141027, 0.002098654, 0.0005487355, 
    0.00055822, 0.06369631,
  0.03572395, 0.003326227, 0.01517266, 0.09214238, -0.001198096, 
    1.340621e-06, 0.05222855, 0.004792522, 0.001033642, 0.04975551, 
    0.08543601, 0.0122242, 0.1178027, 0.1058312, 0.08432914, 0.06279651, 
    0.1464476, 0.2446818, 0.2353259, 0.004296976, 0.03663373, 0.01659278, 
    0.09474181, 0.04676867, 0.128916, 0.06551942, 0.04057136, 0.02828935, 
    0.04666623,
  0.05876298, 0.1604743, 0.1529725, 0.1544488, 0.08783332, 0.06239987, 
    0.1311124, 0.232564, 0.09902436, 0.08384453, 0.1545358, 0.249827, 
    0.1421181, 0.03538425, 0.08340449, 0.2385388, 0.1838923, 0.3687077, 
    0.3459612, 0.1418038, 0.04762599, 0.08733404, 0.2472345, 0.476712, 
    0.1535211, 0.1859045, 0.1509226, 0.0772297, 0.04409578,
  0.09967768, 0.5289468, 0.3334807, 0.3972779, 0.5577818, 0.3263054, 
    0.3573808, 0.4400222, 0.3429376, 0.3079332, 0.307784, 0.5047915, 
    0.2641505, 0.09854179, 0.07994308, 0.3902938, 0.6230149, 0.3691943, 
    0.3893872, 0.2591035, 0.216685, 0.1308012, 0.07762784, 0.356133, 
    0.1712155, 0.1620744, 0.07726373, 0.1199394, 0.1296714,
  0.227277, 0.1087913, 0.3640846, 0.2724423, 0.3400875, 0.2276736, 0.5447321, 
    0.5461646, 0.2821091, 0.484574, 0.379357, 0.3105731, 0.2531164, 
    0.2366671, 0.4184235, 0.3806913, 0.5007764, 0.3280002, 0.200572, 
    0.1491537, 0.3619062, 0.4722344, 0.4231003, 0.3861209, 0.07106789, 
    0.1548094, 0.3925876, 0.09861573, 0.3086969,
  0.355908, 0.1952445, 0.3577788, 0.3391644, 0.3256596, 0.365661, 0.4104172, 
    0.4952285, 0.6056015, 0.5748088, 0.5705632, 0.5070526, 0.524092, 
    0.5094835, 0.481117, 0.5568786, 0.6191752, 0.6876889, 0.675731, 
    0.6730019, 0.5845328, 0.2996371, 0.2691517, 0.6101322, 0.1660968, 
    0.2003681, 0.04692787, 0.2963956, 0.4433075,
  0.1916758, 0.183056, 0.1744362, 0.1658163, 0.1571965, 0.1485767, 0.1399568, 
    0.1105477, 0.1099612, 0.1093747, 0.1087883, 0.1082018, 0.1076154, 
    0.1070289, 0.1095668, 0.1176376, 0.1257084, 0.1337792, 0.1418501, 
    0.1499209, 0.1579917, 0.1785329, 0.1796683, 0.1808038, 0.1819393, 
    0.1830747, 0.1842102, 0.1853456, 0.1985717,
  0.3217882, 0.3519646, 0.2329805, 0.1473613, 0.0508168, -0.001264639, 
    0.003647941, 0.01328611, 0.02873717, 0.03359657, 0.04124446, 0.03278234, 
    0.1165133, -0.0003721526, 0.1384847, 0.2958283, 0.3558269, 0.2450667, 
    0.1669643, 0.2111429, 0.3177315, 0.3697894, 0.2084718, 0.1587764, 
    0.2905149, 0.5354882, 0.112615, 0.08415007, 0.2565246,
  0.3939466, 0.05816627, 0.0796608, 0.008934479, 0.01624894, 0.08399283, 
    0.00376038, 0.03750653, 0.06591957, 0.09498348, 0.08478942, 0.08279867, 
    0.06019184, 0.08367199, 0.2418926, 0.2701819, 0.2732566, 0.3249527, 
    0.2992163, 0.2934331, 0.2769578, 0.3564659, 0.2382936, 0.3023461, 
    0.1405425, 0.4003028, 0.3705885, 0.3931373, 0.4518498,
  0.3773195, 0.3144782, 0.3245072, 0.1223676, 0.06493104, 0.1102933, 
    0.190942, 0.2422422, 0.2806453, 0.1796955, 0.172107, 0.125065, 0.1587301, 
    0.1478228, 0.06182119, 0.1288299, 0.1836663, 0.2841351, 0.3009969, 
    0.2266479, 0.1279564, 0.08643901, 0.1320246, 0.1382862, 0.2153723, 
    0.3038931, 0.3723585, 0.3917949, 0.39372,
  0.2734613, 0.1989717, 0.1415565, 0.08064408, 0.1024154, 0.1010679, 
    0.1159609, 0.138647, 0.1652218, 0.1131753, 0.09688802, 0.03110815, 
    0.02010367, 0.02934282, 0.03357236, 0.1188468, 0.2053578, 0.1632561, 
    0.2031908, 0.2231272, 0.1547236, 0.08312068, 0.0581106, 0.08429381, 
    0.01040806, 0.1572754, 0.3899392, 0.2786421, 0.3978317,
  0.08309031, 0.04710423, 0.0120932, 0.04424816, 0.05212852, 0.03975873, 
    0.07498761, 0.0630626, 0.09304731, 0.05328458, 0.01830715, 0.006964727, 
    0.006460387, 0.0418243, 0.1541539, 0.09483723, 0.09809692, 0.076065, 
    0.1104906, 0.09884834, 0.0854762, 0.1259344, 0.06071803, 0.2887163, 
    0.05424495, 0.06164384, 0.09678629, 0.06341507, 0.1152152,
  0.0227283, 0.008814172, 0.0002067184, 0.01597072, 0.02251005, 0.06077346, 
    0.01671213, 0.009184399, 0.0180971, 0.001633024, 0.0006063334, 
    7.327923e-08, 0.01333986, 0.01279049, 0.01497785, 0.0213358, 0.02862932, 
    0.02116145, 0.0706988, 0.00418696, 0.01203962, 0.002720243, 0.01365832, 
    0.0001303668, 0.01977673, 0.05165802, 0.0444724, 0.00496705, 0.04438677,
  0.01651811, 0.0007691341, -8.462368e-08, 0.001092638, -0.0006058835, 
    0.001596999, 0.0005142418, 0.001070147, 0.002275232, 0.0004589966, 
    1.33289e-08, -2.90747e-08, 0.0047133, 0.00236114, 0.003184227, 
    0.007016949, 0.0002391695, 0.00188919, 0.003186132, 0.003356345, 
    0.00169397, 0.005472523, 0.01754626, 0.005899549, 0.001842545, 
    0.08733524, 0.001620968, 0.00190117, 0.02530913,
  0.06538634, 0.01664765, 3.478233e-06, 0.08162678, 0.0003564244, 
    0.0005591376, 0.002685783, 0.0001115276, 0.001127408, 0.003908263, 
    0.0007498704, 0.0005916053, 0.004856349, 0.0008182814, 0.001045288, 
    1.898459e-05, 9.017698e-05, 0.0003336626, 0.0002250506, 0.0003570626, 
    0.004037845, 0.01319687, 0.04919498, 0.01344837, 0.0001371967, 
    -2.70628e-06, 0.001850744, 0.005810376, 0.02441349,
  0.005612474, 0.102713, 0.009386773, 0.01052387, 0.006972603, 0.0002115329, 
    0.001676294, 0.002887133, 0.04124014, 0.007079591, 0.0004009002, 
    0.001438686, 0.0004424438, 0.0001581611, 0.0005529911, 0.001641238, 
    0.0005491815, 0.0002753326, 6.364599e-05, 0.0008184666, 0.004719807, 
    0.05827975, 0.0654663, 0.000562282, 4.646009e-05, 0.00177302, 
    0.0002537198, 0.000603338, 0.01251144,
  5.0662e-07, 6.284583e-06, 9.873461e-06, 0.02048614, 0.01194632, 
    0.0009496551, 0.02142102, 0.0001851554, 0.00106949, 0.0001786875, 
    4.26564e-05, 0.0002999347, 0.001278779, 0.001578955, 0.001839225, 
    0.000389435, 0.0009031346, 0.01060909, 0.01362264, 0.001928799, 
    0.00462871, 0.002048669, 0.1594842, 0.01432513, 0.0009724763, 
    0.0004039371, 0.000962691, 0.0008937176, -0.0003659208,
  2.737235e-07, 3.265527e-09, 5.879072e-10, -6.721478e-06, -4.004424e-08, 
    0.0008130253, 0.004659743, 0.0003814998, 0.01081554, 0.001324389, 
    0.003473565, 0.0006272739, 7.212296e-05, 0.0005299317, 0.0003293705, 
    0.0006956777, 0.0002280542, 0.001741082, 0.005124885, 0.03970927, 
    0.002889062, 0.07341449, 0.000241124, -0.0008563491, 8.963658e-05, 
    8.253624e-05, 0.000407652, 0.00251695, 4.082114e-07,
  -9.287454e-06, -1.872759e-06, -3.418133e-05, 1.212741e-06, -0.0006006359, 
    5.925671e-08, -0.0002978644, 0.002607619, 0.1464759, 0.00448505, 
    0.03136431, 0.06661088, 0.005558781, 0.006906981, 0.005471375, 
    0.02185999, 0.0008948223, 0.004156096, 0.009606781, 0.1324064, 
    0.02198533, 0.006060278, 0.008557919, 0.01771372, 0.004022335, 
    0.001276672, 0.0003867809, 0.0003688487, 0.05020649,
  0.02443162, 0.001677528, 0.01167418, 0.08764891, -0.0009645533, 
    1.147618e-06, 0.03762339, 0.003889688, 0.0006195257, 0.03769214, 
    0.07455358, 0.008922412, 0.1002193, 0.06979097, 0.0565283, 0.03953586, 
    0.10648, 0.1722531, 0.1607075, 0.004500622, 0.02785121, 0.01033296, 
    0.06381813, 0.04121148, 0.08518416, 0.03495623, 0.02443174, 0.01388046, 
    0.02594557,
  0.03776899, 0.1423534, 0.1413144, 0.2043172, 0.07403705, 0.04896878, 
    0.09739025, 0.1949023, 0.07673962, 0.0803812, 0.1289573, 0.2177973, 
    0.09557324, 0.02209699, 0.04856624, 0.1693898, 0.1215505, 0.2979177, 
    0.2948099, 0.1295311, 0.03718395, 0.06731397, 0.195721, 0.421424, 
    0.1129654, 0.1545641, 0.1141454, 0.05417781, 0.0275236,
  0.05774578, 0.4850605, 0.2545254, 0.3662409, 0.5134385, 0.2758421, 
    0.292584, 0.3589689, 0.2810365, 0.245744, 0.2400312, 0.4425765, 
    0.2186932, 0.0745513, 0.06274723, 0.3194099, 0.5801033, 0.3235476, 
    0.3474569, 0.2354467, 0.1858734, 0.09265286, 0.05947464, 0.3165676, 
    0.1422253, 0.1376621, 0.04873063, 0.08582514, 0.08352201,
  0.169846, 0.07120416, 0.3139033, 0.1929909, 0.2878824, 0.1878321, 
    0.5315598, 0.4688058, 0.2366761, 0.4343773, 0.3594569, 0.2647117, 
    0.2410156, 0.2348462, 0.3924226, 0.3409779, 0.4034825, 0.2814007, 
    0.1725486, 0.1058815, 0.3132755, 0.414817, 0.4346492, 0.3747126, 
    0.05791067, 0.1173567, 0.4354697, 0.07058691, 0.2481072,
  0.3609563, 0.1654555, 0.3773958, 0.2974596, 0.2612306, 0.3255517, 
    0.4194621, 0.5240006, 0.5654632, 0.4858616, 0.5171703, 0.4471731, 
    0.4774881, 0.4576621, 0.4109626, 0.4945709, 0.5462567, 0.627538, 
    0.5961452, 0.5745552, 0.5203026, 0.274417, 0.2500713, 0.6623439, 
    0.1382584, 0.1494234, 0.05748178, 0.2803285, 0.377091,
  0.1450771, 0.1399068, 0.1347365, 0.1295663, 0.124396, 0.1192257, 0.1140554, 
    0.09328189, 0.09239095, 0.09150001, 0.09060907, 0.08971813, 0.0888272, 
    0.08793626, 0.09448988, 0.09930926, 0.1041286, 0.108948, 0.1137674, 
    0.1185868, 0.1234062, 0.134139, 0.1353809, 0.1366227, 0.1378645, 
    0.1391064, 0.1403482, 0.1415901, 0.1492133,
  0.2666386, 0.2702276, 0.1631273, 0.0950949, 0.02821552, 0.0002410492, 
    0.004735288, 0.01182858, 0.02681756, 0.03425533, 0.02957552, 0.01250773, 
    0.0463785, -0.0002636056, 0.2295888, 0.2602369, 0.3392835, 0.2470767, 
    0.1313448, 0.2362663, 0.3353011, 0.3947441, 0.1777362, 0.1255442, 
    0.2622779, 0.5522221, 0.09942926, 0.06831055, 0.2159703,
  0.3367965, 0.04192925, 0.07061903, 0.005956918, 0.009705982, 0.07361044, 
    0.002009052, 0.03013029, 0.03982295, 0.08392555, 0.07145581, 0.07076834, 
    0.0551658, 0.0762437, 0.2165436, 0.2178804, 0.2354166, 0.2847053, 
    0.2664791, 0.2478518, 0.2311326, 0.3048382, 0.2048404, 0.2698382, 
    0.1325419, 0.3626038, 0.3109876, 0.3371708, 0.3978944,
  0.327417, 0.2598218, 0.26756, 0.1001734, 0.0512054, 0.08925804, 0.1574672, 
    0.1967696, 0.2364801, 0.1459799, 0.1411352, 0.09997175, 0.1321924, 
    0.1192779, 0.04671658, 0.104924, 0.1511192, 0.2453301, 0.2520995, 
    0.1782074, 0.09978953, 0.07270622, 0.1056551, 0.1056257, 0.1663031, 
    0.2343368, 0.3216631, 0.3481429, 0.3563714,
  0.2393945, 0.1691534, 0.1158878, 0.06410249, 0.08651372, 0.07914273, 
    0.1042773, 0.1075749, 0.1253295, 0.08373673, 0.06957674, 0.02101968, 
    0.01477716, 0.0178311, 0.0210397, 0.08070526, 0.1438413, 0.1142772, 
    0.1430606, 0.1675504, 0.1091486, 0.05856847, 0.03871736, 0.07205746, 
    0.00629351, 0.1170113, 0.3226529, 0.2312885, 0.3263368,
  0.05583838, 0.02913878, 0.007538743, 0.03005516, 0.03605896, 0.02651372, 
    0.05152381, 0.03923964, 0.0649056, 0.03608731, 0.01287895, 0.00414733, 
    0.003601967, 0.02711089, 0.1235276, 0.05755602, 0.06470881, 0.05329658, 
    0.07154105, 0.07389132, 0.05749207, 0.09210116, 0.0379022, 0.2592733, 
    0.05322812, 0.04195154, 0.06137937, 0.04572759, 0.07418044,
  0.01656235, 0.005169056, -1.704205e-05, 0.007968306, 0.01236555, 
    0.03421665, 0.009068327, 0.006675553, 0.01370047, 0.001297239, 
    0.0004338328, 9.918821e-08, 0.01314852, 0.007147536, 0.007620513, 
    0.01211179, 0.0146837, 0.01334167, 0.04408397, 0.002064049, 0.005931705, 
    0.002170365, 0.01031405, 9.931091e-05, 0.01677048, 0.02964641, 
    0.01899563, 0.002519407, 0.02705264,
  0.01169984, -3.15384e-05, 9.555869e-09, 0.0006618807, -0.0009240531, 
    0.0007162756, 0.0003861239, 0.0007784114, 0.001719889, 0.0003677386, 
    1.325703e-08, 1.944565e-08, 0.003270282, 0.001698516, 0.00228149, 
    0.003368855, 0.0001626256, 0.0008637466, 0.001406672, 0.001600021, 
    0.001236328, 0.003968006, 0.01326541, 0.004338145, 0.001539643, 
    0.07775329, 0.0007285754, 0.001374945, 0.01761862,
  0.04659648, 0.01151379, 9.295974e-06, 0.0665364, 0.0001776366, 0.000341953, 
    0.0009421125, 7.793523e-05, 0.0008352592, 0.003106748, 0.0005227652, 
    0.0004111393, 0.002112882, 0.0003946547, 0.0006057587, 3.682205e-05, 
    0.0001544344, 0.00024818, 0.0001694933, 0.0002648392, 0.002989166, 
    0.009575715, 0.03558382, 0.01329679, 0.0004695029, -8.62115e-06, 
    0.001515831, 0.004149194, 0.01688862,
  0.003169856, 0.07624681, 0.00751129, 0.007137256, 0.004971662, 
    0.0001430395, 0.001187532, 0.001394009, 0.03053145, 0.01099062, 
    0.0002927437, 0.001032825, 0.0003122622, 0.0001186895, 0.0004044748, 
    0.001174634, 0.0003770724, 0.0001878423, 4.40396e-05, 0.0005815099, 
    0.003290518, 0.04044024, 0.04932489, 0.0003955374, 8.25057e-05, 
    0.001231933, 0.0001882751, 0.0004095919, 0.008529133,
  4.843827e-05, 6.153101e-06, -5.396832e-06, 0.01819805, 0.006590484, 
    0.0006788684, 0.01753132, 0.0001346438, 0.0005978865, 0.0001478968, 
    4.100499e-05, 0.0001855902, 0.0006329569, 0.000761901, 0.0009675469, 
    0.0001713166, 0.0005420293, 0.005060473, 0.006437693, 0.0009814481, 
    0.002168967, 0.001026328, 0.1286811, 0.01792893, 0.0005376687, 
    0.0002640334, 0.0006072763, 0.0005655593, -0.0003253057,
  2.672091e-07, 3.12738e-09, 5.819785e-10, -1.429305e-06, 6.45145e-08, 
    0.0005728548, 0.002932065, 0.0002915677, 0.01805098, 0.00104878, 
    0.001560581, 0.000307763, 4.988958e-05, 0.000372402, 0.0001782491, 
    0.0005170829, 0.0001697929, 0.00102955, 0.003719046, 0.0263308, 
    0.001867607, 0.06311021, 0.0001823995, -0.001278308, 6.358884e-05, 
    5.7836e-05, 0.0002881623, 0.001826703, 4.105756e-07,
  -6.604114e-06, 1.797772e-06, 5.78016e-05, 1.173532e-06, -0.0005972859, 
    5.556763e-08, -0.0004239786, 0.002940426, 0.1336291, 0.002341069, 
    0.01754011, 0.04447448, 0.002151206, 0.003445176, 0.003638608, 
    0.01117572, 0.0005702479, 0.002062361, 0.00621023, 0.1134959, 0.01898739, 
    0.004964612, 0.007482474, 0.004577232, 0.002540398, 0.000929424, 
    0.0002977371, 0.0002786877, 0.03957236,
  0.01892638, 0.0008683454, 0.008583497, 0.08397796, -0.0008115627, 
    1.049151e-06, 0.02839907, 0.003343404, 0.0004453833, 0.02944719, 
    0.06480727, 0.005229144, 0.08103034, 0.04545356, 0.03931586, 0.02498729, 
    0.07584134, 0.1151346, 0.1204114, 0.003845007, 0.02209491, 0.006150467, 
    0.04707021, 0.03214094, 0.05676188, 0.01947116, 0.01340144, 0.007074955, 
    0.01786544,
  0.02636811, 0.132355, 0.1313976, 0.2042139, 0.0666201, 0.04226164, 
    0.07936638, 0.1692485, 0.06807028, 0.07373452, 0.1137112, 0.1984519, 
    0.06591316, 0.01634044, 0.03044342, 0.1158159, 0.07696804, 0.2247486, 
    0.2429641, 0.1182993, 0.03158622, 0.05510344, 0.1662072, 0.3804539, 
    0.09020051, 0.1315943, 0.0871161, 0.03693495, 0.01702601,
  0.03742779, 0.4410405, 0.2075138, 0.3271264, 0.4717986, 0.2556799, 
    0.249434, 0.3024826, 0.2357764, 0.2105654, 0.1984896, 0.3947447, 
    0.1963739, 0.06820314, 0.05393925, 0.2575963, 0.5306668, 0.282758, 
    0.3138117, 0.2163795, 0.1644783, 0.07267734, 0.0486874, 0.2843544, 
    0.1184564, 0.1217025, 0.03351127, 0.05794166, 0.05568545,
  0.1105122, 0.04485044, 0.2710573, 0.1308258, 0.2413522, 0.159564, 
    0.4849744, 0.4052806, 0.2167584, 0.3668453, 0.3496704, 0.2168351, 
    0.214749, 0.183025, 0.322174, 0.314079, 0.3563786, 0.2428461, 0.1422758, 
    0.07566065, 0.2797647, 0.3587637, 0.3983201, 0.4022223, 0.04848752, 
    0.09577822, 0.5173379, 0.05431551, 0.1992969,
  0.3425989, 0.1465676, 0.3512646, 0.2445603, 0.221528, 0.2605468, 0.3197008, 
    0.4418309, 0.4542563, 0.3369473, 0.3761163, 0.331755, 0.3661325, 
    0.3289419, 0.2895608, 0.3583616, 0.3779941, 0.4303399, 0.424073, 
    0.446384, 0.4375142, 0.229377, 0.2511006, 0.7089525, 0.1288943, 
    0.1309497, 0.08881734, 0.2296103, 0.3486348,
  0.1148572, 0.1120314, 0.1092055, 0.1063797, 0.1035539, 0.100728, 
    0.09790219, 0.0886993, 0.08827149, 0.08784369, 0.08741588, 0.08698808, 
    0.08656027, 0.08613247, 0.08542802, 0.08857436, 0.09172071, 0.09486706, 
    0.0980134, 0.1011597, 0.1043061, 0.1181829, 0.1182902, 0.1183975, 
    0.1185048, 0.1186121, 0.1187194, 0.1188267, 0.1171179,
  0.2275236, 0.1835084, 0.1124453, 0.06560344, 0.02572574, 0.01040247, 
    0.005971111, 0.01297857, 0.02504399, 0.03443964, 0.02523353, 0.006703308, 
    0.02876401, 0.00129987, 0.2868323, 0.2105265, 0.3051422, 0.2683051, 
    0.1281934, 0.2421194, 0.3600459, 0.4057689, 0.1683508, 0.1167942, 
    0.2571289, 0.5395383, 0.09481393, 0.05929774, 0.1977943,
  0.3144908, 0.03769628, 0.0741586, 0.004517409, 0.009175724, 0.0697417, 
    0.001795327, 0.02817399, 0.04891618, 0.08244053, 0.07201464, 0.06625804, 
    0.05765997, 0.07389435, 0.1958826, 0.1931015, 0.2240266, 0.2639551, 
    0.2502565, 0.2287827, 0.2019344, 0.2718116, 0.1874912, 0.2463149, 
    0.1270892, 0.3355467, 0.2847499, 0.3098446, 0.3667446,
  0.3030265, 0.2356138, 0.2438195, 0.0899016, 0.04491774, 0.07953227, 
    0.1414617, 0.1769458, 0.2196624, 0.1292237, 0.1239637, 0.08827604, 
    0.1111361, 0.1022857, 0.03987286, 0.09084586, 0.1319588, 0.2107466, 
    0.2153513, 0.1518145, 0.08623314, 0.06295853, 0.09009543, 0.08843251, 
    0.1364162, 0.2043713, 0.2963045, 0.3220621, 0.3337009,
  0.1871125, 0.1461033, 0.09866693, 0.05638086, 0.07240677, 0.06738731, 
    0.08909384, 0.08755285, 0.1039017, 0.07064465, 0.05545734, 0.01643516, 
    0.01155045, 0.01346481, 0.01636071, 0.06071268, 0.1052247, 0.0897563, 
    0.1118458, 0.1281193, 0.08392191, 0.04668458, 0.02974408, 0.07985205, 
    0.004647697, 0.091662, 0.2678879, 0.2019966, 0.2659689,
  0.04337506, 0.02004641, 0.005804365, 0.02272788, 0.02788019, 0.01998162, 
    0.03545004, 0.02709883, 0.04613109, 0.02746103, 0.008061307, 0.002797188, 
    0.002915164, 0.01939486, 0.1078033, 0.04020424, 0.04849, 0.04057566, 
    0.05067548, 0.05672048, 0.04204862, 0.06888485, 0.02586349, 0.2514599, 
    0.04020089, 0.02943515, 0.0429119, 0.03048577, 0.05088559,
  0.01289121, 0.003998871, -0.0001321902, 0.005318767, 0.007478536, 
    0.02150427, 0.005987123, 0.005504313, 0.01153734, 0.001122652, 
    0.0003308352, 1.002551e-07, 0.01573081, 0.004815855, 0.004740036, 
    0.007749696, 0.008829172, 0.008762775, 0.02997071, 0.001168796, 
    0.003974294, 0.001976359, 0.008666245, 8.867282e-05, 0.02699324, 
    0.0197077, 0.009457033, 0.001690994, 0.01947539,
  0.009434316, -0.0001119247, 5.401942e-08, 0.0005181877, -0.001247508, 
    0.0004292393, 0.0003278039, 0.0006484115, 0.001453096, 0.0003188809, 
    1.253971e-08, 6.395176e-08, 0.002629239, 0.001382317, 0.001858912, 
    0.002101882, 0.0001308879, 0.0006129973, 0.0009288372, 0.001075465, 
    0.001016678, 0.003277369, 0.01124668, 0.003478057, 0.0146402, 0.08570705, 
    0.0004755616, 0.001144812, 0.0140338,
  0.03754952, 0.009093536, 0.0005493229, 0.07059684, 0.0001227323, 
    0.0002613507, 0.0005587317, 6.422067e-05, 0.0006959939, 0.002470255, 
    0.0004199614, 0.0003318771, 0.001558653, 0.0002923284, 0.0004540569, 
    3.893468e-05, 0.0001562498, 0.0002066968, 0.0001417068, 0.0002208763, 
    0.002497197, 0.007873799, 0.02896381, 0.07675862, 0.004341473, 
    0.0004602743, 0.001203439, 0.0033787, 0.01343347,
  0.002340382, 0.09022201, 0.01172686, 0.00685345, 0.003981578, 0.0001103978, 
    0.0009421101, 0.0009440698, 0.04693691, 0.03785008, 0.0002417194, 
    0.0008095755, 0.0002499421, 9.934242e-05, 0.0003320315, 0.000944545, 
    0.0002976442, 0.0001512057, 3.617438e-05, 0.0004734643, 0.002633231, 
    0.0320094, 0.04086027, 0.008413951, 0.002079254, 0.0009936941, 
    0.0001595477, 0.000322569, 0.006678816,
  0.00106712, 0.0001243363, -0.0001059127, 0.01365743, 0.00427095, 
    0.0005473539, 0.01156796, 0.0001104521, 1.789271e-05, 0.0001288161, 
    3.88382e-05, 0.0001340056, 0.0004489961, 0.0004908354, 0.0006874714, 
    0.0001202296, 0.0004178755, 0.003265024, 0.003599721, 0.0007025382, 
    0.001410982, 0.0007098879, 0.1929687, 0.03312383, 0.0003804338, 
    0.0002071454, 0.0004727411, 0.0004533248, 0.004602252,
  2.692685e-07, 3.123852e-09, 5.872728e-10, -2.110033e-07, 7.52668e-08, 
    0.0004558509, 0.003722445, 0.0001816611, 0.03122176, 0.0006642638, 
    0.0009842498, 0.0002100959, 4.126709e-05, 0.0002998224, 0.0001275259, 
    0.0004263442, 0.0001414097, 0.000775286, 0.003058426, 0.01847417, 
    0.00142163, 0.05998581, 0.0001538627, -0.002287161, 5.044287e-05, 
    4.751321e-05, 0.0002357814, 0.001511708, 4.151867e-07,
  -4.83921e-06, 2.709657e-06, 0.0004063698, 1.165704e-06, -0.0002947316, 
    5.315402e-08, 0.0001857975, 0.009303202, 0.1372637, 0.001814993, 
    0.01160044, 0.02693775, 0.001336888, 0.002219109, 0.002871503, 
    0.007073794, 0.0004482766, 0.001366145, 0.004949592, 0.1019818, 
    0.01803239, 0.02483481, 0.01151742, 0.002281931, 0.002000897, 
    0.0007580654, 0.0002306873, 0.0002347695, 0.03412094,
  0.01588899, 0.0002315744, 0.007206303, 0.0889897, -0.0007702659, 
    9.974241e-07, 0.02402467, 0.002899379, 0.0003353616, 0.02547703, 
    0.07230451, 0.003061822, 0.06300259, 0.03262535, 0.02681208, 0.01780359, 
    0.05411011, 0.06887695, 0.09826196, 0.003227384, 0.02029381, 0.004613212, 
    0.04361898, 0.02531456, 0.03961326, 0.01065737, 0.008784557, 0.004601385, 
    0.01448448,
  0.01960849, 0.141954, 0.1391166, 0.1988378, 0.06139865, 0.03798229, 
    0.07336389, 0.1700522, 0.07464091, 0.07218129, 0.1210959, 0.1998073, 
    0.05045483, 0.01379543, 0.02320415, 0.08001926, 0.05175721, 0.1670144, 
    0.2035378, 0.1245476, 0.03344787, 0.05185183, 0.1705296, 0.3956879, 
    0.08422016, 0.1081412, 0.06918492, 0.02758285, 0.01109993,
  0.02764055, 0.4501102, 0.2086305, 0.3273067, 0.471325, 0.2488216, 
    0.2417137, 0.2920272, 0.2470481, 0.2215959, 0.2005016, 0.3887757, 
    0.1960899, 0.09817198, 0.05035035, 0.2219887, 0.5377855, 0.2739043, 
    0.3374504, 0.211865, 0.1721844, 0.07580965, 0.04222283, 0.2867485, 
    0.09929136, 0.1087917, 0.0266023, 0.03920185, 0.04117603,
  0.08599441, 0.03446462, 0.2939194, 0.1020569, 0.2055997, 0.1410729, 
    0.4706522, 0.3824696, 0.2217622, 0.3512412, 0.4119214, 0.222714, 
    0.2052329, 0.1511523, 0.2693366, 0.3015147, 0.3516908, 0.2285372, 
    0.1163851, 0.05786064, 0.2453677, 0.3107182, 0.3777584, 0.4280698, 
    0.03892134, 0.09690797, 0.5880013, 0.05517634, 0.1676404,
  0.3293134, 0.1332178, 0.3282363, 0.2147776, 0.1946496, 0.2316261, 
    0.2553374, 0.3571357, 0.3617134, 0.2493993, 0.2883559, 0.2410494, 
    0.2652721, 0.2290161, 0.1996144, 0.2630488, 0.2941378, 0.3457967, 
    0.3479673, 0.3760552, 0.3936873, 0.2172264, 0.2716382, 0.711871, 
    0.1226922, 0.1512974, 0.1191882, 0.2188384, 0.3307973,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0002440453, 0.0004155463, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 4.266566e-07, -5.580489e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, -1.397395e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, -2.173573e-05, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, -1.092543e-05, 0, 0, 0.0008720229, 0.0003618316, 
    -6.710902e-05, 0, 2.657368e-05, 0, 0, -1.203781e-05, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2.934569e-06, 0, -3.586625e-05, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -3.911105e-05, 0, 0, 0,
  0, 0, -7.886582e-06, -0.0001454141, -1.90556e-06, 0, 0, 0, 0, 0, 0, 0, 0, 
    8.075333e-07, -1.104076e-05, 0.00393435, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -2.579026e-05, 0, 0, 0,
  0, 0.001009976, 1.680938e-05, 0, -1.061939e-05, 0, 0, 0, -1.706336e-06, 0, 
    0, 0, 0, 3.768605e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0007393617, 
    -3.657608e-05, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, -0.0001155509, 0, -1.09318e-05, 0.002537977, 
    0.0009053955, 0.0008951779, 0.002172753, 1.388955e-05, 0, 0.00116237, 
    -4.570588e-05, 0, 0, 0, 0, 0, -6.126465e-06, 0, -8.539599e-06, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, -6.655159e-06, 4.627523e-05, 0, -7.121073e-05, 
    0.0001488225, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2.460009e-05, 0, 0, 0, 0, 
    0, 0, 0, 0, -6.074974e-05, 0, 0, 0,
  0, 0, 0.0005685939, -4.407767e-05, 0.000171381, -4.346728e-06, 
    -7.624858e-06, 0, 0, 0, 0, 0, 0, 0.0006513351, 0.003529301, 0.005217134, 
    0, 0, 0, 0, 0, 0, 0, -7.931319e-06, -3.771099e-06, -5.994646e-05, 0, 0, 0,
  0, 0.002363423, 8.465659e-06, 0, -7.209826e-05, 0, 0, 0, 1.328772e-05, 0, 
    0, 0, 0, -1.228383e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.000805977, 
    -6.889108e-05, 0, 0.0002421083, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0.001745693, -2.893791e-05, -5.921533e-05, 
    0.004055782, 0.0009166794, 0.002477263, 0.004443524, -2.242988e-05, 
    -7.372283e-06, 0.001555428, 0.00120193, 0.001234475, -3.999038e-05, 
    0.0001401254, 0, 0, -6.454226e-05, 0, 0.0004721639, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, -5.989643e-05, 0.003949693, 0, -0.0001787008, 
    0.004517681, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.008911253, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, -3.187162e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0009342927, 0, -3.032959e-05, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0001939473, 
    -2.989771e-05, 0, 0, 0, 0, 0, 0, 0, -0.0001091091, 0.000973811, 0, 0,
  0, -3.490283e-05, 0.002185281, 0.002674634, 0.0001904906, 4.998212e-05, 
    -0.0001088375, 0, 0, 0, 0, -4.548292e-05, 0, 0.009959997, 0.009115256, 
    0.00681699, 0.001244814, 0, 0, 0, 0, 0, 0, 0.0001374317, 4.320898e-05, 
    -8.884956e-05, 0, 0, 0,
  0, 0.004925863, 0.0003700269, 0, -0.0001524986, 0, 0, 0, 0.0004451533, 0, 
    -1.490287e-05, -2.419787e-05, -6.091396e-07, 0.0002598021, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.0008315154, -5.506168e-05, 0, 0.00203351, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0.004474666, -8.844726e-05, -0.0001666039, 
    0.005925538, 0.001820327, 0.006812559, 0.008231418, -7.618484e-05, 
    -1.145422e-05, 0.004796765, 0.003711542, 0.004141059, 0.001480117, 
    0.001125382, 0, -7.968488e-06, -0.0001292902, -3.172671e-05, 
    0.0006111814, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, -9.317223e-05, 0.01326941, -8.283371e-05, 
    0.0006662451, 0.01324745, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01283252, 0, 0, 0, 
    0, 0,
  0, 0, 0, 0, -1.818945e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, -1.831888e-05, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -2.473362e-05, -1.266748e-05, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, -2.865726e-05, 0, 0, 0, 0, 0, 0, 0, 0, -5.766806e-07, 0, 0, 0, 
    0, 0.0005776687, 0, 0, 0, 0, 0, 0.001854798, 0, 0, 0, 0,
  0, 0, 0, -2.146829e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -3.148739e-05, 
    0, -1.967653e-05, 0, 0, 0, 0, 0, 0.002159495, 0, 0.0003126549, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.000108399, -1.118932e-05, 0, 
    0.004763357, 0.0002272904, 0, 0, 0, 0, 0, 0, 0.0001689562, -9.237786e-05, 
    0.003423538, 0, 0,
  0, -9.799196e-05, 0.00293086, 0.004931384, 0.0002528698, -6.315537e-05, 
    -0.000221417, 0, -3.885973e-05, 0, 0, -8.632464e-05, -6.779077e-05, 
    0.01761575, 0.01508638, 0.01113783, 0.006652525, 0, 0, 0, 0, 0, 0, 
    4.342123e-05, 1.776326e-05, -0.0001516575, 0, 0, 0,
  -5.074746e-06, 0.008368881, 0.004074507, 0, 0.0006405406, -6.656837e-06, 
    -8.061976e-06, 0, 0.008045668, -6.083902e-06, -0.0001776419, 
    -8.03846e-05, -8.699815e-07, 0.001027355, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0008552884, -6.268333e-06, -4.678502e-05, 0.005330778, 0, 0,
  0, 0, 0, 0, -1.587328e-06, 0, 0, 0.009127958, 0.00113923, -0.0002243902, 
    0.01025386, 0.006094719, 0.01134437, 0.02036252, 0.000881449, 
    0.0008940165, 0.01126297, 0.01748969, 0.007418744, 0.003351537, 
    0.002837576, -0.0001724648, -4.723229e-05, -0.0001561846, -0.0001045616, 
    0.003010146, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, -0.0001622767, 0.03026855, -0.0002636894, 
    0.002584249, 0.02980274, 0, 0, 0, 0, 0, 0, 0.0005726349, 0, 0, 0.0148278, 
    -1.760481e-05, 0.001046788, 0, 0, 0,
  0, 0, 0, 0, -0.0001012767, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0006591894, 
    -2.50705e-05, 0, 0, 0, 0, 0, 0, 0, 2.685829e-08, 0, 0.001483457, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.002436892, 0, 0, 0, 0, 
    0, 0, 0.0008531575, -6.370882e-05, 2.888695e-05, -3.106963e-06, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0003913539, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0008097178, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 3.775357e-05, 5.356846e-05, -1.386089e-05, 0, 0, 0, 0, 0, 0, 0, 
    1.842277e-05, 0, 0, 0, 0, 0.003505494, 0, 0, 0, 0, 0, 0.004352283, 
    0.001222783, 0, 0, 0,
  0, 0, 0, 0.001390799, 0, 0, 0, 0, 0, 0, 0, 0, 0, -8.197431e-05, 0, 0, 
    0.005658449, 4.060432e-06, 0.001120792, 0, -1.1141e-06, 0, 0, 0, 
    0.004896586, -1.811987e-05, 0.00140363, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.002438122, -5.92344e-05, 0, 
    0.0102823, 0.0003208097, -3.085803e-06, 0, 0, 0, 0, -9.287453e-08, 
    0.001356502, -0.0001163367, 0.005664409, 0, 0,
  0, -0.0002296995, 0.003555409, 0.008386916, 0.0007873134, 0.00103744, 
    -0.0003319276, -8.292765e-06, 0.0004387535, 0, 0, -0.0001565866, 
    -0.0003222412, 0.02811295, 0.02165913, 0.01714922, 0.01355612, 0, 0, 0, 
    0, 0, 0, -0.0001087223, 0.0002764579, -0.000197537, 0.003935363, 0, 0,
  -8.951227e-05, 0.01401709, 0.007778207, 0, 0.002481332, -1.242921e-05, 
    -8.061976e-06, -9.806692e-06, 0.02021842, -1.545755e-05, 0.000138159, 
    -0.0001799783, 0.003705739, 0.00118344, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.008534447, 8.328418e-05, -0.0001167532, 0.009279553, 0, 0,
  0, 0, 0, 0, 1.365609e-05, 0, 0, 0.01349821, 0.006098887, 0.001225965, 
    0.02188949, 0.01745724, 0.02170665, 0.04022959, 0.002273865, 0.003750033, 
    0.02225393, 0.03300764, 0.01014962, 0.008114519, 0.008634877, 
    -0.0004027265, -0.0003120649, 0.0004357678, 0.0002908785, 0.006949409, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 3.018409e-05, 0, 8.340162e-05, 0.05248897, 
    -0.0004775838, 0.006665227, 0.05763189, -4.856278e-05, 0, -3.375357e-05, 
    -2.258896e-05, 0, 0, 0.0009611068, 0, -1.078253e-05, 0.01840845, 
    9.634609e-06, 0.006315681, 0, 0, 0,
  0, 0, 0, 0, -9.263463e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001152359, 
    0.0001336227, 0, 0, 0, 0, 0, 0, 0, 0.002052897, 0.001236945, 0.003625826, 
    0, 0, 0,
  0, 0, 0, 0, -2.293612e-05, 0, 0, 0, 0, 0, 0, 0, -2.856716e-05, 
    9.520261e-06, 0, 0.0001584694, -6.063387e-05, 0.008779778, 0, 0, 0, 0, 0, 
    -4.052185e-06, 0.003113586, 0.0006835302, 0.003848509, -7.532645e-05, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0008801354, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.003582535, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  -4.185187e-07, 0, 0, 0.0006003164, 0.002188307, 0.0007630375, 0, 0, 0, 0, 
    0, -1.666773e-07, 0, 0.001869295, 0.0001009252, 0, 0, 0, 0.004864963, 
    -2.949944e-05, 0, 0, 0, 0, 0.007521208, 0.0114219, 0, 0, -1.077152e-05,
  0, 0, 0, 0.01012119, 0.0002591156, 0, 0, 0, 0, 0, 0, 0, -1.019991e-05, 
    0.00195699, 0, 0, 0.01695674, 0.001892371, 0.01196544, -5.015193e-06, 
    0.0005876061, 0, 0, 0, 0.007906216, 0.001095717, 0.004195622, 
    -2.644398e-07, 0,
  0, 0.0002312079, 0.0003762548, 0, -2.601693e-05, 0, -6.326762e-05, 
    0.001479769, 0, 0, 2.043773e-10, 0, 0, 0.006175743, -0.0003003488, 
    -0.0004148457, 0.01796905, 0.005871839, 0.001600538, 0, 0, 0, 0, 
    -3.714981e-07, 0.005090437, 0.001584651, 0.008108177, 0, 0,
  0, 0.0009595202, 0.004556596, 0.01709203, 0.01280185, 0.008490996, 
    -8.702373e-05, -6.040886e-05, 0.003130525, -8.535376e-06, -1.264213e-09, 
    0.0003045498, 0.002064267, 0.04475073, 0.03290631, 0.02802943, 
    0.03089889, 0, 0, 0, 0, 0, 0, 0.001983662, 0.003290962, 0.002274634, 
    0.008366544, 0, 0,
  0.0001183356, 0.02668799, 0.01176774, -1.653015e-05, 0.004752836, 
    6.007907e-05, -2.703687e-05, -5.703585e-05, 0.04270187, -5.434079e-05, 
    0.001284159, -0.0005163419, 0.006158968, 0.007317816, 0, 0.0009917178, 0, 
    -5.115798e-06, 0, 0, 0, 0, -2.45184e-08, 0.01305181, 0.0005555419, 
    0.001371669, 0.01792403, -1.246134e-05, 0,
  0, 0, 7.022102e-05, 0, -1.755526e-05, 0, -5.650578e-06, 0.01693289, 
    0.01212222, 0.002910496, 0.04302636, 0.03344912, 0.0412599, 0.06763509, 
    0.006484502, 0.01013453, 0.03839047, 0.04613888, 0.01481945, 0.01434537, 
    0.02735517, -0.000425032, 0.002128122, 0.004461371, 0.001136933, 
    0.01640177, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0.002698736, -5.462414e-05, 0.004515881, 0.07604823, 
    0.0006102713, 0.01785107, 0.07538486, -4.761626e-05, 0, 0.0003049125, 
    3.71101e-05, 0, 0, 0.001852468, -1.723297e-05, -7.089111e-05, 0.03376165, 
    1.365056e-05, 0.01016504, 0, 0, 0,
  0, 0, 0, 0.001863572, 0.0009992243, 0, 0, 0, -1.444917e-07, 0, 
    -7.497937e-06, 0, 0.001702966, -2.809452e-08, 0.004682661, 0.003159589, 
    0, 0, 0, 0, 0, -0.0002062582, 0.000102406, 0.006125308, 0.004144168, 
    0.008483405, -3.421426e-05, 0, 0,
  0, 0, 0, 0, 0.0002658076, 0, 0, 0, 0, 0, 0, 3.021898e-09, 0.002205839, 
    0.002423963, 4.566245e-05, 0.002135257, 0.001532076, 0.01182368, 0, 0, 0, 
    0, 0.0003503492, 0.005334367, 0.01149127, 0.002387584, 0.005295664, 
    -0.0001854238, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.004556863, 0, 0, 0, 0, 
    -1.620069e-06, 0, 0, 0, 0, 0, 0, -9.637613e-05, -1.95001e-05, 
    -7.280772e-06, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.001790809, 0,
  0, 0, 0, 0, 0, 0, 0.0002098225, -8.951107e-06, 0, 0, 0, 0, 0, 0, 
    0.004311728, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.227866e-05, 0,
  0.0008533139, -2.61781e-05, 0, 0.002112468, 0.01024797, 0.005052563, 
    0.002308398, -1.748454e-05, 0, 0, -4.782893e-06, -0.0001089735, 0, 
    0.003566333, 0.0008377308, 0, -1.172428e-06, 0.003776185, 0.01060708, 
    0.001031569, 0, 0, 0, 0, 0.01086504, 0.0224502, 0.00148316, 
    -5.825792e-06, 0.001609437,
  0, 0, 0.0003644419, 0.0292026, 0.0009917325, 0, 0, 0, 0, 0, 1.155357e-05, 
    0, 6.661312e-05, 0.004291837, -3.836095e-05, -7.430003e-06, 0.03105378, 
    0.004884696, 0.03420154, -0.0001159746, 0.001050398, 0, 0, 0, 0.01642995, 
    0.009933171, 0.0166248, 0.001654052, 0,
  0, 0.0006256954, 0.0004413008, 0, 0.0001080424, 1.229243e-05, 
    -0.0001084732, 0.002734053, 0, 0, 8.823264e-07, -9.990669e-09, 
    1.433551e-07, 0.01708439, 0.0007262888, 0.002312546, 0.03609782, 
    0.009919955, 0.00942198, -1.340881e-08, -9.555196e-07, 0, 0, 
    -1.145128e-05, 0.01036346, 0.01375915, 0.01210383, 0, 0,
  0, 0.005629796, 0.01113113, 0.04629212, 0.02727093, 0.02525379, 
    0.002824517, 0.0009612984, 0.007509382, 5.140114e-05, 0.0009390241, 
    0.005292627, 0.02073509, 0.08173247, 0.04791878, 0.05194962, 0.05170664, 
    0, 0, 0, 0, 0, 0, 0.02213839, 0.04512138, 0.0138921, 0.0110139, 0, 0,
  0.01035715, 0.04624914, 0.04030578, 0.0001690879, 0.03218371, 0.005307198, 
    0.003068603, 0.0004019627, 0.06830542, 0.0002577346, 0.01788406, 
    0.006709528, 0.03092931, 0.01015278, -3.513364e-05, 0.00194208, 0, 
    -7.279358e-05, 0, 0.002688721, -0.0001556442, 0, 1.228796e-05, 
    0.03428496, 0.02033698, 0.003891579, 0.02675158, -7.363526e-06, 
    1.849796e-09,
  0, 0, 0.0002033314, -1.416004e-08, 0.003323031, -2.534368e-05, 
    -3.342597e-05, 0.0195278, 0.02683356, 0.01127878, 0.06331655, 0.06516846, 
    0.08275299, 0.1147913, 0.03139395, 0.02581234, 0.06177139, 0.0613837, 
    0.02075711, 0.02479993, 0.04353866, 0.00303446, 0.02923288, 0.0182036, 
    0.009557357, 0.02857651, -1.753062e-06, -1.625658e-06, 4.114267e-07,
  0, 0, 0, 1.058984e-07, 0, 0, -6.965986e-05, 0.01820435, 0.004944021, 
    0.01295374, 0.1021501, 0.004094883, 0.02879283, 0.09148262, 0.002664915, 
    0.000631562, 0.001345614, 0.005303461, 0.001107539, -5.599885e-05, 
    0.004296022, 0.0002268974, 0.0005397032, 0.04458178, 0.001587489, 
    0.02022827, 0.0008393396, 0, -0.0001008954,
  0, 0, 0, 0.003245535, 0.005351978, 0, 0, 0, -3.086939e-05, 3.423897e-05, 
    -1.358531e-06, 8.956346e-06, 0.005542288, -3.99949e-06, 0.01088596, 
    0.01522503, 0.0004772469, 5.491735e-05, 1.186895e-05, 0, 0, 0.008777819, 
    0.006390339, 0.008818756, 0.0113569, 0.01717503, -0.0001355402, 0, 
    -3.843951e-05,
  0, 0, 0, 0, 0.0006579827, 0, 0, 0, 0, 0, 0, 5.56327e-05, 0.005828421, 
    0.009448292, 0.005907423, 0.009206202, 0.007519037, 0.01669238, 
    0.0003843115, 0, 0, 0, 0.0003371852, 0.01609482, 0.03061039, 0.007538982, 
    0.01010219, 0.0002515179, 0.0001101573,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2.680881e-05, 0.008081416, 
    0.002114825, -1.780016e-05, 0, 0.0009762705, 0.0002458466, 0, 0, 0, 0, 0, 
    0.006889176, 7.78352e-06, 0.0008049367, 3.890189e-05, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.898303e-06, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.00273398, 0, -1.284701e-05, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -4.968161e-07, 0, 0, 0, 0, 0, 
    0, -1.968125e-05, 0, 0, 0, 0, 0.002325105, 0,
  0, 1.531047e-05, 0, 0, 0, 9.275068e-05, 0.003438642, -7.674372e-05, 0, 
    -3.963848e-05, -9.129271e-06, 0, 0, 0, 0.006407732, -8.740925e-06, 0, 0, 
    0, -0.0001204025, -8.71548e-06, 0, 0.001342568, -6.31136e-09, 
    -1.198031e-08, 0.001364156, 0.004842142, 0.00281366, 0,
  0.0028777, 0.000204956, 5.547377e-05, 0.004997342, 0.02653132, 0.009675602, 
    0.006592997, 0.001632132, -6.511388e-07, 0, 9.201045e-06, 0.0006170053, 
    -2.204794e-05, 0.01812931, 0.004673836, 0.003247989, -6.712967e-05, 
    0.01187435, 0.03073593, 0.008408245, 0.001653901, -3.3032e-05, 0, 
    -5.893882e-06, 0.01282773, 0.03859258, 0.01035574, -0.0001496284, 
    0.007036483,
  -7.695762e-07, -2.015892e-09, 0.0005426778, 0.04680926, 0.004723831, 
    3.627802e-05, 0, 5.165047e-06, 1.770571e-05, 4.330853e-08, -5.523908e-06, 
    6.13027e-10, 0.0008967293, 0.006269502, 0.001463366, -0.0002257712, 
    0.04125025, 0.007585557, 0.06330242, 0.004401097, 0.002784343, 0, 
    -5.413706e-10, -2.749303e-09, 0.02611575, 0.01862407, 0.03113891, 
    0.005613518, 3.265328e-05,
  3.650028e-08, 0.003101487, 0.002669731, 0.0001024944, 0.0007464117, 
    0.0007510026, -0.0002069595, 0.00522538, -4.810452e-09, -4.642074e-06, 
    0.0001490984, -8.247212e-06, 9.376727e-05, 0.03859461, 0.00143285, 
    0.008008054, 0.06169191, 0.03010768, 0.02232595, 0.0004119622, 
    0.0007088711, 1.676909e-05, 0, 0.003298101, 0.08184618, 0.02960259, 
    0.02716647, -4.172362e-05, -5.693825e-06,
  -1.105841e-05, 0.1752227, 0.02190333, 0.07791632, 0.06177722, 0.05353752, 
    0.02309882, 0.04782963, 0.01175826, 0.0007614404, 0.005957081, 
    0.03177416, 0.1373795, 0.1949356, 0.09204993, 0.1339755, 0.08236376, 
    -2.710389e-06, 0.0004144793, 0, 0, 5.546969e-08, 5.597974e-06, 0.1483787, 
    0.2222472, 0.0765797, 0.03892229, 0.001939051, 0.0001615494,
  0.01135063, 0.1030238, 0.1240697, 0.001203791, 0.05107465, 0.01151961, 
    0.02495497, 0.01714459, 0.114847, 0.04407483, 0.07086244, 0.07459296, 
    0.1894952, 0.08110113, -0.0001418409, 0.02443183, 6.728944e-07, 
    -0.0001536823, -2.125393e-05, 0.009524162, 0.002029855, -1.003268e-06, 
    0.0001816053, 0.1187077, 0.1587963, 0.0140106, 0.06153038, 6.631942e-05, 
    3.750314e-07,
  -1.070944e-08, -1.773916e-05, 0.0009351966, -1.507964e-06, 0.01123205, 
    0.002660622, -0.0001756057, 0.0311285, 0.04011958, 0.08986658, 0.1764277, 
    0.2287837, 0.2490885, 0.2281699, 0.1399145, 0.0502567, 0.08169641, 
    0.08383483, 0.02599158, 0.0564678, 0.05031554, 0.01391564, 0.03947363, 
    0.06625126, 0.07001086, 0.05333705, 0.0002902853, 0.0005034658, 
    -5.892245e-05,
  -5.869474e-10, 0, -2.935203e-06, 1.165271e-05, 5.778124e-05, 1.71013e-05, 
    0.0008205834, 0.03630566, 0.008340884, 0.02885117, 0.1428073, 0.0336825, 
    0.02836228, 0.1063634, 0.06046748, 0.01009849, 0.009386136, 0.03066781, 
    0.0148938, 0.0004898928, 0.01089292, 0.01010533, 0.01392884, 0.05598518, 
    0.01296427, 0.0361973, 0.003361522, 2.347595e-05, -0.0001404924,
  0, -1.264521e-06, -1.000434e-07, 0.007340891, 0.01568922, 0, -0.0001261217, 
    0, 0.001482579, 0.00779035, 0.000273419, 0.002130997, 0.01021552, 
    0.01025633, 0.02063055, 0.02651582, 0.007255356, 0.005337832, 
    0.008620854, 0.0005081282, -0.0001190505, 0.02577072, 0.01577883, 
    0.012994, 0.02707504, 0.02919151, 0.001009678, -2.893043e-06, 
    -0.0002218104,
  0, 0.0007588434, -1.130499e-07, 0.002002589, 0.00134472, 0, 0, 0, 0, 0, 0, 
    0.01562452, 0.01976954, 0.02548322, 0.01718672, 0.02088472, 0.02067134, 
    0.02476834, 0.009633041, 0, 0, -4.191184e-05, 0.00109474, 0.02769278, 
    0.04892277, 0.02632773, 0.03777657, 0.003006133, 0.0002466378,
  -1.060931e-05, 0, -1.705601e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0004928769, 
    0.01354054, 0.008795573, 0.004170736, 0.000980375, 0.005743729, 
    0.0078297, -1.284363e-05, -5.898054e-09, 0, 0, -3.513795e-05, 0.01143378, 
    0.006311843, 0.007389747, 0.0007755866, 0.003319258,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6.627972e-06, 0, 0, 0, 
    -1.236083e-05, 0, 0.0008196677, 0, 0, 0, 0, 0.003469146, -8.951566e-06, 
    -4.58482e-05, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, -3.47465e-06, -1.335541e-05, -3.9372e-06, 0, 0, 0, 0, 0, 
    0, 0.000971713, 0, 0, 0, 0, 0, 0, -3.277353e-05, -2.784391e-06, 0, 0, 0, 
    0.002361737, 1.849301e-05,
  0.0009337123, 0.001579389, -1.708208e-06, 0, -1.381574e-06, 0.0002463756, 
    0.01233674, -0.0001468978, -5.713543e-08, 0.002775195, -3.660949e-05, 
    9.676614e-05, -2.619307e-10, 0.0005101973, 0.008475699, 0.002808361, 0, 
    0.003031448, 0.001141675, 0.002130747, 0.0009518105, -5.414452e-05, 
    0.004231491, 0.003047485, 6.148566e-05, 0.006649566, 0.01409959, 
    0.01170564, 0.005440996,
  0.008511612, 0.001885332, 5.498078e-06, 0.01484824, 0.05583433, 0.04071526, 
    0.01828319, 0.01037807, 7.100915e-05, -2.899397e-07, 0.001284602, 
    0.00229093, -7.086302e-05, 0.02881422, 0.01897629, 0.00641206, 
    -0.0003283648, 0.02506772, 0.05770744, 0.01505416, 0.003939659, 
    0.001491863, 0.0002302576, 3.453505e-05, 0.0214966, 0.05608162, 
    0.02620514, 0.01244136, 0.01310368,
  0.000547113, 1.055269e-05, 0.003043428, 0.1731537, 0.06045713, 0.01410192, 
    0.009735546, 0.002019219, 0.01717728, 0.0177875, 0.009818497, 
    4.451307e-06, 0.008041875, 0.01057388, 0.02212777, 0.0003004558, 
    0.06165625, 0.03429075, 0.111978, 0.04714852, 0.01999164, 0.002164744, 
    0.0003110968, 0.0004729622, 0.05031824, 0.07914028, 0.09386116, 
    0.05303772, 0.02031064,
  0.0003324918, 0.0307795, 0.05994547, 0.07334867, 0.02056975, 0.007590095, 
    0.0005566417, 0.03613533, 0.005380071, 0.02397018, 0.004917935, 
    -7.314481e-05, 0.005023948, 0.09649983, 0.02975656, 0.02538371, 
    0.1713408, 0.2786905, 0.1959624, 0.04237043, 0.03281733, 0.002665052, 
    4.645422e-08, 0.02666583, 0.1324997, 0.1486437, 0.1265198, 0.05051101, 
    0.005405762,
  0.001809348, 0.2385228, 0.1940213, 0.1552051, 0.1402685, 0.093853, 
    0.0546018, 0.07160358, 0.0187841, 0.005487701, 0.03372842, 0.03681706, 
    0.1230981, 0.1898709, 0.132179, 0.2019391, 0.1176386, 0.003277213, 
    0.0005952652, 1.461071e-06, 3.242991e-07, 6.513039e-07, 0.006958769, 
    0.3008218, 0.3532405, 0.2998261, 0.1069173, 0.0731338, 0.0003983085,
  0.01791914, 0.3836679, 0.4877965, 0.02585453, 0.06305045, 0.02841317, 
    0.04119355, 0.03826446, 0.2919722, 0.2988757, 0.1774015, 0.156425, 
    0.2040485, 0.07252486, 0.001011686, 0.00537825, 0.0001288911, 0.00416389, 
    9.695663e-05, 0.01683794, 0.003091141, 3.651899e-07, 0.03372313, 
    0.4078711, 0.2737241, 0.02650088, 0.1326301, 0.02301525, 9.21072e-06,
  0.01226048, 0.00882713, 0.04730554, 0.004791712, 0.06394621, 0.03677694, 
    0.009372196, 0.07623743, 0.07649457, 0.1529208, 0.1605259, 0.217065, 
    0.2044539, 0.2105427, 0.1172717, 0.1396037, 0.1292061, 0.1399453, 
    0.03931483, 0.1084529, 0.0716425, 0.05989055, 0.09975193, 0.1609113, 
    0.1262072, 0.07878752, 0.06895576, 0.1349968, 0.0263889,
  0.03825092, -0.0001479452, 0.001217075, 0.02216314, 0.03761204, 0.050254, 
    0.008328185, 0.04465886, 0.01068052, 0.02791273, 0.1215049, 0.04532043, 
    0.02496896, 0.1053237, 0.09427361, 0.1198898, 0.09864737, 0.1045751, 
    0.1143085, 0.03289313, 0.0565262, 0.06289126, 0.02986092, 0.122123, 
    0.06120778, 0.09226627, 0.02523351, 0.05278289, 0.03148573,
  -5.341174e-06, -1.469738e-05, 5.140867e-06, 0.01131088, 0.02443876, 
    1.066415e-05, 0.0002860814, -1.663197e-05, 0.004283048, 0.01258014, 
    0.0001761034, 0.01123861, 0.04122265, 0.0358839, 0.05861348, 0.04490551, 
    0.04236407, 0.07592244, 0.02445398, 0.01117678, 0.006756907, 0.0767298, 
    0.04366603, 0.03250943, 0.1235001, 0.09556768, 0.01867723, -5.830704e-06, 
    -0.0006649783,
  7.269002e-05, 0.003697064, -8.439732e-05, 0.00605127, 0.004778884, 0, 0, 0, 
    0, 0, 2.238068e-05, 0.04321833, 0.03508825, 0.05599169, 0.03693585, 
    0.0570519, 0.03911742, 0.05228537, 0.04017353, 5.37721e-05, 0, 
    0.0001449372, 0.003805168, 0.05824246, 0.0756935, 0.0508674, 0.09036588, 
    0.02053452, 0.00434779,
  0.008005774, 1.08084e-05, 0.000266777, 0.001128474, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0009171981, 0.01555945, 0.01454195, 0.0154277, 0.006816434, 
    0.009019735, 0.02005767, 0.002168663, 0.0004168823, -2.030264e-06, 
    -8.974315e-05, 0.001284624, 0.01957362, 0.01737517, 0.01702876, 
    0.006938831, 0.02030476,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.056087e-06, -8.018456e-08, 
    0.0005129931, 0, 0, 0.001123637, -1.289273e-05, 0.002687122, 
    -5.714482e-05, 0, 0, 0, 0.007062329, 0.0009214929, 0.002551033, 
    -1.645255e-05,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  -1.175625e-05, -2.3476e-06, 0, -2.732541e-06, 0, 0, -1.365897e-05, 
    0.002115103, 0.0002435755, 0, 2.055118e-16, 0, 0, -3.066528e-06, 0, 
    0.001902851, 0.004132765, 0, 0, 0, 0, -1.802372e-05, 0.002752126, 
    -3.513843e-06, 0, -1.04418e-05, 0, 0.004305325, 0.0003279301,
  0.006870858, 0.004929577, 0.003080152, 0.001976364, 0.002121908, 
    0.003724144, 0.01731463, 0.01174909, 0.006229713, 0.0118142, 0.004513261, 
    0.0005034528, -1.465765e-05, 0.003869578, 0.01273216, 0.01100557, 
    9.483349e-06, 0.00453576, 0.006419457, 0.007330477, 0.007182417, 
    0.001561236, 0.01922236, 0.005848145, -6.040098e-06, 0.01102814, 
    0.02573694, 0.03195352, 0.01150799,
  0.03728846, 0.02321468, 0.04708084, 0.07753804, 0.1123658, 0.08891765, 
    0.08035519, 0.07853381, 0.04701509, 0.04270032, 0.0507653, 0.03204484, 
    0.01160024, 0.04602771, 0.03944842, 0.04590052, 0.0107613, 0.04337101, 
    0.1069749, 0.06048033, 0.05468055, 0.02157575, 0.03467459, 0.002518445, 
    0.03019453, 0.1131427, 0.06364801, 0.09357031, 0.04882362,
  0.05840775, 0.005369095, 0.0407311, 0.1810579, 0.09323951, 0.08623373, 
    0.03240002, 0.05965858, 0.04314677, 0.02306282, 0.06042907, 0.01186908, 
    0.01875165, 0.03196071, 0.06433152, 0.04108445, 0.1049777, 0.06133074, 
    0.183629, 0.1446775, 0.1205046, 0.07715248, 0.0250807, 0.01781387, 
    0.0623391, 0.08310195, 0.1812958, 0.1611221, 0.1131606,
  0.003448932, 0.0295247, 0.06579242, 0.05449722, 0.01529191, 0.002686637, 
    0.0003178881, 0.02548763, 0.0001627659, 0.005086443, 0.005450435, 
    -3.968877e-05, 0.006617574, 0.1144378, 0.05533674, 0.02660893, 0.152693, 
    0.2698331, 0.1885647, 0.03774215, 0.03683225, 0.001453148, -4.810525e-09, 
    0.01793209, 0.08661576, 0.14356, 0.1430712, 0.08681971, 0.001418618,
  0.002669894, 0.1733512, 0.138523, 0.1325339, 0.1155461, 0.071748, 
    0.04544434, 0.05854835, 0.01236282, 0.003464457, 0.01587046, 0.03362888, 
    0.07997887, 0.149337, 0.1221931, 0.16101, 0.09121788, 0.001207641, 
    1.258008e-05, 3.750048e-07, 4.043346e-07, 6.743984e-07, 0.002043182, 
    0.2823807, 0.2951477, 0.2655149, 0.08715806, 0.05356241, -1.141317e-06,
  0.01547695, 0.3483624, 0.3732401, 0.02106159, 0.0416072, 0.01744167, 
    0.02837868, 0.02383246, 0.236982, 0.2256426, 0.126807, 0.1062857, 
    0.1516412, 0.04330144, 0.000369298, 0.0004149171, 0.000146572, 
    8.299355e-05, -5.413587e-05, 0.002440749, 0.00126392, -4.32566e-05, 
    0.03060469, 0.3036744, 0.2261074, 0.03540152, 0.09765181, 0.01585328, 
    6.945122e-06,
  0.004911098, 2.280317e-05, 0.0373595, 0.0470644, 0.04132321, 0.02703724, 
    0.004490189, 0.05413807, 0.06133074, 0.1107432, 0.1292281, 0.1709971, 
    0.1873251, 0.1805044, 0.07987929, 0.1204818, 0.1308015, 0.09988014, 
    0.03100696, 0.08974284, 0.06367894, 0.02924667, 0.06781062, 0.1117678, 
    0.113895, 0.07735036, 0.03864409, 0.1022584, 0.0249371,
  0.09453663, 0.002242996, 0.001344254, 0.009406778, 0.05501613, 0.04722015, 
    0.0278138, 0.04104434, 0.01308578, 0.02305132, 0.1055622, 0.04084048, 
    0.0201671, 0.1028973, 0.08973379, 0.08700204, 0.08226559, 0.07664239, 
    0.09968368, 0.02935713, 0.03765453, 0.05663804, 0.02272925, 0.1124129, 
    0.05382121, 0.08263801, 0.1162216, 0.1435351, 0.2679816,
  0.0414147, 0.03472803, 0.07241975, 0.03089282, 0.04606179, 0.02446642, 
    0.09658296, -6.838945e-05, 0.01442488, 0.03684719, 0.02585745, 
    0.02820216, 0.04293737, 0.04671568, 0.1135876, 0.159531, 0.08119157, 
    0.1244339, 0.1145504, 0.07710586, 0.02724306, 0.1427586, 0.102898, 
    0.07285701, 0.2132226, 0.168883, 0.1146808, 0.03207893, 0.012048,
  0.0008412028, 0.008272881, 0.001494967, 0.01160406, 0.008264279, 
    -2.238834e-05, -1.899879e-05, -1.246117e-06, 1.608656e-06, -4.321228e-07, 
    0.004931862, 0.05401313, 0.04944022, 0.08273928, 0.07729874, 0.1051763, 
    0.1237418, 0.13963, 0.1203743, 0.004260708, -6.420361e-12, 0.0007396783, 
    0.009642424, 0.09912504, 0.1133787, 0.1021223, 0.1705648, 0.08241028, 
    0.0274777,
  0.02621275, 0.004205208, 0.005865517, 0.001986528, -6.953619e-06, 
    -4.128701e-07, 0, -3.07193e-06, 0, 0, 0, 0, 0.005618033, 0.02156112, 
    0.02594685, 0.03530132, 0.03021534, 0.03012457, 0.0652658, 0.01361281, 
    0.004019985, 0.0001144938, 0.00457065, 0.007619814, 0.03717327, 
    0.03339788, 0.02986541, 0.02230744, 0.06365622,
  -0.0001285653, 0, 0.001843411, 0, -5.038997e-05, 0, 0, 0, 0, 0, 0, 0, 0, 
    -4.180584e-06, 0.00126197, 0.00284763, -0.0001470307, 0.0008896702, 
    0.003391216, -4.699394e-05, 0.002215659, -0.0002017645, 0, 4.136826e-05, 
    0.0001445243, 0.01185049, 0.009971753, 0.004620789, 0.0008314641,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0001754747, -1.580943e-05, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, -3.085784e-06, -4.347651e-06, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  -3.526874e-05, -4.810633e-05, 0, -8.667537e-05, -7.051001e-05, 
    2.466891e-06, -1.140926e-05, 0.01381577, 0.0210615, 0.01162161, 
    0.0001736338, 7.495387e-09, 0, 0.001511777, 0.01075957, 0.01051156, 
    0.01373732, 0.0002498174, 0.0004161781, -3.531009e-05, 2.905556e-09, 
    0.0001006375, 0.003331088, 0.003093089, 4.591438e-05, 9.241178e-05, 
    -2.673377e-05, 0.005995864, 0.003616532,
  0.03938416, 0.02312445, 0.009249701, 0.03168991, 0.02547195, 0.02987745, 
    0.05260944, 0.06924225, 0.08097276, 0.0746044, 0.05359736, 0.02996968, 
    0.02390172, 0.05428242, 0.03363496, 0.08648131, 0.03832271, 0.03555495, 
    0.06675917, 0.09617671, 0.07322044, 0.02635419, 0.05120966, 0.01613362, 
    0.02208641, 0.09438, 0.1452663, 0.1255189, 0.07244946,
  0.09030972, 0.06295499, 0.07048011, 0.1013884, 0.1375364, 0.1268482, 
    0.1506887, 0.1832568, 0.1322517, 0.1121932, 0.1176447, 0.1132856, 
    0.0326667, 0.08676706, 0.108231, 0.1273734, 0.1231619, 0.08256033, 
    0.1697185, 0.1230134, 0.1490185, 0.1516524, 0.1008985, 0.03681692, 
    0.1016437, 0.1408524, 0.09185316, 0.09165642, 0.08149515,
  0.04126621, 0.0006539692, 0.06524274, 0.1607345, 0.09333928, 0.06461005, 
    0.02285402, 0.04323747, 0.02953316, 0.01051935, 0.05173919, 0.008452525, 
    0.02808145, 0.01512857, 0.09396869, 0.0444667, 0.1076878, 0.09458864, 
    0.1788258, 0.134291, 0.1489888, 0.09042667, 0.01780571, 0.01014956, 
    0.0929132, 0.08269749, 0.1848058, 0.1298723, 0.07854087,
  -1.346066e-05, 0.0252104, 0.04246886, 0.0177494, 0.009518898, 
    -8.610565e-06, 0.002143137, 0.02999377, 3.590891e-06, 0.000616221, 
    0.005638701, -4.385424e-06, 0.0167311, 0.1518375, 0.06287213, 0.03592634, 
    0.1342557, 0.2337024, 0.1762306, 0.03091497, 0.04097401, 0.001398061, 
    -8.079298e-07, 0.01420004, 0.06531651, 0.1507912, 0.1335532, 0.08267086, 
    -2.638819e-05,
  0.001587284, 0.1484261, 0.08508274, 0.132896, 0.09147974, 0.06433112, 
    0.04835996, 0.04053552, 0.01422902, 0.001050907, 0.01054765, 0.03667525, 
    0.06070541, 0.1362084, 0.1124323, 0.1342677, 0.08315396, 0.0003701804, 
    2.273397e-05, 1.617928e-07, 9.69875e-08, 3.785498e-07, 0.0003615658, 
    0.2439396, 0.270875, 0.2468775, 0.08357092, 0.040266, 4.310711e-07,
  0.01637326, 0.3117107, 0.2958718, 0.01870368, 0.04300089, 0.01403684, 
    0.02242377, 0.02390149, 0.1920476, 0.1553807, 0.09901903, 0.08793375, 
    0.1320263, 0.0191058, 0.0003395093, 0.00072581, 5.086243e-05, 
    -0.0001688704, -1.102001e-07, 1.858969e-06, -0.0001200946, -1.72547e-06, 
    0.02778791, 0.2377794, 0.1888269, 0.054302, 0.1031604, 0.01414734, 
    0.000297502,
  0.004210352, -2.362788e-05, 0.03119612, 0.02519925, 0.02053751, 0.01517954, 
    0.003793472, 0.06129721, 0.05784003, 0.0846509, 0.1172071, 0.1452815, 
    0.1750752, 0.165949, 0.06874842, 0.09536363, 0.1324111, 0.1004464, 
    0.03253356, 0.08392549, 0.06083252, 0.0207777, 0.05228101, 0.09957951, 
    0.1012404, 0.08262128, 0.02959337, 0.08766518, 0.02931987,
  0.06895397, 0.0002049826, 0.0002985731, 0.005131995, 0.04965984, 
    0.05288864, 0.03424935, 0.04120086, 0.0201837, 0.01878479, 0.09667657, 
    0.03565551, 0.01839162, 0.1028206, 0.08255461, 0.06921967, 0.075386, 
    0.0678346, 0.0669831, 0.008937312, 0.03111935, 0.03191066, 0.02224313, 
    0.1096757, 0.04674186, 0.07343164, 0.1041629, 0.1248145, 0.2373754,
  0.04470244, 0.05889222, 0.1077847, 0.1343289, 0.1212086, 0.09728184, 
    0.1533797, 0.0004948113, 0.02299352, 0.07327154, 0.03691113, 0.04392751, 
    0.03429617, 0.03977009, 0.1070436, 0.1192323, 0.07330025, 0.09947474, 
    0.1215416, 0.07662016, 0.07958917, 0.1428442, 0.09168639, 0.06530491, 
    0.1429125, 0.1454173, 0.1127409, 0.03287887, 0.02724925,
  0.08310273, 0.09120432, 0.07519444, 0.03087654, 0.0774316, 0.04026401, 
    2.243082e-05, -9.033419e-06, 2.586886e-05, -7.881597e-05, 0.01961591, 
    0.1016436, 0.07353129, 0.163446, 0.1668984, 0.1950272, 0.2087442, 
    0.2236892, 0.1563033, 0.04247506, -2.245658e-05, 0.01359241, 0.09919003, 
    0.1611761, 0.1281269, 0.1788509, 0.2322929, 0.1587385, 0.08254452,
  0.09650803, 0.01700683, 0.02557494, 0.003022601, 0.00979393, 0.01079562, 
    0.002439815, -3.282642e-05, 0, 0, 0, 0, 0.007827047, 0.02584014, 
    0.03139232, 0.03772428, 0.08729131, 0.0937221, 0.2244554, 0.03447158, 
    0.01871267, 0.01175056, 0.01041348, 0.02085795, 0.082222, 0.06534164, 
    0.07335375, 0.08007651, 0.1269122,
  0.01510566, -0.0001413919, 0.002358494, -5.165745e-06, -0.0003279835, 
    0.003591891, 0, 5.872782e-05, 0, 0, 0, 0, 0, -2.395262e-05, 0.007708594, 
    0.008097909, 0.001365852, 0.003444593, 0.01209085, 0.002329827, 
    0.004505525, -0.0004549477, -5.220421e-09, 0.01178202, 0.003822202, 
    0.02647957, 0.02860838, 0.0110771, 0.005149638,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.006332856, 0.0002735714, -5.83845e-07, 0.0003703115, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  -0.00017978, -0.000204056, 0.003316446, 0, 0, 0, 0, -4.100167e-05, 
    -8.17496e-05, -6.220874e-09, 0, 0, 0, 0, -0.0002656059, -0.0004784028, 
    -7.874722e-05, -4.414643e-05, -1.915694e-05, -1.024669e-06, 0, 
    -5.19909e-06, 0, -4.938303e-06, 0, -1.142462e-05, 0.0003229301, 
    0.002191882, 0.002305656,
  0.02543387, 0.0126509, 0.003764756, 0.00179969, 0.005256293, 0.01254279, 
    0.008110463, 0.04400955, 0.05100789, 0.04807, 0.03339845, 0.01194902, 
    0.0127452, 0.03450217, 0.07741268, 0.06560323, 0.08301956, 0.04698677, 
    0.04055136, 0.02810447, 0.05342754, 0.0915067, 0.08851985, 0.06898649, 
    0.04590793, 0.04945337, 0.05433793, 0.05575642, 0.03656079,
  0.08845105, 0.09765305, 0.08092285, 0.09454028, 0.07722189, 0.09905886, 
    0.1469489, 0.1248732, 0.1037531, 0.1073009, 0.1158283, 0.1009914, 
    0.07124888, 0.1094887, 0.07740249, 0.152588, 0.1031417, 0.1710585, 
    0.1582303, 0.2042408, 0.1455455, 0.131368, 0.129961, 0.05804141, 
    0.07054365, 0.1498518, 0.229571, 0.1697455, 0.1137362,
  0.09910221, 0.06364413, 0.04383876, 0.08983539, 0.1121164, 0.1143912, 
    0.132358, 0.1691004, 0.1481247, 0.1242579, 0.09778231, 0.1269798, 
    0.05951482, 0.1015297, 0.1040038, 0.1584613, 0.1544297, 0.1033488, 
    0.164461, 0.1440495, 0.1792555, 0.1800616, 0.1055293, 0.06011447, 
    0.1092912, 0.1505253, 0.09983422, 0.08011649, 0.09171313,
  0.0200491, 0.0002746021, 0.04816313, 0.1551419, 0.08041468, 0.06041989, 
    0.01336198, 0.02666268, 0.02025204, 0.001156715, 0.05119724, 0.009295767, 
    0.02002615, 0.01368859, 0.09724849, 0.03637071, 0.1055261, 0.09511222, 
    0.155153, 0.1073135, 0.1237339, 0.0735494, 0.01503386, 0.006546053, 
    0.1004887, 0.07916686, 0.1591882, 0.1128666, 0.0578731,
  7.455552e-06, 0.0226574, 0.04102341, 0.01092477, 0.006512451, 2.860054e-06, 
    -2.309007e-05, 0.04691749, -6.125978e-06, 8.343228e-06, 0.005204483, 
    0.0003538285, 0.009785354, 0.1535594, 0.07447983, 0.04794616, 0.115329, 
    0.1896736, 0.1566294, 0.01872291, 0.0528605, -1.557359e-05, 3.760551e-08, 
    0.006877783, 0.0486467, 0.1453292, 0.1339963, 0.06916983, 1.33052e-05,
  0.0002565182, 0.1487178, 0.06068811, 0.1312792, 0.06194771, 0.06888793, 
    0.04182762, 0.01749067, 0.01713551, 0.001178316, 0.004971015, 0.04051698, 
    0.04871754, 0.1225562, 0.12177, 0.1113385, 0.07580242, 0.0006052587, 
    9.997416e-07, 1.998214e-08, -5.244776e-10, 4.504947e-08, 0.0009300562, 
    0.1899079, 0.2286211, 0.1931694, 0.07934137, 0.01967652, 1.103391e-07,
  0.01675591, 0.2669134, 0.2206542, 0.01554195, 0.05302477, 0.008015459, 
    0.01126346, 0.01851934, 0.1372337, 0.09732608, 0.06578602, 0.07755823, 
    0.1007744, 0.01288092, 0.002356447, 0.0010377, -5.553632e-07, 
    -6.458002e-05, 6.717772e-07, 3.456621e-06, -0.0002663218, 7.180477e-07, 
    0.006255381, 0.1720318, 0.1455483, 0.06308142, 0.1099722, 0.009319381, 
    5.6662e-05,
  0.002424622, 3.479415e-05, 0.01625868, 0.01287077, 0.02824406, 0.007823032, 
    0.008505782, 0.06086633, 0.05791375, 0.05287473, 0.09699241, 0.1200048, 
    0.1523865, 0.1461302, 0.05858222, 0.07534565, 0.1350837, 0.08819638, 
    0.03387595, 0.0777643, 0.06814494, 0.01369122, 0.04403344, 0.08245888, 
    0.08669117, 0.08301172, 0.02173937, 0.07659961, 0.0319899,
  0.05169459, 8.692248e-05, -3.770394e-05, 0.00196955, 0.03852547, 
    0.03052442, 0.02190237, 0.04470434, 0.02278274, 0.0149113, 0.09067529, 
    0.02996228, 0.01777544, 0.09964243, 0.06794816, 0.04643926, 0.07311287, 
    0.05642724, 0.05021417, 0.0008556088, 0.02994952, 0.01829896, 0.01869412, 
    0.1163201, 0.04344365, 0.0686096, 0.08420619, 0.09448767, 0.1939282,
  0.02815626, 0.05847146, 0.09365695, 0.1233796, 0.1613656, 0.1022738, 
    0.1425646, 0.002540492, 0.03517762, 0.08130534, 0.01472737, 0.05659572, 
    0.02862764, 0.04824705, 0.09970533, 0.07826895, 0.06339485, 0.09534919, 
    0.1195042, 0.05924239, 0.1118284, 0.1117387, 0.07755315, 0.07659932, 
    0.09359949, 0.1323327, 0.08528253, 0.02872156, 0.02697029,
  0.09546658, 0.1206378, 0.1099384, 0.1192247, 0.09615169, 0.09914594, 
    0.0009052432, 0.03509708, 0.01515415, 0.02165312, 0.1013836, 0.200593, 
    0.1566496, 0.2151272, 0.2059446, 0.1892513, 0.213207, 0.2061485, 
    0.1611285, 0.0808023, 0.00490963, 0.04941713, 0.1443698, 0.1741686, 
    0.1676229, 0.1701931, 0.2251079, 0.1612698, 0.09687844,
  0.1657574, 0.1514759, 0.1624863, 0.1619707, 0.187592, 0.1079693, 
    0.04612542, 4.856292e-05, 9.234172e-05, -2.375953e-06, -1.047137e-05, 
    -3.248151e-05, 0.02527616, 0.03937786, 0.06193236, 0.07370424, 0.1605891, 
    0.139221, 0.2818021, 0.08779085, 0.0337272, 0.07141848, 0.05206405, 
    0.05517117, 0.1438359, 0.1207119, 0.1167065, 0.1269827, 0.2052712,
  0.02987423, 0.01777745, 0.01975124, 0.008172342, 0.02719544, 0.01882317, 
    0.01244727, 0.009838602, -6.264239e-06, 0, 0, 0, 0, 0.009392839, 
    0.01950301, 0.01234725, 0.01659293, 0.01387592, 0.01868502, 0.02217793, 
    0.01316968, 0.01067926, 0.0006655034, 0.02853743, 0.07658342, 0.07768109, 
    0.07805014, 0.04459526, 0.02883013,
  0.0002298686, 0, 6.714185e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, -7.88148e-07, 0.01057211, 0.006221407, -4.630969e-05, 
    0.01155544, -0.0001441075,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -1.17589e-05, -1.463445e-05, 0, 0,
  0.01156008, 0.02236223, 0.01918714, 0.004312627, -8.211828e-06, 0, 
    0.01041648, 1.249364e-05, 2.69288e-05, -2.798919e-06, 0, -3.257227e-06, 
    -0.0002348545, 0.009570437, 0.01397278, 0.03494149, 0.0446514, 
    0.05091717, 0.02993839, 0.02454761, 0.004770984, -2.858006e-05, 
    -3.114e-06, 0.004281865, 0.02287496, 0.03723583, 0.01979156, 0.03199981, 
    0.0276974,
  0.1337862, 0.1078099, 0.0941682, 0.0917474, 0.03746254, 0.06964337, 
    0.1191565, 0.08374178, 0.06382969, 0.09130887, 0.08074977, 0.05471414, 
    0.08358052, 0.0958157, 0.1662853, 0.1975143, 0.1723929, 0.1785313, 
    0.1365934, 0.1605266, 0.1224183, 0.1319932, 0.1323295, 0.1537063, 
    0.1975483, 0.1545403, 0.1489512, 0.1561077, 0.1442521,
  0.1143011, 0.1021147, 0.1210548, 0.140877, 0.1287847, 0.1559653, 0.2195547, 
    0.193637, 0.1332391, 0.11421, 0.1211775, 0.1408883, 0.1097245, 0.1480746, 
    0.1254842, 0.1688387, 0.1124894, 0.1479485, 0.164484, 0.1830068, 
    0.1598746, 0.135673, 0.1615906, 0.0845783, 0.07077026, 0.1664447, 
    0.1968487, 0.1652061, 0.1292184,
  0.1194626, 0.07605439, 0.03483119, 0.07215478, 0.09231949, 0.1037256, 
    0.1207902, 0.1501049, 0.1276107, 0.1090949, 0.0858927, 0.1076323, 
    0.05423564, 0.1214687, 0.1005745, 0.1343256, 0.1446514, 0.1098996, 
    0.1342333, 0.1351383, 0.1676217, 0.1854254, 0.1036731, 0.06469338, 
    0.09407522, 0.1443908, 0.09758316, 0.06977172, 0.08900717,
  0.005229584, 0.0003130773, 0.04713175, 0.1719887, 0.07888526, 0.04626743, 
    0.007577785, 0.02031737, 0.0194824, -2.531723e-06, 0.05341483, 
    0.01336297, 0.01687175, 0.01846668, 0.1017279, 0.03273201, 0.09035948, 
    0.09301662, 0.1276184, 0.09699591, 0.1427408, 0.04708992, 0.008711482, 
    0.001184401, 0.09592824, 0.07354862, 0.151985, 0.1002967, 0.02409262,
  7.122046e-06, 0.01836395, 0.0374028, 0.006551865, 0.004507159, 
    1.120503e-06, -0.000272028, 0.02961221, -4.759752e-06, -0.0001720372, 
    0.004444381, 0.0003158836, 0.01232733, 0.1671051, 0.0817422, 0.05230834, 
    0.1109052, 0.1338076, 0.1409814, 0.01152787, 0.04339293, -1.185092e-05, 
    1.118153e-09, 0.0007653552, 0.03126291, 0.1521372, 0.1236415, 0.05058407, 
    8.864135e-06,
  3.396048e-06, 0.1285803, 0.04837088, 0.1257063, 0.04534243, 0.07078391, 
    0.02787411, 0.00647119, 0.02077796, 0.0008646058, 0.008146198, 
    0.03507775, 0.03901128, 0.1069713, 0.09421255, 0.1053523, 0.07669845, 
    0.0008366731, 1.091326e-06, 2.43783e-08, 0, 1.148091e-08, 0.0004509676, 
    0.1501966, 0.184265, 0.1287872, 0.06585435, 0.008740127, 8.98717e-08,
  0.0220579, 0.2533486, 0.1720464, 0.01498376, 0.05010597, 0.005930227, 
    0.006414072, 0.0134239, 0.1008157, 0.06645195, 0.03614196, 0.06587891, 
    0.07182689, 0.013209, 0.004748911, 0.001053463, -2.807505e-06, 
    0.006641622, 3.913471e-07, 1.57879e-07, -0.0001697964, 2.924627e-06, 
    7.74423e-05, 0.1309941, 0.09425115, 0.06190443, 0.1324494, 0.01907878, 
    2.177319e-05,
  0.000727018, 0.000280151, 0.006969154, 0.01263603, 0.03868899, 0.005412353, 
    0.0235967, 0.05758753, 0.05394009, 0.02990623, 0.06813413, 0.1085703, 
    0.1287034, 0.1161956, 0.04590115, 0.07064262, 0.1301284, 0.08390933, 
    0.03676622, 0.06273314, 0.0653012, 0.008620146, 0.04027508, 0.06791372, 
    0.06536283, 0.08732823, 0.01561139, 0.06175152, 0.02689336,
  0.0163457, 0.003332158, -3.983729e-05, 0.001943046, 0.03314749, 0.0111123, 
    0.01351194, 0.03981144, 0.01601297, 0.01038669, 0.07418732, 0.01523206, 
    0.01764873, 0.09891069, 0.04767702, 0.02422768, 0.06639583, 0.04135987, 
    0.01692021, 0.005198318, 0.03112204, 0.01683101, 0.01192489, 0.1150421, 
    0.03769754, 0.06966287, 0.08406383, 0.06350588, 0.1385011,
  0.0236029, 0.06673758, 0.06399649, 0.08909401, 0.1546383, 0.09830259, 
    0.1228239, 0.007071834, 0.06018695, 0.07802982, 0.01465294, 0.03638138, 
    0.01858682, 0.03017544, 0.06823243, 0.05760905, 0.06422563, 0.09451865, 
    0.09330444, 0.02854785, 0.08628157, 0.09337828, 0.0716019, 0.07582323, 
    0.06972317, 0.1193091, 0.0699113, 0.01727915, 0.02534158,
  0.09155575, 0.1301268, 0.09090858, 0.153778, 0.07412881, 0.100604, 
    0.006137389, 0.08248591, 0.03069924, 0.05408125, 0.1569346, 0.1987548, 
    0.216834, 0.2264153, 0.2107455, 0.1763358, 0.2068592, 0.2211744, 
    0.2125146, 0.1020498, 0.01945205, 0.03983613, 0.1248686, 0.1601043, 
    0.1751177, 0.1605691, 0.2050968, 0.1399413, 0.1082551,
  0.203894, 0.2158332, 0.2507496, 0.2370652, 0.2332261, 0.2363753, 0.1540614, 
    0.002989264, 0.001127939, 0.004127227, 0.007112542, 0.002937696, 
    0.04132483, 0.08835234, 0.09088627, 0.1035183, 0.1646867, 0.1870941, 
    0.3156216, 0.1783297, 0.05827343, 0.1291109, 0.109361, 0.1310782, 
    0.1651519, 0.1426831, 0.1104963, 0.129754, 0.2225207,
  0.1468914, 0.08522789, 0.07798856, 0.0846599, 0.1395499, 0.1837588, 
    0.1074368, 0.0918185, 0.02814003, -3.103333e-05, 0, 0, -0.0002380084, 
    0.0427393, 0.04176123, 0.01915984, 0.02707155, 0.02021413, 0.06291053, 
    0.1211433, 0.07855008, 0.04614992, 0.007358751, 0.09520403, 0.1356041, 
    0.1236775, 0.1840212, 0.07213596, 0.09624884,
  0.009908199, 1.9161e-05, 0.0001074874, 0.0009573026, 0.03216712, 
    0.03710885, 0.01664493, -2.287581e-07, 0, 0, 0, 0, 0, 0, -2.440381e-05, 
    0.0001063161, 0.001056598, 0.007530954, 0.006967816, 0.001919645, 
    0.0102822, 0.004676544, -0.00110078, -0.003539287, 0.03398779, 
    0.01925153, -0.0002584474, 0.03560962, 0.02034982,
  0, 0, -4.234663e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5.497586e-06, 4.076722e-05, 
    0.0004117214, 0.02170673, 0.008798834, 0.0002548091, 0, 0, 0, 0, 
    0.03905908, 7.918218e-05, -0.0007119414, -0.001011041, 0, 0,
  0.03764333, 0.04634277, 0.05049202, 0.04596369, -0.001030141, -0.001649905, 
    0.07578607, -0.0002151128, -0.0002081937, -0.0002661711, 2.4934e-05, 
    0.0001578671, -0.003225184, 0.035858, 0.04097785, 0.08271537, 0.09556142, 
    0.1120871, 0.09461912, 0.05415532, 0.04068347, 0.03703814, 0.04114874, 
    0.04842562, 0.08841789, 0.08421687, 0.1351351, 0.07001803, 0.04996168,
  0.1806255, 0.1456479, 0.144738, 0.1230503, 0.1038066, 0.1467233, 0.2484502, 
    0.1857118, 0.1354548, 0.1485356, 0.1465028, 0.1071409, 0.1701044, 
    0.1482071, 0.218746, 0.1880754, 0.2051378, 0.2311478, 0.1900885, 
    0.1748082, 0.1680821, 0.1965075, 0.2220667, 0.2096953, 0.2405663, 
    0.1884332, 0.1663047, 0.1840672, 0.2237224,
  0.1216774, 0.1136813, 0.1274264, 0.1701108, 0.1621283, 0.162298, 0.2371236, 
    0.1994997, 0.1569282, 0.1241568, 0.1310792, 0.1545258, 0.1269233, 
    0.1503915, 0.1463246, 0.172174, 0.117044, 0.1449315, 0.1344973, 
    0.1728247, 0.1656312, 0.1573841, 0.1629181, 0.08871237, 0.07693448, 
    0.136445, 0.178635, 0.1412252, 0.1334178,
  0.1074291, 0.07103572, 0.02880109, 0.05024811, 0.08398969, 0.08479589, 
    0.1233629, 0.1433435, 0.1166854, 0.0875949, 0.08125964, 0.0860124, 
    0.05056692, 0.1288258, 0.09861552, 0.1196568, 0.1206907, 0.1037656, 
    0.1112471, 0.124122, 0.168394, 0.1794413, 0.06980827, 0.05058544, 
    0.07661923, 0.1540349, 0.09010407, 0.05560832, 0.08569105,
  0.0005865246, 0.0008909264, 0.05007576, 0.1972249, 0.06944048, 0.03887875, 
    0.008065241, 0.01466267, 0.02215618, 4.979533e-05, 0.06262282, 
    0.01571098, 0.0169235, 0.02416313, 0.1039521, 0.03569232, 0.07700876, 
    0.0851753, 0.1085042, 0.07800139, 0.131829, 0.02419372, 0.001089138, 
    -3.711895e-05, 0.0843283, 0.06985659, 0.1060692, 0.07971784, 0.01533056,
  4.001442e-06, 0.01399085, 0.03284395, 0.005340176, 0.001603535, 
    2.906867e-07, -0.0002529004, 0.02487038, -3.968135e-07, 0.0005812792, 
    0.003947451, 0.0003016572, 0.009234241, 0.1902012, 0.08455152, 
    0.05306837, 0.1098363, 0.08048943, 0.1151967, 0.01365218, 0.03012104, 
    -2.304602e-07, 1.436865e-08, -3.469717e-05, 0.01922728, 0.1454581, 
    0.1023064, 0.04748035, 1.96144e-05,
  0.0004330147, 0.1109929, 0.03920432, 0.1261619, 0.0550863, 0.0809868, 
    0.01562986, 0.003303544, 0.02664501, 0.0008438826, 0.004698996, 
    0.02191036, 0.03864892, 0.08611645, 0.08465668, 0.09859673, 0.07365998, 
    0.0009308334, 1.127384e-07, -1.508615e-09, 0, 5.165748e-11, 0.001627197, 
    0.1110989, 0.146804, 0.08294787, 0.04801983, 0.0016479, 3.354349e-08,
  0.02605247, 0.2403721, 0.1227053, 0.02708536, 0.05098863, 0.005849005, 
    0.01006744, 0.01372604, 0.06476357, 0.05508611, 0.02036953, 0.05042892, 
    0.05538189, 0.0185165, 0.004359476, 0.001471726, -3.097016e-06, 
    0.002422248, -2.88191e-06, -1.392385e-09, 0.0008696973, 5.823358e-06, 
    0.0007367076, 0.1054908, 0.05780366, 0.05155186, 0.146914, 0.0138573, 
    0.0001687449,
  0.0004797994, 0.0001500251, 0.005156488, 0.01277302, 0.01615235, 
    0.004028391, 0.02998672, 0.04993882, 0.05966275, 0.01767099, 0.04709184, 
    0.1054763, 0.1163108, 0.09240143, 0.04387495, 0.05557489, 0.1170393, 
    0.08663382, 0.04312212, 0.07060228, 0.0631211, 0.007249844, 0.03215614, 
    0.05394249, 0.04980321, 0.09419985, 0.01113903, 0.04387249, 0.01839637,
  0.002520189, 0.001045543, -8.195991e-07, 0.002731306, 0.03275418, 
    0.002380094, 0.006138443, 0.02890137, 0.01597592, 0.006291474, 
    0.05287954, 0.00946937, 0.0222512, 0.09144954, 0.03521389, 0.01099342, 
    0.07890148, 0.0332863, 0.01471519, 0.01878587, 0.03366594, 0.01745188, 
    0.006967289, 0.1285716, 0.03710913, 0.07323676, 0.07132064, 0.047228, 
    0.08414931,
  0.03074429, 0.07061532, 0.03631394, 0.06102586, 0.1374105, 0.09711532, 
    0.09888429, 0.01430113, 0.1159585, 0.06428194, 0.01600338, 0.02507116, 
    0.01376641, 0.01997984, 0.06191139, 0.05129493, 0.04680197, 0.07773544, 
    0.06509452, 0.02441286, 0.06037333, 0.06646096, 0.06463712, 0.06442291, 
    0.06035783, 0.1018585, 0.0569616, 0.009907926, 0.03012659,
  0.1089717, 0.1257692, 0.07938814, 0.1632462, 0.04967044, 0.07022262, 
    0.02385315, 0.1113558, 0.05443434, 0.07475843, 0.1585768, 0.1682684, 
    0.2263662, 0.2059775, 0.2065705, 0.1653944, 0.2087997, 0.2023899, 
    0.1788514, 0.1201557, 0.06294334, 0.03369521, 0.1074755, 0.1530192, 
    0.1502792, 0.1410874, 0.1792935, 0.1561578, 0.1156689,
  0.2230216, 0.2216687, 0.2626851, 0.2320966, 0.2096225, 0.2226539, 
    0.1548649, 0.01870118, 0.02131764, 0.06102043, 0.07881158, 0.03069619, 
    0.05531984, 0.1263879, 0.134542, 0.1256783, 0.1579733, 0.1976149, 
    0.3167925, 0.1952761, 0.09205947, 0.1536827, 0.1628222, 0.1977001, 
    0.1601662, 0.1527333, 0.1092218, 0.1385968, 0.2273129,
  0.1860982, 0.1729599, 0.2097147, 0.1926426, 0.1987581, 0.2568399, 
    0.1913284, 0.217766, 0.1773315, 0.04898991, 0.01198864, 0.002084094, 
    0.001255011, 0.06778004, 0.06996109, 0.08292005, 0.05677816, 0.05563148, 
    0.1242513, 0.1516403, 0.1375153, 0.1195365, 0.08435785, 0.2631032, 
    0.2329367, 0.2082028, 0.1938767, 0.1412086, 0.1641602,
  0.05017017, 0.04852379, 0.05069181, 0.1920525, 0.1934973, 0.1402717, 
    0.1007541, 0.05367018, 0.005828083, 0.008457493, 0.000150506, 
    -1.118897e-05, 0, 0.007634613, 0.03178418, 0.03481094, 0.03425299, 
    0.01286931, 0.03255152, 0.05761063, 0.05651569, 0.02255163, 0.0452251, 
    0.02665618, 0.1710826, 0.03011956, 0.00184757, 0.06099132, 0.03491776,
  0.01380529, 0.01068199, 0.004078253, 0.0045896, 0.0002818014, 0.0002663803, 
    -3.840732e-07, -7.34501e-08, 0, 0, 0, 0, 0, 0, 0.0005258986, 0.003842548, 
    0.006975011, 0.004058803, -6.209405e-05, -9.030245e-07, 0.0001156494, 
    -3.850879e-07, 0, -5.611059e-08, -2.186506e-08, -1.643453e-05, 0, 
    -0.005104327, 0.02255559,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3.353403e-06, 0.0005902312, 0.029076, 
    0.03751743, 0.03817778, 0.03321038, 0.01246419, 0.0002305893, 0, 0, 
    0.004268645, 0.06389428, 0.02852774, 0.01585803, 0.04111802, 
    9.940142e-05, 1.393584e-07,
  0.06355072, 0.1101023, 0.1526572, 0.1129104, -0.001818964, 0.004010099, 
    0.1151147, -0.001634198, 0.001958104, -0.001493857, 0.0005118824, 
    0.001660481, 0.01804904, 0.1549756, 0.1515667, 0.2013752, 0.1653749, 
    0.1455229, 0.1361403, 0.1292414, 0.1222485, 0.09929132, 0.1103102, 
    0.1466182, 0.2091081, 0.1815886, 0.1932239, 0.09985783, 0.06426994,
  0.2450052, 0.163184, 0.2029361, 0.2337202, 0.2016063, 0.2041236, 0.3071043, 
    0.2467503, 0.1570631, 0.1609241, 0.1883567, 0.2035895, 0.2787887, 
    0.1886251, 0.2938772, 0.2391527, 0.2067251, 0.2291892, 0.1807556, 
    0.1818765, 0.1910032, 0.2673025, 0.2595676, 0.2236311, 0.2883279, 
    0.2442277, 0.2117895, 0.1961364, 0.2644193,
  0.1233097, 0.1085322, 0.1333556, 0.1747778, 0.1580472, 0.1636868, 0.210695, 
    0.2040204, 0.1527243, 0.1268273, 0.1341884, 0.1413114, 0.1211643, 
    0.1363097, 0.1485384, 0.1560627, 0.1030824, 0.1483213, 0.121906, 
    0.1600723, 0.1819493, 0.174136, 0.1695149, 0.1169055, 0.06375838, 
    0.10447, 0.1638011, 0.1413676, 0.134031,
  0.1036699, 0.05753732, 0.02960439, 0.03969233, 0.08216271, 0.07703764, 
    0.1193595, 0.1430447, 0.1291613, 0.07242212, 0.06302618, 0.0889919, 
    0.0561064, 0.1345852, 0.09679269, 0.1149873, 0.1124478, 0.09848347, 
    0.09384261, 0.1102484, 0.1776054, 0.1880561, 0.0837756, 0.04617711, 
    0.06521161, 0.162041, 0.07769704, 0.0460244, 0.07774194,
  8.236249e-05, 0.001398383, 0.03762266, 0.1799861, 0.06990051, 0.03757606, 
    0.008145784, 0.008676318, 0.03118507, 0.0009417789, 0.0699464, 
    0.02100771, 0.01886855, 0.0278238, 0.09970622, 0.03799891, 0.06218426, 
    0.08575577, 0.08043581, 0.05875874, 0.1412892, 0.005596778, 6.802774e-05, 
    -6.823817e-05, 0.07309451, 0.06187405, 0.08277529, 0.08511245, 0.01899786,
  3.652813e-06, 0.01028134, 0.02445912, 0.003673274, 0.0007486996, 
    5.610932e-08, -0.0002236534, 0.02757758, 2.678642e-07, 0.0008574853, 
    0.01346009, 0.0002303904, 0.01211961, 0.1880816, 0.06095721, 0.06063434, 
    0.0951211, 0.05921637, 0.0985728, 0.01927304, 0.006497984, 1.999572e-07, 
    4.975341e-08, 0.0005371512, 0.01361366, 0.1488529, 0.08027048, 
    0.06206792, 8.499263e-06,
  0.001167567, 0.09034543, 0.0302827, 0.1209553, 0.06149033, 0.08844839, 
    0.01412699, 0.003500219, 0.02593607, 0.0005810214, 0.009818201, 
    0.01738604, 0.04876879, 0.07507271, 0.08869696, 0.07930509, 0.06346769, 
    0.00378881, 6.378787e-08, 0, 0, 3.767549e-09, 0.001920951, 0.08371755, 
    0.1250628, 0.06472136, 0.0281314, 3.820587e-05, -4.522515e-08,
  0.04643795, 0.2413551, 0.09328593, 0.02715602, 0.05223935, 0.007066566, 
    0.02184642, 0.0119243, 0.03567672, 0.04709218, 0.02489285, 0.03071873, 
    0.0488876, 0.01517207, 0.004717678, 0.001766482, -3.225301e-06, 
    0.001927474, -0.0001274881, 3.221807e-08, 0.000990991, 2.47362e-06, 
    0.0007417591, 0.09967297, 0.03906828, 0.04456689, 0.1699769, 0.009595281, 
    0.0001680685,
  0.000330643, 0.0001340353, 0.003843289, 0.01317575, 0.01908495, 
    0.003835211, 0.009489124, 0.04724124, 0.06168467, 0.01733007, 0.03462414, 
    0.09461682, 0.1048055, 0.07721241, 0.04248826, 0.05541553, 0.08967517, 
    0.08590364, 0.04722271, 0.07066129, 0.08102321, 0.01633222, 0.02601046, 
    0.05035555, 0.04121192, 0.09406735, 0.009171824, 0.01625577, 0.01793837,
  0.002037967, 4.703281e-05, 4.356889e-06, 0.001663406, 0.02882251, 
    0.0008613601, 0.004091811, 0.0246683, 0.01924751, 0.00426965, 0.04404814, 
    0.008203894, 0.02669486, 0.09398229, 0.02964044, 0.009940811, 0.06107667, 
    0.02538697, 0.02994449, 0.01293478, 0.03284019, 0.02469857, 0.004106442, 
    0.1318413, 0.02716954, 0.07570581, 0.08390687, 0.03438988, 0.07365548,
  0.0367617, 0.06642941, 0.03142321, 0.04455459, 0.1143864, 0.0787062, 
    0.08713498, 0.04541837, 0.1793466, 0.06131215, 0.0108663, 0.02134538, 
    0.01106613, 0.02028215, 0.05112571, 0.05002496, 0.03542952, 0.0753807, 
    0.05184456, 0.01676378, 0.02808854, 0.05025054, 0.06286868, 0.06609526, 
    0.05479512, 0.09845019, 0.04151523, 0.01153195, 0.0323046,
  0.1115871, 0.1096024, 0.07848539, 0.1523575, 0.02854387, 0.04685178, 
    0.05028856, 0.1123362, 0.04688602, 0.06524551, 0.148459, 0.1533567, 
    0.2241376, 0.1925117, 0.2150892, 0.1530307, 0.221487, 0.2181341, 
    0.1391547, 0.1128836, 0.07344324, 0.04052797, 0.1173905, 0.1511189, 
    0.1388179, 0.1332397, 0.1656403, 0.1388282, 0.1210494,
  0.2405555, 0.2000409, 0.2744526, 0.2397979, 0.1857687, 0.2034942, 
    0.1555938, 0.06188932, 0.03426971, 0.09846959, 0.1401411, 0.08075415, 
    0.1245809, 0.1879634, 0.1361901, 0.1465708, 0.1744981, 0.2041363, 
    0.3114471, 0.2263641, 0.1279895, 0.1753454, 0.2110053, 0.2776103, 
    0.1988183, 0.1638631, 0.1137875, 0.1581048, 0.2481944,
  0.2116634, 0.2339372, 0.2691315, 0.2749273, 0.2600435, 0.3134982, 
    0.2297864, 0.2569662, 0.2741708, 0.09680005, 0.06013409, 0.01717843, 
    -0.001513775, 0.09651392, 0.1899826, 0.1382307, 0.1206418, 0.1207244, 
    0.1517571, 0.1909813, 0.1693709, 0.178022, 0.2152514, 0.3116946, 
    0.2814054, 0.2355938, 0.2687463, 0.1924353, 0.2176001,
  0.04413803, 0.1039669, 0.2459088, 0.2722242, 0.2502174, 0.2217655, 
    0.1411412, 0.1093527, 0.02712087, 0.03537881, 0.0095453, 0.009000865, 
    0.02292375, 0.06393687, 0.07146461, 0.06049026, 0.05533586, 0.04335196, 
    0.1027031, 0.1936008, 0.09089998, 0.09362417, 0.1214562, 0.1045053, 
    0.1982882, 0.03734447, 0.005406654, 0.09860854, 0.0585227,
  0.1046323, 0.07772055, 0.06870135, 0.06165988, 0.05911493, 0.02846119, 
    0.00304967, -2.149442e-06, 0, 0, 0.0002623624, 0.0218002, 0.0349529, 
    0.05417113, 0.02115882, 0.006951139, 0.01387708, 0.03597906, 0.04928857, 
    0.05306027, 0.03189938, 0.01850837, -2.55079e-05, -0.001489075, 
    -0.001493436, -2.917801e-05, -0.004217028, 0.02874668, 0.1099856,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  -1.71803e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001145325, 0.06170427, 
    0.08648607, 0.08572701, 0.09092393, 0.07246725, 0.02565772, 0.01790774, 
    0.004147435, -9.688102e-05, 0.01929222, 0.141902, 0.08674253, 0.05854387, 
    0.06466766, 0.032428, 2.868961e-05,
  0.1488932, 0.1665071, 0.2383134, 0.1737665, 0.01329421, 0.03169963, 
    0.1539293, 0.00444952, 0.003478838, 0.005218659, 0.0001230034, 
    0.001117396, 0.03922956, 0.2744746, 0.2163956, 0.2534435, 0.1781208, 
    0.1658084, 0.2419564, 0.1668084, 0.2216879, 0.2462277, 0.1779054, 
    0.2225864, 0.3183974, 0.1982047, 0.2541112, 0.1415964, 0.1206464,
  0.2566718, 0.1833496, 0.1937434, 0.2725813, 0.2286565, 0.2529822, 
    0.3485703, 0.2608556, 0.1812062, 0.1718584, 0.2172854, 0.2746639, 
    0.3418389, 0.2312875, 0.3032087, 0.2541676, 0.2240407, 0.2117442, 0.1697, 
    0.1757835, 0.1985987, 0.2762198, 0.2481252, 0.2736557, 0.2756807, 
    0.251293, 0.2032108, 0.1906704, 0.2963346,
  0.1218421, 0.1046289, 0.1283774, 0.187379, 0.1582183, 0.163661, 0.2105264, 
    0.2074274, 0.1405997, 0.1213277, 0.1323838, 0.1485472, 0.118703, 
    0.1369059, 0.141619, 0.1392596, 0.09488686, 0.1490352, 0.125081, 
    0.1619014, 0.1694819, 0.1642499, 0.1790239, 0.1163238, 0.05763969, 
    0.08635762, 0.1463844, 0.1287055, 0.1341812,
  0.1064321, 0.06253736, 0.03095683, 0.03617457, 0.08876058, 0.0728838, 
    0.1172267, 0.1100167, 0.1157237, 0.06059876, 0.04799915, 0.08820412, 
    0.05943912, 0.1391909, 0.09729874, 0.1154737, 0.1131053, 0.09284513, 
    0.07444464, 0.09780418, 0.163101, 0.1701946, 0.05628411, 0.03427162, 
    0.07093091, 0.1517997, 0.0602567, 0.04235259, 0.07277568,
  8.778835e-05, 0.0008650087, 0.02621817, 0.1761851, 0.07671497, 0.04880464, 
    0.007646917, 0.004183802, 0.01432156, 0.0009446571, 0.08634891, 
    0.01902583, 0.01901895, 0.03649021, 0.07883178, 0.02737265, 0.05226174, 
    0.08412996, 0.06390484, 0.05098358, 0.1523352, 0.003555905, 0.000265885, 
    -0.000130892, 0.07367564, 0.05454329, 0.07506444, 0.08579651, 0.01262375,
  3.384378e-06, 0.008397324, 0.03352739, 0.0007544295, 0.001309412, 
    -2.088358e-08, -0.0001960768, 0.02825572, -9.115264e-08, 0.0001732973, 
    0.02841613, 0.0005173162, 0.01398497, 0.1325679, 0.05417288, 0.06548518, 
    0.07648128, 0.03869294, 0.08333412, 0.01750359, 0.0002706711, 
    1.08099e-08, 2.67518e-08, 0.0009068315, 0.01526919, 0.1221423, 
    0.06623571, 0.05575768, -1.123883e-05,
  0.003448635, 0.0917516, 0.03267665, 0.1095527, 0.06893282, 0.08689766, 
    0.01852975, 0.002963233, 0.02904089, 0.0006625879, 0.01563879, 
    0.01609575, 0.04630081, 0.06989038, 0.07977013, 0.08090502, 0.05360982, 
    0.005134766, -3.174648e-08, -4.251895e-11, 8.519221e-11, 4.870335e-09, 
    0.001140563, 0.06397252, 0.109487, 0.06422744, 0.01327723, -1.769697e-06, 
    -1.611252e-05,
  0.1054104, 0.2555192, 0.08488871, 0.02431287, 0.05636272, 0.01901584, 
    0.03401982, 0.007522381, 0.02628339, 0.04548334, 0.03164129, 0.01655111, 
    0.04562824, 0.01023937, 0.003950455, 0.001781151, 1.681716e-05, 
    0.0005421001, 0.006243477, 4.744074e-08, 0.0008311932, 1.087246e-06, 
    0.00695594, 0.09628429, 0.02699317, 0.03930289, 0.1604959, 0.00678474, 
    0.01484196,
  0.003527986, 0.0002281488, 0.003030211, 0.02886987, 0.0169741, 0.003150621, 
    0.001203459, 0.03944968, 0.06424504, 0.02298163, 0.02551816, 0.08911522, 
    0.09691733, 0.07406713, 0.0476452, 0.06767917, 0.05586633, 0.08322845, 
    0.06061279, 0.07095961, 0.07910869, 0.03487387, 0.02724633, 0.04010859, 
    0.0355405, 0.08221939, 0.008102683, 0.005253883, 0.0271037,
  0.0007532099, 2.792664e-06, 2.309461e-06, 0.00145648, 0.02530246, 
    0.0008232779, 0.004366349, 0.01752417, 0.01578299, 0.002710712, 
    0.03573926, 0.007378275, 0.02864047, 0.09387526, 0.02745143, 0.01086882, 
    0.04945948, 0.01871859, 0.01739069, 0.00526537, 0.02850625, 0.0264364, 
    0.002610361, 0.1283261, 0.02119325, 0.07167891, 0.09090087, 0.0318383, 
    0.04361207,
  0.03929974, 0.0289799, 0.017191, 0.03639557, 0.1065458, 0.04747294, 
    0.0735203, 0.04481661, 0.2195539, 0.05951509, 0.006449367, 0.03726855, 
    0.007312119, 0.02042953, 0.04741255, 0.03750111, 0.02493235, 0.06229436, 
    0.04246224, 0.01623676, 0.01200431, 0.05858372, 0.05345289, 0.07413619, 
    0.04913087, 0.1116632, 0.03800681, 0.01050035, 0.03776925,
  0.1233405, 0.1029118, 0.07087751, 0.134472, 0.01681079, 0.03309323, 
    0.06843662, 0.1062787, 0.03223426, 0.05337987, 0.1436922, 0.1459162, 
    0.2242737, 0.1913562, 0.2147924, 0.1394478, 0.20989, 0.2095183, 
    0.1018534, 0.09485017, 0.07980096, 0.04829901, 0.1222992, 0.139098, 
    0.1437296, 0.1287399, 0.1501229, 0.1416985, 0.1005887,
  0.263356, 0.1895761, 0.2586153, 0.2526152, 0.1706745, 0.1781939, 0.138026, 
    0.09252218, 0.0581289, 0.1305088, 0.1547096, 0.113893, 0.1462964, 
    0.1971589, 0.1442235, 0.1732939, 0.1773764, 0.1942189, 0.2936008, 
    0.2401699, 0.1626694, 0.2037486, 0.2364772, 0.3291555, 0.2293562, 
    0.1781746, 0.1141221, 0.1633255, 0.2679285,
  0.2086928, 0.2757518, 0.2795075, 0.3228299, 0.3143653, 0.3149207, 
    0.2320355, 0.2695629, 0.3381656, 0.1707592, 0.088454, 0.03267933, 
    0.01049328, 0.1400077, 0.2428924, 0.1933682, 0.1974484, 0.193424, 
    0.1917285, 0.26821, 0.1753203, 0.27417, 0.3507352, 0.3589891, 0.2985505, 
    0.2755443, 0.2791526, 0.2098583, 0.2389535,
  0.1248028, 0.1637886, 0.2493119, 0.2700619, 0.2860491, 0.2610267, 
    0.1752909, 0.1784504, 0.1258511, 0.108702, 0.06066335, 0.04726928, 
    0.09585472, 0.1690795, 0.2040475, 0.115849, 0.1281286, 0.1359033, 
    0.2248887, 0.242842, 0.109532, 0.1465348, 0.3324921, 0.2115841, 
    0.1716266, 0.0558287, 0.007900752, 0.1130013, 0.09287741,
  0.1627021, 0.165555, 0.1470632, 0.1394686, 0.1097046, 0.07675504, 
    0.05199794, 0.03366658, 0.01576919, 0.01881302, 0.03755635, 0.04071114, 
    0.04595626, 0.08969187, 0.0935979, 0.03201941, 0.01699275, 0.06463864, 
    0.0901216, 0.07935499, 0.09802246, 0.1343456, 0.05789162, -0.01183918, 
    0.01130135, 0.001848839, 0.01180767, 0.06859295, 0.1572287,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -5.385984e-05, -5.385984e-05, -5.385984e-05, -5.385984e-05, 
    -5.385984e-05, -5.385984e-05, -5.385984e-05, 0,
  0.0005680366, 0.0003388887, -1.075159e-10, 0, 0, 0, 0, 0, 0, 0, 0, 
    1.273549e-05, 0.0007269121, 0.09326658, 0.0781004, 0.0869447, 0.09642301, 
    0.0959446, 0.08537108, 0.05884396, 0.03839676, 0.009574044, 0.024077, 
    0.1833384, 0.1062337, 0.08484442, 0.1556679, 0.05680473, 0.0006289842,
  0.1638448, 0.2191868, 0.214201, 0.1839255, 0.083366, 0.124754, 0.1553796, 
    0.06428409, 0.04466096, 0.07695636, 0.006896044, 0.03418599, 0.06216267, 
    0.2929928, 0.2233576, 0.2167398, 0.1895853, 0.1907207, 0.2752263, 
    0.2001066, 0.2500302, 0.308395, 0.2753029, 0.3124247, 0.309717, 
    0.1831203, 0.2562721, 0.1522362, 0.1221364,
  0.2589748, 0.1991224, 0.2479832, 0.2645929, 0.2338849, 0.26236, 0.3700808, 
    0.2539547, 0.1918216, 0.1952903, 0.2565857, 0.3151182, 0.3462386, 
    0.240362, 0.3120323, 0.2408378, 0.2246666, 0.192148, 0.1501815, 
    0.1739361, 0.2203424, 0.2693307, 0.2389106, 0.2590214, 0.2726742, 
    0.23039, 0.196203, 0.1809821, 0.2861114,
  0.1151903, 0.09697964, 0.1332876, 0.191879, 0.1519209, 0.1635136, 
    0.2131105, 0.2103575, 0.1364375, 0.1275358, 0.1328725, 0.1720932, 
    0.1314389, 0.1621482, 0.1352234, 0.1284982, 0.09463356, 0.137213, 
    0.1337464, 0.1450636, 0.169057, 0.1712247, 0.1982002, 0.112763, 
    0.04813874, 0.07345525, 0.1385729, 0.1349465, 0.1358147,
  0.1001749, 0.06341922, 0.03196704, 0.04821641, 0.1055344, 0.07298926, 
    0.1111488, 0.1015281, 0.1191516, 0.03642423, 0.04638759, 0.08313885, 
    0.06361401, 0.1466619, 0.09760837, 0.1340473, 0.1179089, 0.09681574, 
    0.06163979, 0.08316371, 0.1647858, 0.1354361, 0.07100405, 0.02388146, 
    0.08310045, 0.1389123, 0.06232393, 0.04579595, 0.09339232,
  0.0008454102, 0.0002775009, 0.02571754, 0.1549423, 0.06842213, 0.03413482, 
    0.01129247, 0.004666139, 0.01099726, 0.0009538686, 0.07001939, 0.0107111, 
    0.0233146, 0.02375214, 0.05407649, 0.02351793, 0.05003013, 0.06111361, 
    0.04078333, 0.04275708, 0.1379635, 0.005290116, -5.806549e-06, 
    -1.860356e-05, 0.06694596, 0.0459967, 0.06511796, 0.09632713, 0.00613807,
  2.461278e-06, 0.008374218, 0.08147886, 8.471785e-05, 0.007537235, 
    -3.965089e-09, -0.0002374501, 0.02483957, -4.028978e-08, -4.389886e-05, 
    0.05459925, 0.01187864, 0.01476831, 0.1147069, 0.09003113, 0.06732118, 
    0.05640491, 0.02818636, 0.08333437, 0.007061431, 6.611829e-06, 
    1.361104e-08, 2.084352e-08, 0.001195222, 0.02142911, 0.1249838, 
    0.06703626, 0.03055098, 1.552511e-06,
  0.009504138, 0.1043993, 0.04516312, 0.09912824, 0.07657216, 0.07787651, 
    0.01741876, 0.006184932, 0.0162136, 0.001031484, 0.02745884, 0.01646083, 
    0.04726612, 0.07256602, 0.08243768, 0.08594951, 0.04506649, 0.006591307, 
    5.375572e-08, 3.212766e-09, 1.121458e-09, 9.300471e-08, 0.0007477125, 
    0.05783925, 0.1042901, 0.07706818, 0.007408116, 2.538114e-07, 0.01621646,
  0.2213603, 0.2545656, 0.08754882, 0.0238884, 0.05619972, 0.0112539, 
    0.0405782, 0.005311977, 0.02712755, 0.04866315, 0.05340744, 0.02746287, 
    0.04169768, 0.01252987, 0.004471883, 0.001153089, -2.693624e-05, 
    9.106418e-05, 0.01595412, 1.760979e-07, 0.004453565, 1.28e-06, 
    0.02378509, 0.1197262, 0.03308202, 0.01555784, 0.1485204, 0.005786127, 
    0.03781322,
  0.002047417, 0.0001691107, 0.002672578, 0.03687057, 0.02503761, 
    0.003284678, 0.002415687, 0.04290961, 0.06629153, 0.0405937, 0.02852979, 
    0.0935555, 0.1084676, 0.07895075, 0.05963747, 0.07208195, 0.04677015, 
    0.08566494, 0.07852942, 0.08864939, 0.1066763, 0.03626145, 0.03221153, 
    0.03885162, 0.03597494, 0.07065415, 0.008173874, 0.004216987, 0.02063175,
  -0.0001461317, 1.480116e-06, 2.680051e-06, 0.002070521, 0.01629286, 
    6.805905e-05, 0.006689175, 0.01074207, 0.01902944, 0.003388169, 
    0.03522005, 0.008023885, 0.03239695, 0.09349963, 0.0208847, 0.01339498, 
    0.043313, 0.02235929, 0.003958326, 0.0006966569, 0.02496555, 0.03108769, 
    0.001991692, 0.1194123, 0.01947513, 0.06371359, 0.06940367, 0.007063167, 
    0.02077686,
  0.03696308, 0.0155958, 0.005148908, 0.02780662, 0.1025392, 0.02783774, 
    0.06326206, 0.0595683, 0.2355961, 0.04755165, 0.004083129, 0.05761464, 
    0.009067722, 0.0242622, 0.04916592, 0.03967078, 0.02321723, 0.05990937, 
    0.03485914, 0.009775996, 0.006675255, 0.0631584, 0.05318134, 0.07217864, 
    0.04673865, 0.1162597, 0.04211957, 0.01050138, 0.05324643,
  0.1202966, 0.09994305, 0.06391115, 0.1216944, 0.01318205, 0.0259464, 
    0.0761546, 0.09175343, 0.02190974, 0.04150735, 0.1394598, 0.126221, 
    0.2131305, 0.1855296, 0.2058234, 0.1301801, 0.2102409, 0.1954817, 
    0.09117467, 0.07734381, 0.0662296, 0.05292571, 0.1368291, 0.1437161, 
    0.1348222, 0.121647, 0.1452557, 0.1402765, 0.09769659,
  0.2983781, 0.1799791, 0.2402441, 0.2224676, 0.1610439, 0.1467322, 
    0.1404803, 0.1279328, 0.09417553, 0.1337718, 0.1648888, 0.1229674, 
    0.1484741, 0.1969563, 0.1414673, 0.1567398, 0.1709179, 0.2033669, 
    0.2837012, 0.2595175, 0.1978973, 0.2191894, 0.2302572, 0.3379606, 
    0.205357, 0.192469, 0.1184781, 0.1780035, 0.2564243,
  0.2091798, 0.2680533, 0.2940463, 0.3268133, 0.3121133, 0.3064483, 
    0.2340294, 0.3027816, 0.365568, 0.2375714, 0.1364865, 0.0426969, 
    0.03844559, 0.1829576, 0.2374469, 0.2125461, 0.2231919, 0.219179, 
    0.2374616, 0.286075, 0.2019579, 0.2937401, 0.4302158, 0.3858626, 
    0.2827095, 0.3411087, 0.2398553, 0.1913903, 0.2411764,
  0.1688987, 0.182817, 0.2432531, 0.3002141, 0.3152725, 0.2878808, 0.2183319, 
    0.2106892, 0.2454975, 0.2182494, 0.1270435, 0.06229353, 0.1742657, 
    0.2701812, 0.3399028, 0.2735515, 0.2375655, 0.1853122, 0.2592479, 
    0.2507436, 0.1206292, 0.1802671, 0.3034111, 0.2096038, 0.1397695, 
    0.09990419, 0.02096898, 0.1055693, 0.1101241,
  0.1453684, 0.160835, 0.1633454, 0.177091, 0.1762191, 0.1707425, 0.1345721, 
    0.09474712, 0.05805144, 0.06150602, 0.05780615, 0.07387646, 0.1113927, 
    0.102113, 0.1201063, 0.1273459, 0.1085789, 0.1001032, 0.1159196, 
    0.1383511, 0.1581286, 0.1975684, 0.1248057, 0.007690009, 0.0547138, 
    0.008526702, 0.02782063, 0.0792805, 0.1624708,
  0.005770106, 0.005239251, 0.004708395, 0.00417754, 0.003646685, 0.00311583, 
    0.002584974, 0.001752094, 0.00163948, 0.001526865, 0.001414251, 
    0.001301637, 0.001189023, 0.001076409, -0.00048762, -0.0001075306, 
    0.0002725588, 0.0006526482, 0.001032738, 0.001412827, 0.001792916, 
    0.005041773, 0.005305153, 0.005568533, 0.005831913, 0.006095293, 
    0.006358674, 0.006622054, 0.00619479,
  0.001159403, 0.003063783, 0.001465679, -3.367505e-06, 0, -1.157652e-05, 0, 
    0, 0, 0, -7.156119e-06, 0.000146639, 0.008367135, 0.08731987, 0.07096571, 
    0.085205, 0.1064738, 0.09982274, 0.09420459, 0.1107738, 0.08381867, 
    0.02852341, 0.05762542, 0.1834291, 0.09394246, 0.06591228, 0.13754, 
    0.174534, 0.004300921,
  0.1691433, 0.2334549, 0.1974149, 0.1889373, 0.1773915, 0.1906236, 
    0.1415235, 0.1213804, 0.07654507, 0.1967608, 0.108703, 0.08864998, 
    0.06450576, 0.2842475, 0.2333344, 0.2188838, 0.191833, 0.1980396, 
    0.2614967, 0.2014422, 0.2507464, 0.3188853, 0.281527, 0.3409033, 
    0.2975036, 0.1622067, 0.2551346, 0.1546638, 0.1318543,
  0.2608542, 0.2162642, 0.302288, 0.276332, 0.2400675, 0.2704492, 0.3846963, 
    0.2358249, 0.1923285, 0.2081734, 0.2630024, 0.3175117, 0.3216073, 
    0.2453839, 0.3249506, 0.2652696, 0.2626649, 0.1775999, 0.1583716, 
    0.175994, 0.2247894, 0.2398198, 0.2326968, 0.2754321, 0.2518332, 
    0.2279251, 0.188901, 0.1736542, 0.2732506,
  0.1249102, 0.1105236, 0.1474018, 0.2184197, 0.1615249, 0.1776081, 
    0.2064374, 0.1952379, 0.1609529, 0.1353509, 0.1429474, 0.1872855, 
    0.1457015, 0.1766092, 0.1336233, 0.11188, 0.1187078, 0.1447679, 
    0.1316086, 0.147884, 0.1617397, 0.1661672, 0.1883542, 0.1058121, 
    0.04728057, 0.09058036, 0.1267928, 0.1558245, 0.1408388,
  0.09309638, 0.0690238, 0.02724596, 0.05057769, 0.1157123, 0.07442702, 
    0.1046377, 0.09318903, 0.1185499, 0.02332329, 0.04713516, 0.06555846, 
    0.06440823, 0.1358442, 0.09622838, 0.1380618, 0.08160509, 0.1074911, 
    0.05384149, 0.08679163, 0.1271232, 0.130078, 0.05770069, 0.01899496, 
    0.1042234, 0.1533344, 0.05973788, 0.05712783, 0.1046292,
  0.002450959, 0.0001630036, 0.05149603, 0.1473414, 0.04422205, 0.02886282, 
    0.01659391, 0.007982983, 0.008167785, 0.0001832563, 0.03470711, 
    0.01305267, 0.03329321, 0.00919659, 0.03760825, 0.02977134, 0.05227333, 
    0.05439601, 0.03805987, 0.04371268, 0.1184932, 0.01692214, 0.0001929434, 
    -9.954045e-07, 0.07344577, 0.04231995, 0.05908529, 0.09380563, 
    5.148432e-05,
  6.617481e-06, 0.0129747, 0.1679981, 7.269494e-05, 0.01288624, 9.386028e-07, 
    -0.000191954, 0.02904034, -8.290777e-06, 0.001337792, 0.05522454, 
    0.03950142, 0.02217131, 0.1109191, 0.08828209, 0.07826763, 0.05978785, 
    0.02843017, 0.08107647, 0.004220332, 4.890177e-07, 1.942572e-08, 
    2.635841e-07, 0.00299796, 0.01856854, 0.1326321, 0.07822682, 0.01078798, 
    3.206424e-06,
  0.007790123, 0.1307925, 0.08053264, 0.08655022, 0.08833099, 0.07275219, 
    0.02223452, 0.01202947, 0.01091389, 0.001571016, 0.03093345, 0.02604006, 
    0.05790365, 0.08360431, 0.08978888, 0.09898034, 0.03816463, 0.0061969, 
    3.547294e-06, 1.239756e-07, 9.340015e-09, 1.27289e-06, 0.003091697, 
    0.07198807, 0.1333202, 0.1042388, 0.00114619, 5.923819e-07, 0.002256094,
  0.2770443, 0.290204, 0.1210857, 0.02568667, 0.05690367, 0.005950685, 
    0.0387734, 0.008635839, 0.03338952, 0.07090344, 0.07931642, 0.05761388, 
    0.05767293, 0.01582164, 0.003566011, 0.001189114, 9.449766e-05, 
    0.0006328803, 0.0008025328, 7.524418e-06, -8.320466e-06, 6.836129e-06, 
    0.03351839, 0.1474746, 0.05582193, 0.01138676, 0.1493771, 0.007111709, 
    0.05139539,
  0.0005302961, 0.0003626411, 0.003614476, 0.01996505, 0.03568424, 
    0.004645341, 0.005141877, 0.04708197, 0.07713552, 0.0596692, 0.03245311, 
    0.1059273, 0.1400377, 0.1056073, 0.06814193, 0.08466552, 0.04986412, 
    0.09902089, 0.1126648, 0.1200509, 0.1308877, 0.04209498, 0.05647729, 
    0.04382502, 0.03930301, 0.07872247, 0.01339363, 0.005475566, 0.01725073,
  -7.669418e-05, 1.655598e-06, 2.190884e-06, 0.003511773, 0.0111291, 
    0.000117785, 0.01003172, 0.003920306, 0.02445205, 0.008497479, 
    0.04411598, 0.01604316, 0.03437644, 0.1047528, 0.02189536, 0.01936002, 
    0.03276569, 0.02977995, 0.001115431, 1.804185e-05, 0.02663621, 0.0432989, 
    0.003142758, 0.1070246, 0.02532228, 0.0680197, 0.05581069, 0.003888977, 
    0.01073448,
  0.02420145, 0.01129986, 0.003484115, 0.02636677, 0.0969997, 0.0179136, 
    0.06513179, 0.1172638, 0.2324172, 0.04507675, 0.002209196, 0.08554608, 
    0.02141726, 0.02956272, 0.0533473, 0.04329991, 0.03268371, 0.05732643, 
    0.01694224, 0.008571536, 0.005634274, 0.07205419, 0.05268872, 0.07476488, 
    0.04632444, 0.1162057, 0.05234256, 0.009527073, 0.08849989,
  0.1017378, 0.09997995, 0.03669279, 0.111718, 0.009482794, 0.02085398, 
    0.07566179, 0.0704348, 0.02031216, 0.03770526, 0.133856, 0.1123577, 
    0.1781085, 0.1754575, 0.1834127, 0.1337814, 0.204858, 0.1892616, 
    0.09565005, 0.05993957, 0.06274935, 0.04571736, 0.1428942, 0.1444283, 
    0.1341285, 0.115176, 0.1381418, 0.1362624, 0.08920843,
  0.2610893, 0.1547859, 0.2438102, 0.2096165, 0.1485934, 0.1298991, 
    0.1063527, 0.1609977, 0.1064627, 0.1471837, 0.1630331, 0.1179236, 
    0.1586375, 0.1987295, 0.1512103, 0.1445555, 0.1617084, 0.2260562, 
    0.2648276, 0.2770303, 0.2020972, 0.1849216, 0.2243101, 0.3271208, 
    0.2065637, 0.1847, 0.1139998, 0.205891, 0.2494278,
  0.2021113, 0.285905, 0.269361, 0.3089625, 0.3341911, 0.2918818, 0.2613091, 
    0.3076447, 0.4127649, 0.291314, 0.1927458, 0.05780933, 0.1041212, 
    0.2180017, 0.1979295, 0.1840128, 0.2364652, 0.212142, 0.2794544, 
    0.2691684, 0.189683, 0.3154103, 0.4350773, 0.3561728, 0.2843563, 
    0.3547165, 0.1965344, 0.1962815, 0.2377961,
  0.1434406, 0.1894029, 0.2309896, 0.3737662, 0.4040878, 0.3065571, 
    0.2078559, 0.2082637, 0.2556278, 0.2471615, 0.1855312, 0.1456095, 
    0.2105864, 0.3164947, 0.3557113, 0.2789681, 0.2680774, 0.1924095, 
    0.2716523, 0.2552451, 0.1620418, 0.213609, 0.3105051, 0.221426, 
    0.1306697, 0.1178467, 0.04833527, 0.100418, 0.1752932,
  0.1294551, 0.1368608, 0.1639781, 0.1852863, 0.1897983, 0.1928582, 
    0.2104897, 0.173772, 0.1574793, 0.1470028, 0.1127663, 0.1271477, 
    0.1651676, 0.1248989, 0.1600102, 0.1531726, 0.2142783, 0.2777663, 
    0.2349338, 0.1775163, 0.2347326, 0.2644413, 0.1735243, 0.03185493, 
    0.08846249, 0.01268967, 0.04434698, 0.09138317, 0.1524661,
  0.01464422, 0.01385491, 0.01306559, 0.01227628, 0.01148697, 0.01069765, 
    0.009908339, 0.01062692, 0.01042406, 0.01022121, 0.01001836, 0.009815504, 
    0.009612651, 0.009409797, 0.005776464, 0.006660927, 0.007545391, 
    0.008429855, 0.009314319, 0.01019878, 0.01108325, 0.01865046, 0.01875816, 
    0.01886586, 0.01897356, 0.01908127, 0.01918897, 0.01929667, 0.01527567,
  -9.875018e-05, 0.01295865, 0.02108196, 0.009532487, 0.001689846, 
    -0.0004602962, -0.001189746, -0.0002689318, 5.22606e-05, 0.001386621, 
    -0.0001769821, 0.00812504, 0.0679944, 0.07976026, 0.06472041, 0.08552005, 
    0.12243, 0.1104246, 0.08519616, 0.1091266, 0.1387938, 0.113825, 
    0.08213117, 0.1627819, 0.09625718, 0.06669586, 0.1360099, 0.1577587, 
    0.03350196,
  0.1731038, 0.2296293, 0.1842275, 0.1938644, 0.2299681, 0.1978717, 
    0.1573439, 0.1986524, 0.1719111, 0.3073227, 0.2270809, 0.1001692, 
    0.08466056, 0.2768951, 0.2221838, 0.208315, 0.1726513, 0.1829879, 
    0.2854955, 0.2383747, 0.2579626, 0.319851, 0.2560264, 0.3757925, 
    0.2885125, 0.1447471, 0.2646022, 0.1790434, 0.1383136,
  0.2471749, 0.2269391, 0.3284393, 0.3185305, 0.3173738, 0.2633239, 
    0.3644632, 0.2370586, 0.1938925, 0.198216, 0.285356, 0.3496104, 
    0.3595168, 0.2448138, 0.310622, 0.2454791, 0.1991031, 0.1877314, 
    0.1409695, 0.1508446, 0.2386315, 0.2165134, 0.2382465, 0.2876239, 
    0.256743, 0.2336314, 0.20554, 0.1788984, 0.2575261,
  0.1274028, 0.130444, 0.1754681, 0.221356, 0.162869, 0.1391326, 0.1979879, 
    0.2009844, 0.1957929, 0.1578882, 0.167562, 0.2235915, 0.1868723, 
    0.1679788, 0.1274476, 0.1247062, 0.1095597, 0.1371763, 0.1069625, 
    0.1457789, 0.165262, 0.1483149, 0.1852212, 0.1015269, 0.06022847, 
    0.08734865, 0.1147748, 0.1368617, 0.1274181,
  0.08413045, 0.05059563, 0.01978564, 0.06530026, 0.1174365, 0.08264419, 
    0.0959962, 0.08861732, 0.1079303, 0.01649345, 0.03438044, 0.0533323, 
    0.06738095, 0.1239294, 0.1081685, 0.1424432, 0.06365237, 0.1082049, 
    0.05003875, 0.09433379, 0.1306899, 0.09621596, 0.0612173, 0.01630919, 
    0.09987285, 0.1724278, 0.07473732, 0.06952133, 0.09664784,
  0.005445775, -5.975596e-05, 0.06579756, 0.1586973, 0.03631033, 0.02891964, 
    0.02386324, 0.005164196, 0.003180734, -4.248958e-06, 0.01998921, 
    0.002546388, 0.03091633, 0.008811708, 0.03235204, 0.03042721, 0.05214558, 
    0.05438432, 0.04591454, 0.04527087, 0.1074406, 0.01426658, 0.0001019449, 
    -6.254937e-09, 0.08146252, 0.04135162, 0.07553655, 0.07204498, 
    5.636975e-05,
  7.795543e-06, 0.01491164, 0.2144258, 8.184111e-05, 0.009842121, 
    1.623126e-06, -8.843736e-05, 0.01669845, 0.0002483826, 0.0005336627, 
    0.03950115, 0.04148138, 0.0247338, 0.109989, 0.07168801, 0.08082782, 
    0.06922938, 0.03341623, 0.09841645, 0.00473045, 1.248318e-07, 
    4.365877e-08, 1.338512e-07, 0.002565667, 0.03326858, 0.1424886, 
    0.08984723, 0.001799471, 6.350684e-06,
  0.00681756, 0.1707347, 0.1242822, 0.09359743, 0.09536225, 0.07143096, 
    0.02418966, 0.01905914, 0.006384349, 0.002341622, 0.0286621, 0.03342714, 
    0.06515741, 0.08365706, 0.09497555, 0.1237464, 0.03560985, 0.004366247, 
    8.130796e-06, -2.15308e-07, 3.662888e-08, -4.369864e-07, 0.004506859, 
    0.08044249, 0.1731026, 0.1728153, 0.0002631794, 1.445241e-06, 0.0002530101,
  0.2776839, 0.3524149, 0.1723304, 0.04376959, 0.05764886, 0.003795455, 
    0.04003215, 0.01270472, 0.04893563, 0.1089458, 0.09304868, 0.07352754, 
    0.07054681, 0.01407596, 0.003164657, 0.004645631, 9.602197e-06, 
    0.004820967, -0.0002054249, 0.0001490202, 0.0003438192, 1.232283e-05, 
    0.04924785, 0.173067, 0.07965927, 0.01140835, 0.1625398, 0.01040437, 
    0.03963809,
  0.001878937, 0.0006692291, 0.006090669, 0.0417421, 0.03869546, 0.009308591, 
    0.008289129, 0.05051289, 0.09422696, 0.06527579, 0.04785379, 0.1115918, 
    0.1549063, 0.123739, 0.07765344, 0.08004287, 0.05624084, 0.09498054, 
    0.1174474, 0.1609641, 0.1246699, 0.05623228, 0.08472635, 0.05975955, 
    0.03959375, 0.08264881, 0.03185571, 0.01215601, 0.01138953,
  7.740144e-05, 3.665545e-06, 2.004984e-05, 0.00776383, 0.009231233, 
    0.0001731305, 0.01232593, 0.01156907, 0.03113329, 0.01767332, 0.06060865, 
    0.01497664, 0.03493438, 0.09853734, 0.02696577, 0.03373402, 0.03305029, 
    0.03117615, 0.0008596766, 0.0001891182, 0.04145187, 0.05208936, 
    0.004489824, 0.1131806, 0.0319646, 0.06953762, 0.04768883, 0.01926112, 
    0.02223622,
  0.007482722, 0.01917346, 0.005329006, 0.02488313, 0.09631516, 0.01407874, 
    0.05810339, 0.1529904, 0.229151, 0.06409201, 0.0001076577, 0.08881617, 
    0.04359058, 0.04175851, 0.06400799, 0.04281053, 0.03303538, 0.05766097, 
    0.005539666, 0.0112244, 0.01288818, 0.08318987, 0.05535904, 0.07937589, 
    0.04728007, 0.1187569, 0.05619691, 0.01084179, 0.08773916,
  0.0865605, 0.09728803, 0.02624189, 0.1105171, 0.01687859, 0.0423595, 
    0.07362018, 0.04018957, 0.01829697, 0.03229428, 0.1246844, 0.1088467, 
    0.1519896, 0.1541119, 0.1599047, 0.1437646, 0.2043231, 0.188153, 
    0.09849096, 0.0608892, 0.06372287, 0.05552232, 0.1292718, 0.1410332, 
    0.1348125, 0.09827996, 0.1240137, 0.1276296, 0.0937577,
  0.2476866, 0.1441948, 0.2395684, 0.1909482, 0.1198754, 0.1135634, 
    0.1076006, 0.1736297, 0.1107481, 0.1484221, 0.162355, 0.1135695, 
    0.1554378, 0.2056678, 0.1572076, 0.1322501, 0.151223, 0.2031927, 
    0.2459217, 0.2639818, 0.1867478, 0.1965871, 0.2379276, 0.3151452, 
    0.2178884, 0.1926302, 0.122984, 0.2075843, 0.2343949,
  0.1975435, 0.3070476, 0.2938102, 0.4029061, 0.3791894, 0.3011143, 
    0.2810001, 0.3235162, 0.4375391, 0.3103499, 0.2170934, 0.1031525, 
    0.1258317, 0.21055, 0.1658695, 0.1683701, 0.2479846, 0.2218002, 
    0.2772282, 0.2658098, 0.2096394, 0.2704325, 0.4764637, 0.3936777, 
    0.2930416, 0.3560474, 0.210509, 0.2237963, 0.2029025,
  0.1501023, 0.1420555, 0.2123639, 0.3932302, 0.416577, 0.2914924, 0.2071469, 
    0.2160289, 0.24854, 0.2461914, 0.1929957, 0.1833886, 0.1876613, 0.3181, 
    0.3719217, 0.2791318, 0.2586219, 0.1933668, 0.2703886, 0.2530171, 
    0.1627864, 0.192563, 0.2997584, 0.2390789, 0.1177665, 0.1146647, 
    0.05966383, 0.09780885, 0.1446579,
  0.1403651, 0.1244418, 0.1834632, 0.2154042, 0.1951742, 0.1937594, 
    0.2332801, 0.2012412, 0.1799405, 0.220737, 0.2239692, 0.1793359, 
    0.2022031, 0.1425905, 0.1721332, 0.1697053, 0.2360106, 0.3150368, 
    0.3221145, 0.2183509, 0.3006345, 0.3150798, 0.2007374, 0.08666721, 
    0.1305029, 0.01902305, 0.04552297, 0.08975638, 0.2054775,
  0.02625817, 0.02518668, 0.02411519, 0.0230437, 0.02197221, 0.02090072, 
    0.01982924, 0.01957732, 0.01987235, 0.02016738, 0.02046242, 0.02075745, 
    0.02105249, 0.02134752, 0.02387135, 0.02492017, 0.02596899, 0.0270178, 
    0.02806662, 0.02911543, 0.03016425, 0.03156602, 0.03129366, 0.03102129, 
    0.03074893, 0.03047657, 0.03020421, 0.02993185, 0.02711536,
  0.008766535, 0.02011747, 0.03571406, 0.03134743, 0.02933468, 0.005203595, 
    0.01454042, 0.01549353, 0.01276068, 0.002452903, 0.01278417, 0.071303, 
    0.08625448, 0.07230977, 0.04975931, 0.07135883, 0.1208563, 0.1201441, 
    0.08393741, 0.09357542, 0.1386382, 0.1885837, 0.1049898, 0.1535629, 
    0.101028, 0.0708539, 0.128821, 0.1326885, 0.0779145,
  0.1938301, 0.2327195, 0.2072335, 0.2446202, 0.2773101, 0.1917249, 
    0.1769848, 0.255817, 0.2410646, 0.3267301, 0.2369964, 0.1105832, 
    0.0997633, 0.2741981, 0.2111901, 0.207198, 0.2051322, 0.2300829, 
    0.3158147, 0.2291547, 0.2573516, 0.2976694, 0.276947, 0.4082431, 
    0.2964995, 0.1439901, 0.245488, 0.1985704, 0.1633499,
  0.2279781, 0.2382464, 0.3763911, 0.3645625, 0.3797969, 0.3045032, 
    0.3691292, 0.2347301, 0.2416671, 0.2185058, 0.2745315, 0.3670771, 
    0.3437114, 0.2683276, 0.2924669, 0.2579048, 0.2401948, 0.2004433, 
    0.1680068, 0.1899259, 0.254335, 0.2405968, 0.2403301, 0.2797527, 
    0.2258955, 0.2390992, 0.2149232, 0.1917088, 0.2356746,
  0.1291417, 0.1352308, 0.1833435, 0.2336307, 0.1603184, 0.1601774, 0.191437, 
    0.1723547, 0.1916405, 0.155764, 0.2100306, 0.2452511, 0.1905124, 
    0.1803068, 0.1234257, 0.1177472, 0.1134147, 0.1340849, 0.1232179, 
    0.123658, 0.1481472, 0.1545416, 0.1849105, 0.1037821, 0.06445833, 
    0.08254156, 0.1187984, 0.137545, 0.1238425,
  0.08130601, 0.07190318, 0.02225861, 0.09244746, 0.1220878, 0.0918743, 
    0.09973647, 0.0870565, 0.114668, 0.02269998, 0.02865655, 0.04576048, 
    0.06008868, 0.1015577, 0.1240561, 0.1421807, 0.07850315, 0.1163588, 
    0.05563346, 0.105866, 0.141338, 0.0861541, 0.07359505, 0.01753284, 
    0.09305642, 0.1659252, 0.09165769, 0.07551666, 0.1184527,
  0.006601868, -3.426796e-05, 0.0914808, 0.1773536, 0.02065107, 0.03891401, 
    0.02818422, 0.004403146, 0.004503264, 2.116056e-06, 0.005437169, 
    0.0003342478, 0.03072843, 0.009833364, 0.03413044, 0.03657412, 
    0.05135469, 0.05299169, 0.0530739, 0.05565453, 0.09734424, 0.0189853, 
    4.614598e-06, 1.185945e-07, 0.08176529, 0.04752878, 0.1057428, 
    0.06809583, 0.00046473,
  3.886416e-06, 0.01435853, 0.1556029, 8.582357e-05, 0.007432334, 
    7.056784e-05, -0.0001997782, 0.006291224, 4.328247e-06, 4.163719e-06, 
    0.01424596, 0.01114938, 0.02408797, 0.1105715, 0.05688495, 0.0837829, 
    0.07970133, 0.03864628, 0.1148182, 0.006526096, 2.511528e-07, 
    2.99985e-08, 7.06756e-08, 0.0002030845, 0.04935748, 0.1696721, 0.1123658, 
    0.001714202, 5.816627e-06,
  0.001140172, 0.1347022, 0.1379161, 0.09786474, 0.09571868, 0.07145407, 
    0.02804668, 0.01785284, 0.005059727, 0.006014952, 0.02939202, 0.020792, 
    0.05203455, 0.068136, 0.08133956, 0.1146164, 0.04094742, 0.005522656, 
    0.0001524883, -1.288948e-05, 4.559666e-08, 0.0003099786, 0.002139097, 
    0.09027739, 0.1566833, 0.1970933, 0.006282711, 1.240976e-06, 4.162617e-05,
  0.2753032, 0.4103115, 0.1860399, 0.06791169, 0.05879742, 0.005001712, 
    0.03901462, 0.0167133, 0.05822906, 0.1287694, 0.09167572, 0.06658486, 
    0.0542509, 0.01223394, 0.002905537, 0.00317947, 0.0001633422, 
    0.001331703, -5.394809e-05, 0.0001692864, 0.009026742, 0.0009945057, 
    0.06035317, 0.160813, 0.09404832, 0.009186212, 0.1178988, 0.01615676, 
    0.0410389,
  0.002108671, 0.000582272, 0.01324313, 0.04857027, 0.0430163, 0.006949132, 
    0.01847651, 0.04929968, 0.1036036, 0.04858305, 0.04712694, 0.09133349, 
    0.1162545, 0.1108475, 0.08192687, 0.07043115, 0.05679471, 0.08658855, 
    0.1290783, 0.1395467, 0.1307701, 0.05404813, 0.1112806, 0.06972194, 
    0.03842471, 0.07401707, 0.05787593, 0.01091388, 0.002739068,
  1.388928e-05, 2.898906e-06, 0.001675478, 0.01394087, 0.01326618, 
    0.0001887122, 0.01390991, 0.02485208, 0.03793095, 0.01956389, 0.04838441, 
    0.01754024, 0.03549482, 0.09633726, 0.02229955, 0.03843627, 0.0388295, 
    0.03403481, 0.001017367, 0.001930358, 0.05292687, 0.06406865, 
    0.002711703, 0.1218498, 0.03179318, 0.0741569, 0.05034442, 0.02171928, 
    0.01706963,
  0.002947257, 0.009531152, 0.01304185, 0.01936012, 0.1009103, 0.01172432, 
    0.0389008, 0.1512111, 0.2302617, 0.07308275, 0.004482095, 0.0932462, 
    0.05576488, 0.07441215, 0.1072115, 0.05018797, 0.03372438, 0.06357332, 
    0.002256084, 0.005876024, 0.02126475, 0.08398017, 0.06701534, 0.08280499, 
    0.05709391, 0.1204453, 0.06368992, 0.01425213, 0.07325275,
  0.0702256, 0.1000176, 0.02887601, 0.1177669, 0.01289629, 0.02749847, 
    0.08196189, 0.02531189, 0.01530503, 0.02598857, 0.1140285, 0.1102877, 
    0.1321272, 0.1293673, 0.1454777, 0.1581749, 0.2074058, 0.1858109, 
    0.1130235, 0.05909897, 0.06938451, 0.04973675, 0.1212633, 0.137032, 
    0.1439517, 0.1046205, 0.1245942, 0.1328324, 0.1051031,
  0.2472834, 0.11728, 0.2175778, 0.1879146, 0.1466641, 0.1332064, 0.1077583, 
    0.1835554, 0.1122913, 0.1509423, 0.1596863, 0.1048262, 0.1430475, 
    0.2071888, 0.1743145, 0.1264212, 0.1449215, 0.2110967, 0.2582405, 
    0.2566487, 0.1735208, 0.1968147, 0.2722222, 0.3094431, 0.2236473, 
    0.1896085, 0.1467148, 0.2006758, 0.2269803,
  0.2085442, 0.3185565, 0.2553453, 0.349321, 0.385676, 0.3288248, 0.2740127, 
    0.3294853, 0.4344124, 0.3133315, 0.2370938, 0.1293637, 0.154704, 
    0.2024366, 0.154722, 0.1704866, 0.2540633, 0.2472827, 0.2653721, 
    0.2642656, 0.2435674, 0.3460848, 0.4467039, 0.3837039, 0.2546805, 
    0.3431121, 0.2011597, 0.223159, 0.2252418,
  0.1705345, 0.1830408, 0.2745239, 0.3961009, 0.4414858, 0.2552527, 
    0.2055195, 0.226942, 0.2485369, 0.2407835, 0.1932619, 0.203567, 
    0.1718165, 0.3051864, 0.3771004, 0.2728598, 0.2613955, 0.2093167, 
    0.2606702, 0.2762427, 0.1685483, 0.1932213, 0.259239, 0.273093, 
    0.1168816, 0.1271147, 0.07593136, 0.09672488, 0.1300743,
  0.1223415, 0.1286936, 0.202818, 0.2257251, 0.2216194, 0.2014535, 0.2460398, 
    0.222642, 0.1738674, 0.2101164, 0.2026091, 0.169766, 0.1840097, 
    0.1340646, 0.1590476, 0.1513507, 0.2003666, 0.2695848, 0.2798056, 
    0.2773343, 0.3065831, 0.3335655, 0.2314352, 0.1212541, 0.1542618, 
    0.05861815, 0.05322568, 0.1240918, 0.2129599,
  0.06238401, 0.06150869, 0.06063338, 0.05975807, 0.05888276, 0.05800745, 
    0.05713214, 0.04692703, 0.04506294, 0.04319885, 0.04133476, 0.03947067, 
    0.03760657, 0.03574248, 0.03143785, 0.03328687, 0.03513588, 0.0369849, 
    0.03883392, 0.04068293, 0.04253195, 0.03889273, 0.03978312, 0.0406735, 
    0.04156389, 0.04245427, 0.04334466, 0.04423504, 0.06308425,
  0.02986054, 0.03213101, 0.06922974, 0.07223701, 0.08205822, 0.03766213, 
    0.03023827, 0.01609951, 0.02142962, 0.01418855, 0.07356397, 0.08581904, 
    0.08640483, 0.07141785, 0.05177034, 0.08752821, 0.1038194, 0.1211966, 
    0.07797191, 0.07882993, 0.1319425, 0.211484, 0.1346104, 0.1626775, 
    0.1140444, 0.07512788, 0.1267203, 0.1246591, 0.06562714,
  0.2185583, 0.2460579, 0.2252961, 0.2621909, 0.3068281, 0.1955882, 
    0.2099989, 0.2758732, 0.2769132, 0.3131555, 0.2373144, 0.1256912, 
    0.1027754, 0.293807, 0.2177276, 0.2052382, 0.2399668, 0.2559941, 
    0.3274536, 0.2244374, 0.278385, 0.3427209, 0.2978263, 0.4277261, 
    0.2788549, 0.1505583, 0.2661681, 0.195486, 0.1915085,
  0.2691246, 0.2360057, 0.3910638, 0.4715219, 0.3172377, 0.2615655, 
    0.3183721, 0.2906325, 0.2435066, 0.2413056, 0.3167457, 0.4105032, 
    0.3761421, 0.263693, 0.3119867, 0.2321829, 0.2123777, 0.2102673, 
    0.1411359, 0.1729975, 0.2781722, 0.2793033, 0.2653534, 0.3019707, 
    0.2413454, 0.2181691, 0.2382103, 0.1991698, 0.2652898,
  0.1277184, 0.155808, 0.2098962, 0.2593834, 0.175071, 0.1674455, 0.2011018, 
    0.2073552, 0.2351325, 0.1898306, 0.2234441, 0.2436879, 0.1776282, 
    0.1587892, 0.1129148, 0.1528416, 0.1277689, 0.1252483, 0.1356093, 
    0.1380357, 0.1489605, 0.1572024, 0.184533, 0.1121636, 0.07595982, 
    0.07557049, 0.1044951, 0.1459485, 0.1184835,
  0.08497608, 0.07720471, 0.03400706, 0.1007868, 0.1333565, 0.09924192, 
    0.1192116, 0.07522155, 0.1124565, 0.05149481, 0.02471547, 0.02803028, 
    0.05300685, 0.1119585, 0.1107488, 0.1583426, 0.09451193, 0.1211343, 
    0.05984421, 0.1088707, 0.1539868, 0.0865247, 0.05703122, 0.02030981, 
    0.09182651, 0.182609, 0.08910133, 0.08818551, 0.1263674,
  0.008228998, -1.850648e-06, 0.07539415, 0.1461599, 0.02584581, 0.03427633, 
    0.01845405, 0.002970782, 0.0168543, 2.063547e-06, 0.001972024, 
    0.0007733807, 0.03077189, 0.01484906, 0.03749281, 0.04823541, 0.06192597, 
    0.0534119, 0.06527895, 0.07713502, 0.09185833, 0.02630662, 5.352294e-06, 
    1.120939e-07, 0.06900574, 0.06249214, 0.1087291, 0.08643259, 0.003011255,
  9.412843e-07, 0.009882675, 0.06921515, 4.935007e-05, 0.003308418, 
    0.0003355787, -0.0001383185, 0.0007590399, -2.336737e-07, 2.807691e-07, 
    0.002057847, 0.006122958, 0.01692705, 0.0849955, 0.05144346, 0.07837655, 
    0.09124365, 0.03838377, 0.1102434, 0.0388231, 6.031076e-08, 
    -2.166891e-07, 3.042403e-08, 6.154407e-06, 0.07133707, 0.1997594, 
    0.1059335, 0.001166516, 4.121274e-06,
  0.002388909, 0.09288085, 0.09903832, 0.0859639, 0.0914775, 0.06461722, 
    0.03688597, 0.02585767, 0.003255918, 0.002464631, 0.02880646, 0.01597053, 
    0.04900041, 0.05477557, 0.07463688, 0.09455731, 0.03927106, 0.01124989, 
    0.001030337, 0.0003102668, 8.040738e-08, 1.327931e-05, 0.0001116859, 
    0.05493117, 0.09323999, 0.1539199, 0.01065075, 8.978548e-07, -2.024816e-05,
  0.244588, 0.3722147, 0.1097986, 0.0892733, 0.05056029, 0.007638549, 
    0.04119743, 0.01461423, 0.06383345, 0.1223252, 0.08189186, 0.06110855, 
    0.04342111, 0.01269076, 0.00366324, 0.001652165, 5.353393e-05, 
    5.999675e-05, -0.0001210404, 0.0006602888, 0.005403675, 0.01211411, 
    0.02807397, 0.1144635, 0.1120929, 0.004085501, 0.09476738, 0.01993051, 
    0.0423763,
  0.001955125, 0.002228906, 0.0272492, 0.06239711, 0.03975758, 0.007274278, 
    0.01749147, 0.04767033, 0.09572292, 0.03556117, 0.05286239, 0.07280221, 
    0.09139238, 0.1003683, 0.08548548, 0.06895137, 0.05040479, 0.07457327, 
    0.1403238, 0.135369, 0.1516349, 0.04847096, 0.1127832, 0.07377712, 
    0.03746189, 0.05999639, 0.04372068, 0.009047484, 0.001117189,
  1.772564e-05, 1.815398e-06, 0.01377478, 0.01609911, 0.03003592, 
    0.0001585603, 0.01510716, 0.02772585, 0.04143964, 0.02962918, 0.03667158, 
    0.02490045, 0.03375057, 0.1021052, 0.02404678, 0.04483218, 0.03529315, 
    0.03006927, 0.002157368, 0.001374163, 0.03636216, 0.08011319, 0.00299896, 
    0.1049335, 0.03447906, 0.07600099, 0.04374301, 0.02323489, 0.004791828,
  0.008610184, 0.006927602, 0.01804146, 0.02235137, 0.1087822, 0.008094118, 
    0.0256065, 0.1462445, 0.2378205, 0.08260217, 0.01474801, 0.1048538, 
    0.07758035, 0.1073224, 0.1334145, 0.06383536, 0.03328684, 0.0658415, 
    0.003128679, 0.003027589, 0.02690672, 0.09134066, 0.0811877, 0.07009586, 
    0.06048092, 0.1219772, 0.07769533, 0.014579, 0.07254839,
  0.05964967, 0.1035849, 0.02981468, 0.1407222, 0.01781217, 0.0192618, 
    0.0973516, 0.02225847, 0.01571892, 0.0161547, 0.1152228, 0.1071492, 
    0.1226193, 0.1084849, 0.147577, 0.1633285, 0.2085232, 0.1705661, 
    0.1235018, 0.05401086, 0.0790112, 0.03877966, 0.1193251, 0.153112, 
    0.1535541, 0.122854, 0.1358573, 0.1501632, 0.1186041,
  0.2305614, 0.1132417, 0.2450515, 0.1900219, 0.1161317, 0.1008447, 
    0.09070281, 0.1890149, 0.1046191, 0.150407, 0.1515746, 0.09466194, 
    0.1454673, 0.2094922, 0.2138406, 0.1325841, 0.1436485, 0.1917063, 
    0.2587679, 0.2542632, 0.1840338, 0.2346278, 0.2398194, 0.3930292, 
    0.2288247, 0.2059337, 0.1671822, 0.2037818, 0.215878,
  0.2242691, 0.3437475, 0.2719187, 0.3422589, 0.4247276, 0.3276815, 
    0.3585487, 0.387305, 0.4914173, 0.373209, 0.2637046, 0.1349293, 0.164933, 
    0.1996722, 0.1671732, 0.1744955, 0.2452288, 0.2791169, 0.2516632, 
    0.2642228, 0.3295555, 0.3282822, 0.4900862, 0.3816169, 0.2710908, 
    0.3229989, 0.1663599, 0.2290229, 0.2248913,
  0.1904763, 0.2188449, 0.2954362, 0.3895774, 0.4191012, 0.2324064, 
    0.1984578, 0.2304615, 0.2598507, 0.2420469, 0.2130013, 0.2121198, 
    0.1736501, 0.2784961, 0.3606317, 0.256192, 0.2779781, 0.2346446, 
    0.2765385, 0.2454074, 0.1663556, 0.2773986, 0.2802455, 0.2526931, 
    0.1279393, 0.146036, 0.090216, 0.1072355, 0.1381177,
  0.1341227, 0.1684354, 0.2310709, 0.2241556, 0.2331677, 0.2058038, 0.254123, 
    0.2400284, 0.1721787, 0.2061796, 0.1970269, 0.1620311, 0.1590439, 
    0.113825, 0.1500938, 0.1329895, 0.1594531, 0.2411309, 0.3030529, 
    0.3028955, 0.2902941, 0.304781, 0.2387192, 0.149043, 0.1691437, 
    0.07936495, 0.05379794, 0.1323989, 0.2163091,
  0.1222565, 0.1170061, 0.1117558, 0.1065054, 0.1012551, 0.0960047, 
    0.09075434, 0.05865664, 0.05612886, 0.05360109, 0.05107331, 0.04854554, 
    0.04601776, 0.04348999, 0.04007557, 0.04671767, 0.05335977, 0.06000187, 
    0.06664397, 0.07328607, 0.07992817, 0.09886214, 0.09999818, 0.1011342, 
    0.1022702, 0.1034063, 0.1045423, 0.1056783, 0.1264568,
  0.02774042, 0.07342289, 0.05243254, 0.1131813, 0.09486811, 0.0883972, 
    0.06474633, 0.0560258, 0.05594335, 0.06837817, 0.08229741, 0.08445932, 
    0.0860155, 0.07079843, 0.04459367, 0.06967424, 0.08566198, 0.1097321, 
    0.08766949, 0.06474835, 0.1270775, 0.2201479, 0.1651324, 0.2068579, 
    0.1782137, 0.1012004, 0.1282152, 0.1184753, 0.05607907,
  0.2380551, 0.2486452, 0.2354105, 0.2842177, 0.2977932, 0.2210643, 0.211121, 
    0.2658297, 0.2495825, 0.3077008, 0.2499646, 0.1416144, 0.133969, 
    0.3282054, 0.2172547, 0.1838133, 0.2076693, 0.2203797, 0.2950016, 
    0.2343109, 0.3611182, 0.3820772, 0.3478541, 0.455937, 0.2669273, 
    0.1711447, 0.2422611, 0.2709613, 0.2510243,
  0.2456031, 0.2759803, 0.3044814, 0.4760338, 0.3179361, 0.2658844, 
    0.3833241, 0.3135099, 0.2293174, 0.2227128, 0.3274166, 0.3565802, 
    0.3986938, 0.2870985, 0.298699, 0.2361646, 0.2016587, 0.2182613, 
    0.191325, 0.2191876, 0.3176902, 0.2896663, 0.2645859, 0.3084238, 
    0.2391258, 0.2381794, 0.2585367, 0.2131056, 0.2470539,
  0.1438802, 0.1804622, 0.2219297, 0.3101234, 0.1796401, 0.1925591, 
    0.2386781, 0.2282873, 0.2201726, 0.2133512, 0.2358877, 0.2431259, 
    0.168621, 0.1967453, 0.1209997, 0.131518, 0.1371377, 0.1662995, 
    0.1416832, 0.1512021, 0.1670037, 0.1600353, 0.1858062, 0.111837, 
    0.07292573, 0.08988925, 0.1098335, 0.1368074, 0.1407759,
  0.0960763, 0.0832089, 0.04473285, 0.1146689, 0.1396271, 0.1068323, 
    0.1360305, 0.08150912, 0.1284518, 0.05441773, 0.05582162, 0.0283491, 
    0.05455723, 0.1192146, 0.1181401, 0.1508763, 0.10075, 0.1269994, 
    0.08082327, 0.1319661, 0.1737646, 0.1064844, 0.05559326, 0.01968541, 
    0.09547532, 0.1969414, 0.1003935, 0.1057894, 0.1510769,
  0.006193973, 9.391944e-06, 0.04325869, 0.1000186, 0.03529753, 0.03123367, 
    0.02916255, 0.003013142, 0.01545358, 3.185631e-06, 0.002412165, 
    0.001969988, 0.02106991, 0.01977129, 0.04652091, 0.04936818, 0.09485021, 
    0.06724224, 0.06127958, 0.0964537, 0.1017568, 0.03861302, 3.977297e-05, 
    1.801613e-07, 0.03840818, 0.06054827, 0.1038873, 0.08661351, 0.006116194,
  8.092138e-07, 0.004905929, 0.03434353, 0.0001291964, 0.002436238, 
    0.0005406614, 0.004995508, -1.878528e-05, -2.436672e-07, 8.474388e-08, 
    0.0002516965, 0.0003737859, 0.01963971, 0.0811694, 0.06041009, 
    0.06574652, 0.09053645, 0.03830603, 0.1070054, 0.06406871, 0.001654786, 
    -4.645001e-06, 2.053892e-08, -3.017361e-05, 0.07234084, 0.1831268, 
    0.1092023, 6.863565e-05, 9.902724e-06,
  0.006210579, 0.07573115, 0.06031934, 0.08283222, 0.08529335, 0.06837974, 
    0.04601019, 0.04178202, 0.00355683, 0.001761732, 0.01964456, 0.01146999, 
    0.04872936, 0.04771062, 0.06832993, 0.08071209, 0.04527028, 0.02658378, 
    0.004497977, 0.003214461, 7.404952e-08, 1.360009e-06, 2.731492e-05, 
    0.03890844, 0.08176459, 0.1457792, 0.01360917, 7.027667e-07, 1.751834e-07,
  0.1899064, 0.3348518, 0.07962551, 0.1070741, 0.03973204, 0.0110064, 
    0.03799575, 0.01935431, 0.07267188, 0.1326586, 0.06909809, 0.04561728, 
    0.03387339, 0.01369686, 0.005375961, 0.002914474, 8.988553e-06, 
    0.0002556002, -1.065971e-05, 1.912487e-05, 0.01680275, 0.0199947, 
    0.02117776, 0.09583981, 0.1503291, 0.002547241, 0.08315404, 0.03108096, 
    0.03672715,
  0.001585403, 0.001982733, 0.02943246, 0.09289239, 0.03226904, 0.00891128, 
    0.02009828, 0.05895355, 0.1005658, 0.02976266, 0.05540492, 0.06515657, 
    0.08118609, 0.09586932, 0.07713472, 0.05728396, 0.04166314, 0.08571775, 
    0.1500521, 0.1247913, 0.1774553, 0.04456626, 0.1171085, 0.0776448, 
    0.03792315, 0.04840553, 0.03538712, 0.002962271, 0.0008370655,
  2.011601e-05, 7.391674e-07, 0.0008513725, 0.01733807, 0.0334713, 
    0.0003819644, 0.01633528, 0.01964309, 0.0352876, 0.03363549, 0.02705536, 
    0.02840392, 0.0393492, 0.1048805, 0.03301581, 0.05185495, 0.04246531, 
    0.02293051, 0.008750392, 0.001105098, 0.03081238, 0.1053216, 0.006126371, 
    0.1061211, 0.04528654, 0.08293153, 0.03089382, 0.02295576, -2.661356e-05,
  0.001852379, 0.005436526, 0.01683537, 0.02468155, 0.1225455, 0.00366348, 
    0.02008226, 0.1347175, 0.2263856, 0.07391053, 0.01060893, 0.103181, 
    0.07504673, 0.1195535, 0.1537313, 0.07249393, 0.0482863, 0.06638376, 
    0.005848273, 0.00434467, 0.0311215, 0.09982602, 0.1082824, 0.06673985, 
    0.05164966, 0.123059, 0.07550083, 0.01929332, 0.05747438,
  0.05354584, 0.1118607, 0.03690975, 0.1222576, 0.02284755, 0.0185807, 
    0.100689, 0.02549461, 0.01433677, 0.009233519, 0.120159, 0.1018678, 
    0.1199037, 0.09394952, 0.1563501, 0.1676171, 0.2088142, 0.1689196, 
    0.1268811, 0.0602963, 0.0831755, 0.03034905, 0.1228326, 0.1666571, 
    0.164115, 0.1501741, 0.1377098, 0.1702701, 0.1319185,
  0.2404473, 0.1297962, 0.2391375, 0.1705117, 0.1562741, 0.1038184, 
    0.08927844, 0.19804, 0.09759105, 0.1539506, 0.1485283, 0.08432656, 
    0.1682109, 0.2367299, 0.2315325, 0.1405987, 0.1516819, 0.1845313, 
    0.2455457, 0.2566238, 0.1796743, 0.1598254, 0.231538, 0.4319043, 
    0.2248509, 0.2226834, 0.1717422, 0.2257767, 0.2115271,
  0.2424681, 0.3597241, 0.3251423, 0.3427573, 0.4111638, 0.3370935, 
    0.3487895, 0.4026597, 0.4554904, 0.3632328, 0.2912267, 0.1349927, 
    0.1685334, 0.1817039, 0.1679396, 0.1819365, 0.252885, 0.3145438, 
    0.2592917, 0.2671444, 0.248968, 0.3216107, 0.4663061, 0.3599135, 
    0.2915048, 0.2800521, 0.1915665, 0.2358499, 0.2362747,
  0.2348175, 0.2673441, 0.3438864, 0.3833617, 0.4507723, 0.2324538, 
    0.2047646, 0.3021866, 0.2866348, 0.2585632, 0.2391763, 0.2184711, 
    0.1679442, 0.2561426, 0.33995, 0.218298, 0.2774091, 0.2398122, 0.2279584, 
    0.250866, 0.1965066, 0.3203503, 0.2509341, 0.2501447, 0.1264217, 
    0.184674, 0.09835291, 0.102294, 0.1350205,
  0.1524399, 0.2042586, 0.272076, 0.2620557, 0.2463679, 0.2281621, 0.2562078, 
    0.2570188, 0.1885215, 0.2018402, 0.1956768, 0.1465748, 0.1442723, 
    0.1138076, 0.1451286, 0.1460167, 0.1612492, 0.2547457, 0.373138, 
    0.4029633, 0.3428952, 0.3154032, 0.280439, 0.1611025, 0.184075, 
    0.1441251, 0.08104779, 0.1370462, 0.2174968,
  0.1194098, 0.1170025, 0.1145953, 0.1121881, 0.1097808, 0.1073736, 
    0.1049664, 0.1044088, 0.1013008, 0.09819283, 0.09508482, 0.09197681, 
    0.0888688, 0.08576079, 0.09112316, 0.09702349, 0.1029238, 0.1088241, 
    0.1147245, 0.1206248, 0.1265251, 0.1238118, 0.1234267, 0.1230416, 
    0.1226565, 0.1222714, 0.1218863, 0.1215012, 0.1213355,
  0.02739816, 0.08381601, 0.055105, 0.127203, 0.09289663, 0.1077588, 
    0.0902291, 0.07884832, 0.06169525, 0.0934343, 0.08304182, 0.08404589, 
    0.101288, 0.07328848, 0.06273138, 0.07034101, 0.07195608, 0.09436719, 
    0.09443433, 0.05864207, 0.1328455, 0.2202306, 0.2120356, 0.2281283, 
    0.245993, 0.181562, 0.1376615, 0.1055081, 0.05950882,
  0.2150936, 0.2241228, 0.2150263, 0.2646244, 0.2953944, 0.2559888, 0.168471, 
    0.2578926, 0.2363216, 0.3252968, 0.2492676, 0.140089, 0.1755085, 
    0.3002414, 0.1574139, 0.1946713, 0.191815, 0.2084217, 0.2998023, 
    0.2579876, 0.2510328, 0.3487569, 0.3057977, 0.45045, 0.2350959, 
    0.1960068, 0.324708, 0.3716992, 0.2946412,
  0.2678669, 0.3236526, 0.3688117, 0.4316668, 0.3686836, 0.2673889, 
    0.4298676, 0.2453779, 0.2171601, 0.2562277, 0.3398216, 0.3720139, 
    0.3785445, 0.2900886, 0.2975263, 0.2468801, 0.2617418, 0.267181, 
    0.2009271, 0.2460316, 0.3322488, 0.290222, 0.2845019, 0.3450643, 
    0.2548255, 0.2265656, 0.249182, 0.2137941, 0.2785342,
  0.1484743, 0.2156941, 0.2448714, 0.3284775, 0.2039669, 0.1703699, 
    0.2271429, 0.2426616, 0.2341724, 0.2376519, 0.2773816, 0.2156541, 
    0.175154, 0.1962347, 0.1100785, 0.1369132, 0.1714439, 0.1794647, 
    0.1684856, 0.1823335, 0.186001, 0.2003502, 0.2266596, 0.114354, 
    0.05374373, 0.08856659, 0.1196621, 0.1552086, 0.1414168,
  0.1113324, 0.1006164, 0.06644027, 0.1331401, 0.1543744, 0.1189628, 
    0.1531382, 0.1158445, 0.1265828, 0.05353199, 0.05973251, 0.04432458, 
    0.06175973, 0.1246744, 0.1528823, 0.1459177, 0.1457549, 0.1344019, 
    0.09990027, 0.1413872, 0.1784994, 0.1203877, 0.07335057, 0.02644018, 
    0.08656495, 0.205346, 0.1029729, 0.1227282, 0.1793432,
  0.007650028, 0.0003300166, 0.02114675, 0.05985891, 0.0421783, 0.03614617, 
    0.03459787, 0.007363089, 0.02420424, 1.907041e-06, 0.0004191264, 
    0.004045466, 0.01736665, 0.02710532, 0.04223281, 0.0580757, 0.1093238, 
    0.06988811, 0.05883917, 0.08190932, 0.1026446, 0.04960051, 0.0005528321, 
    6.244376e-07, 0.0293038, 0.05992541, 0.09934638, 0.09180587, 0.01265072,
  -5.704744e-09, 0.001983336, 0.01513167, 0.0002101868, 0.007716755, 
    0.003058465, 0.01175108, 0.0008562895, -1.597214e-05, 9.701382e-08, 
    4.051151e-05, 5.796831e-05, 0.02115915, 0.09998997, 0.06612258, 
    0.0592711, 0.09061869, 0.04025896, 0.1025495, 0.07390735, 0.008905104, 
    -2.240155e-05, 1.492227e-08, -1.913034e-05, 0.06339581, 0.1690416, 
    0.1147914, 0.001760392, 4.67676e-05,
  0.004998802, 0.07136729, 0.04142978, 0.09391323, 0.08963195, 0.0723964, 
    0.05161901, 0.0557804, 0.006637202, 0.001197023, 0.007458481, 0.00979147, 
    0.04925863, 0.04394558, 0.06493713, 0.06435307, 0.05504117, 0.04210131, 
    0.01720639, 0.006515697, -5.459862e-06, 2.603219e-07, 1.136564e-05, 
    0.0349051, 0.06750023, 0.08809198, 0.01376158, 3.66676e-06, 4.441031e-07,
  0.1311664, 0.3111572, 0.06906845, 0.1455869, 0.03184874, 0.01265466, 
    0.04038936, 0.02031362, 0.08792026, 0.1305092, 0.04747339, 0.03967561, 
    0.02648003, 0.01400151, 0.006354629, 0.005991719, 8.833732e-05, 
    7.947829e-05, -1.19059e-05, 0.001246053, 0.01388445, 0.02338774, 
    0.02152263, 0.08239855, 0.1374026, 0.004178312, 0.08203737, 0.05476746, 
    0.03886884,
  0.0005143778, 0.0008768498, 0.005372741, 0.1172891, 0.03854739, 0.01779773, 
    0.03203669, 0.07060348, 0.1125832, 0.02545357, 0.0656823, 0.05801234, 
    0.07478997, 0.09099934, 0.06869291, 0.05463885, 0.04053183, 0.08973022, 
    0.1570238, 0.1264811, 0.1814297, 0.04921446, 0.1389393, 0.08665442, 
    0.04138502, 0.04378641, 0.03157693, 0.0004281822, 0.0003145972,
  1.437759e-05, 4.692234e-07, 0.01827333, 0.01951734, 0.03346888, 
    0.002437865, 0.01769594, 0.02080732, 0.03823796, 0.04161246, 0.03640568, 
    0.02793484, 0.04659098, 0.09868535, 0.03687885, 0.04267072, 0.04620137, 
    0.0215684, 0.01415563, 0.007441932, 0.02765499, 0.1323854, 0.02057407, 
    0.09483222, 0.05234215, 0.0785531, 0.02387198, 0.01661009, -4.597262e-07,
  0.0003059314, 0.005385902, 0.01796263, 0.02526172, 0.1254296, 0.00203007, 
    0.01214686, 0.1216279, 0.1967155, 0.07484831, 0.03078157, 0.1016937, 
    0.06979468, 0.1117117, 0.1683362, 0.09301275, 0.0636178, 0.08038653, 
    0.0099404, 0.005743853, 0.02471272, 0.08815432, 0.1226392, 0.06385175, 
    0.05660108, 0.1360554, 0.07178632, 0.04815513, 0.03709527,
  0.04569163, 0.1162316, 0.04655055, 0.106896, 0.01453276, 0.018925, 
    0.09715687, 0.01393951, 0.009342131, 0.00829933, 0.1240064, 0.1001422, 
    0.1345717, 0.1087095, 0.1773662, 0.1680377, 0.2147604, 0.190582, 
    0.1342838, 0.0678536, 0.07948823, 0.0264101, 0.1115522, 0.1666601, 
    0.1735138, 0.1544906, 0.1606019, 0.1837, 0.1436375,
  0.2402028, 0.134995, 0.2514313, 0.206445, 0.1926866, 0.07972912, 
    0.09777243, 0.2171883, 0.08585058, 0.1398968, 0.137893, 0.09120011, 
    0.196126, 0.2688466, 0.2557692, 0.1812232, 0.164961, 0.1828724, 0.242355, 
    0.2660089, 0.1560635, 0.155069, 0.2675093, 0.4236402, 0.2485987, 
    0.2381604, 0.1849808, 0.2613417, 0.2056109,
  0.2295662, 0.3743916, 0.2734185, 0.4088396, 0.3959017, 0.3118435, 0.323393, 
    0.3869242, 0.4089434, 0.3526042, 0.3038538, 0.1485294, 0.1671038, 
    0.1698884, 0.180102, 0.2392541, 0.2559487, 0.2974337, 0.2751487, 
    0.256672, 0.2477008, 0.3303438, 0.4090804, 0.3552606, 0.2629378, 
    0.2646144, 0.2245271, 0.2427124, 0.2256894,
  0.2738362, 0.2638887, 0.3407604, 0.349907, 0.4421449, 0.224286, 0.1823329, 
    0.3490734, 0.3133357, 0.2790984, 0.2833562, 0.2089629, 0.1633625, 
    0.2507378, 0.3288678, 0.2158346, 0.2902105, 0.263337, 0.2076898, 
    0.2480356, 0.1932085, 0.2302354, 0.2015149, 0.2258935, 0.1399924, 
    0.2255488, 0.1084914, 0.1311728, 0.1679937,
  0.1707373, 0.2186752, 0.2823791, 0.2506472, 0.258708, 0.2614085, 0.2454437, 
    0.2485405, 0.203633, 0.2190563, 0.1889694, 0.1379043, 0.1304696, 
    0.1119049, 0.1538302, 0.1327659, 0.1616334, 0.2461651, 0.3491917, 
    0.3388154, 0.3173188, 0.3198994, 0.2793251, 0.2111213, 0.2159077, 
    0.1746227, 0.08649266, 0.1400817, 0.232549,
  0.1272156, 0.125129, 0.1230423, 0.1209557, 0.118869, 0.1167824, 0.1146957, 
    0.1223653, 0.1185689, 0.1147726, 0.1109762, 0.1071798, 0.1033834, 
    0.09958705, 0.09867837, 0.1051499, 0.1116213, 0.1180928, 0.1245643, 
    0.1310358, 0.1375073, 0.1331786, 0.1325902, 0.1320017, 0.1314133, 
    0.1308248, 0.1302363, 0.1296479, 0.1288849,
  0.03114708, 0.08020636, 0.06092149, 0.120553, 0.09835419, 0.1303844, 
    0.09722545, 0.07920668, 0.06695497, 0.126033, 0.0771331, 0.08959151, 
    0.1043361, 0.06759194, 0.06081874, 0.07046209, 0.0723139, 0.08289383, 
    0.07932461, 0.05395007, 0.1195931, 0.212124, 0.2567227, 0.1887006, 
    0.2027766, 0.2246905, 0.07637979, 0.09053306, 0.06423847,
  0.23374, 0.2455349, 0.2290642, 0.2442826, 0.3086951, 0.2907915, 0.1853487, 
    0.2437394, 0.247664, 0.3472877, 0.2370214, 0.1261514, 0.1891172, 
    0.2577819, 0.1662585, 0.1558587, 0.1788694, 0.1820603, 0.2741089, 
    0.2525816, 0.2659453, 0.3685585, 0.3195099, 0.4282953, 0.2203475, 
    0.2171687, 0.3608164, 0.3071584, 0.2948208,
  0.3196544, 0.3293115, 0.40676, 0.3785826, 0.3642265, 0.3765928, 0.3836581, 
    0.2291263, 0.2275069, 0.2243102, 0.3452913, 0.3705584, 0.3220134, 
    0.2676956, 0.3056721, 0.2460221, 0.2512941, 0.2346788, 0.2165939, 
    0.2525072, 0.3196172, 0.295348, 0.3018706, 0.33769, 0.2394532, 0.2436051, 
    0.301081, 0.2516187, 0.2722803,
  0.1656608, 0.2388244, 0.2550235, 0.3169062, 0.2051356, 0.1955686, 
    0.2270623, 0.2437126, 0.2614878, 0.2738458, 0.2823408, 0.2239089, 
    0.1880261, 0.2026016, 0.1152867, 0.1473465, 0.1811523, 0.1756474, 
    0.1811919, 0.215031, 0.2195789, 0.2561022, 0.2220646, 0.1102481, 
    0.04116056, 0.08656768, 0.1293617, 0.1423958, 0.1536154,
  0.1011754, 0.1300338, 0.09545326, 0.1459143, 0.1663196, 0.1599724, 
    0.1879837, 0.1584325, 0.147411, 0.05348669, 0.05196984, 0.06854043, 
    0.06979634, 0.1408305, 0.171289, 0.1666083, 0.1597939, 0.149325, 
    0.1090042, 0.1230946, 0.1722624, 0.1245108, 0.08990149, 0.02993531, 
    0.06756122, 0.2165819, 0.1048975, 0.1321202, 0.1567851,
  0.01528866, 0.002004739, 0.01772604, 0.04227612, 0.07502805, 0.05558402, 
    0.0398953, 0.02059996, 0.02569241, 6.078474e-07, 0.000155839, 
    0.004011898, 0.01362767, 0.02987466, 0.04316722, 0.04297654, 0.1079544, 
    0.07028036, 0.06794506, 0.09558564, 0.09432328, 0.05279683, 0.01004326, 
    2.843999e-07, 0.02483295, 0.05618415, 0.08569551, 0.1056289, 0.03274108,
  -1.578982e-05, 0.0003690242, 0.008081191, 5.825143e-05, 0.0195807, 
    0.009866188, 0.01190272, 0.01610521, 0.0002261222, 1.433715e-07, 
    3.905082e-06, 6.863105e-06, 0.01813852, 0.07938996, 0.07178697, 
    0.05702196, 0.08436053, 0.04062365, 0.08616745, 0.08941098, 0.03252918, 
    0.0006305975, 2.964108e-08, -9.786704e-06, 0.06265547, 0.1713163, 
    0.106964, 0.04176023, 0.002494884,
  0.0007966438, 0.05987159, 0.03423985, 0.102444, 0.09096275, 0.07427329, 
    0.05150077, 0.06833322, 0.009290368, 0.001480669, 0.004951966, 
    0.00933819, 0.05213324, 0.03738281, 0.06241689, 0.05014992, 0.05321271, 
    0.04237195, 0.03276009, 0.01963411, 0.0004225023, 6.704392e-07, 
    6.149036e-06, 0.03460026, 0.05792875, 0.04865727, 0.02106989, 
    2.447049e-05, 1.388426e-06,
  0.09275065, 0.2946326, 0.06898114, 0.1883089, 0.0290333, 0.0144002, 
    0.03855206, 0.02049887, 0.1050825, 0.1268739, 0.03071594, 0.02507023, 
    0.0215269, 0.01408143, 0.009056994, 0.009843844, 0.000780142, 0.00105992, 
    -6.5279e-06, 0.01930629, 0.01019309, 0.01767823, 0.01590924, 0.0734227, 
    0.1023811, 0.00582343, 0.08408253, 0.07591614, 0.04970145,
  0.0001836316, 4.416287e-05, 0.002901947, 0.127579, 0.04854861, 0.02115002, 
    0.05079171, 0.06244315, 0.08682572, 0.02801877, 0.0738074, 0.04591443, 
    0.06766879, 0.07618921, 0.06801049, 0.05134298, 0.04320415, 0.09160336, 
    0.164431, 0.1238409, 0.1734542, 0.04201258, 0.1641507, 0.08376254, 
    0.03961417, 0.0393388, 0.03002024, 0.0002521136, 0.000181595,
  5.540877e-06, 2.139153e-07, 0.01188632, 0.02156834, 0.02321174, 0.01163251, 
    0.01983431, 0.01843676, 0.06798577, 0.07472067, 0.04933486, 0.03048152, 
    0.0596657, 0.09884342, 0.03974281, 0.04558194, 0.06857247, 0.02720541, 
    0.01644341, 0.01102205, 0.02405972, 0.1747278, 0.03566634, 0.0921412, 
    0.05596471, 0.06525577, 0.02013277, 0.01200424, 4.770971e-06,
  2.478031e-05, 0.008313328, 0.01895473, 0.02192314, 0.1113587, 0.007997471, 
    0.005822523, 0.09616105, 0.1837967, 0.04832661, 0.06525861, 0.1035982, 
    0.07390123, 0.09902897, 0.1607186, 0.09921864, 0.08707415, 0.09010306, 
    0.01201457, 0.006343561, 0.01793607, 0.06086706, 0.1132503, 0.06642903, 
    0.0659854, 0.1239249, 0.05699423, 0.07222713, 0.01719105,
  0.03877667, 0.1128583, 0.05852851, 0.1029553, 0.009348528, 0.02828719, 
    0.08721209, 0.001401562, 0.005383696, 0.01513499, 0.1263845, 0.110738, 
    0.147339, 0.1513147, 0.2175816, 0.1833807, 0.2168985, 0.2163532, 
    0.1406882, 0.06938661, 0.06601663, 0.02702498, 0.09219671, 0.1577049, 
    0.1853923, 0.142566, 0.1742895, 0.220803, 0.165241,
  0.2594101, 0.1204903, 0.2597773, 0.2172355, 0.2037812, 0.07751051, 
    0.07705548, 0.2361405, 0.07572604, 0.1298369, 0.1235522, 0.09718905, 
    0.2365447, 0.3135613, 0.2574708, 0.2128382, 0.1828099, 0.1938614, 
    0.2450419, 0.2790453, 0.1518305, 0.1728884, 0.2667558, 0.4034171, 
    0.2464405, 0.2304471, 0.2084997, 0.2778181, 0.2243904,
  0.2346454, 0.3581448, 0.3083932, 0.4302606, 0.3309472, 0.3230714, 
    0.3102579, 0.356772, 0.3903767, 0.3521752, 0.3226099, 0.1756161, 
    0.1574317, 0.2105659, 0.2155144, 0.2572129, 0.2808602, 0.3171483, 
    0.2841884, 0.2352443, 0.2850001, 0.3120908, 0.4426493, 0.4068879, 
    0.2748275, 0.2364831, 0.2565957, 0.2750016, 0.2521778,
  0.2952574, 0.2707208, 0.3632419, 0.3317675, 0.4299868, 0.2394451, 
    0.1897439, 0.3014788, 0.3050343, 0.3453785, 0.3247664, 0.2133692, 
    0.1663246, 0.283507, 0.3400616, 0.2068447, 0.2811055, 0.288219, 0.182586, 
    0.3102662, 0.1727924, 0.1785976, 0.2085537, 0.1838351, 0.1176093, 
    0.2595752, 0.1160892, 0.1566764, 0.2455728,
  0.2013038, 0.2405825, 0.3026279, 0.2654548, 0.2580631, 0.2907651, 
    0.2478526, 0.2381412, 0.2233103, 0.221131, 0.1840963, 0.1466685, 
    0.1402068, 0.1270754, 0.1458972, 0.1226039, 0.1837472, 0.2734006, 
    0.360387, 0.4491473, 0.3918971, 0.269297, 0.224587, 0.2336661, 0.243958, 
    0.206877, 0.09094582, 0.1467755, 0.2570782,
  0.1474065, 0.1454343, 0.1434621, 0.1414899, 0.1395177, 0.1375455, 
    0.1355733, 0.1391989, 0.134971, 0.1307431, 0.1265152, 0.1222873, 
    0.1180595, 0.1138316, 0.1100528, 0.1172644, 0.1244761, 0.1316878, 
    0.1388994, 0.1461111, 0.1533228, 0.1460105, 0.1449989, 0.1439873, 
    0.1429757, 0.1419641, 0.1409525, 0.1399409, 0.1489843,
  0.04245842, 0.07979512, 0.07252863, 0.1281791, 0.1350376, 0.1810837, 
    0.1557955, 0.09430139, 0.09133627, 0.1356137, 0.07579324, 0.09469955, 
    0.1032645, 0.06433763, 0.09135246, 0.1055466, 0.08441751, 0.05805849, 
    0.0607439, 0.0562952, 0.1117449, 0.2115187, 0.2909361, 0.1977399, 
    0.2584827, 0.1718803, 0.06957401, 0.07882144, 0.07596405,
  0.2330677, 0.2620808, 0.2421497, 0.1954727, 0.308796, 0.3062466, 0.1704384, 
    0.2153751, 0.2557675, 0.325984, 0.2276084, 0.09366689, 0.1610152, 
    0.2807469, 0.2599983, 0.1900167, 0.2218162, 0.1940726, 0.2918733, 0.2705, 
    0.3446285, 0.3957123, 0.319516, 0.4290535, 0.2190607, 0.2989442, 
    0.3894641, 0.2472345, 0.2489983,
  0.3362288, 0.3244083, 0.4145598, 0.4270686, 0.31272, 0.305009, 0.4312296, 
    0.2683965, 0.3467063, 0.3056413, 0.3982226, 0.3487227, 0.3355115, 
    0.3402479, 0.2971763, 0.267644, 0.2687983, 0.3006705, 0.2348577, 
    0.3162649, 0.3440603, 0.3258796, 0.3138991, 0.3494951, 0.2334592, 
    0.2554285, 0.3250638, 0.2852442, 0.3028232,
  0.1967656, 0.2740009, 0.2822792, 0.3136361, 0.23104, 0.2606289, 0.2822006, 
    0.2939433, 0.3001772, 0.2599169, 0.2994598, 0.269334, 0.2503093, 
    0.2053545, 0.123982, 0.1694767, 0.2149921, 0.2140996, 0.2127686, 
    0.2379977, 0.2481082, 0.2392071, 0.2095435, 0.1203558, 0.0344143, 
    0.08911226, 0.1283939, 0.1265554, 0.16213,
  0.1092781, 0.1738679, 0.1203474, 0.1834823, 0.2130001, 0.2296775, 
    0.2407583, 0.1994988, 0.1920916, 0.09291925, 0.06838542, 0.07677961, 
    0.07193696, 0.1550176, 0.1991567, 0.1736445, 0.2224733, 0.1466386, 
    0.1487284, 0.1316691, 0.2093872, 0.1567496, 0.1157385, 0.03731428, 
    0.0753779, 0.2554962, 0.1060956, 0.158177, 0.1561131,
  0.05061866, 0.01908627, 0.02266174, 0.06984144, 0.09706736, 0.07960859, 
    0.04482215, 0.03599729, 0.03283873, 0.0003554049, 0.000155354, 
    0.0005085737, 0.01202953, 0.03191205, 0.05116517, 0.04744586, 0.107745, 
    0.08785397, 0.06874874, 0.106915, 0.1011559, 0.07401364, 0.01187062, 
    4.422568e-07, 0.0145643, 0.07515638, 0.09049056, 0.1320888, 0.06734002,
  0.001047143, 5.961092e-05, 0.003182585, 0.0001031916, 0.0407238, 
    0.02453258, 0.02251831, 0.03796329, 0.001088014, 1.247912e-07, 
    -1.107476e-06, -3.386291e-07, 0.02489386, 0.0562474, 0.07475687, 
    0.06500468, 0.05127048, 0.03874046, 0.06264415, 0.08784803, 0.05283962, 
    0.01677359, 1.289991e-06, -7.06224e-06, 0.07886872, 0.1848512, 
    0.09431984, 0.128948, 0.03829296,
  5.364002e-05, 0.04060768, 0.02952558, 0.1073368, 0.0746192, 0.0719079, 
    0.04577519, 0.0742887, 0.01333268, 0.003099761, 0.004641218, 0.009775297, 
    0.05673156, 0.03708222, 0.05901337, 0.04189494, 0.0455612, 0.03863936, 
    0.03943021, 0.05184831, 0.01011036, 0.0002863779, 4.515093e-06, 
    0.03539353, 0.04809552, 0.02928625, 0.04124376, 0.001784699, 1.362915e-05,
  0.08697043, 0.2529262, 0.0682366, 0.2079925, 0.02909919, 0.01621999, 
    0.03402037, 0.02006368, 0.1151154, 0.1471304, 0.02828561, 0.0197777, 
    0.02144681, 0.0136222, 0.01237315, 0.01423023, 0.004514285, 0.00295753, 
    0.0003016075, 0.01143341, 0.0131612, 0.004909613, 0.0185428, 0.06317479, 
    0.07358644, 0.008895428, 0.07854968, 0.0743144, 0.05249091,
  6.090982e-05, 9.061923e-06, 0.0005425983, 0.1145899, 0.07133304, 
    0.02380896, 0.06536776, 0.05665193, 0.0771313, 0.02939795, 0.06720343, 
    0.0346218, 0.05882409, 0.06543776, 0.06260248, 0.04972101, 0.05872358, 
    0.08929663, 0.1685578, 0.1110644, 0.1516788, 0.03867671, 0.1593081, 
    0.09188122, 0.03656248, 0.03687065, 0.02876626, 0.0003393516, 0.0001828775,
  1.90131e-06, 5.74437e-08, 7.589115e-05, 0.02107995, 0.01452965, 0.06570969, 
    0.02208072, 0.01831151, 0.1050569, 0.07777374, 0.08520224, 0.03383363, 
    0.06306408, 0.1071796, 0.04783311, 0.07853253, 0.0521412, 0.03703716, 
    0.05096509, 0.008375823, 0.02167059, 0.2123234, 0.06046812, 0.0968286, 
    0.05494863, 0.04977299, 0.02227187, 0.002547334, 2.8478e-06,
  7.802412e-06, 0.02213522, 0.03960752, 0.02750926, 0.1095437, 0.000898275, 
    0.004207716, 0.07296859, 0.1858656, 0.02035714, 0.1201202, 0.1371599, 
    0.09837945, 0.09890635, 0.1802448, 0.1636479, 0.1300756, 0.1022327, 
    0.02260395, 0.006238485, 0.01561307, 0.06368569, 0.1198081, 0.0784443, 
    0.08965357, 0.1155786, 0.0557296, 0.09254888, 0.01055367,
  0.03160305, 0.1062615, 0.06850868, 0.1046861, 0.0194987, 0.008513947, 
    0.08642802, 0.0005804688, 0.002255577, 0.01433797, 0.1221441, 0.1403656, 
    0.1945792, 0.21052, 0.2897309, 0.2038737, 0.2507422, 0.247502, 0.1520358, 
    0.0810002, 0.06289513, 0.03779596, 0.1157845, 0.1682402, 0.214181, 
    0.1668584, 0.1920695, 0.263516, 0.1840938,
  0.2777224, 0.1342201, 0.2691334, 0.2263845, 0.1676617, 0.06585748, 
    0.08892114, 0.2595935, 0.07880246, 0.1463286, 0.1195958, 0.1047316, 
    0.2836165, 0.3579807, 0.2641156, 0.23027, 0.2043889, 0.2490975, 
    0.2583733, 0.3024895, 0.1635993, 0.2321646, 0.2944554, 0.4115195, 
    0.2891073, 0.2422308, 0.2401619, 0.3124282, 0.239758,
  0.222351, 0.3479211, 0.3348254, 0.388427, 0.3648364, 0.2784784, 0.3213745, 
    0.4000395, 0.4379789, 0.4127655, 0.4165899, 0.2166593, 0.1430073, 
    0.2510241, 0.3688958, 0.2786544, 0.3035966, 0.3019951, 0.302779, 
    0.250916, 0.3478673, 0.3033067, 0.4619421, 0.4270187, 0.3705186, 
    0.2151662, 0.2797663, 0.3023002, 0.2484335,
  0.2595683, 0.2614719, 0.3915575, 0.3858172, 0.4574845, 0.2530344, 
    0.2432764, 0.298362, 0.3017483, 0.3472725, 0.3492617, 0.2248175, 
    0.2171603, 0.3317963, 0.3797354, 0.235939, 0.2871063, 0.3534793, 
    0.2033689, 0.3789047, 0.2362929, 0.1758497, 0.1996852, 0.182313, 
    0.108632, 0.2647523, 0.1178687, 0.1680469, 0.3322865,
  0.2319258, 0.2745499, 0.2833222, 0.294044, 0.2537478, 0.2664128, 0.2143883, 
    0.2287416, 0.2500876, 0.259316, 0.2162714, 0.1466438, 0.1595042, 
    0.1748692, 0.2208793, 0.1728488, 0.294889, 0.2849629, 0.4166034, 
    0.4579858, 0.3291449, 0.3045498, 0.185547, 0.2638496, 0.2780113, 
    0.2548174, 0.1098379, 0.1606326, 0.2885329,
  0.1521569, 0.1505543, 0.1489517, 0.147349, 0.1457464, 0.1441438, 0.1425412, 
    0.1596004, 0.155659, 0.1517176, 0.1477762, 0.1438348, 0.1398934, 
    0.1359521, 0.131679, 0.1391655, 0.1466521, 0.1541386, 0.1616251, 
    0.1691116, 0.1765981, 0.1623636, 0.1604211, 0.1584786, 0.1565361, 
    0.1545936, 0.1526511, 0.1507086, 0.153439,
  0.05448104, 0.07823371, 0.08407517, 0.1425514, 0.1613826, 0.2252872, 
    0.1874029, 0.1078086, 0.1215342, 0.1428491, 0.0815879, 0.09446125, 
    0.1190912, 0.04895883, 0.06724662, 0.2069418, 0.1958911, 0.1118817, 
    0.05791043, 0.0465344, 0.116339, 0.2050286, 0.3212503, 0.3532622, 
    0.26678, 0.1772057, 0.09225591, 0.05501755, 0.08138749,
  0.2652793, 0.2578764, 0.2398157, 0.1471252, 0.301384, 0.3139065, 0.1390354, 
    0.2185733, 0.2588651, 0.3187372, 0.2153024, 0.0802016, 0.1485059, 
    0.2720847, 0.2907271, 0.2300213, 0.2523651, 0.2044192, 0.3213035, 
    0.2481704, 0.2777543, 0.4104565, 0.3144749, 0.4483352, 0.218405, 
    0.3024103, 0.4405645, 0.3034699, 0.313757,
  0.3861384, 0.3659057, 0.4248647, 0.4325051, 0.420459, 0.337067, 0.4915985, 
    0.3584969, 0.4373852, 0.3675991, 0.4291393, 0.4425295, 0.4913707, 
    0.4377481, 0.334897, 0.3548258, 0.3442137, 0.3553481, 0.2706515, 
    0.3629509, 0.343895, 0.3512118, 0.3280001, 0.371551, 0.2574317, 
    0.3072763, 0.3378622, 0.3129762, 0.3370399,
  0.2391731, 0.3260583, 0.3264346, 0.3667649, 0.3406853, 0.3148558, 0.36623, 
    0.3820717, 0.3461255, 0.3350163, 0.3338717, 0.2622749, 0.2669137, 
    0.2734404, 0.1446575, 0.2422101, 0.3697795, 0.2500797, 0.2481154, 
    0.303337, 0.2641768, 0.259358, 0.2491676, 0.1388542, 0.02975521, 
    0.0859552, 0.1400235, 0.1291842, 0.2324453,
  0.1819833, 0.2148959, 0.2001204, 0.2103747, 0.2930877, 0.2487126, 
    0.2544343, 0.2168854, 0.2211718, 0.1733187, 0.1031255, 0.1146234, 
    0.07531437, 0.1682636, 0.2259305, 0.2199744, 0.3245946, 0.2424863, 
    0.2009884, 0.1573006, 0.2871506, 0.2422861, 0.1885054, 0.04569467, 
    0.06115146, 0.2792194, 0.1231523, 0.1891422, 0.2380597,
  0.07409919, 0.02620651, 0.02722979, 0.07274564, 0.131407, 0.1788711, 
    0.08045834, 0.09941163, 0.05831877, 0.006606318, 4.117649e-06, 
    0.0001341943, 0.00983148, 0.04382339, 0.06999823, 0.0626476, 0.1371715, 
    0.1027893, 0.09174955, 0.1543916, 0.1018562, 0.1272851, 0.08097244, 
    1.057204e-06, 0.009297688, 0.07503304, 0.0980894, 0.1554189, 0.1446334,
  0.0528474, -7.18138e-05, 0.001443389, 0.002904114, 0.03925875, 0.0535537, 
    0.05860348, 0.03976129, 0.007985329, 8.910429e-08, -1.242521e-07, 
    -1.461766e-06, 0.02550965, 0.05271973, 0.06761758, 0.05950359, 
    0.06047351, 0.03959534, 0.05143755, 0.08126877, 0.1910085, 0.07066, 
    0.0001012723, 3.085893e-06, 0.08068243, 0.2107456, 0.08455967, 0.1397681, 
    0.3559434,
  0.0002451642, 0.0359799, 0.02596394, 0.113222, 0.05394323, 0.06721193, 
    0.04038043, 0.06044034, 0.02461281, 0.004599735, 0.007703998, 0.01254561, 
    0.05361898, 0.03678058, 0.05402967, 0.04941563, 0.04045148, 0.03824749, 
    0.03699437, 0.0503906, 0.1045012, 0.0105086, 0.0001923662, 0.03306079, 
    0.04191398, 0.01821238, 0.05164782, 0.03432361, 0.003818048,
  0.09190901, 0.2313584, 0.06213501, 0.2129677, 0.03258064, 0.02226566, 
    0.03221342, 0.02144898, 0.1237605, 0.1526372, 0.03116601, 0.02016666, 
    0.024139, 0.01647162, 0.01682901, 0.01939104, 0.01065023, 0.005964763, 
    0.007202453, 0.001722563, 0.02300173, 0.001260989, 0.01020942, 
    0.06263001, 0.05005256, 0.01733692, 0.06747788, 0.06569836, 0.06265592,
  4.093114e-05, 3.328293e-06, 0.0001634083, 0.07569043, 0.07528365, 
    0.02267967, 0.05662212, 0.05718658, 0.09629704, 0.03992459, 0.06022314, 
    0.03489815, 0.05015458, 0.05759117, 0.05603324, 0.04583225, 0.06352696, 
    0.08596398, 0.1657931, 0.09939651, 0.1351789, 0.04845976, 0.1558295, 
    0.1008503, 0.03708611, 0.03489826, 0.03394777, 0.000506184, 4.582543e-05,
  6.677167e-07, 1.468518e-08, 8.760482e-06, 0.02759288, 0.003667641, 
    0.07463156, 0.02492639, 0.0339492, 0.1202077, 0.1075483, 0.1229896, 
    0.05711986, 0.06276805, 0.1019959, 0.07328951, 0.06798097, 0.0483649, 
    0.04235403, 0.1103233, 0.05182134, 0.02728887, 0.2422015, 0.07738026, 
    0.09497033, 0.05205157, 0.04612127, 0.03674258, 0.001818335, 1.779597e-06,
  2.130972e-06, 0.02477477, 0.05623871, 0.02534238, 0.1128363, 7.600066e-05, 
    0.002829141, 0.05622884, 0.1794147, 0.004918796, 0.2007729, 0.1778706, 
    0.1234216, 0.1296429, 0.2052235, 0.2048699, 0.1396133, 0.1465181, 
    0.05503552, 0.02329694, 0.0200641, 0.07048766, 0.1420823, 0.1665235, 
    0.1287124, 0.1201926, 0.06036057, 0.1224431, 0.01465249,
  0.02266836, 0.09946555, 0.08385289, 0.1048967, 0.03369742, 0.0104716, 
    0.06634021, -0.0002233257, 0.0006033987, 0.01410586, 0.1146274, 
    0.3109147, 0.3376026, 0.3255272, 0.3157348, 0.2354949, 0.306044, 
    0.2371697, 0.1813665, 0.09025564, 0.05841312, 0.05785872, 0.1536741, 
    0.1742796, 0.2462031, 0.1957413, 0.2348449, 0.2682827, 0.2037636,
  0.2902476, 0.1841883, 0.2574653, 0.2402688, 0.1588549, 0.06764345, 
    0.106783, 0.2624343, 0.075538, 0.1478819, 0.1330062, 0.1068272, 
    0.3380414, 0.3708196, 0.2677121, 0.2196151, 0.2159818, 0.2827951, 
    0.2916687, 0.3281749, 0.1627744, 0.2834851, 0.332226, 0.47275, 0.3140225, 
    0.2970766, 0.2652381, 0.2877452, 0.2339679,
  0.2233204, 0.3687583, 0.3274192, 0.4025781, 0.4415684, 0.2851508, 
    0.3779151, 0.4195248, 0.4777853, 0.4841643, 0.4848364, 0.2817102, 
    0.1342706, 0.2514044, 0.4906317, 0.3146321, 0.3379172, 0.3102113, 
    0.3398573, 0.2659462, 0.4000835, 0.3223069, 0.5881739, 0.4559112, 
    0.3931001, 0.220636, 0.3232389, 0.3584287, 0.2559204,
  0.2519829, 0.2503772, 0.3865713, 0.4223847, 0.4783415, 0.2686574, 
    0.2797596, 0.3040714, 0.326537, 0.3687484, 0.3721293, 0.2479023, 
    0.2187884, 0.3500105, 0.3846745, 0.2486615, 0.3274772, 0.3731492, 
    0.2083164, 0.4214556, 0.2743293, 0.2236744, 0.2480651, 0.2036988, 
    0.1427373, 0.2727655, 0.1214548, 0.2188997, 0.3380274,
  0.2188489, 0.3061242, 0.3160746, 0.2652597, 0.2207772, 0.2789567, 
    0.2290342, 0.237553, 0.2782357, 0.2868074, 0.2471019, 0.1691487, 
    0.1640353, 0.2192427, 0.3008763, 0.2855028, 0.3527515, 0.3749554, 
    0.4537727, 0.4318605, 0.3171679, 0.2972034, 0.2100511, 0.2648145, 
    0.3192897, 0.3125101, 0.1121279, 0.1789552, 0.2957455,
  0.162397, 0.1620773, 0.1617576, 0.1614379, 0.1611182, 0.1607985, 0.1604788, 
    0.1834445, 0.1792567, 0.175069, 0.1708812, 0.1666935, 0.1625058, 
    0.158318, 0.1660247, 0.1740641, 0.1821036, 0.1901431, 0.1981826, 
    0.2062221, 0.2142616, 0.1839682, 0.1804362, 0.1769042, 0.1733721, 
    0.1698401, 0.166308, 0.162776, 0.1626528,
  0.05930302, 0.07474802, 0.09163346, 0.1537362, 0.1783323, 0.2380045, 
    0.2264332, 0.1234273, 0.1526391, 0.1561434, 0.09362803, 0.09035978, 
    0.1221262, 0.03722353, 0.1112523, 0.15412, 0.1897607, 0.09395782, 
    0.04887998, 0.02876394, 0.1261386, 0.1860376, 0.343789, 0.2943387, 
    0.2496454, 0.2013168, 0.1019878, 0.03927164, 0.07544729,
  0.2665395, 0.2601295, 0.1939873, 0.1204507, 0.2694932, 0.3361999, 
    0.1174109, 0.2289353, 0.2700478, 0.3088554, 0.2045141, 0.06979811, 
    0.1421742, 0.2513591, 0.2850461, 0.2624615, 0.2763421, 0.2946889, 
    0.3992369, 0.2566776, 0.2845638, 0.4219241, 0.3366659, 0.5172843, 
    0.2070278, 0.340424, 0.4758942, 0.3762201, 0.3858643,
  0.4691316, 0.4081674, 0.4497264, 0.4465411, 0.564693, 0.4193745, 0.4827472, 
    0.4264486, 0.4116363, 0.4082093, 0.4426356, 0.5405588, 0.4308419, 
    0.3950866, 0.3518121, 0.4086558, 0.4247658, 0.3817382, 0.3384799, 
    0.3641428, 0.4116063, 0.3441071, 0.3192896, 0.3728756, 0.3065142, 
    0.3174478, 0.4111756, 0.3528286, 0.3743785,
  0.2982926, 0.3655796, 0.4028401, 0.3335596, 0.3398343, 0.3976401, 0.395231, 
    0.4402498, 0.3956096, 0.3733369, 0.3072077, 0.270905, 0.2442578, 
    0.2999628, 0.1862635, 0.2709249, 0.4195056, 0.3063478, 0.2721661, 
    0.3350045, 0.2648022, 0.3678871, 0.2627528, 0.1464882, 0.01791377, 
    0.1049556, 0.1794422, 0.1735056, 0.278278,
  0.254561, 0.2449223, 0.1891186, 0.1813116, 0.2990642, 0.2483763, 0.218166, 
    0.2292912, 0.3196006, 0.2360162, 0.1766893, 0.09340791, 0.04605445, 
    0.153023, 0.2610763, 0.3166517, 0.3402959, 0.3604299, 0.2323013, 
    0.3345012, 0.3298744, 0.3128829, 0.1927192, 0.05482632, 0.05085336, 
    0.3114988, 0.2054791, 0.2566761, 0.336962,
  0.2150007, 0.07277842, 0.03143242, 0.1098487, 0.1440964, 0.157296, 
    0.1966535, 0.1941604, 0.1013973, 0.04119044, -2.674111e-05, 4.410286e-05, 
    0.008668985, 0.07668279, 0.1285264, 0.1003599, 0.1499021, 0.1387804, 
    0.124289, 0.2462558, 0.1580367, 0.1516066, 0.2648645, 3.715443e-06, 
    0.009999012, 0.08889315, 0.1190514, 0.2131213, 0.228459,
  0.3606304, -5.690857e-05, 0.0006735608, 0.01479278, 0.05700769, 0.07200707, 
    0.07420726, 0.07296102, 0.06451356, 2.71943e-07, 3.98682e-08, 
    -6.759558e-07, 0.05849495, 0.0944358, 0.09323263, 0.1074793, 0.1272522, 
    0.06690005, 0.05650563, 0.1118198, 0.170503, 0.3023695, 0.03593208, 
    0.0001891963, 0.05842885, 0.2219941, 0.1001633, 0.1658752, 0.4450241,
  0.01360312, 0.05165443, 0.0189277, 0.1055754, 0.06215929, 0.07756852, 
    0.04435827, 0.06374113, 0.09185594, 0.009653385, 0.01199275, 0.01569388, 
    0.06785493, 0.03887435, 0.06922724, 0.06923179, 0.04788174, 0.06485355, 
    0.05092231, 0.0509227, 0.1538523, 0.1607414, 0.004222057, 0.02582866, 
    0.0310582, 0.01279689, 0.08324245, 0.07731541, 0.05646255,
  0.09098917, 0.2041612, 0.04959938, 0.2024725, 0.04052833, 0.02952555, 
    0.05110502, 0.02618988, 0.1238373, 0.1418556, 0.06365592, 0.024678, 
    0.06829636, 0.05810815, 0.0400365, 0.070021, 0.04285061, 0.03595193, 
    0.01765092, 0.01676823, 0.01788191, 0.0006088183, 0.00144642, 0.04528629, 
    0.03016748, 0.02410414, 0.06932168, 0.0662314, 0.06583103,
  2.006608e-05, 3.016374e-06, 7.297917e-05, 0.03809636, 0.06520366, 
    0.1220061, 0.02672987, 0.08169817, 0.16438, 0.07838483, 0.07761921, 
    0.071179, 0.04919342, 0.05832563, 0.07235057, 0.05318072, 0.06742411, 
    0.09911246, 0.1526459, 0.08768737, 0.121905, 0.05283262, 0.1546647, 
    0.08706504, 0.05390691, 0.1042439, 0.1275667, 0.001413022, 2.319991e-05,
  2.44482e-07, 2.45991e-09, 4.610236e-06, 0.02670783, 0.001900404, 0.111273, 
    0.02228765, 0.05278889, 0.1284778, 0.1424587, 0.1061816, 0.07809618, 
    0.07158653, 0.117198, 0.0821114, 0.06040528, 0.07160331, 0.04725865, 
    0.1787818, 0.169286, 0.03997885, 0.2721223, 0.07202177, 0.1008114, 
    0.05674127, 0.06524447, 0.0918098, 0.01229263, 7.986817e-07,
  6.443464e-07, 0.03474782, 0.03844761, 0.0210786, 0.115627, 8.975465e-06, 
    0.00221714, 0.03332683, 0.1621733, 0.001775657, 0.2015252, 0.1692062, 
    0.1363098, 0.1663673, 0.2863837, 0.1727195, 0.164118, 0.1371881, 
    0.2479633, 0.01504056, 0.01411626, 0.07740459, 0.1460598, 0.1483529, 
    0.1520656, 0.1210289, 0.06970245, 0.149315, 0.01409091,
  0.03009623, 0.1166582, 0.09256301, 0.1143816, 0.0406378, 0.007251482, 
    0.06270938, -0.0002211092, 1.134983e-05, 0.01229648, 0.1422379, 
    0.2723408, 0.3808033, 0.3001693, 0.2876656, 0.3015924, 0.3450398, 
    0.2494523, 0.2918555, 0.08996783, 0.04975436, 0.06300952, 0.195328, 
    0.1929857, 0.2334423, 0.1719826, 0.2325276, 0.2664067, 0.2436517,
  0.2728377, 0.2309757, 0.2661135, 0.2883037, 0.2087097, 0.1435855, 
    0.1439091, 0.2607018, 0.08615121, 0.1582733, 0.1556166, 0.1710004, 
    0.3604743, 0.3104116, 0.2676837, 0.2121434, 0.2503811, 0.2686725, 
    0.2872529, 0.3640269, 0.1557382, 0.3472819, 0.3852313, 0.5644287, 
    0.3120112, 0.342876, 0.2184163, 0.2241221, 0.2085152,
  0.2001953, 0.4357019, 0.3968448, 0.4406841, 0.5126405, 0.463451, 0.450671, 
    0.491485, 0.485425, 0.5050694, 0.4676629, 0.327486, 0.1367583, 0.2319003, 
    0.5301495, 0.254283, 0.4002883, 0.3130717, 0.4233503, 0.2533253, 
    0.4358007, 0.3962938, 0.5335691, 0.4707083, 0.3736725, 0.2057381, 
    0.2740401, 0.3269613, 0.2109882,
  0.1722371, 0.2304821, 0.3633392, 0.3720812, 0.4785096, 0.395248, 0.248843, 
    0.3612238, 0.3613179, 0.4604011, 0.3715339, 0.2842665, 0.2314643, 
    0.3722363, 0.4106958, 0.2385194, 0.299681, 0.3661479, 0.2613827, 
    0.4408737, 0.2946542, 0.3011878, 0.3132861, 0.2207205, 0.2284154, 
    0.275613, 0.1244148, 0.2084052, 0.2693848,
  0.2241564, 0.3615384, 0.3003735, 0.2289128, 0.2165646, 0.2791118, 
    0.2572027, 0.2631548, 0.2674295, 0.3128125, 0.2653872, 0.2421222, 
    0.2002736, 0.2774918, 0.3686748, 0.3935023, 0.418463, 0.4273402, 0.50506, 
    0.4218536, 0.3530492, 0.3401458, 0.2611378, 0.3036373, 0.3357922, 
    0.3351339, 0.1192209, 0.2060676, 0.2905618,
  0.190781, 0.1941935, 0.197606, 0.2010184, 0.2044309, 0.2078433, 0.2112558, 
    0.2405453, 0.2338377, 0.2271301, 0.2204225, 0.2137149, 0.2070073, 
    0.2002997, 0.2133704, 0.2202584, 0.2271464, 0.2340344, 0.2409225, 
    0.2478105, 0.2546985, 0.209535, 0.2059422, 0.2023493, 0.1987564, 
    0.1951636, 0.1915707, 0.1879779, 0.1880511,
  0.04880956, 0.07337786, 0.08815006, 0.1918407, 0.2051746, 0.2440125, 
    0.2425863, 0.1352908, 0.1870826, 0.1764255, 0.1091226, 0.09086669, 
    0.1138479, 0.03067797, 0.04377697, 0.05883656, 0.06838977, 0.1218304, 
    0.06759429, 0.03046084, 0.1782272, 0.191101, 0.368536, 0.2363301, 
    0.2766718, 0.242178, 0.09599607, 0.03286926, 0.04872895,
  0.289377, 0.1801077, 0.1590603, 0.096932, 0.2340581, 0.3327309, 0.07741738, 
    0.2083242, 0.2654222, 0.3026756, 0.1694111, 0.06707539, 0.1246436, 
    0.2412813, 0.3009491, 0.2914326, 0.3026005, 0.3266243, 0.40116, 
    0.2557406, 0.2630194, 0.3060711, 0.3450097, 0.5599841, 0.1899379, 
    0.330628, 0.368184, 0.3789178, 0.3642868,
  0.4228758, 0.4158004, 0.4691305, 0.4584853, 0.5277701, 0.427095, 0.4388431, 
    0.4770205, 0.4065886, 0.3695216, 0.4617776, 0.5404812, 0.4437761, 
    0.4186162, 0.3474597, 0.4445644, 0.4398484, 0.5088575, 0.4093558, 
    0.3816579, 0.3528779, 0.2724189, 0.2953911, 0.3981785, 0.3526332, 
    0.3442101, 0.4427994, 0.3963017, 0.4641365,
  0.3787045, 0.3950878, 0.4081561, 0.3440489, 0.3585821, 0.4111345, 
    0.3852306, 0.3744127, 0.3463125, 0.3622519, 0.2772094, 0.286113, 
    0.181932, 0.2877543, 0.2516798, 0.3358632, 0.4241105, 0.440134, 
    0.3416771, 0.3574269, 0.292915, 0.3735982, 0.3631358, 0.1352717, 
    0.01383813, 0.1583564, 0.282696, 0.262152, 0.2775086,
  0.3504226, 0.2762821, 0.1232338, 0.2102501, 0.2224583, 0.1862496, 
    0.2076243, 0.2426165, 0.3049322, 0.330597, 0.2873585, 0.131248, 
    0.0283222, 0.1677242, 0.2929631, 0.3544484, 0.3127365, 0.3694189, 
    0.2927936, 0.4379562, 0.3625003, 0.2895482, 0.2228659, 0.08589959, 
    0.06101299, 0.3430304, 0.3168086, 0.3103453, 0.3403369,
  0.3135318, 0.09371501, 0.02930219, 0.1415647, 0.2310071, 0.1806977, 
    0.2084597, 0.2064613, 0.2330964, 0.06908882, -2.851519e-05, 3.078618e-05, 
    0.007096996, 0.1037636, 0.1542837, 0.2175905, 0.1219543, 0.137521, 
    0.133432, 0.181076, 0.1424691, 0.1733029, 0.3917694, 0.0002513271, 
    0.01505439, 0.08161429, 0.1168057, 0.1782281, 0.1875149,
  0.4293165, -0.000213918, 0.0003494954, 0.04445046, 0.1157947, 0.1058223, 
    0.118651, 0.1734263, 0.2122536, 4.817576e-07, 4.438964e-08, 
    -3.249361e-07, 0.05029586, 0.08458097, 0.1460662, 0.1239722, 0.08704136, 
    0.0622199, 0.07036583, 0.0768972, 0.1153152, 0.366426, 0.5561478, 
    0.003141768, 0.03644977, 0.2197621, 0.08777217, 0.09236097, 0.345778,
  0.2061845, 0.09801022, 0.0134877, 0.1174217, 0.07378306, 0.0857994, 
    0.07389897, 0.07845264, 0.1909177, 0.1367879, 0.03366333, 0.04065588, 
    0.06518304, 0.05921062, 0.07875551, 0.0772054, 0.07042403, 0.08949019, 
    0.08507872, 0.09758735, 0.1748923, 0.4206886, 0.03809553, 0.01820364, 
    0.01946091, 0.006149219, 0.1092136, 0.07881268, 0.321263,
  0.08153152, 0.1856517, 0.02660529, 0.170095, 0.1034414, 0.1460307, 
    0.1682507, 0.05765903, 0.1122904, 0.1152444, 0.05760821, 0.1029697, 
    0.1232865, 0.1112065, 0.1186557, 0.1054343, 0.08765301, 0.1002253, 
    0.08294982, 0.08023862, 0.06852913, 0.01610574, 0.01315109, 0.02950016, 
    0.01281501, 0.04497405, 0.08783074, 0.07409769, 0.07205067,
  1.080268e-05, 8.562167e-07, 3.866836e-05, 0.02184077, 0.09043121, 
    0.1830886, 0.01606234, 0.07758623, 0.1162089, 0.104537, 0.06241464, 
    0.04359413, 0.06877555, 0.0699101, 0.06327718, 0.05983197, 0.08803447, 
    0.1045404, 0.1509113, 0.09503246, 0.1107247, 0.06534989, 0.184496, 
    0.09521402, 0.08190119, 0.06970077, 0.0996584, 0.05888768, 7.600668e-06,
  1.482062e-07, 1.046023e-09, 3.089941e-06, 0.02345505, 0.00147307, 
    0.06032289, 0.01602399, 0.09180228, 0.1027121, 0.1225461, 0.07978476, 
    0.09348506, 0.1073091, 0.09377971, 0.06358446, 0.0605999, 0.1119448, 
    0.04617068, 0.2147851, 0.2779691, 0.1642769, 0.2692019, 0.0444256, 
    0.08065043, 0.06221273, 0.06490017, 0.1234469, 0.03898744, 3.465132e-07,
  2.293804e-07, 0.03332004, 0.03775731, 0.01365009, 0.09912997, 
    -1.911018e-06, 0.001348204, 0.01993943, 0.1594265, 0.0004066185, 
    0.1445986, 0.1812924, 0.1228625, 0.1509281, 0.2308692, 0.1455201, 
    0.103011, 0.1012165, 0.2433723, 0.02004014, 0.0189029, 0.09466015, 
    0.1585966, 0.08814979, 0.1345957, 0.1925253, 0.05918713, 0.1071153, 
    0.0217162,
  0.03004856, 0.1364688, 0.1420109, 0.1248777, 0.03717986, 0.003899954, 
    0.07899368, -0.000288501, -0.0001201636, 0.0124267, 0.1491055, 0.1740248, 
    0.2632088, 0.2299102, 0.2716771, 0.2725584, 0.3264894, 0.2928947, 
    0.2671545, 0.09050226, 0.04009044, 0.08013789, 0.2134002, 0.2132649, 
    0.1671248, 0.1845439, 0.1982037, 0.2599402, 0.179399,
  0.2597176, 0.2525588, 0.2754101, 0.3863901, 0.2771071, 0.1511612, 
    0.1454174, 0.2761122, 0.08923105, 0.1927019, 0.1196321, 0.2097316, 
    0.2124058, 0.2287975, 0.2229144, 0.2047145, 0.2173323, 0.2802788, 
    0.2837237, 0.3704588, 0.1660628, 0.270713, 0.3534398, 0.650496, 
    0.3592169, 0.3023963, 0.2247321, 0.1855891, 0.1807171,
  0.1634806, 0.4209051, 0.5170417, 0.4934573, 0.5882007, 0.4884327, 
    0.5092632, 0.6010332, 0.5023066, 0.543608, 0.4999258, 0.3431715, 
    0.119799, 0.289173, 0.4311135, 0.2004625, 0.4113443, 0.3154665, 
    0.4428983, 0.2368757, 0.4867495, 0.4551339, 0.489049, 0.5077343, 
    0.3183669, 0.1781614, 0.2296732, 0.2414264, 0.1563242,
  0.1138945, 0.1761146, 0.3795331, 0.2775418, 0.3950996, 0.4872497, 
    0.2748864, 0.4112325, 0.3642887, 0.4710271, 0.404016, 0.3209463, 
    0.2775109, 0.4571579, 0.4205756, 0.2412018, 0.3348244, 0.407654, 
    0.3037484, 0.4609791, 0.3813571, 0.3030066, 0.3245704, 0.2635901, 
    0.2570894, 0.2880118, 0.134405, 0.1600324, 0.1873149,
  0.268272, 0.5120638, 0.3068324, 0.2359336, 0.2240548, 0.3039728, 0.2438401, 
    0.2837857, 0.282858, 0.3534938, 0.3341526, 0.2794846, 0.2764504, 
    0.3443344, 0.4176628, 0.428198, 0.4538462, 0.438563, 0.516733, 0.4547789, 
    0.3755865, 0.3000127, 0.291212, 0.2710522, 0.3272742, 0.3742971, 
    0.1618411, 0.2337219, 0.303638,
  0.2558433, 0.2643838, 0.2729243, 0.2814648, 0.2900054, 0.2985459, 
    0.3070864, 0.3289601, 0.3162582, 0.3035564, 0.2908546, 0.2781528, 
    0.2654509, 0.2527491, 0.2492965, 0.2550429, 0.2607893, 0.2665357, 
    0.2722821, 0.2780285, 0.2837749, 0.2406986, 0.2391135, 0.2375284, 
    0.2359434, 0.2343583, 0.2327732, 0.2311881, 0.2490109,
  0.0318316, 0.06975681, 0.08236156, 0.2150936, 0.2430999, 0.2474438, 
    0.2520626, 0.14738, 0.2611336, 0.2272843, 0.135636, 0.1047588, 0.1158179, 
    0.03176184, 0.0437469, 0.09609058, 0.1020394, 0.129717, 0.1342559, 
    0.04523441, 0.1719009, 0.2102116, 0.4012753, 0.2399632, 0.2292892, 
    0.2423115, 0.06623251, 0.02047713, 0.03428934,
  0.2811963, 0.1352475, 0.1599903, 0.07859481, 0.2028234, 0.3044968, 
    0.05260462, 0.1510987, 0.2209456, 0.2547028, 0.1424323, 0.06479447, 
    0.09493928, 0.2058583, 0.2889509, 0.2885985, 0.3003783, 0.2937131, 
    0.3854867, 0.2792642, 0.2680044, 0.2750033, 0.3103606, 0.503661, 
    0.1606744, 0.2610527, 0.3388537, 0.3448009, 0.3149896,
  0.3800154, 0.333992, 0.4279095, 0.4613453, 0.4558374, 0.4124752, 0.4159946, 
    0.4590128, 0.4305158, 0.3330149, 0.4504832, 0.4896975, 0.4701074, 
    0.3834891, 0.3799975, 0.5040168, 0.4995955, 0.5990197, 0.4964253, 
    0.3096398, 0.2844057, 0.2374975, 0.2847863, 0.396941, 0.3466529, 
    0.3648674, 0.4246086, 0.4171261, 0.4963175,
  0.4725956, 0.4298022, 0.417266, 0.369908, 0.335566, 0.3490815, 0.3856727, 
    0.3258829, 0.3136519, 0.345918, 0.2565065, 0.2488987, 0.1408625, 
    0.2154711, 0.2339815, 0.3510408, 0.3652693, 0.4464863, 0.5770345, 
    0.3589244, 0.3665595, 0.3687146, 0.3928922, 0.1213318, 0.01530091, 
    0.1978946, 0.3596176, 0.2999452, 0.3164952,
  0.3294131, 0.1895282, 0.09008819, 0.1631666, 0.1847242, 0.1467986, 
    0.1751432, 0.2534487, 0.3106178, 0.2498452, 0.2611896, 0.06823, 
    0.02051916, 0.1414515, 0.3180986, 0.3112797, 0.3036533, 0.3201698, 
    0.3118429, 0.310325, 0.3563816, 0.3023516, 0.2281303, 0.1096806, 
    0.06239314, 0.3136487, 0.3370987, 0.3361131, 0.3580929,
  0.1213817, 0.05427961, 0.02378277, 0.1415463, 0.2707085, 0.1433432, 
    0.1640254, 0.1372609, 0.3095637, 0.04813952, 0.001031795, 8.040795e-06, 
    0.004116355, 0.1749671, 0.1283012, 0.08785793, 0.07808746, 0.0725335, 
    0.09970287, 0.1183812, 0.1028307, 0.06282309, 0.2611741, 0.01255437, 
    0.01735859, 0.09275142, 0.1291288, 0.1196161, 0.06768653,
  0.2682249, -0.000717651, 0.000113236, 0.06514568, 0.06017106, 0.0718549, 
    0.07766528, 0.1092994, 0.2361498, -0.0001793051, -2.022897e-09, 
    3.153282e-08, 0.117913, 0.08977076, 0.05976372, 0.0918096, 0.0345365, 
    0.06778127, 0.03380755, 0.03476271, 0.03745023, 0.1281161, 0.4986686, 
    0.1092594, 0.0236764, 0.2001107, 0.05831566, 0.02296604, 0.1416386,
  0.421395, 0.1617633, 0.004688811, 0.1469151, 0.03725724, 0.04194357, 
    0.0486978, 0.02848387, 0.07681151, 0.1595341, 0.03450545, 0.067749, 
    0.07252114, 0.02686658, 0.03318295, 0.03361156, 0.03320219, 0.04593736, 
    0.01952183, 0.02381232, 0.08034184, 0.2193415, 0.6206231, 0.008037572, 
    0.009951299, 0.002312594, 0.03391186, 0.04182001, 0.1974007,
  0.08254441, 0.1654664, 0.01521151, 0.1740631, 0.06089524, 0.1469371, 
    0.1174833, 0.2054581, 0.107596, 0.08036286, 0.01600737, 0.02191604, 
    0.02206765, 0.01857411, 0.06320351, 0.04135491, 0.04123003, 0.05664244, 
    0.08642738, 0.1451177, 0.3710656, 0.252931, 0.2101753, 0.02277005, 
    0.003885591, 0.05813793, 0.09485302, 0.07062253, 0.1412681,
  3.789859e-06, -2.413605e-08, 1.948431e-05, 0.0238402, 0.09924003, 
    0.0487275, 0.01516798, 0.02787673, 0.04451715, 0.01788131, 0.03549127, 
    0.02513261, 0.02933435, 0.04366883, 0.03077625, 0.03849667, 0.06895579, 
    0.08088532, 0.1268822, 0.08257824, 0.1025143, 0.128732, 0.2054369, 
    0.08550764, 0.03301773, 0.02642053, 0.03097325, 0.09085936, 7.007091e-06,
  1.447017e-07, 7.786695e-10, 2.400551e-06, 0.0124924, 0.0006266041, 
    0.03393682, 0.02378375, 0.03008947, 0.06378734, 0.07252665, 0.03919361, 
    0.02748695, 0.04344816, 0.05670998, 0.02659531, 0.02374407, 0.03977795, 
    0.06307818, 0.1018454, 0.1712004, 0.08075812, 0.199343, 0.00638578, 
    0.04275296, 0.02624681, 0.020838, 0.02871072, 0.004946875, 2.073869e-07,
  -2.857177e-07, 0.02877179, 0.0163858, 0.03055592, 0.08794595, 
    -1.211871e-06, 0.001362347, 0.01015503, 0.1487858, 0.0019701, 0.1056817, 
    0.1539713, 0.1137292, 0.1284572, 0.1593774, 0.1033354, 0.07312609, 
    0.07393655, 0.1158665, 0.02324285, 0.01981632, 0.08600593, 0.1608623, 
    0.05449584, 0.06581741, 0.1313655, 0.02456804, 0.03969743, 0.01839996,
  0.04023586, 0.09978914, 0.1364102, 0.129234, 0.01364717, 0.002519478, 
    0.0976494, -0.0003893836, -0.000164559, 0.02094154, 0.1827602, 0.1197168, 
    0.1735694, 0.1513112, 0.2189099, 0.2035423, 0.2430699, 0.2447227, 
    0.2409495, 0.09180892, 0.03061514, 0.07289492, 0.1904346, 0.1814932, 
    0.130553, 0.1425453, 0.169695, 0.2035855, 0.1269511,
  0.2238483, 0.2858055, 0.304095, 0.4610581, 0.2785563, 0.1695226, 0.1267941, 
    0.2888836, 0.08962367, 0.1980666, 0.07388819, 0.2157807, 0.1356488, 
    0.1904703, 0.1740714, 0.1535404, 0.150407, 0.2540223, 0.2498991, 
    0.3841211, 0.1979041, 0.2266946, 0.2638806, 0.6693771, 0.3383306, 
    0.2536051, 0.2019509, 0.1598953, 0.1534929,
  0.09867002, 0.4372928, 0.524788, 0.630405, 0.7356972, 0.428051, 0.5397798, 
    0.6272338, 0.5991264, 0.4805842, 0.4883914, 0.4151385, 0.1206914, 
    0.340782, 0.3079396, 0.1788981, 0.3580921, 0.3062031, 0.4415085, 
    0.2489104, 0.5717039, 0.4094955, 0.3235638, 0.5050614, 0.2779087, 
    0.1338129, 0.1568633, 0.1857107, 0.1129203,
  0.0794246, 0.114872, 0.3897064, 0.153167, 0.3134567, 0.4405341, 0.3441235, 
    0.3933943, 0.3802282, 0.4734018, 0.4116018, 0.3455459, 0.3217059, 
    0.5327531, 0.4522329, 0.2697409, 0.3704029, 0.4052956, 0.3121484, 
    0.4389127, 0.42484, 0.3432096, 0.3464497, 0.3159981, 0.2625101, 
    0.3006898, 0.1620534, 0.140322, 0.1052569,
  0.2611012, 0.5169445, 0.3289842, 0.2311536, 0.2176276, 0.3003675, 0.295589, 
    0.3000943, 0.3430224, 0.4247666, 0.3575238, 0.3307886, 0.3517661, 
    0.4369728, 0.5039864, 0.4706558, 0.4750983, 0.4804062, 0.5378641, 
    0.4614469, 0.3950603, 0.2705919, 0.2842103, 0.2639116, 0.2887168, 
    0.3862371, 0.1913185, 0.2425428, 0.2912957,
  0.4036934, 0.4097953, 0.4158973, 0.4219992, 0.4281011, 0.434203, 0.440305, 
    0.4314605, 0.416173, 0.4008855, 0.3855979, 0.3703104, 0.3550228, 
    0.3397353, 0.3469823, 0.3536994, 0.3604166, 0.3671338, 0.3738509, 
    0.3805681, 0.3872852, 0.3479839, 0.3504524, 0.3529209, 0.3553893, 
    0.3578578, 0.3603262, 0.3627947, 0.3988118,
  0.02305798, 0.05787795, 0.0735241, 0.2246489, 0.2882428, 0.2436381, 
    0.2655916, 0.1646001, 0.3195255, 0.3060731, 0.199746, 0.1253335, 
    0.1017622, 0.01598345, 0.09816016, 0.1664654, 0.1438326, 0.08596198, 
    0.1453971, 0.07419693, 0.1542565, 0.2149902, 0.4103943, 0.2068085, 
    0.1672785, 0.2735538, 0.03493136, 0.01571605, 0.02800309,
  0.2071263, 0.1016685, 0.1212541, 0.05553212, 0.155883, 0.2537637, 
    0.02901744, 0.08498897, 0.1696152, 0.17704, 0.1069099, 0.05460056, 
    0.07364924, 0.1816902, 0.256666, 0.2569469, 0.2789403, 0.2758707, 
    0.3805759, 0.269749, 0.2707033, 0.2610339, 0.291313, 0.4110748, 
    0.1153837, 0.2556433, 0.3211581, 0.3058524, 0.2681078,
  0.3526775, 0.2872086, 0.3831422, 0.4322774, 0.4013743, 0.3989562, 
    0.4476885, 0.4513082, 0.4219854, 0.2845862, 0.4092672, 0.465297, 
    0.4661174, 0.3396774, 0.389697, 0.5035984, 0.5596081, 0.6134724, 
    0.4878764, 0.270812, 0.241868, 0.2120285, 0.2770402, 0.3744627, 
    0.3500454, 0.4052277, 0.4491308, 0.475022, 0.5015956,
  0.4298042, 0.4098666, 0.3753072, 0.3284605, 0.3139752, 0.3082941, 
    0.3614405, 0.3061143, 0.2924875, 0.3223518, 0.2236792, 0.2120077, 
    0.1138949, 0.2041688, 0.1910561, 0.3072594, 0.3672693, 0.3810194, 
    0.4959038, 0.402396, 0.3271475, 0.3596938, 0.3245564, 0.09979389, 
    0.01588444, 0.2379599, 0.3555382, 0.281677, 0.38424,
  0.2431064, 0.1226826, 0.03807713, 0.1330855, 0.1520022, 0.133806, 
    0.1438856, 0.2205302, 0.2670961, 0.1637358, 0.135442, 0.03560878, 
    0.01077119, 0.1268018, 0.3166704, 0.2976236, 0.3031028, 0.2644664, 
    0.2654083, 0.2248295, 0.3262662, 0.2519871, 0.1584117, 0.1174732, 
    0.05886239, 0.2730182, 0.3065089, 0.3348809, 0.2895415,
  0.03945137, 0.05577973, 0.01721984, 0.1649397, 0.2478645, 0.09017179, 
    0.09619434, 0.08128231, 0.177702, 0.01400546, 0.0007318135, 2.073648e-06, 
    0.003500488, 0.2129218, 0.1019774, 0.06147986, 0.04862794, 0.04898384, 
    0.05786034, 0.07878949, 0.05950933, 0.02946104, 0.09697368, 0.02012869, 
    0.01526453, 0.05844283, 0.1348276, 0.08266452, 0.02469693,
  0.1031487, 0.00327213, -4.606273e-05, 0.01697823, 0.01207485, 0.01304339, 
    0.02598927, 0.04689718, 0.08129332, -6.927593e-05, 3.328686e-08, 
    3.891462e-08, 0.06088041, 0.03061358, 0.01891814, 0.03824605, 0.0130135, 
    0.04086537, 0.01740797, 0.01572888, 0.008277652, 0.04063127, 0.1893636, 
    0.1594746, 0.01746926, 0.1843941, 0.03938907, 0.004114592, 0.04029494,
  0.2482932, 0.1631505, 0.002546435, 0.1953181, 0.009560497, 0.01555528, 
    0.01185811, 0.003781212, 0.0197119, 0.04066261, 0.01274543, 0.02169886, 
    0.02839607, 0.008400477, 0.01884515, 0.0134901, 0.005185422, 0.00575677, 
    0.004156491, 0.004890351, 0.02034868, 0.07008881, 0.3970475, 0.004927973, 
    0.006036161, 0.001235407, 0.0001537838, 0.004803142, 0.1013097,
  0.1029289, 0.1412447, 0.007791462, 0.1684596, 0.02096714, 0.02386604, 
    0.02255862, 0.02759985, 0.09827639, 0.04350124, 0.005975265, 0.004210236, 
    0.005412901, 0.005436392, 0.01396265, 0.008190383, 0.008128247, 
    0.01349642, 0.02819007, 0.06226308, 0.2083401, 0.5131905, 0.3256511, 
    0.01284021, 0.001395898, 0.02254126, 0.04297356, 0.04155524, 0.1033501,
  5.308671e-06, 3.849763e-07, 1.066358e-05, 0.0202199, 0.08010495, 
    0.01246821, 0.003024495, 0.009431365, 0.01852046, 0.00824327, 0.01708963, 
    0.007367871, 0.01315224, 0.02169368, 0.01326098, 0.01031098, 0.0177781, 
    0.04408306, 0.08531972, 0.07088025, 0.05714531, 0.03136528, 0.2483867, 
    0.06004342, 0.01207298, 0.01351085, 0.005592263, 0.01471492, 3.590337e-06,
  1.42429e-07, 6.718746e-10, 2.066222e-06, 0.006378571, 0.0002229472, 
    0.009399266, 0.01602538, 0.007680899, 0.0484153, 0.03417205, 0.01588853, 
    0.0077492, 0.015234, 0.02742699, 0.01236924, 0.006425455, 0.02087454, 
    0.03295627, 0.04844581, 0.0637176, 0.03342715, 0.1387551, 0.001509911, 
    0.02769478, 0.006007756, 0.008644837, 0.007612283, 0.0009927996, 
    1.604712e-07,
  -7.5782e-07, 0.02623178, 0.003879207, 0.02181885, 0.07891893, 
    -9.025433e-06, 0.0008965675, 0.005405839, 0.1278403, 0.004218898, 
    0.03261495, 0.08720025, 0.07743285, 0.0646771, 0.1211497, 0.05574542, 
    0.04362976, 0.07434303, 0.08660108, 0.0071064, 0.02111292, 0.07048128, 
    0.1495693, 0.02785244, 0.02809123, 0.06144951, 0.007973104, 0.01064657, 
    0.01861214,
  0.01878016, 0.04901749, 0.1035644, 0.1248073, 0.03268562, 0.002060359, 
    0.09477193, 6.274543e-05, -0.0001234208, 0.01549834, 0.2033246, 
    0.08259207, 0.1294969, 0.1095753, 0.1604456, 0.1446461, 0.1910015, 
    0.1824073, 0.2100967, 0.09539273, 0.02211207, 0.06362791, 0.1460655, 
    0.1529195, 0.101683, 0.1164856, 0.1422596, 0.1536658, 0.08795899,
  0.1849158, 0.2621482, 0.2940629, 0.4295003, 0.218434, 0.1819184, 0.1118605, 
    0.2774733, 0.0677197, 0.1558875, 0.0570053, 0.2081175, 0.09797965, 
    0.1513102, 0.1278445, 0.1066837, 0.108839, 0.2173442, 0.2046813, 
    0.4083476, 0.1852155, 0.186825, 0.2158854, 0.7086793, 0.2864156, 
    0.2080987, 0.1684976, 0.1369169, 0.1436918,
  0.06569979, 0.4390446, 0.4441612, 0.7620544, 0.7624621, 0.4268385, 
    0.5957512, 0.5987832, 0.6052508, 0.4556936, 0.4665901, 0.4791968, 
    0.1189086, 0.2700657, 0.2229449, 0.1552462, 0.3300911, 0.273246, 
    0.3805803, 0.2641039, 0.718173, 0.3188803, 0.2105258, 0.4729537, 
    0.2315925, 0.1029677, 0.1184925, 0.1255461, 0.07499411,
  0.05408363, 0.07245994, 0.3497815, 0.0797988, 0.2052671, 0.3795967, 
    0.5098826, 0.3652104, 0.3734147, 0.5191264, 0.4154044, 0.3753974, 
    0.3536984, 0.5600542, 0.4598994, 0.2866096, 0.3903547, 0.3993921, 
    0.3620052, 0.4142174, 0.432114, 0.4215511, 0.3865401, 0.382046, 
    0.1654243, 0.3085646, 0.1776189, 0.1247265, 0.0530843,
  0.3032326, 0.427956, 0.3587398, 0.2693928, 0.2478954, 0.340494, 0.3611872, 
    0.3867516, 0.4535021, 0.4781828, 0.4033092, 0.3797445, 0.439742, 
    0.5144865, 0.5744557, 0.5525329, 0.5498325, 0.5503082, 0.6210444, 
    0.4880634, 0.4256192, 0.2580482, 0.3183176, 0.2520061, 0.2486738, 
    0.4074059, 0.2100187, 0.2646982, 0.3147159,
  0.5170724, 0.5234949, 0.5299174, 0.5363398, 0.5427623, 0.5491847, 
    0.5556072, 0.5267663, 0.5169966, 0.5072268, 0.4974571, 0.4876874, 
    0.4779177, 0.468148, 0.5229923, 0.5266818, 0.5303714, 0.534061, 
    0.5377506, 0.5414402, 0.5451298, 0.4830944, 0.482752, 0.4824097, 
    0.4820673, 0.481725, 0.4813827, 0.4810404, 0.5119345,
  0.01807222, 0.05745756, 0.06921196, 0.211994, 0.3235233, 0.246678, 
    0.2632977, 0.2092868, 0.352765, 0.3169978, 0.212726, 0.1113537, 
    0.09429233, 0.01062896, 0.1208737, 0.1774042, 0.1542437, 0.1142547, 
    0.1527882, 0.08432839, 0.1288766, 0.2033441, 0.377753, 0.1538913, 
    0.1164439, 0.2036687, 0.02001869, 0.01127581, 0.02293336,
  0.1320179, 0.07671699, 0.07590725, 0.04157032, 0.1196267, 0.1898858, 
    0.01044056, 0.05217276, 0.1227725, 0.1028382, 0.06054855, 0.05018963, 
    0.04526681, 0.1585635, 0.2409546, 0.2586733, 0.2595892, 0.2414743, 
    0.3786103, 0.2551283, 0.2580852, 0.2298952, 0.262284, 0.35867, 
    0.09928152, 0.2608756, 0.2725756, 0.2105289, 0.2126453,
  0.3138655, 0.2338804, 0.3506104, 0.3562461, 0.345949, 0.3674947, 0.430355, 
    0.3837114, 0.3992146, 0.2543712, 0.3403563, 0.4175001, 0.4170902, 
    0.2925041, 0.3470571, 0.4488973, 0.5385705, 0.5745878, 0.4263961, 
    0.2341769, 0.2062742, 0.186371, 0.239755, 0.3440558, 0.3597715, 
    0.4439031, 0.4887026, 0.4756926, 0.4314667,
  0.353025, 0.3662895, 0.3313945, 0.2879388, 0.2735797, 0.270414, 0.326091, 
    0.2623951, 0.2600749, 0.2905469, 0.1680267, 0.1695407, 0.08468554, 
    0.1729232, 0.1949751, 0.2567802, 0.3301164, 0.320288, 0.3586522, 
    0.332683, 0.2696764, 0.3353889, 0.2562411, 0.07695082, 0.01391438, 
    0.2815359, 0.3472196, 0.3073888, 0.4228275,
  0.155035, 0.06965542, 0.01633906, 0.09697043, 0.1247547, 0.1133911, 
    0.1144979, 0.1768204, 0.1945198, 0.1071105, 0.05791431, 0.02013727, 
    0.006163427, 0.1148443, 0.2979921, 0.2846111, 0.2697927, 0.2357458, 
    0.2483946, 0.1515793, 0.2912516, 0.1790213, 0.1314527, 0.114429, 
    0.04519525, 0.2352638, 0.2644941, 0.3150179, 0.2020299,
  0.01952599, 0.02595978, 0.01289152, 0.1694219, 0.1721215, 0.04320806, 
    0.06031046, 0.03150215, 0.08724742, 0.005433119, 0.0004326485, 
    7.235387e-07, 0.003669631, 0.1473017, 0.05760042, 0.03429899, 0.03773715, 
    0.03871711, 0.03922172, 0.05069814, 0.02415685, 0.01130487, 0.04248423, 
    0.02518843, 0.009692388, 0.03131819, 0.1146532, 0.05345212, 0.01083199,
  0.04452902, 0.008239628, -4.889644e-05, 0.01115007, 0.002797466, 
    0.004527789, 0.006663275, 0.01172221, 0.04341751, -2.951975e-05, 
    2.834076e-08, 3.665932e-08, 0.01675223, 0.01069822, 0.01078951, 
    0.01967976, 0.002771358, 0.01145158, 0.005059312, 0.007517871, 
    0.00265359, 0.01596216, 0.07966637, 0.058734, 0.01111377, 0.181977, 
    0.02129675, 0.001279637, 0.01412255,
  0.0913302, 0.04256099, 0.0009786258, 0.1982787, 0.001731738, 0.003752663, 
    0.002240211, 0.0004792013, 0.006713178, 0.01159944, 0.004292193, 
    0.007752737, 0.01091267, 0.001332312, 0.01072432, 0.00867664, 
    0.0005294197, 0.001141676, 0.001698501, 0.002080026, 0.008024968, 
    0.02627126, 0.1658377, 0.006585647, 0.002697853, 0.000482921, 
    -0.001670554, 0.001088822, 0.03066595,
  0.03151078, 0.1441106, 0.009904286, 0.1418976, 0.004092105, 0.005941727, 
    0.005098188, 0.006465957, 0.1071328, 0.02549435, 0.002368096, 
    0.001053717, 0.001967233, 0.001591717, 0.004825801, 0.002795054, 
    0.001965373, 0.002647904, 0.006410638, 0.01477892, 0.05952598, 0.2075087, 
    0.1303744, 0.008119494, 0.0007188009, 0.003418141, 0.0359043, 
    0.003586546, 0.01007394,
  7.63377e-06, 9.339807e-08, 5.75149e-06, 0.01195357, 0.06587555, 
    0.004687021, -0.0009628023, 0.004050895, 0.007021004, 0.002072443, 
    0.0062949, 0.001114798, 0.002763049, 0.008676931, 0.004282316, 
    0.002317502, 0.007556725, 0.01450891, 0.05377251, 0.02158443, 0.03135787, 
    0.006652848, 0.2339174, 0.04713363, 0.004995236, 0.006003979, 
    0.001500609, 0.00544259, 1.510199e-08,
  1.392134e-07, 6.398661e-10, 1.54285e-06, 0.003347982, 0.002177356, 
    0.004121319, 0.007259873, 0.003627406, 0.0370377, 0.01337572, 0.0035915, 
    0.002136925, 0.007066079, 0.01197863, 0.001559115, 0.001180441, 
    0.003444052, 0.01297573, 0.02130605, 0.02897397, 0.0163952, 0.09653617, 
    0.0006008316, 0.009198776, 0.0008403151, 0.003948208, 0.00343767, 
    0.0004183347, 1.510222e-07,
  -7.563699e-06, 0.01986444, 0.0008267103, 0.01754344, 0.06582906, 
    -8.268415e-06, 0.001163226, 0.003670984, 0.1127221, 0.004770802, 
    0.01312355, 0.05930295, 0.05144041, 0.0193563, 0.08493094, 0.0279124, 
    0.0203476, 0.04544555, 0.05548082, 0.006036842, 0.0186546, 0.05500958, 
    0.1359167, 0.02095246, 0.01428393, 0.03499004, 0.002462011, 0.004035129, 
    0.01206997,
  0.01113027, 0.0175754, 0.06199561, 0.1216928, 0.01357182, 0.001436952, 
    0.08915095, 0.001737905, -9.024872e-05, 0.01040122, 0.2075995, 
    0.05904552, 0.1030012, 0.08436875, 0.1209929, 0.1096054, 0.1576632, 
    0.1476362, 0.1520342, 0.08884066, 0.0144983, 0.06391218, 0.1156012, 
    0.1239333, 0.07481883, 0.09655405, 0.09098758, 0.1056888, 0.05411223,
  0.1417609, 0.2424365, 0.2868903, 0.3919372, 0.2611153, 0.1866017, 
    0.0828132, 0.256435, 0.05389892, 0.1201001, 0.04682169, 0.2072302, 
    0.07637081, 0.1152151, 0.08980501, 0.08143657, 0.07852019, 0.1808536, 
    0.1749244, 0.4353419, 0.1651362, 0.1517634, 0.1910509, 0.6909576, 
    0.2240767, 0.182055, 0.1361132, 0.1119962, 0.1298838,
  0.04196582, 0.4413915, 0.4041454, 0.7521293, 0.7399291, 0.4045545, 
    0.6390129, 0.5722325, 0.6103994, 0.4446713, 0.4628735, 0.5002702, 
    0.1027444, 0.2290987, 0.166321, 0.1269937, 0.3468936, 0.2330256, 
    0.3105778, 0.29113, 0.7961084, 0.2696386, 0.1395696, 0.4050821, 
    0.1784782, 0.09152855, 0.09384485, 0.07718318, 0.05075845,
  0.0379543, 0.03240044, 0.3579492, 0.04544342, 0.1465091, 0.2807558, 
    0.5712069, 0.3160528, 0.3597573, 0.4942759, 0.4333235, 0.4070133, 
    0.4027653, 0.5947416, 0.4671496, 0.3150438, 0.4266126, 0.3898056, 
    0.3907559, 0.3842528, 0.4881113, 0.515349, 0.3955016, 0.4642824, 
    0.138636, 0.3050954, 0.1764902, 0.1036939, 0.03185603,
  0.4186095, 0.3712187, 0.4097867, 0.3113168, 0.2757092, 0.417524, 0.4708964, 
    0.4927526, 0.4779411, 0.5407276, 0.4799243, 0.4533557, 0.5571993, 
    0.590549, 0.6015978, 0.6132125, 0.5842729, 0.6689127, 0.6888292, 
    0.609286, 0.4474809, 0.2380734, 0.3584931, 0.2690894, 0.2345999, 
    0.3963959, 0.2114609, 0.2807726, 0.4489134,
  0.5832077, 0.5919046, 0.6006016, 0.6092986, 0.6179956, 0.6266926, 
    0.6353896, 0.5531633, 0.5515543, 0.5499452, 0.5483361, 0.546727, 
    0.5451179, 0.5435088, 0.6579689, 0.6558507, 0.6537325, 0.6516144, 
    0.6494962, 0.647378, 0.6452599, 0.5956612, 0.5906914, 0.5857217, 
    0.580752, 0.5757823, 0.5708126, 0.5658429, 0.5762501,
  0.01817741, 0.07435265, 0.05348718, 0.1959299, 0.3522601, 0.2216547, 
    0.2452363, 0.255787, 0.3005215, 0.2403078, 0.1610994, 0.07935011, 
    0.07654684, 0.006797125, 0.1584587, 0.2138886, 0.1884959, 0.1291978, 
    0.1077568, 0.108835, 0.1030353, 0.192271, 0.3182235, 0.09703585, 
    0.1053334, 0.1784346, 0.01206634, 0.01090358, 0.01262981,
  0.1157111, 0.06131002, 0.06686924, 0.0322125, 0.09282902, 0.1324972, 
    0.002981488, 0.03512384, 0.09041659, 0.06301153, 0.03729506, 0.04630097, 
    0.02894228, 0.1257585, 0.2480718, 0.227746, 0.2294541, 0.2213826, 
    0.3483595, 0.229288, 0.2776699, 0.2141939, 0.2181465, 0.3203303, 
    0.07983416, 0.2303355, 0.2078886, 0.1436817, 0.1719959,
  0.2631725, 0.2131721, 0.3030171, 0.2729458, 0.2846628, 0.2761163, 
    0.3357675, 0.3089306, 0.3417187, 0.1953503, 0.2837501, 0.3465705, 
    0.3449378, 0.2541155, 0.2994038, 0.3861038, 0.4746358, 0.4847118, 
    0.3458765, 0.1954967, 0.173837, 0.1448794, 0.1851212, 0.2938867, 
    0.3163615, 0.4364627, 0.4413853, 0.3970696, 0.3316344,
  0.3083839, 0.3034305, 0.269074, 0.2322476, 0.2120855, 0.2100855, 0.2656164, 
    0.2094049, 0.2208102, 0.2392504, 0.1219408, 0.1138064, 0.05248362, 
    0.12142, 0.2031628, 0.21187, 0.2619185, 0.2433543, 0.2824745, 0.2380908, 
    0.1874491, 0.2682463, 0.1971477, 0.05987057, 0.04229439, 0.2708418, 
    0.3399112, 0.3017358, 0.3816066,
  0.09391388, 0.03616125, 0.008959132, 0.0683134, 0.09532169, 0.08481573, 
    0.08397368, 0.1218541, 0.1338716, 0.06381508, 0.0300298, 0.01057135, 
    0.004132201, 0.1044356, 0.2607394, 0.2228914, 0.2284372, 0.2266864, 
    0.2085684, 0.1238518, 0.2725055, 0.1158682, 0.107382, 0.104997, 
    0.04120146, 0.1972501, 0.1986683, 0.263203, 0.1730181,
  0.01218499, 0.01372011, 0.008047873, 0.1305654, 0.1119349, 0.01955572, 
    0.03333058, 0.01240538, 0.03946765, 0.003130565, 0.000214253, 
    3.320657e-07, 0.002276036, 0.06845251, 0.03017116, 0.01403397, 
    0.02657033, 0.02857985, 0.0273897, 0.02639955, 0.01129055, 0.00461016, 
    0.02504361, 0.02115587, 0.006908188, 0.01577606, 0.08052942, 0.03010583, 
    0.005095008,
  0.02369638, 0.00684544, -3.575861e-05, 0.005875653, 0.0009982579, 
    0.002424735, 0.002622371, 0.005493823, 0.02274234, 2.167834e-05, 
    2.550516e-08, 3.290992e-08, 0.005466346, 0.003635373, 0.008769206, 
    0.007911996, 0.0005508211, 0.003412828, 0.001746334, 0.003157117, 
    0.001182456, 0.008650879, 0.04131927, 0.02915088, 0.007045995, 0.1654837, 
    0.00894089, 0.0006386756, 0.006253063,
  0.04540952, 0.01332656, 0.0005250893, 0.1567915, 0.0004879987, 0.001012537, 
    0.0009768882, 0.0001873871, 0.00354482, 0.006240201, 0.001456042, 
    0.004941873, 0.003674543, 9.552891e-05, 0.006766213, 0.004077494, 
    0.0001758762, 0.0005344882, 0.000973767, 0.001172121, 0.004367027, 
    0.0134428, 0.08593509, 0.009595154, 0.002109074, 0.0001379818, 
    -0.0006790681, 0.0005076843, 0.01470968,
  0.008794845, 0.1395696, 0.006182254, 0.1227314, 0.001636063, 0.002614343, 
    0.001902343, 0.002965938, 0.09269403, 0.02452903, 0.001177197, 
    0.0004638744, 0.0008956824, 0.0007854693, 0.002596807, 0.00147445, 
    0.001001121, 0.001144089, 0.002744536, 0.005393128, 0.02136523, 
    0.08684611, 0.06533761, 0.007957246, 0.0005000154, 0.001249012, 
    0.02039708, 0.0003157798, 0.002265553,
  3.708039e-06, -4.513516e-08, 9.001725e-06, 0.01084349, 0.04095326, 
    0.002674954, -0.002788359, 0.001599717, 0.002579093, 0.0008478342, 
    0.002482732, 0.0002557851, 0.0007918002, 0.002869311, 0.001343599, 
    0.0006313947, 0.003341363, 0.004951128, 0.02933027, 0.007738843, 
    0.01284839, 0.002185584, 0.1882889, 0.04562528, 0.001962075, 0.002567902, 
    0.0008841756, 0.00291577, 4.941654e-07,
  1.359159e-07, 5.959805e-10, 1.459945e-06, 0.002174589, 0.00234837, 
    0.002423905, 0.008722234, 0.002222739, 0.02914846, 0.006250423, 
    0.001170512, 0.0008929145, 0.002871776, 0.00394817, 0.0003975024, 
    0.0005456924, 0.001103185, 0.004313671, 0.008919697, 0.01715208, 
    0.008812527, 0.07754613, 0.0003906843, 0.003038665, 0.0001785244, 
    0.001793665, 0.001994702, 0.0002374658, 1.542056e-07,
  -1.68055e-05, 0.0138856, 0.0006219922, 0.01270404, 0.0524888, 
    -6.757641e-06, 0.001557591, 0.005038592, 0.09782966, 0.00295029, 
    0.007852804, 0.03944457, 0.03272425, 0.005353861, 0.05468575, 0.0130226, 
    0.009617585, 0.02415512, 0.03073853, 0.003587519, 0.01372379, 0.04613099, 
    0.1207372, 0.01432812, 0.005514939, 0.02170352, 0.0009514263, 
    0.002274072, 0.01007039,
  0.00692313, 0.008169807, 0.03733281, 0.11087, 0.007741392, 0.0004884826, 
    0.08697148, 0.00211222, -6.435355e-05, 0.009093613, 0.2010384, 
    0.04016827, 0.08416977, 0.06525015, 0.08617543, 0.08420128, 0.1245254, 
    0.1242038, 0.1007763, 0.08096237, 0.01121669, 0.05997565, 0.09351522, 
    0.09541458, 0.05301047, 0.06579216, 0.05198367, 0.05829467, 0.03389382,
  0.1023161, 0.1910729, 0.23024, 0.3728947, 0.2308555, 0.1600063, 0.0568054, 
    0.2257378, 0.04995482, 0.09298459, 0.03918251, 0.1883772, 0.06099598, 
    0.08802646, 0.06350003, 0.0574657, 0.05239075, 0.1422319, 0.1255421, 
    0.4329532, 0.1409539, 0.1126594, 0.1550494, 0.6408596, 0.1706872, 
    0.1612034, 0.1070826, 0.0825121, 0.1102982,
  0.01980263, 0.4465335, 0.3712858, 0.6747268, 0.6861616, 0.3495342, 
    0.5779703, 0.5607006, 0.554359, 0.4139777, 0.4459967, 0.4897353, 
    0.09410699, 0.2022998, 0.1312031, 0.09446278, 0.3833461, 0.191108, 
    0.2613348, 0.2825403, 0.7895228, 0.2193311, 0.0859374, 0.3355862, 
    0.1360146, 0.08390943, 0.07012707, 0.04845893, 0.02880582,
  0.02747811, 0.01606841, 0.3292477, 0.025654, 0.1089664, 0.2139778, 
    0.5679839, 0.3003798, 0.348956, 0.5177178, 0.4938309, 0.4395183, 
    0.3977499, 0.6160576, 0.4333076, 0.3685608, 0.3571355, 0.334594, 
    0.3863567, 0.320621, 0.5079765, 0.6073003, 0.3670456, 0.5355252, 
    0.1146505, 0.2959741, 0.1924813, 0.07841257, 0.02205944,
  0.4654299, 0.3454972, 0.4610058, 0.3360422, 0.304699, 0.4923871, 0.5478718, 
    0.5569605, 0.6021491, 0.6361788, 0.5627686, 0.488355, 0.5743584, 
    0.6135158, 0.6162519, 0.6469944, 0.6186415, 0.6453228, 0.6781994, 
    0.6464298, 0.4648548, 0.2025831, 0.4134836, 0.3138914, 0.2055477, 
    0.3833747, 0.2177672, 0.305369, 0.4446163,
  0.5544297, 0.5636647, 0.5728997, 0.5821348, 0.5913698, 0.6006048, 
    0.6098399, 0.4714868, 0.4733148, 0.4751428, 0.4769708, 0.4787988, 
    0.4806268, 0.4824548, 0.6844622, 0.6782088, 0.6719555, 0.6657021, 
    0.6594487, 0.6531954, 0.646942, 0.5911862, 0.5863765, 0.5815669, 
    0.5767572, 0.5719475, 0.5671378, 0.5623282, 0.5470416,
  0.02246189, 0.07595833, 0.0390124, 0.186293, 0.3499193, 0.1897414, 
    0.1995258, 0.2441196, 0.2190179, 0.1671209, 0.09694728, 0.04711133, 
    0.06365385, 0.006817487, 0.1969266, 0.2101898, 0.176468, 0.1349124, 
    0.07494012, 0.1358184, 0.0765213, 0.1892529, 0.2594839, 0.06639899, 
    0.08462636, 0.1621045, 0.006329128, 0.01022132, 0.005100579,
  0.08119521, 0.04964827, 0.06484248, 0.02566019, 0.07239655, 0.0923994, 
    0.001222357, 0.02809473, 0.0654726, 0.04273695, 0.02660564, 0.04988976, 
    0.02018799, 0.1010998, 0.234267, 0.1923272, 0.1970744, 0.1840312, 
    0.2822008, 0.2070433, 0.2390831, 0.1785271, 0.1652915, 0.2631976, 
    0.07775919, 0.1769188, 0.1458615, 0.09709952, 0.1312223,
  0.1934417, 0.1727396, 0.2276973, 0.1831721, 0.1936719, 0.1963439, 
    0.2361363, 0.2387859, 0.269297, 0.139773, 0.213537, 0.2693874, 0.2583728, 
    0.2126966, 0.2335361, 0.2973718, 0.3806832, 0.3713422, 0.269969, 
    0.1570914, 0.1375842, 0.1016716, 0.1279277, 0.2110128, 0.2603898, 
    0.3713804, 0.3509876, 0.3137971, 0.2405997,
  0.2649574, 0.2334734, 0.2076715, 0.1714478, 0.1479714, 0.163285, 0.2048424, 
    0.1511184, 0.1690015, 0.1881765, 0.08195023, 0.06751952, 0.02928937, 
    0.07586135, 0.1600478, 0.1517377, 0.1830815, 0.1717641, 0.2106242, 
    0.1615221, 0.1161562, 0.2005469, 0.1323759, 0.04702426, 0.03704577, 
    0.2332236, 0.2943433, 0.263533, 0.3366373,
  0.04825415, 0.01785272, 0.006159612, 0.04566111, 0.06097695, 0.05861915, 
    0.05635406, 0.07525143, 0.07351518, 0.03577693, 0.01759744, 0.006531809, 
    0.002642805, 0.08938262, 0.2296926, 0.1479671, 0.1588285, 0.197694, 
    0.1628141, 0.09695584, 0.2370831, 0.07528318, 0.07372328, 0.09320031, 
    0.03030456, 0.1487018, 0.120503, 0.1903542, 0.1289992,
  0.008694062, 0.009240652, 0.005186544, 0.06611015, 0.05773666, 0.005888149, 
    0.01412103, 0.006208047, 0.02279597, 0.00216111, 8.910603e-05, 
    1.978401e-07, 0.0006928452, 0.03611215, 0.01818641, 0.007157695, 
    0.0156655, 0.01763179, 0.01859391, 0.01490352, 0.005769683, 0.002470322, 
    0.01754063, 0.01390039, 0.004843927, 0.008036632, 0.04067435, 0.01363941, 
    0.00330785,
  0.01526794, 0.005905137, -2.447813e-05, 0.003556834, 0.0006855731, 
    0.001587309, 0.001493503, 0.003432208, 0.01442298, -6.957599e-06, 
    2.366908e-08, 2.69275e-08, 0.002768441, 0.001684721, 0.004509383, 
    0.003412743, 0.0002395339, 0.00141959, 0.0006351457, 0.00139517, 
    0.000667981, 0.005626905, 0.02618414, 0.01888229, 0.005658725, 0.1425782, 
    0.00326971, 0.0003968573, 0.003560376,
  0.02799381, 0.00226025, 0.0004611652, 0.1183316, 0.0002265929, 
    0.0004665749, 0.0006131624, 0.0001133523, 0.002284511, 0.004255579, 
    0.0006408815, 0.002502095, 0.001541482, -2.425435e-06, 0.003557252, 
    0.001661398, 0.0001198399, 0.000333291, 0.0006506369, 0.0007826617, 
    0.002851512, 0.008490631, 0.05359628, 0.01122808, 0.001253875, 
    5.751532e-06, -0.0002058387, 0.0003082087, 0.009028568,
  0.003168178, 0.1123628, 0.005554353, 0.09746917, 0.0009222876, 0.001601555, 
    0.001147431, 0.001780133, 0.08648103, 0.02466155, 0.0005534173, 
    0.0002829533, 0.0005435614, 0.0005031898, 0.001670998, 0.0009594288, 
    0.0006442092, 0.000686431, 0.001672132, 0.002978545, 0.01115229, 
    0.04954597, 0.04015774, 0.008291307, 0.0002442927, 0.0006970527, 
    0.009861254, 9.770406e-05, 0.001159659,
  -2.912556e-06, -1.571631e-07, 3.858363e-06, 0.01170572, 0.0275178, 
    0.001803275, -0.002707454, 0.0005627008, 0.0006437468, 0.0005544729, 
    0.0008531389, 0.0001047929, 0.000416523, 0.001096857, 0.0005138669, 
    0.0002211826, 0.00143816, 0.001974552, 0.01233028, 0.003914854, 
    0.004822489, 0.001327456, 0.1496208, 0.04100558, 0.0008719739, 
    0.00107369, 0.000619789, 0.001850699, 2.156208e-07,
  1.315274e-07, 5.97277e-10, 1.323323e-06, 0.001314736, 0.0008161277, 
    0.001667496, 0.01421822, 0.001535121, 0.01702643, 0.003466197, 
    0.0006726215, 0.0005711046, 0.001295895, 0.00130295, 0.0002272414, 
    0.0003093999, 0.0006137908, 0.002308228, 0.004863173, 0.01195089, 
    0.005072565, 0.05957036, 0.0002849912, -0.0002985057, 0.0001085339, 
    0.000996289, 0.001336604, 0.0001581172, 1.567645e-07,
  -1.464873e-05, 0.007319819, 0.0007309491, 0.009305967, 0.03814709, 
    -2.744933e-06, 0.0008218344, 0.009996264, 0.0874696, 0.001278521, 
    0.005639288, 0.02123174, 0.0139318, 0.002596172, 0.02792208, 0.006384313, 
    0.005507697, 0.008924023, 0.01741171, 0.002175223, 0.01014532, 
    0.04021192, 0.1001966, 0.003460194, 0.002545251, 0.01011969, 
    0.0004890896, 0.001602181, 0.007719534,
  0.005244329, 0.004157863, 0.02351871, 0.1076357, 0.004980452, 0.000261565, 
    0.08280392, 0.002061747, -4.560662e-05, 0.007200086, 0.1819839, 
    0.02730448, 0.06303272, 0.04875363, 0.05576453, 0.05664218, 0.09457535, 
    0.09639163, 0.06089089, 0.07363555, 0.01074925, 0.05033657, 0.07493152, 
    0.07416955, 0.03197301, 0.03671431, 0.02562941, 0.02869123, 0.02048289,
  0.06641612, 0.1574326, 0.178649, 0.3133422, 0.1898681, 0.141644, 
    0.04111348, 0.1940595, 0.05806513, 0.07267112, 0.03664774, 0.1645334, 
    0.04772573, 0.06696898, 0.04496614, 0.03866694, 0.03619726, 0.09966629, 
    0.07455085, 0.4104302, 0.1183837, 0.0892961, 0.1159559, 0.5728034, 
    0.1323665, 0.1409506, 0.07590315, 0.0509092, 0.0768658,
  0.01021955, 0.4348211, 0.3545808, 0.5797157, 0.6187788, 0.2944569, 
    0.4942597, 0.4819915, 0.4562206, 0.3819059, 0.3903591, 0.4802857, 
    0.1302797, 0.2075818, 0.1058912, 0.07413501, 0.4099853, 0.1551548, 
    0.2070788, 0.2770539, 0.7343352, 0.1644842, 0.05823364, 0.2907928, 
    0.1043841, 0.07609943, 0.05280848, 0.03122763, 0.01683846,
  0.02046916, 0.01011062, 0.3035629, 0.01710585, 0.08347437, 0.1720479, 
    0.5425104, 0.3332469, 0.3432842, 0.5051317, 0.5604313, 0.4082356, 
    0.4192411, 0.5019594, 0.3184173, 0.3064428, 0.3070415, 0.2727225, 
    0.3972804, 0.2753262, 0.4979254, 0.6638804, 0.3677015, 0.569623, 
    0.09522738, 0.2856444, 0.2658542, 0.05754118, 0.01683443,
  0.4366187, 0.314071, 0.4987378, 0.3182368, 0.3781623, 0.5079358, 0.5513912, 
    0.5434912, 0.5623794, 0.6246262, 0.6112482, 0.5376732, 0.6077569, 
    0.5968577, 0.5342801, 0.628857, 0.5550236, 0.5659806, 0.6284083, 
    0.5978205, 0.457542, 0.1713106, 0.441497, 0.3876595, 0.1942701, 
    0.3286824, 0.2088003, 0.303412, 0.3879924,
  0.404533, 0.4135377, 0.4225424, 0.4315471, 0.4405518, 0.4495565, 0.4585612, 
    0.3401125, 0.3388367, 0.3375608, 0.336285, 0.3350092, 0.3337334, 
    0.3324575, 0.5034011, 0.4985001, 0.4935992, 0.4886982, 0.4837973, 
    0.4788963, 0.4739954, 0.4302703, 0.4274424, 0.4246144, 0.4217865, 
    0.4189586, 0.4161307, 0.4133028, 0.3973292,
  0.03188274, 0.06713018, 0.03659197, 0.1509768, 0.3281984, 0.1597642, 
    0.1510459, 0.1974344, 0.1639421, 0.1191126, 0.06420071, 0.02785518, 
    0.05470951, 0.00674881, 0.2413464, 0.1950635, 0.1533296, 0.1315202, 
    0.06500079, 0.1452391, 0.06359366, 0.1726727, 0.2221684, 0.05544571, 
    0.07793046, 0.1411013, 0.007372138, 0.009599404, 0.0002188764,
  0.06706166, 0.04378051, 0.06741818, 0.01977738, 0.05827097, 0.07755157, 
    0.0008414881, 0.02259564, 0.05779364, 0.03262698, 0.02228944, 0.04661413, 
    0.01149946, 0.09009903, 0.2073101, 0.1690461, 0.1613018, 0.1553947, 
    0.219212, 0.1804331, 0.194268, 0.1347047, 0.1304697, 0.2156948, 
    0.06915869, 0.1357173, 0.1101427, 0.0763473, 0.0990373,
  0.1466497, 0.1370502, 0.1831759, 0.1411507, 0.144585, 0.1549208, 0.1832546, 
    0.1837213, 0.2103316, 0.1125515, 0.1662828, 0.2189145, 0.1948278, 
    0.175773, 0.1847427, 0.2358539, 0.3047852, 0.3103886, 0.2176115, 
    0.1246937, 0.1132808, 0.07663516, 0.09579049, 0.1582497, 0.2103201, 
    0.3038816, 0.2835127, 0.2596179, 0.1962615,
  0.2187418, 0.1892859, 0.173785, 0.1315875, 0.1137077, 0.1387644, 0.1658788, 
    0.1137889, 0.1270907, 0.1367025, 0.0535459, 0.04581372, 0.01914598, 
    0.04992234, 0.117756, 0.1064277, 0.1292593, 0.1213021, 0.1559974, 
    0.1068547, 0.08001175, 0.1458231, 0.09692596, 0.04046657, 0.03019756, 
    0.1865498, 0.2467259, 0.2145505, 0.2914737,
  0.02933352, 0.01083577, 0.004788053, 0.03024083, 0.03907651, 0.04177129, 
    0.03475795, 0.04812154, 0.04384641, 0.02197507, 0.01106975, 0.004790679, 
    0.001899376, 0.06542332, 0.2007662, 0.09830962, 0.1124946, 0.1346416, 
    0.1214958, 0.0696544, 0.1753852, 0.04916226, 0.05082614, 0.0795755, 
    0.02592652, 0.1078717, 0.07430502, 0.1331181, 0.08233918,
  0.006850641, 0.007145641, 0.003586566, 0.03756024, 0.0333703, 0.003009193, 
    0.008345575, 0.004038579, 0.01614451, 0.001657629, 4.682222e-05, 
    1.394226e-07, -0.0003207821, 0.02192799, 0.009735853, 0.004408262, 
    0.008960699, 0.009680714, 0.01215869, 0.008822349, 0.003243128, 
    0.001812987, 0.0136367, 0.01010495, 0.003786349, 0.003715898, 0.02171823, 
    0.009904654, 0.002659391,
  0.01126724, 0.003310863, -1.566166e-05, 0.002420822, 0.0006560787, 
    0.001182232, 0.001073858, 0.00249737, 0.01061631, -6.802119e-06, 
    2.098745e-08, 2.604963e-08, 0.001843033, 0.001194336, 0.002198278, 
    0.002078404, 0.0001730579, 0.0008891128, 0.0003098454, 0.0007356027, 
    0.0004485093, 0.004167117, 0.01905478, 0.01415192, 0.004088365, 
    0.1211192, 0.001154734, 0.0002861261, 0.00242623,
  0.02012276, -0.002201175, 0.001121991, 0.08873373, 0.0001549521, 
    0.0002657344, 0.0004478758, 8.155359e-05, 0.001678173, 0.00321461, 
    0.0004161029, 0.00131377, 0.0009246432, 3.558837e-05, 0.001646803, 
    0.0008648385, 8.944501e-05, 0.0002414435, 0.000488203, 0.0005886804, 
    0.002112376, 0.006177582, 0.03903573, 0.0128109, 0.0009586613, 
    1.222852e-05, -6.83739e-05, 0.000219103, 0.006497455,
  0.001619787, 0.09426372, 0.003476867, 0.08570544, 0.0005803449, 
    0.001136246, 0.000834277, 0.00123955, 0.07817541, 0.02533756, 
    0.0003502168, 0.0002025236, 0.0003822338, 0.0003643123, 0.001216795, 
    0.0006852203, 0.0004754346, 0.0004773871, 0.001191275, 0.00201718, 
    0.007312767, 0.03439371, 0.02875775, 0.005701315, 0.0001106563, 
    0.0004744474, 0.004410287, 6.621493e-05, 0.0007847404,
  -9.462729e-07, -8.785594e-06, 6.510388e-07, 0.0148011, 0.02517045, 
    0.001366718, -0.002327098, 0.0002891427, 0.0003863132, 0.000420074, 
    0.0004882732, 9.294844e-05, 0.0002879105, 0.0006464255, 0.0002498697, 
    0.0001352853, 0.0007123747, 0.001055136, 0.005411985, 0.001878647, 
    0.00190165, 0.001028012, 0.1349533, 0.03356479, 0.0004685599, 
    0.0004833925, 0.0004685602, 0.001344319, 5.338657e-07,
  1.29191e-07, 6.069862e-10, 1.172905e-06, 0.0006999778, 0.0003487031, 
    0.00125193, 0.02139477, 0.001152872, 0.01194376, 0.002276846, 
    0.0004800904, 0.000434585, 0.0007502236, 0.0005640467, 0.0001687835, 
    0.0002193374, 0.0004419717, 0.001579067, 0.003475186, 0.009224323, 
    0.003301557, 0.04972483, 0.000228982, -0.0009677981, 8.600362e-05, 
    0.0006533641, 0.001006345, 0.0001187655, 1.56153e-07,
  -1.087677e-05, 0.005172332, 0.0002400264, 0.005796495, 0.0282837, 
    -6.973285e-07, 0.0002179206, 0.01340206, 0.08334005, 0.0008032696, 
    0.004477432, 0.01308781, 0.006390987, 0.001903691, 0.01493865, 
    0.003678672, 0.003787993, 0.00403876, 0.01135555, 0.001553959, 
    0.007882804, 0.03799202, 0.0812788, 0.00165964, 0.001644387, 0.004810876, 
    0.000338169, 0.001227757, 0.006829056,
  0.006925646, 0.002490929, 0.01503617, 0.1079308, 0.0037626, 0.0001769008, 
    0.07722668, 0.001244718, -3.532243e-05, 0.005575574, 0.1580679, 
    0.02020578, 0.04693687, 0.03357638, 0.03444315, 0.03809154, 0.07640561, 
    0.06245998, 0.04036403, 0.06857237, 0.009526072, 0.04537985, 0.05794509, 
    0.06002061, 0.0204322, 0.0200899, 0.01434991, 0.01505091, 0.01338965,
  0.04642345, 0.1414535, 0.1493881, 0.2784774, 0.1640832, 0.1360612, 
    0.03254369, 0.1865059, 0.08857883, 0.05966653, 0.03060155, 0.1583725, 
    0.03584456, 0.055343, 0.03404408, 0.02794567, 0.02753848, 0.07351257, 
    0.04640635, 0.4004728, 0.1051124, 0.07116041, 0.09503862, 0.5060599, 
    0.1092418, 0.1211013, 0.05424815, 0.03144028, 0.05132399,
  0.006761482, 0.3986066, 0.3352476, 0.5092816, 0.570246, 0.2613828, 
    0.4388475, 0.4233055, 0.3699217, 0.3343331, 0.3336272, 0.4875947, 
    0.1888204, 0.2298891, 0.08985828, 0.06291916, 0.4197384, 0.1484655, 
    0.1845854, 0.267057, 0.6652436, 0.164816, 0.04480045, 0.2703451, 
    0.0905833, 0.06783628, 0.04141039, 0.0236161, 0.01198128,
  0.01548113, 0.007338319, 0.3083523, 0.01318096, 0.06785716, 0.1454544, 
    0.5104456, 0.3968716, 0.3413801, 0.4603032, 0.5729623, 0.381197, 
    0.3818927, 0.3909759, 0.2211774, 0.244179, 0.2853287, 0.2231371, 
    0.3608851, 0.2378479, 0.4226423, 0.6016153, 0.4109909, 0.5736012, 
    0.07886291, 0.2696677, 0.3997082, 0.05081422, 0.01403492,
  0.424664, 0.2904213, 0.522965, 0.3057417, 0.3526709, 0.4665697, 0.4541669, 
    0.4078532, 0.4367971, 0.4926053, 0.3954844, 0.364894, 0.4055783, 
    0.4735698, 0.4150126, 0.4761184, 0.3825057, 0.4246656, 0.4782689, 
    0.447173, 0.3581946, 0.1565607, 0.4390189, 0.4736615, 0.1980376, 
    0.2951558, 0.2134119, 0.2911451, 0.3077126,
  0.2443429, 0.2501571, 0.2559713, 0.2617855, 0.2675997, 0.2734139, 
    0.2792281, 0.2261515, 0.2273843, 0.2286171, 0.2298499, 0.2310827, 
    0.2323155, 0.2335483, 0.3322822, 0.3274045, 0.3225267, 0.3176489, 
    0.3127711, 0.3078934, 0.3030156, 0.3251198, 0.3229506, 0.3207814, 
    0.3186122, 0.3164429, 0.3142737, 0.3121045, 0.2396916,
  0.0532366, 0.06128776, 0.0398071, 0.1250742, 0.2909491, 0.1535531, 
    0.1342438, 0.1902721, 0.1287282, 0.09677317, 0.05515045, 0.02004647, 
    0.04091067, 0.006785051, 0.2933979, 0.1809669, 0.1557664, 0.1510083, 
    0.06016261, 0.1695102, 0.06361301, 0.1601085, 0.195864, 0.04995645, 
    0.09173868, 0.1322234, 0.01099657, 0.01124761, -0.00259487,
  0.06169213, 0.04297743, 0.07459426, 0.01755147, 0.05333743, 0.07499524, 
    0.0007857122, 0.01810555, 0.05099572, 0.02620659, 0.02142322, 0.04887532, 
    0.008915183, 0.09512974, 0.212312, 0.158364, 0.1419391, 0.1391152, 
    0.1884309, 0.158859, 0.1755357, 0.1187096, 0.1135668, 0.187467, 
    0.06574107, 0.1206938, 0.09535076, 0.06638724, 0.08256303,
  0.1242331, 0.1199672, 0.1569718, 0.1221987, 0.1184502, 0.1287582, 
    0.1498856, 0.1574039, 0.1768544, 0.09428657, 0.1420497, 0.1857009, 
    0.1569906, 0.1478868, 0.1551551, 0.1955709, 0.2537073, 0.2716862, 
    0.188359, 0.1071438, 0.09637419, 0.06395038, 0.07977621, 0.1308254, 
    0.1761732, 0.2603143, 0.2495002, 0.2292218, 0.1716581,
  0.1875257, 0.1626128, 0.150116, 0.1109491, 0.09380273, 0.1222665, 
    0.1365181, 0.09214523, 0.1068561, 0.110198, 0.03902065, 0.03600474, 
    0.01449673, 0.03874881, 0.09397846, 0.07944535, 0.09324894, 0.08863141, 
    0.1249366, 0.07983185, 0.06187729, 0.1152244, 0.08081143, 0.04410493, 
    0.02722074, 0.1516973, 0.2013667, 0.179665, 0.2478598,
  0.02173607, 0.008053299, 0.004097063, 0.02144384, 0.02841607, 0.03089008, 
    0.02319545, 0.03467642, 0.03056956, 0.01575977, 0.008193732, 0.004006009, 
    0.001556005, 0.04907605, 0.2010106, 0.0704044, 0.08005912, 0.093849, 
    0.0934998, 0.04898118, 0.1309652, 0.03446699, 0.04094863, 0.0743534, 
    0.02198446, 0.07617696, 0.05015851, 0.09626435, 0.05814627,
  0.005893665, 0.006055109, 0.009882268, 0.02711299, 0.02083876, 0.002318462, 
    0.006034258, 0.003489769, 0.01297462, 0.001384129, 3.133016e-05, 
    1.08171e-07, 0.001600673, 0.01589314, 0.005738727, 0.003369611, 
    0.005514916, 0.00579965, 0.007989654, 0.006042797, 0.00208736, 
    0.001487971, 0.01153634, 0.008718658, 0.00409742, 0.002513412, 
    0.01401106, 0.006089248, 0.002313859,
  0.009361136, 0.002711187, -1.772196e-05, 0.0018615, 0.0004236709, 
    0.0009836507, 0.0008240542, 0.002061494, 0.008783706, -5.983387e-06, 
    2.051829e-08, 2.542479e-08, 0.001453258, 0.0009713486, 0.001444358, 
    0.001549903, 0.0001421337, 0.0006916429, 0.0002134135, 0.0005174191, 
    0.0003526611, 0.003475395, 0.01571602, 0.01172187, 0.007332616, 
    0.1529544, 0.0006782598, 0.0002358118, 0.001947833,
  0.01634846, -0.003748025, 0.008365578, 0.0822876, 0.0001273642, 
    0.0001958433, 0.0003668468, 6.69517e-05, 0.001391335, 0.002182561, 
    0.0003282056, 0.0008408975, 0.0006850889, 4.495444e-05, 0.001006501, 
    0.0005841076, 7.313497e-05, 0.0001963388, 0.0004063711, 0.00049221, 
    0.001754754, 0.005080597, 0.03186605, 0.02947309, 0.001452239, 
    0.001956219, -2.120259e-05, 0.0001793955, 0.005317023,
  0.001130306, 0.1058394, 0.00354729, 0.0897412, 0.0004570062, 0.000908024, 
    0.0006758761, 0.0009773723, 0.105731, 0.05169579, 0.0002794745, 
    0.0001624874, 0.0002877639, 0.0002941311, 0.0009853655, 0.000560291, 
    0.0003926378, 0.0003819742, 0.000958218, 0.001597412, 0.005584589, 
    0.02717886, 0.02318778, 0.03849442, 0.002203133, 0.000370413, 
    0.002504595, 5.568388e-05, 0.0006185493,
  -4.414467e-05, -0.0001101804, -3.738338e-07, 0.03035745, 0.02198724, 
    0.001153632, -0.00204086, 0.0002143014, 0.0002612804, 0.0003527743, 
    0.0003801237, 8.523659e-05, 0.0002112134, 0.0004825712, 0.0001809048, 
    0.0001029383, 0.000527061, 0.0007514991, 0.002976231, 0.001084158, 
    0.00111237, 0.0008650143, 0.1724851, 0.03457468, 0.0003580239, 
    0.000332947, 0.0003389265, 0.001093843, 8.406123e-06,
  1.294102e-07, 6.14266e-10, -1.284601e-07, 0.0004523542, 0.0002009987, 
    0.001037468, 0.02787185, 0.0009215206, 0.01200716, 0.001447451, 
    0.0004291077, 0.000369393, 0.0005533769, 0.0003627505, 0.0001428394, 
    0.0001793541, 0.0003646353, 0.001257447, 0.002859107, 0.007800385, 
    0.002593784, 0.04696348, 0.0002020418, -0.001257083, 7.208325e-05, 
    0.0005028471, 0.0008475562, 0.0001004961, 1.5817e-07,
  -7.111457e-06, 0.004309462, 0.0006068107, 0.004426989, 0.02751585, 
    -3.554725e-07, -0.0001023532, 0.02045641, 0.09012705, 0.0006212911, 
    0.003886989, 0.009486783, 0.003997087, 0.001607456, 0.008293062, 
    0.002530377, 0.003034842, 0.002541749, 0.008196411, 0.001265657, 
    0.006191751, 0.03819336, 0.08406493, 0.001359684, 0.001295224, 
    0.003043072, 0.0002757231, 0.0009925768, 0.008790764,
  0.008995301, 0.001404461, 0.01137801, 0.1107869, 0.003113347, 0.0001335818, 
    0.07193965, 0.0008769089, -3.083806e-05, 0.004810564, 0.1577183, 
    0.01710678, 0.03878052, 0.02564951, 0.02455177, 0.02850339, 0.06239842, 
    0.04358158, 0.02988699, 0.06655622, 0.007938032, 0.04453583, 0.05874689, 
    0.04955391, 0.01481522, 0.01388662, 0.009583133, 0.01002723, 0.01239045,
  0.03486748, 0.1540816, 0.1532716, 0.2764867, 0.1554303, 0.1338982, 
    0.03015554, 0.2652683, 0.1439227, 0.05781233, 0.05762097, 0.1937949, 
    0.0299318, 0.05032621, 0.0290354, 0.02324338, 0.02318229, 0.06027338, 
    0.03480409, 0.4231735, 0.1053851, 0.06353797, 0.1111523, 0.4985421, 
    0.106374, 0.1012292, 0.04279355, 0.02201814, 0.03680339,
  0.005462385, 0.4124967, 0.3269178, 0.4886603, 0.5704494, 0.3037868, 
    0.441274, 0.4157863, 0.3598391, 0.3169014, 0.3103376, 0.524078, 
    0.2745871, 0.2770107, 0.08108909, 0.0571683, 0.4602936, 0.1563197, 
    0.2226393, 0.3094741, 0.6416934, 0.1954063, 0.03823333, 0.2995856, 
    0.08113042, 0.06131968, 0.03519276, 0.02056199, 0.009961819,
  0.01291262, 0.006267574, 0.3463863, 0.01098452, 0.05971183, 0.1316055, 
    0.4854892, 0.4414091, 0.3888857, 0.4513902, 0.6008368, 0.4393789, 
    0.402495, 0.3033208, 0.1796658, 0.2151967, 0.3058158, 0.198599, 
    0.3242067, 0.202765, 0.3573073, 0.5430873, 0.4143606, 0.5570827, 
    0.07069146, 0.2488125, 0.5197003, 0.0491881, 0.01268002,
  0.4492614, 0.2810862, 0.4854694, 0.2753496, 0.3165487, 0.3683237, 
    0.3542752, 0.3222934, 0.3473453, 0.3350908, 0.2736023, 0.2494418, 
    0.2922454, 0.3716282, 0.3345514, 0.391594, 0.3055272, 0.3257338, 
    0.3732746, 0.352824, 0.2888708, 0.1513844, 0.4583878, 0.5381601, 
    0.1991666, 0.2598725, 0.2268116, 0.3028871, 0.2682506,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2.035369e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0004559944, -3.937145e-05, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 1.800889e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, -3.287091e-05, 0.0005168325, 0, 0, 0, 0, 0, 2.70987e-05, 0, 0, 
    0, -1.742014e-05, 0, 0, 0, 0, 0, 0, 0, 0, -3.880469e-05, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0008951412, -0.0001154514, 0, 
    -2.539627e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -6.055576e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 8.061308e-05, 0, -3.402034e-05, 0, 0, 0, 0, 0, 0, -8.058232e-06, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0002229527, 0, 0, 0,
  0, 0, 0, 0, 0.0001095764, 0.002595317, -7.57428e-05, -9.854371e-06, 0, 0, 
    0, 0.0001798783, 0, 0, -2.195077e-06, -2.334628e-05, 0, 0, 0, 0, 0, 0, 0, 
    0, -0.0001018995, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -3.714435e-06, -1.960992e-05, 
    -1.90404e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0008584302, 4.143742e-05, 
    0.0004394028, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001258824, -0.0002863811, 0, -5.086977e-05, 
    0, 0, 0, 0, -1.568458e-05, 0, 0.001049196, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -3.122739e-05, 0, 0, 0, 0, 0, 0, 0, 0, 
    -7.587672e-06, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, -7.806105e-06, 0, 0,
  0, 0, 6.821541e-05, 0, -0.0001416483, 0, 0, 0, 0, 0, 0, -8.058232e-06, 0, 
    0, -2.539555e-06, 0, -6.958488e-06, 0, 0, 0, 0, 0, 0, 0, -3.980906e-05, 
    0.003846079, 0, 0, 0,
  0, 0, -2.430001e-05, 0, 0.000274413, 0.01108279, -9.910921e-05, 
    0.0001298263, 0, 0, 0, 0.0004897209, -1.123539e-05, 0, -4.172014e-06, 
    0.001269813, 0, -1.625438e-05, 0, 0, 0, 0, 0, 0, 0.0006697606, 0, 0, 0, 0,
  0, 0, 0, 0, -6.819164e-07, -1.691663e-05, 0.001872647, -7.493085e-05, 
    -2.923306e-05, -2.375209e-06, 0, 0, 1.800066e-05, -3.921985e-05, 
    -1.525024e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.002727781, 0.0002293094, 
    0.002692553, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001012976, 0.003587988, 0.003148673, 
    -9.081009e-06, -0.0002706352, -0.0001199609, -6.346301e-05, 0, 
    0.0005789567, -7.838094e-05, -7.904969e-05, 0.003816813, 0, 0, 0, 0, 0, 
    0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.43409e-05, 0.0004274588, 0, 0, 0, 0, 0, 0, 
    0, 0, -8.016109e-05, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -1.71915e-05, 0.0002404974, 0, 0,
  0, 0.0005525416, 0.0006223523, 0, -0.0003654164, 0, 0, 0, 0, 0, 0, 
    -8.058232e-06, 0, 0, -2.961557e-06, 0, -4.182822e-05, 0, 0, 0, 0, 0, 0, 
    0, 0.0001794857, 0.008232606, 0, 0, 0,
  0, 0, 0.002726616, 0, 0.0006574962, 0.0200262, 0.002039794, 0.001356715, 0, 
    0, 0, 0.002710771, -6.005486e-05, -5.989786e-05, -2.195733e-05, 
    0.002300579, 0.0003108154, -1.858428e-07, 0, 0, 0, 0, 0, -1.812667e-05, 
    0.005393077, 0, 0, 0, 0,
  0, 0, -1.545226e-10, 0, -6.765424e-06, -2.645253e-05, 0.00246748, 
    -0.0002227389, -0.0001023138, 0.0001476208, 0, -5.416658e-06, 
    -9.212796e-06, -5.882977e-05, 0.0005079589, 0, -1.009916e-05, 0, 0, 0, 0, 
    0, 0.0008913795, 3.580267e-05, 0.005559081, 0.0002099831, 0.005467258, 0, 0,
  0, 0, 0, 0, 0, 0, 0, -4.665813e-06, 0, 0.003580335, 0.005912163, 
    0.01064888, 0.0003680014, -0.000271607, -0.0001791132, -0.0002345868, 
    -0.0001429918, 0.001379275, -0.000124437, 0.001394716, 0.01678577, 0, 0, 
    0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6.425977e-05, 0.0006405271, 0, 0, 0, 0, 0, 0, 
    0.0008771936, 0, -0.0001559014, 0, -4.885277e-05, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0004695607, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.0001208151, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -9.907733e-06, -2.492103e-05, 0, 0, 
    -6.24009e-06, 0.0005132896, 0, -2.390788e-05, 0, 0, 0, 0, 0, 0, 
    -7.010981e-05, 0.003043511, 0, 0,
  0, 0.0007738483, 0.0009609332, 0, 0.0007542617, 2.375044e-05, 0, 0, 0, 0, 
    0, -3.944665e-05, -2.795559e-05, 0, -2.198378e-05, 0, -4.874172e-05, 0, 
    0, 0, 0, 0, 0, 0, 0.0006456791, 0.01133252, 0, 0, 0,
  0, 0, 0.002493368, -1.004786e-05, 0.003025208, 0.03936836, 0.008358356, 
    0.004015384, 0, 0, 0, 0.01054648, 0.0001375097, -0.0001201399, 
    4.758646e-06, 0.00713515, 0.002035847, 0.0003020327, 0, 0, 0, 0, 0, 
    -5.063819e-05, 0.006932309, -2.388576e-06, 0, 0, 0,
  0, 0, -8.491455e-07, 0, -2.798568e-05, -1.760308e-05, 0.005130193, 
    -0.0003729422, -0.0001594388, 0.000267692, 4.672314e-06, -6.116576e-05, 
    -0.0001007182, -9.208807e-05, 0.001008068, 0, -5.997354e-05, 0, 0, 0, 0, 
    0, 0.00382456, 0.0003939229, 0.00664996, 0.002705722, 0.0122306, 0, 0,
  0, 0, 0, 0, 0, 0, 0, -5.225099e-05, 0, 0.007273513, 0.01443017, 0.01948995, 
    0.002981839, -0.0005246954, -0.0001311444, -0.0001197091, 0.001236126, 
    0.002608887, 0.002516086, 0.002722668, 0.04508179, 0, 0, 0, 0, 
    -1.65284e-05, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.002189284, 0.002622165, 0, 0, 0, 0, 
    -6.554586e-06, 0, 0.00246087, -1.995355e-06, 0.001182912, 0, 
    -7.013187e-05, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3.847141e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, -4.73234e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, -9.816469e-06, -5.227466e-06, 0, 0, 0,
  0, 0, 0, 0, 0.001443719, 3.012697e-06, 0, 0, 0, 0, -5.675969e-05, 0, 0, 
    0.003281212, 0, -2.680297e-05, 0, 0, 0.001480213, 0, 0, 0, 0, 0, 
    0.002568404, 0, -3.957727e-05, 0, 0,
  0, 0, 0, 0.001674686, 0, 0.0001157191, -1.521656e-05, 0, 0, 0, 
    0.0002170751, 0.0004129252, 0.0001511878, 0.002143348, 0, 0.004109432, 
    0.001551095, -6.365958e-06, 0.001125165, 0, -8.706382e-06, 0, 0, 0, 
    -4.177781e-07, 0.004164485, 0.006256554, 0, 0,
  0, 0.002356931, 0.001441412, 0, 0.001792122, 5.704816e-05, -0.0001071897, 
    0, 0, 0, 0.0001498005, 1.776444e-05, -9.842323e-05, 0, 0.0009039291, 
    -2.861002e-05, 8.106139e-05, 0, 0, 0, 0, 0, 0, 0, 0.001766497, 
    0.01951364, -3.252182e-05, 0, 0,
  0, -4.064097e-05, 0.003129896, -0.0001014253, 0.01114463, 0.06205584, 
    0.01563371, 0.009883877, 0, -6.306319e-06, 0, 0.01315059, 4.020454e-05, 
    -0.0001259665, 0.0005546919, 0.01518941, 0.004407702, 0.000855968, 0, 0, 
    0, 0, 0, 0.000452741, 0.01240968, -2.465021e-05, 0, 0, 0,
  0, 0, 2.537962e-06, 0, -3.89958e-05, 0.0003065836, 0.007764616, 
    -0.0003743553, -0.0001245555, 0.006422822, 0.0003645304, -9.23471e-05, 
    -6.559455e-05, -0.0001891238, 0.002041267, 0, 0.0006379107, 0, 0, 0, 0, 
    0, 0.00838727, 0.0004535811, 0.007757646, 0.004831776, 0.02013155, 0, 0,
  0, 0, 0, 0, 0, 0, 0, -0.0002713485, 0, 0.01225354, 0.03331949, 0.03518049, 
    0.00558418, -0.000614011, 0.001886479, 0.0002041374, 0.004801897, 
    0.007329891, 0.01183228, 0.006894059, 0.08040992, 0, 3.591376e-05, 0, 0, 
    -5.350062e-05, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.02527078, 0.004434943, 0, 0, 0, 0, 
    -6.918953e-05, 7.591023e-05, 0.006266023, 3.959412e-05, 0.005317878, 0, 
    0.000394008, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -5.451076e-09, 0.0002019622, 0.0001753983, 0, 
    -2.027281e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.10388e-05, 0, 0.00100121, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.00126603, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.252192e-05, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0.0002437, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2.217836e-05, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, -4.879832e-05, 0.001305953, 0, 0, 0,
  0, 0, 0, -5.711585e-05, 0.006451403, 9.642785e-06, -9.201442e-05, 0, 0, 0, 
    0.001273173, 0.0002341638, 0.0002573402, 0.01998055, 0.0002123029, 
    -7.147458e-05, 0, -1.419561e-05, 0.003381266, 0.0004306634, 3.878123e-05, 
    0, 0, 0, 0.004729534, 0.000128713, 0.001207374, -1.131546e-05, 
    -7.14206e-06,
  0, 0, 0.0002084504, 0.01142471, 0, 0.01094928, 0.0004096995, 0, 0, 0, 
    0.005827912, 0.008770349, 0.0009179353, 0.003597739, 0, 0.01610036, 
    0.007660621, 0.002072755, 0.002175724, 0, -0.0001603738, 0, 0, 0, 
    -0.0001632382, 0.0134915, 0.01489016, 0, 0.002717857,
  0, 0.005525683, 0.004530138, 1.97734e-05, 0.01300323, 0.000793835, 
    -0.0002710394, -7.250292e-05, 0, 0, 0.0002207796, 0.001640703, 
    0.002240175, -9.361489e-06, 0.005866764, -0.0001290849, 0.0002969365, 
    -2.150435e-05, -8.212277e-06, 0, 0, 0, 0, -9.93175e-05, 0.00659831, 
    0.028082, 0.0009616418, 0, 0,
  0, -0.0003670656, 0.004745374, 2.58266e-05, 0.01852967, 0.09099255, 
    0.03068985, 0.02170069, -1.08114e-05, -5.625495e-05, -2.323653e-06, 
    0.02323578, 0.003933433, 0.0006917875, 0.00430538, 0.02362449, 
    0.01214412, 0.002993929, 0, 0, 0, 0, 0, 0.001974324, 0.01845776, 
    -1.708261e-06, 0, 0, 0,
  0, 0.0002650213, 0.0001689472, 0, 5.316757e-05, 0.004126392, 0.0153378, 
    0.00351911, 0.0002809282, 0.01357007, 0.002589279, 0.0006747541, 
    0.008470355, 0.001081327, 0.01065773, -4.431267e-07, 0.007872494, 
    -9.446329e-06, 0, 0, 0, 0, 0.01690506, 0.002047802, 0.009974284, 
    0.00793968, 0.02664783, -1.913837e-05, -7.728248e-06,
  0, 0, 0, 0, 0, 0, 0, 0.001113472, 0, 0.02274909, 0.0546671, 0.05868977, 
    0.009485868, 0.004490828, 0.006117046, 0.004000097, 0.01289352, 
    0.01514791, 0.03969996, 0.01902056, 0.118942, -3.618628e-05, 
    0.0001257387, 0, -6.925569e-06, 0.001272578, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, -0.0001078651, 0.05596312, 0.005698379, 
    -1.93346e-05, -2.432098e-06, 0, -1.506299e-05, 0.001581008, 0.003910638, 
    0.01386389, 0.0008260311, 0.01008068, 0, 0.001716196, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4.237156e-06, 0.003838469, 0.005207187, 0, 
    0.0003805698, 0.003860643, 0.000106466, 0, 0, -1.1255e-05, 0, 0, 0, 0, 0, 
    0, -4.209e-05, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9.245885e-05, 2.016102e-05, -5.963665e-09, 
    0.00314593, 0.0005945713, 0.003662794, 0, 0, 0, 0, 0, 0, -6.838588e-06, 
    0.002455595, -2.857404e-05, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.24165e-06, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.004631095, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001319711, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  -1.071902e-05, 0.0003104234, 0, 0, 0.003985148, 0.0009183214, 0, 0, 0, 0, 
    0, 0, 0, 0, -8.624535e-05, -3.212061e-05, 0, 0, 0, -1.601272e-05, 0, 0, 
    0.0005265421, 0, -2.764706e-05, 0.003516892, 0.001082256, -2.677388e-06, 0,
  -1.710659e-05, 0, 0, 0.0004445918, 0.0107999, -5.344901e-05, 0.003792807, 
    -9.705276e-06, -1.304825e-05, 0, 0.004152217, 0.004010295, 0.001653608, 
    0.04273355, 0.00136338, 0.0001959943, 0, 0.0002503181, 0.005740532, 
    0.005184408, 0.0008234375, 0.001474289, 0, 0, 0.005946141, 0.009186662, 
    0.01018728, 1.926962e-05, 8.569416e-05,
  0, -1.211316e-08, 0.003576165, 0.01751742, -1.813928e-05, 0.03133665, 
    0.001334026, -2.817731e-05, 0, 0.0001301101, 0.008060237, 0.0301805, 
    0.00302785, 0.00802448, -1.319406e-06, 0.03486002, 0.02305472, 
    0.01345193, 0.01198118, -1.054535e-05, -0.0003408901, 0, 0, 5.048402e-07, 
    0.0006663553, 0.01795491, 0.0256762, -1.630522e-05, 0.003923317,
  0, 0.01309418, 0.00933286, 0.0004530372, 0.01647745, 0.01189321, 
    0.0001647077, 0.0004072068, -5.766939e-06, 0, 0.0003850897, 0.01520489, 
    0.02601611, 0.0001519483, 0.01853394, 0.003993249, 0.0008514334, 
    7.265022e-06, -1.933235e-05, -3.149181e-09, 0, 0, 0, 0.001353263, 
    0.05434966, 0.04778849, 0.009864794, 0, 0,
  0, 0.006413547, 0.0156058, 0.001878137, 0.05229056, 0.1103154, 0.05469188, 
    0.03886306, 0.0006145977, -0.0001431286, -2.805345e-05, 0.05307472, 
    0.01539576, 0.004258135, 0.0222337, 0.04379997, 0.02055378, 0.007192855, 
    0, -3.805121e-08, 0, 0, -5.154201e-07, 0.02184298, 0.05318718, 
    0.002025311, -0.000106964, -1.377754e-10, 0,
  0.0008707473, 0.002071158, 0.006228382, -1.753302e-05, 0.003017906, 
    0.01433534, 0.05267559, 0.01891467, 0.01325723, 0.03161201, 0.004898778, 
    0.006271528, 0.02712894, 0.01754393, 0.01233344, -1.66771e-05, 
    0.008690462, -7.365897e-05, 0, -6.466485e-09, 0, 1.605772e-06, 
    0.02272521, 0.0272568, 0.01644002, 0.01552915, 0.03776956, -6.959793e-05, 
    9.328658e-05,
  0, 0, 0, -1.628012e-05, 0.00104567, 6.183302e-05, 0, 0.008701912, 
    -4.431028e-08, 0.03803796, 0.07894669, 0.1007564, 0.01890872, 0.03125632, 
    0.01356323, 0.01772618, 0.02499225, 0.02237327, 0.08270354, 0.0427014, 
    0.154461, -0.0002072583, 0.0003374349, -9.773536e-06, -4.921604e-05, 
    0.003127988, -2.759485e-07, -2.911865e-09, 0,
  0, 0, -1.566449e-07, 0, 0, 0, 0.0003769825, 5.832989e-06, 0, -7.798889e-06, 
    0.08230487, 0.007306145, -0.0002375652, -1.677341e-05, 0.002306567, 
    0.00277603, 0.0146308, 0.0168736, 0.03097507, 0.001746924, 0.01915432, 
    0.001305323, 0.006737057, 0, 0, 1.184739e-06, 0, 0, 0,
  0, 0, 0, 0, -8.708702e-07, 0, 0, 0, 0, 0, 0.001113895, 0.01079374, 
    0.01286473, 0.0002827033, 0.008774512, 0.02056255, 0.001959188, 0, 
    0.0005141585, 0.0002506266, -3.289374e-05, -5.43822e-05, 0.0002865411, 
    -4.221799e-05, -1.002602e-05, 0, 7.455992e-05, 0, 0,
  0, 0, 0, 0, -1.711844e-06, 0, 0, 0, 0, 0, 0, 0.001419681, 0.0007514321, 
    0.0002696218, 0.009019515, 0.007927594, 0.01116594, -7.34804e-07, 0, 
    0.0001761168, 0, 0, 0, 0.001266385, 0.01171861, 0.003481978, 
    -1.068491e-06, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.002192522, 0, 0, 0, 0, 0, 
    0, 0, -7.664561e-06, 0.008063523, 0.003395772, -6.449562e-05, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, -6.191959e-05, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0002081825, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.00533515, 0, 0, 0.001286464, 0, 0, 
    0, 0, 7.105446e-05, 0, 0, 0, 0, 0, 0, 0,
  0.0001398612, 0.005587675, 0.0001036509, 9.808793e-05, 0.01468475, 
    0.009525413, -5.690532e-07, 0, 0, 0, -2.650433e-05, 0, 0, -9.937902e-05, 
    0.004223273, -4.418451e-05, 0.0001596142, 0, 0.0006102083, 0.003206418, 
    3.70709e-05, -9.912927e-06, 0.003032451, 0.0005253585, 0.0003506916, 
    0.005481086, 0.004821521, -9.582433e-05, 0.001703612,
  0.001453956, 9.609547e-09, 1.83578e-08, 0.01157135, 0.01988744, 
    0.002070092, 0.01011437, 0.003817846, -8.853643e-05, 0, 0.005690647, 
    0.01216396, 0.003128693, 0.05732026, 0.002816682, 0.004092608, 0, 
    0.008739803, 0.01612315, 0.01222105, 0.008457737, 0.005418535, 0, 0, 
    0.01319823, 0.0215646, 0.03115743, 0.008400056, 0.001469355,
  7.586092e-07, 0.0001531978, 0.0210789, 0.03628554, 0.002228296, 0.07092244, 
    0.006741264, 0.002239123, 1.990292e-05, 0.004156885, 0.01726194, 
    0.07039057, 0.01063513, 0.01596943, -3.272992e-05, 0.05576539, 
    0.04837219, 0.04155124, 0.0313115, 0.0007471567, 0.00144208, 0, 
    3.88441e-05, 0.0001626651, 0.01390155, 0.03369245, 0.04552605, 
    0.001631113, 0.00722171,
  -1.112065e-06, 0.0524854, 0.05922394, 0.006522651, 0.06752689, 0.1326414, 
    0.01145134, 0.007952131, 0.0001610426, 4.476382e-09, 0.01303747, 
    0.04723231, 0.1203928, 0.0586522, 0.09081013, 0.03901257, 0.005422938, 
    0.008990459, 0.001878839, -1.973598e-06, 0, -1.775838e-06, -3.990554e-06, 
    0.07635562, 0.2866382, 0.06931593, 0.02983839, -6.364968e-05, 
    -8.506891e-10,
  -4.347116e-05, 0.1176216, 0.05818296, 0.01403497, 0.1549126, 0.2080474, 
    0.1005078, 0.1074601, 0.04103789, 0.005147557, 0.01463525, 0.1687052, 
    0.08936292, 0.04785482, 0.0594158, 0.0704408, 0.02599204, 0.01127508, 
    -3.651595e-07, 5.281111e-06, 0, 0, 0.001052512, 0.1592866, 0.289002, 
    0.01332857, -8.113085e-06, -2.632532e-05, -1.073471e-10,
  0.004564492, 0.01207183, 0.02597537, 0.0002040143, 0.02487735, 0.05188342, 
    0.09505875, 0.1516001, 0.08126158, 0.06880455, 0.09050976, 0.1029031, 
    0.1435882, 0.06831305, 0.04134732, 0.003376791, 0.008499911, 0.003430911, 
    -1.127992e-05, 0.001181333, -1.585739e-05, 2.803474e-05, 0.02930727, 
    0.1336362, 0.1304835, 0.03758568, 0.05403275, -4.710578e-05, 8.416439e-05,
  0, -1.700739e-06, -1.300201e-06, -2.819628e-05, 0.001186485, 0.004850541, 
    -1.532354e-05, 0.03637607, 0.0001672712, 0.09444425, 0.2144659, 
    0.1868099, 0.07939381, 0.07675353, 0.05294319, 0.05608237, 0.03279647, 
    0.0316762, 0.1169069, 0.07027894, 0.1791254, -0.0008144027, 0.0008557719, 
    -2.286589e-05, -9.576002e-05, 0.009549589, -0.0002327689, 0.0001113881, 
    7.798612e-14,
  0, 0, 0.000366339, 4.247332e-06, -5.876957e-06, 0, 0.003849557, 
    0.0006317876, 8.82103e-05, 0.002138266, 0.130278, 0.02383723, 0.03383298, 
    0.00476246, 0.003884088, 0.02480915, 0.03925991, 0.03274747, 0.05591096, 
    0.01270825, 0.03942813, 0.01100682, 0.01156167, 1.170332e-05, 
    -4.072976e-10, 0.0001204864, 9.526497e-05, -5.552007e-06, -1.530561e-05,
  0, 0, 0, -7.283662e-06, 0.0006052134, -7.666988e-06, -2.644073e-06, 0, 0, 
    0.008141057, 0.01039456, 0.0303311, 0.02339978, 0.003771063, 0.02088764, 
    0.0351829, 0.00908877, -5.144954e-05, 0.004718713, 0.008206009, 
    0.0001307594, 0.004803488, 0.0048586, 0.0001395754, 0.0007652071, 
    0.0001584277, 0.002081596, -3.94959e-12, 0,
  0, 0, 0, -1.933855e-05, 0.0002226822, 0, 0, 0, 0, 0, -2.554187e-07, 
    0.006881827, 0.00819505, 0.008000206, 0.0174137, 0.03277215, 0.0319296, 
    0.00631179, -1.144464e-05, 0.0004004457, 0, -3.503417e-06, 0.0002486621, 
    0.01849776, 0.03530812, 0.01873638, 0.009622197, -7.291191e-05, 0,
  -2.609787e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -4.442318e-05, 0, 
    0.0002455968, 0.004001081, -2.013022e-05, -1.369795e-05, 0, 0, 0, 0, 
    -9.889526e-06, 0.001871811, 0.0180217, 0.01910972, 0.00165562, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0006057986, 0, 0, 0, 
    0, 0, 0, 0, 0.0002189474, 0.001576098, 0.001477555, -1.166276e-05,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -4.726047e-05, 0.003422793, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, -1.919122e-06, 0, 0, 0, 0.005731489, 
    -2.997124e-05, -6.254108e-05, 0.005819083, -5.42979e-06, -1.95149e-05, 0, 
    0, 0.0005391448, 0, 0.0007973321, -1.05277e-05, 0.001093463, 0, 
    0.0004442194, 0,
  0.001908154, 0.0121145, 0.005351612, 0.002939467, 0.02526363, 0.01789797, 
    0.003341118, -6.653954e-06, 0.0001887862, 9.726064e-05, -0.0002025081, 0, 
    -1.39656e-05, -0.0003019554, 0.01868838, 0.0002399077, 0.006700934, 
    0.0003092765, 0.008441142, 0.007402618, 0.000722524, 0.002284466, 
    0.0150012, 0.005777288, 0.00167821, 0.009741641, 0.01874631, 0.006544385, 
    0.003345912,
  0.02340213, 0.003026205, 0.0001660842, 0.02327967, 0.05059176, 0.009821986, 
    0.01595527, 0.01053824, 0.02484589, 0.003923869, 0.007440844, 0.02179891, 
    0.009118103, 0.07823017, 0.01055395, 0.00822765, 9.072627e-05, 
    0.02389879, 0.02838807, 0.03874205, 0.01912724, 0.01298174, 
    -3.059214e-06, -1.045053e-05, 0.02597345, 0.04405312, 0.07285275, 
    0.01790113, 0.02078089,
  2.51563e-05, 0.001791902, 0.1050702, 0.1065486, 0.07785663, 0.1850078, 
    0.08409295, 0.07113841, 0.01301233, 0.01358641, 0.05046283, 0.1324733, 
    0.04111, 0.05388906, 0.05285615, 0.1501965, 0.1302482, 0.1682122, 
    0.2330956, 0.08098606, 0.01142704, 0.0004994519, 0.01362038, 0.001554963, 
    0.07087907, 0.1079461, 0.1287355, 0.05189316, 0.01526594,
  0.0001653278, 0.1475928, 0.3565799, 0.02993811, 0.06403036, 0.1704267, 
    0.07364188, 0.02312243, 0.01003759, 8.103339e-06, 0.02850391, 0.1244228, 
    0.1653884, 0.0937136, 0.2002797, 0.2097094, 0.09640541, 0.204834, 
    0.111211, 0.01345152, 8.089401e-06, -0.000147713, 0.00226461, 0.1030964, 
    0.2553302, 0.3235347, 0.2128928, 0.02172003, 2.488036e-05,
  0.003811068, 0.1986995, 0.3296514, 0.07588031, 0.1754802, 0.2168125, 
    0.1317279, 0.1275346, 0.03815747, 0.005012012, 0.009929243, 0.1447671, 
    0.06783637, 0.09512407, 0.07678176, 0.07844801, 0.02860117, 0.03721521, 
    -4.909246e-05, 1.641227e-06, 3.193629e-07, 5.138706e-06, 0.004605309, 
    0.2733543, 0.3249125, 0.1763989, 0.009966782, 0.04586242, -1.072544e-05,
  0.02258368, 0.102898, 0.1774148, 0.07101619, 0.1090582, 0.1091392, 
    0.1796924, 0.1880915, 0.1795742, 0.2457787, 0.1163518, 0.09746027, 
    0.1386162, 0.0598234, 0.06398146, 0.0002569488, 0.007489754, 0.01545637, 
    0.0001628307, 0.001555794, 9.969302e-06, 0.0008454663, 0.0349821, 
    0.3983206, 0.2790926, 0.09530878, 0.1450543, 0.01872221, 0.000863074,
  -2.458448e-06, 0.009551242, 0.000283015, -3.1072e-05, 0.005327721, 
    0.02172074, -0.0001635406, 0.04777613, 0.0003416239, 0.09112976, 
    0.199374, 0.1777223, 0.06737635, 0.05210428, 0.07046289, 0.06161212, 
    0.04349359, 0.1250239, 0.2068056, 0.1792944, 0.2447936, 0.07174002, 
    0.01560085, 0.004097199, 0.005351121, 0.02403375, 0.03011373, 0.1067752, 
    -6.513264e-05,
  -5.322508e-06, 1.628021e-07, 0.003439163, 0.004209374, 1.392981e-05, 
    3.388632e-07, 0.006953846, 0.0007911169, 0.008791359, 0.00234301, 
    0.1307227, 0.02458223, 0.02457312, 0.009185486, 0.04885628, 0.0751009, 
    0.1209685, 0.08783705, 0.1302017, 0.1288726, 0.1254354, 0.0488761, 
    0.03708439, 0.01435291, 0.008672191, 0.003241311, 0.007449537, 
    0.05940805, 0.006790535,
  -2.046452e-06, 0, 0, -4.654288e-05, -6.803263e-05, -0.000142756, 
    -0.000304501, -1.249697e-07, 0, 0.01812878, 0.0301616, 0.1057232, 
    0.05580833, 0.004185109, 0.1167281, 0.1227314, 0.03255797, 0.01548509, 
    0.01744752, 0.05266121, 0.01085177, 0.04514053, 0.02429152, 0.04615691, 
    0.01867235, 0.005449638, 0.008723295, 7.433572e-05, -5.568027e-05,
  4.88729e-05, 0, 0, 0.0001853261, 0.002042931, 0.0006470896, 0, 0, 0, 0, 
    -5.62571e-07, 0.02107896, 0.01276774, 0.01973477, 0.03407079, 0.06917807, 
    0.09317485, 0.03911242, 0.01614054, 0.001492579, 0, 0.002031503, 
    0.009797464, 0.04473901, 0.06590834, 0.05611365, 0.02779301, 0.001734698, 0,
  0.002943919, 0.0001725653, 0, 0, 0, -7.277134e-08, 0, 0, 0, 0, 0, 0, 
    -6.121177e-05, 0.005830853, 0.001150323, 0.002496981, 0.01645861, 
    0.002674036, 0.001005197, -2.172558e-06, 0, 0, 0, -6.383645e-05, 
    0.01064776, 0.04239945, 0.04534465, 0.02317015, -0.0002299365,
  0.0007464107, -1.0421e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.001028761, 0.003310637, -2.841786e-05, 0, 0, 0, 0, 0, 0, 0.007569211, 
    0.007705164, 0.003707675, 0.001290087,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, -2.662068e-06, 0, 0, 0, 0, 0, 0, -1.029833e-05, 
    0.005932055, 7.542806e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  -1.901586e-05, 0, 0, 0, -1.81492e-05, 0.001714205, 0.0004007616, 
    0.0006998566, -4.586653e-05, -2.679231e-05, 0, 0.0001456876, 
    -7.803325e-05, 0.008084945, 0.0001159344, 0.0002500857, 0.009305312, 
    0.0006870979, 0.0001534425, -3.072124e-05, 7.754233e-05, 0.002000153, 
    -2.904232e-05, 0.001206105, 0.002813366, 0.009058621, 0.002081837, 
    0.00130426, 0.0004287907,
  0.01142963, 0.02224564, 0.01419463, 0.01466715, 0.03462054, 0.04099932, 
    0.01949493, 0.0029629, 0.00467039, 0.01646046, 0.03031767, 0.004527489, 
    0.001943879, 0.008002862, 0.03144777, 0.02338636, 0.02066894, 
    0.008842385, 0.02622917, 0.01587643, 0.01584283, 0.008795068, 0.02352053, 
    0.01627608, 0.00938161, 0.03494918, 0.04298929, 0.03269239, 0.01059589,
  0.1151065, 0.06405952, 0.02165892, 0.04853499, 0.086937, 0.06642821, 
    0.07822977, 0.05622886, 0.05998809, 0.04105842, 0.04975182, 0.0510329, 
    0.04423829, 0.1124828, 0.06477332, 0.04939068, 0.03348857, 0.0855604, 
    0.08269213, 0.1764342, 0.1510011, 0.09198923, 0.02539507, 0.002892753, 
    0.06748476, 0.1164909, 0.130588, 0.1111142, 0.1200228,
  0.001368467, -8.329317e-07, 0.1077652, 0.1025368, 0.07392313, 0.1671701, 
    0.0901672, 0.1099354, 0.02205928, 0.05808983, 0.1543782, 0.2252256, 
    0.1475084, 0.2001092, 0.1500345, 0.1937458, 0.1257953, 0.2455056, 
    0.405803, 0.1683661, 0.1277909, 0.02343374, 0.01144159, 0.002622318, 
    0.08966592, 0.106183, 0.1523556, 0.0971127, 0.01109696,
  0.0001454678, 0.1068396, 0.2902131, 0.02097565, 0.0572355, 0.1441091, 
    0.06562505, 0.01629365, 0.002369327, 2.603995e-06, 0.02753555, 0.1093661, 
    0.1143283, 0.07618546, 0.1529876, 0.1698065, 0.07150665, 0.1587945, 
    0.0854945, 0.01281121, 1.414076e-05, 0.0004580762, 0.0009618875, 
    0.1055793, 0.2156225, 0.3238079, 0.1411151, 0.004627617, 9.872958e-06,
  0.0001752683, 0.1517271, 0.2844132, 0.04117705, 0.1432582, 0.1787435, 
    0.1187089, 0.1168741, 0.0255026, 0.00351304, 0.003722063, 0.1318364, 
    0.05915999, 0.05830112, 0.05228776, 0.06262667, 0.03067979, 0.02508239, 
    -0.0001008931, 9.696572e-06, 1.774539e-08, 7.875857e-08, 0.002596772, 
    0.2589178, 0.2881474, 0.1387949, 0.003406148, 0.01282977, -1.306894e-05,
  0.009562742, 0.06928481, 0.1051499, 0.03769215, 0.06456578, 0.07957281, 
    0.1382412, 0.1353562, 0.1167937, 0.1938933, 0.08739351, 0.07703893, 
    0.1089969, 0.03798101, 0.03861583, 5.143086e-05, 0.006181237, 
    0.006402013, 1.516113e-05, 5.065903e-05, 2.383632e-06, 0.002441358, 
    0.03774498, 0.2994148, 0.2139578, 0.06581421, 0.08802979, 0.004365318, 
    0.0004126458,
  2.900651e-05, 0.003928058, 0.001043724, 0.004055744, 0.002389623, 
    0.01565106, -0.0001353159, 0.03982681, 0.0001534384, 0.07274936, 
    0.1743942, 0.1555102, 0.05015249, 0.0361312, 0.05285237, 0.04941673, 
    0.03102815, 0.104884, 0.1565063, 0.1514094, 0.2240165, 0.03834879, 
    0.00575388, 0.000499133, 0.003982353, 0.02221212, 0.05021431, 0.048165, 
    0.002233237,
  0.05016483, -2.053399e-05, 0.0006861027, 0.003613806, 3.360325e-05, 
    1.163305e-06, 0.005288825, 0.002130582, 0.01423304, 0.006140465, 
    0.1220205, 0.02293711, 0.006353118, 0.007450047, 0.04757706, 0.07715881, 
    0.08525109, 0.08827456, 0.1331258, 0.1759181, 0.09556849, 0.03580914, 
    0.0222565, 0.008596373, 0.006696675, 0.02036925, 0.06993356, 0.1846278, 
    0.1066195,
  0.01348539, 7.582578e-05, 0.01231424, 0.00250609, 0.003794477, 0.01132955, 
    0.0110601, -0.0001349411, -6.094808e-06, 0.03546334, 0.06538939, 
    0.1312526, 0.06181962, 0.01159008, 0.1630997, 0.1823445, 0.1016762, 
    0.04382547, 0.04067038, 0.1039977, 0.04591009, 0.1200021, 0.1007791, 
    0.1284679, 0.09219787, 0.05677931, 0.05353846, 0.04228936, 0.009478355,
  0.00116072, -2.758645e-05, -1.3326e-08, 0.002887174, 0.0121632, 
    0.003360762, -2.865267e-05, 0, 0, 0, -4.007553e-05, 0.04159372, 
    0.02806095, 0.04121225, 0.07424431, 0.1090353, 0.1588304, 0.1094835, 
    0.06512304, 0.007617167, 0.001226046, 0.01347605, 0.03876429, 0.101734, 
    0.1178419, 0.1299205, 0.09075584, 0.01400443, 4.848094e-06,
  0.0103719, 0.005859364, -3.648319e-05, 0, 0, -2.030416e-05, -1.435071e-06, 
    0, 0, 0, 0, 0, 0.0002493188, 0.01156843, 0.004371879, 0.01017629, 
    0.04600737, 0.02176461, 0.01156269, -0.0001520192, -3.639783e-07, 0, 0, 
    -9.333677e-05, 0.02464715, 0.06526954, 0.09678202, 0.05989046, 0.007635064,
  0.003438483, 0.0010117, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0003511727, 0.007250898, 0.01671128, 0.009136763, -4.040964e-08, 0, 0, 
    0, 0, -8.937569e-06, 0.009074206, 0.02119, 0.01704867, 0.009045721,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -3.81627e-06, 0, 0, 
    0, 0, 0, 0, 0, 0, -2.983107e-05, -3.844158e-05,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, -6.094946e-06, -1.424419e-06, 0, 0, 0, 0, 0, 0.001106188, 
    0.009705536, 0.006499229, 4.912584e-10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  -0.0002868673, -6.815611e-06, 0, 0, 1.123179e-05, 0.01036526, 0.01652833, 
    0.01789152, 0.01105501, 0.0003139969, -3.202385e-05, 0.001043246, 
    0.002252914, 0.0146022, 0.006672292, 0.01147062, 0.03497741, 0.01450571, 
    0.005041346, -8.478646e-05, 0.004749029, 0.007307538, 0.003152293, 
    0.003688381, 0.0147472, 0.01955244, 0.005905141, 0.011424, 0.002377851,
  0.09197451, 0.0949404, 0.0738435, 0.1012766, 0.1001146, 0.08710361, 
    0.1033979, 0.08336588, 0.07497632, 0.09959862, 0.08814792, 0.0549089, 
    0.06914808, 0.05321976, 0.1030931, 0.1125585, 0.105279, 0.1186442, 
    0.1541879, 0.1137161, 0.093607, 0.08333542, 0.1002909, 0.04488153, 
    0.09817537, 0.1294612, 0.154369, 0.1075568, 0.09421709,
  0.1259066, 0.05554068, 0.02640932, 0.06406953, 0.1171582, 0.1228273, 
    0.1433567, 0.1562447, 0.1060238, 0.04343037, 0.0575146, 0.06067006, 
    0.1027362, 0.2358906, 0.1505944, 0.1267882, 0.1039945, 0.09688715, 
    0.1326018, 0.1994226, 0.1762168, 0.1297622, 0.05774855, 0.02587741, 
    0.08491794, 0.1128362, 0.1731865, 0.1515661, 0.1317896,
  0.0006252906, 1.023819e-06, 0.1151838, 0.08934467, 0.0443693, 0.1403935, 
    0.1264313, 0.093881, 0.01310943, 0.03562033, 0.1319878, 0.1978698, 
    0.1269817, 0.1497265, 0.1345593, 0.2032318, 0.1107867, 0.2427622, 
    0.3921664, 0.166361, 0.1071467, 0.009419943, 0.001416743, 0.005948441, 
    0.08596368, 0.08425727, 0.1389683, 0.07238337, 0.009146529,
  3.673298e-05, 0.0952056, 0.2439385, 0.01863482, 0.04799736, 0.1284586, 
    0.07179634, 0.02758957, 0.0001429008, 8.766143e-07, 0.03862071, 
    0.09383783, 0.06435048, 0.07411858, 0.1210424, 0.1337681, 0.04431577, 
    0.1416536, 0.0627032, 0.009022051, -6.787718e-06, -0.0001142446, 
    7.811843e-05, 0.09840237, 0.1780882, 0.2807607, 0.1007861, 7.720815e-05, 
    4.857132e-06,
  0.0001054011, 0.1055805, 0.260382, 0.03441165, 0.1278602, 0.1813077, 
    0.1063575, 0.1064953, 0.01772044, 0.00446788, 0.005740837, 0.1165546, 
    0.06001026, 0.03996907, 0.04638299, 0.0577907, 0.0357849, 0.0203437, 
    0.001000088, 6.797608e-07, -5.034916e-08, 6.835273e-07, 0.003028347, 
    0.238069, 0.2871214, 0.1209182, 0.003251868, 0.00135285, -1.572424e-07,
  0.007196001, 0.0584383, 0.0657573, 0.0187656, 0.04527261, 0.07088921, 
    0.1235906, 0.1057299, 0.07789361, 0.1674749, 0.06009582, 0.05906432, 
    0.1001653, 0.03807387, 0.03139474, 1.625382e-05, 0.005717706, 
    0.0006789223, 4.603563e-06, 4.354047e-05, 1.669369e-06, 0.001282995, 
    0.04049577, 0.22863, 0.1940164, 0.07019823, 0.07657754, 0.002805693, 
    0.002241282,
  2.79913e-06, 0.0008009752, 0.0006162809, 0.002583542, 0.001372259, 
    0.01754667, -3.588069e-05, 0.03607485, 0.00178721, 0.06682096, 0.1487978, 
    0.1388106, 0.04948596, 0.03203336, 0.03123035, 0.0495077, 0.03016452, 
    0.08807414, 0.1374347, 0.1407663, 0.2253725, 0.02581982, 0.005227736, 
    0.001108352, 0.003890505, 0.02639163, 0.06179029, 0.02612925, 
    -0.0002309865,
  0.02629518, -1.207237e-05, 0.0001957765, 0.0004577146, 2.162135e-05, 
    1.743463e-06, 0.01300596, 0.005164115, 0.01059068, 0.01971993, 0.1160618, 
    0.02389687, 0.001351709, 0.01036163, 0.03274616, 0.06153743, 0.07069468, 
    0.09275249, 0.1314924, 0.1138962, 0.07632811, 0.02157116, 0.01683223, 
    0.00545845, 0.001125956, 0.01691623, 0.0790195, 0.1518438, 0.103,
  0.08131375, 0.007806376, 0.01483979, 0.0008690649, 0.003173514, 
    0.008176032, 0.04135125, -0.0001586106, -6.559349e-06, 0.0507533, 
    0.07606438, 0.1299967, 0.07959835, 0.02002706, 0.166922, 0.188992, 
    0.08651868, 0.06198167, 0.04280181, 0.1043569, 0.1136239, 0.1272008, 
    0.1362425, 0.1214052, 0.1050324, 0.07655532, 0.0784066, 0.08116825, 
    0.04130096,
  0.02088437, 0.003701875, 0.009100812, 0.00757209, 0.05650784, 0.02037849, 
    0.0003834743, 0, -1.188994e-06, -3.529768e-10, 0.0001957834, 0.07005568, 
    0.05887791, 0.08923622, 0.09805149, 0.1486831, 0.2652128, 0.1851641, 
    0.1443952, 0.03843367, 0.006363504, 0.03349944, 0.06317665, 0.1666456, 
    0.1901713, 0.2547203, 0.1827113, 0.09750997, 0.05147888,
  0.05495629, 0.0234534, 0.001007126, 9.834195e-05, -7.737725e-08, 
    -3.469914e-05, 0.001176541, 0, 0, 0, 0, 0, 0.0006002226, 0.01608155, 
    0.008980452, 0.02631729, 0.09674097, 0.04289445, 0.03898941, 0.002030944, 
    0.00532734, 0.002080717, 0, 0.001708979, 0.04581957, 0.1192325, 
    0.1863948, 0.1918696, 0.09956414,
  0.01857012, 0.009735387, 0.0004095069, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -0.0001491006, 0.0009364106, 0.01967697, 0.05024751, 0.01789252, 
    0.0004181534, -1.85072e-05, 0, 0, 0, 0.007858081, 0.02121186, 0.0513931, 
    0.07346015, 0.05296008,
  0.003099, 0.0001201568, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -7.885298e-06, 0.002465308, 0.00430367, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.001880184, 0.002013508,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -4.59428e-06, 0, 0, 0, 0,
  0, 0, 0, -3.249954e-05, 0, -1.698221e-09, 0.005460706, -4.197158e-05, 0, 0, 
    0, 0, 0, 0.01584138, 0.01067818, 0.01889271, 0.01989738, 0.01219042, 
    -6.432715e-05, -4.300774e-06, -7.779593e-05, 0, 0, 0.0001862743, 
    0.0197203, 0.01472025, 0.002025225, 0, 0,
  0.02547653, 0.009295185, 0.007296623, 0.008929819, 0.008721753, 0.03245248, 
    0.06396259, 0.04561326, 0.08209498, 0.03919426, 0.04196751, 0.03208495, 
    0.02409627, 0.05109736, 0.03524782, 0.04716493, 0.0961014, 0.0741436, 
    0.06015656, 0.03701052, 0.03438605, 0.0360883, 0.04154474, 0.05381426, 
    0.06005673, 0.07220604, 0.02745783, 0.03473355, 0.01643123,
  0.1436075, 0.1097564, 0.1522356, 0.1915677, 0.1720982, 0.1552516, 
    0.1803119, 0.1432742, 0.1841343, 0.1938248, 0.1698557, 0.114909, 
    0.1801781, 0.1127346, 0.2189157, 0.1888368, 0.2214061, 0.1301532, 
    0.1695585, 0.1850175, 0.1618101, 0.1616193, 0.1649506, 0.07100093, 
    0.1122998, 0.1607043, 0.1899913, 0.1295418, 0.145732,
  0.1169527, 0.04252744, 0.02337765, 0.0653582, 0.1100286, 0.113404, 
    0.1401264, 0.1352086, 0.07971467, 0.04902141, 0.04682493, 0.0474906, 
    0.07510126, 0.2030383, 0.1618469, 0.1119337, 0.09590234, 0.08482348, 
    0.1223275, 0.196129, 0.1699732, 0.1411695, 0.04484573, 0.04711319, 
    0.07571872, 0.08922988, 0.171312, 0.1346016, 0.1283351,
  0.003146082, -1.4278e-05, 0.1187914, 0.08297238, 0.03728338, 0.1142097, 
    0.1320367, 0.07863089, 0.007974376, 0.01461981, 0.1209955, 0.1782342, 
    0.09958599, 0.1183315, 0.1106198, 0.1961378, 0.1164986, 0.218794, 
    0.3933768, 0.1659198, 0.09043495, 0.003244778, 0.0001449251, 0.008109195, 
    0.07437263, 0.07455491, 0.1321137, 0.05017627, 0.008264027,
  6.748502e-06, 0.09401757, 0.2180347, 0.01822713, 0.04436829, 0.1068452, 
    0.0673626, 0.03267172, 0.0004267668, 4.00424e-07, 0.0279641, 0.06139623, 
    0.0487555, 0.06498472, 0.1128266, 0.1126607, 0.02961371, 0.1073889, 
    0.02675748, 0.00385319, -5.423974e-05, -0.0001014334, 6.609083e-05, 
    0.1009778, 0.1310777, 0.2423987, 0.08885267, 1.676748e-05, 3.350521e-06,
  0.0006669417, 0.06222742, 0.2052378, 0.02423336, 0.1227285, 0.1727593, 
    0.09159996, 0.0950454, 0.01245558, 0.007453822, 0.007838983, 0.09560084, 
    0.05199482, 0.02857981, 0.04241732, 0.05172309, 0.04227513, 0.01365349, 
    0.001265911, -4.156497e-09, 6.577376e-09, 1.071296e-06, 0.001119231, 
    0.1793997, 0.2677626, 0.09423921, 0.0005539457, -1.069041e-05, 
    9.924125e-09,
  0.005242407, 0.05493346, 0.05936663, 0.0133354, 0.02270146, 0.06268305, 
    0.1048213, 0.06897274, 0.03926662, 0.1142979, 0.03631118, 0.04879523, 
    0.07669337, 0.03555617, 0.02792621, 2.285037e-05, 0.005239934, 
    -7.25754e-05, 6.626e-06, 0.0003575497, 1.780855e-07, -5.00631e-05, 
    0.05173839, 0.1564048, 0.1684151, 0.09107715, 0.06921194, 0.001766903, 
    0.01440804,
  1.836132e-07, 4.612059e-05, -3.251482e-05, 0.002266471, 0.0005669365, 
    0.01152475, 4.852263e-05, 0.03576064, 0.0112759, 0.06765916, 0.1255586, 
    0.1390068, 0.04503051, 0.03430652, 0.02049503, 0.06322211, 0.03568304, 
    0.08088433, 0.1237315, 0.1282714, 0.2283453, 0.01882058, 0.004937041, 
    0.0009342074, 0.004089135, 0.03463717, 0.09267496, 0.04017891, 
    9.371958e-05,
  0.02076794, -1.959606e-06, 4.305793e-06, 7.90183e-06, 1.606179e-05, 
    -1.183448e-05, 0.01862613, 0.007714559, 0.02885833, 0.01899658, 
    0.1082341, 0.02537544, 0.0003718048, 0.008375586, 0.01625453, 0.07592642, 
    0.05824165, 0.09287877, 0.1171325, 0.07519047, 0.0445391, 0.0106632, 
    0.01616614, 0.0002601332, 0.0009338508, 0.01940065, 0.06773586, 
    0.1129021, 0.1038615,
  0.07997609, 0.01780204, 0.02061075, 0.01011372, 0.009238216, 0.01033376, 
    0.05133347, -0.0003375515, -0.0001157761, 0.04939545, 0.06804404, 
    0.1047452, 0.07930718, 0.04471196, 0.1552374, 0.1521502, 0.1115799, 
    0.04332501, 0.06732146, 0.08699322, 0.1169829, 0.1224645, 0.09307916, 
    0.1013456, 0.0882872, 0.0561333, 0.06754684, 0.07638459, 0.06785072,
  0.07031554, 0.03167731, 0.0479941, 0.02437558, 0.0837328, 0.06049588, 
    0.005295715, 0.00661522, 0.0007662604, -1.055479e-05, 0.02719492, 
    0.1325198, 0.06607838, 0.1256841, 0.1120459, 0.1653466, 0.2920876, 
    0.1805287, 0.1612169, 0.1071289, 0.02284375, 0.03912793, 0.08186851, 
    0.1781197, 0.1637784, 0.2588654, 0.1711351, 0.1129583, 0.09767032,
  0.1446468, 0.06985079, 0.0222628, 0.017296, 0.02760136, -5.510615e-05, 
    0.003162392, 0, 0, 0, 0, -2.139563e-06, 0.003437675, 0.03230201, 
    0.03900636, 0.07288827, 0.1514807, 0.09169731, 0.1309368, 0.007979001, 
    0.02455472, 0.04197433, 0.02933692, 0.01827011, 0.04924958, 0.1328506, 
    0.2411726, 0.2721581, 0.1560425,
  0.1297489, 0.04216384, 0.004354456, -9.512171e-07, 0, 2.178444e-06, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.007604989, 0.01450092, 0.04922482, 0.1024477, 
    0.0224661, 0.002859073, 0.0003824009, -4.196522e-05, -3.364724e-05, 
    -7.009313e-06, 0.01033714, 0.03732684, 0.1075748, 0.1446002, 0.1549947,
  0.01275104, 0.001869212, -2.924651e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0001786749, -4.770072e-05, 0.0004138214, 0.007715863, 0.00735914, 
    0.005164474, 0, 0, 0, 0, 0, 0, -0.0001279253, 0.01610473, 0.01087213,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -3.324147e-05, 0, 0, 0, 0, 
    0, 0, 0.02987806, 0.02122088, 0.01471384, -0.002218735, 0, 0,
  0.02914923, 0.0289526, -0.0004596857, 0.006037111, -0.0001162519, 
    0.001931111, 0.08285295, -0.001359823, 0, -9.983028e-10, 0, 0, 
    -0.000836689, 0.04535022, 0.04964364, 0.05747541, 0.04164422, 0.04348707, 
    0.03591025, 0.001800814, 0.001655006, 0, 1.303506e-05, 0.02920064, 
    0.02677373, 0.01543493, 0.05154642, 0.04101207, 0.02151701,
  0.06383995, 0.05914366, 0.09015208, 0.05365247, 0.042876, 0.0432443, 
    0.08358654, 0.08621489, 0.1194893, 0.07749721, 0.09727593, 0.0683291, 
    0.0913616, 0.1511728, 0.06941511, 0.07229643, 0.1422217, 0.1553848, 
    0.151371, 0.1236169, 0.1339841, 0.1326344, 0.1275686, 0.09243017, 
    0.1408453, 0.1574225, 0.1106883, 0.07889606, 0.05659917,
  0.1738014, 0.1226666, 0.1619689, 0.1966944, 0.2057608, 0.1648118, 
    0.1876189, 0.1701811, 0.1705833, 0.1691969, 0.1595137, 0.1199724, 
    0.1885651, 0.1236909, 0.2096989, 0.1775567, 0.2044358, 0.1258035, 
    0.1784008, 0.1845164, 0.167724, 0.1679127, 0.1891059, 0.1028779, 
    0.1121979, 0.1759988, 0.2168848, 0.1590063, 0.168404,
  0.1028434, 0.0381673, 0.02294128, 0.06430004, 0.102112, 0.09406603, 
    0.1323373, 0.1214969, 0.0722556, 0.04937608, 0.03004934, 0.03585874, 
    0.06474898, 0.1531622, 0.1382915, 0.09852906, 0.09035922, 0.08112808, 
    0.1148914, 0.1699905, 0.1555004, 0.1336214, 0.0380301, 0.05179028, 
    0.05881532, 0.07068626, 0.1688284, 0.1247223, 0.1261607,
  0.002476709, -9.838611e-05, 0.1226575, 0.07077935, 0.02813956, 0.09943622, 
    0.1261314, 0.06825212, 0.001792501, 0.004172266, 0.0969709, 0.1626531, 
    0.07653178, 0.09742824, 0.08659813, 0.1660288, 0.115708, 0.2273493, 
    0.4062284, 0.1329906, 0.08508382, 4.924604e-05, 0.0007580851, 
    0.005798343, 0.05844956, 0.06864267, 0.1143258, 0.03111179, 0.008161681,
  2.748238e-06, 0.09562935, 0.1812766, 0.01813539, 0.03756078, 0.07465975, 
    0.05641496, 0.03179882, 0.00644088, 1.5579e-08, 0.01980085, 0.04314023, 
    0.03817594, 0.03409256, 0.1086876, 0.07783682, 0.02468678, 0.08720479, 
    0.01453601, 0.0007708819, -1.726752e-05, -3.973112e-05, 7.100341e-06, 
    0.09186457, 0.09366945, 0.2035402, 0.0672664, 1.652675e-06, 1.874547e-06,
  1.853098e-05, 0.03040227, 0.1700549, 0.01919468, 0.1115738, 0.1651287, 
    0.07537988, 0.08045208, 0.0100559, 0.007297249, 0.005790362, 0.07272502, 
    0.03926067, 0.01866275, 0.03213217, 0.04817267, 0.04761085, 0.008313044, 
    4.706179e-05, -6.436571e-11, 6.337488e-09, 6.274171e-07, 0.0001664776, 
    0.1145051, 0.2384046, 0.06355304, 0.001317678, -9.837145e-05, 5.825767e-08,
  0.01132309, 0.03835338, 0.06684536, 0.008753813, 0.0101778, 0.05555176, 
    0.08209526, 0.04159965, 0.02566625, 0.07787874, 0.02366212, 0.03363438, 
    0.05049167, 0.02864179, 0.01892502, 0.0001840581, 0.007570922, 
    -5.996425e-06, 1.738961e-05, 0.001013616, -9.775025e-08, 0.0001187975, 
    0.04327338, 0.1188326, 0.1563767, 0.09615891, 0.0695468, 0.006734618, 
    0.03498788,
  5.637845e-08, 2.726393e-05, 0.0001711381, 0.004708452, 0.0003793449, 
    0.006091232, 0.000121322, 0.03726683, 0.01364571, 0.06418577, 0.1004094, 
    0.1331566, 0.03862136, 0.03159408, 0.02699094, 0.07349268, 0.04986175, 
    0.06709594, 0.1179395, 0.1294783, 0.2166685, 0.01398471, 0.004665732, 
    0.001164149, 0.007235008, 0.04287063, 0.08007336, 0.04490414, 
    -9.451629e-07,
  0.02157606, 1.843411e-06, 2.459596e-07, 1.236292e-06, 1.502578e-05, 
    -4.493056e-05, 0.01866398, 0.005615357, 0.03204066, 0.02144994, 
    0.1119512, 0.0252007, 6.790984e-05, 0.005995024, 0.006765902, 0.0724423, 
    0.0477579, 0.08421136, 0.1194536, 0.06514362, 0.03306, 0.004622968, 
    0.01471325, 0.001141088, 0.001574146, 0.0192409, 0.05668, 0.08769834, 
    0.0662348,
  0.07090508, 0.01539071, 0.02435942, 0.005240472, 0.00543645, 0.01202493, 
    0.04677914, 0.001818508, -0.0001954341, 0.03528943, 0.06205501, 
    0.08688377, 0.07938059, 0.05214057, 0.126411, 0.1205795, 0.09886593, 
    0.04893643, 0.07004393, 0.05783924, 0.09214924, 0.09882147, 0.06712295, 
    0.07811379, 0.0533895, 0.03852157, 0.05867689, 0.06157695, 0.07050473,
  0.06706586, 0.04480844, 0.09265155, 0.06764343, 0.2133361, 0.176263, 
    0.0143985, 0.06875466, 0.01375536, 0.001653379, 0.07784974, 0.1399265, 
    0.09358831, 0.1518526, 0.1242169, 0.1822281, 0.2816945, 0.1621739, 
    0.1554205, 0.1472249, 0.05952503, 0.06555784, 0.1148023, 0.1716461, 
    0.1636464, 0.2608436, 0.1312968, 0.1008647, 0.08976018,
  0.1891545, 0.1239623, 0.1133058, 0.1156827, 0.1036248, 0.05259333, 
    0.00413439, -3.344545e-06, 0, 0, 0.0004769088, 0.001006023, 0.02145334, 
    0.04374215, 0.1230259, 0.1302507, 0.1885178, 0.1177734, 0.1550081, 
    0.05634949, 0.05571372, 0.07450598, 0.08417587, 0.04072691, 0.0852157, 
    0.1519042, 0.2624709, 0.2909842, 0.1348114,
  0.1847512, 0.1325329, 0.06077209, 0.00559985, 0.03564175, 0.05876775, 
    0.04038369, 2.257606e-05, 1.344479e-05, 0, 0, 0, 0, -1.736775e-05, 
    0.03333199, 0.04922961, 0.1236912, 0.1265642, 0.0411433, 0.02853344, 
    0.03983017, 0.05368035, 0.03368028, 0.0001861445, 0.01428537, 0.05053763, 
    0.1371043, 0.1916681, 0.2268243,
  0.05682876, 0.02825416, 0.000438487, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.007087566, 0.009682808, 0.03359229, 0.05491679, 0.03167392, 
    0.009773458, -6.09793e-05, 0, 0, 0, -2.005184e-06, -1.888924e-06, 
    -0.0003216186, 0.06233579, 0.06089,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2.886677e-06, -9.113041e-06, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -3.444591e-05, -1.895172e-05, 
    -5.541787e-05, -1.114945e-05, 0, 0, 0, 0, 0.006405809, 0.03960893, 
    0.0436826, 0.01606392, 0.02755736, -0.001965381, 0,
  0.05746908, 0.09945945, 0.08593798, 0.09078772, -0.00144454, 0.001516707, 
    0.170823, 0.01049207, 0.0009148781, -0.001863641, -7.344904e-05, 0, 
    -0.0008791218, 0.07220011, 0.09473284, 0.09131405, 0.06095061, 0.1297469, 
    0.06649379, 0.0982566, 0.05475348, 0.04961023, 0.05461142, 0.1219549, 
    0.1411359, 0.0923823, 0.161509, 0.1186001, 0.05466755,
  0.1320883, 0.1546843, 0.1471955, 0.1419287, 0.08965293, 0.09454751, 
    0.1389918, 0.1255683, 0.149, 0.116303, 0.1295423, 0.09760074, 0.1608948, 
    0.1884177, 0.1226552, 0.1273527, 0.1635705, 0.1771057, 0.1789254, 
    0.1474532, 0.1954385, 0.1930426, 0.2003016, 0.1754312, 0.256425, 
    0.2457711, 0.1711685, 0.129755, 0.1241766,
  0.1723072, 0.1207111, 0.1682972, 0.2118965, 0.2133102, 0.1496849, 
    0.1717679, 0.1676961, 0.1605252, 0.1430592, 0.1419267, 0.1069926, 
    0.1846197, 0.1177158, 0.2027517, 0.1660421, 0.1769299, 0.1300837, 
    0.1781811, 0.1593266, 0.163239, 0.1672552, 0.1877775, 0.1327596, 
    0.1048401, 0.1607523, 0.1953475, 0.1645066, 0.1677877,
  0.08461191, 0.0315323, 0.02352075, 0.07390233, 0.0827483, 0.06802282, 
    0.1125761, 0.1120182, 0.06261058, 0.05247179, 0.02869818, 0.03045035, 
    0.06491274, 0.13425, 0.1268172, 0.07195184, 0.08368297, 0.08344308, 
    0.08607313, 0.1517853, 0.1559862, 0.1427033, 0.02527736, 0.03605253, 
    0.04979838, 0.06045144, 0.1615615, 0.1126195, 0.1089602,
  -7.57311e-05, -3.208662e-05, 0.1044792, 0.06018608, 0.02186996, 0.09064373, 
    0.1244767, 0.05175849, 0.0004045916, 0.0008286599, 0.08141667, 0.140782, 
    0.05961345, 0.08428748, 0.06447595, 0.1358245, 0.1072954, 0.2329732, 
    0.4079922, 0.09447842, 0.07878871, 0.001895475, 0.0005496424, 
    0.007043959, 0.05596242, 0.06280062, 0.1198312, 0.03190459, 0.005356198,
  1.826166e-06, 0.08895063, 0.1511952, 0.01623934, 0.0340419, 0.0454097, 
    0.04997062, 0.02582741, 0.0001966642, 4.287869e-10, 0.01360651, 
    0.02923835, 0.03020702, 0.0218411, 0.1089719, 0.05609203, 0.03667356, 
    0.05861178, 0.008382281, 1.260103e-05, 0.0007486808, -1.060908e-05, 
    2.240858e-06, 0.07979342, 0.08395144, 0.1940235, 0.06864554, 
    6.109841e-06, 7.274582e-07,
  1.048868e-05, 0.02168752, 0.1260127, 0.0137156, 0.1265804, 0.1711846, 
    0.06941599, 0.07508662, 0.007850649, 0.006070138, 0.004423358, 
    0.05944563, 0.02427298, 0.01538593, 0.0349553, 0.04040193, 0.06309145, 
    0.006307207, 6.295685e-05, 0, 0, -4.273471e-06, 0.0003654642, 0.073475, 
    0.2170812, 0.03978995, 0.0004035945, -1.761498e-05, -1.12352e-07,
  0.02862468, 0.02052988, 0.05953119, 0.007249748, 0.009827883, 0.05466889, 
    0.0598221, 0.03492087, 0.03242123, 0.06206966, 0.02312733, 0.02782205, 
    0.03585367, 0.01989107, 0.02083509, 0.01051789, 0.009691617, 
    -1.595376e-06, 5.356238e-06, -2.728479e-06, -5.458743e-05, 0.005555946, 
    0.04367362, 0.0955262, 0.1507635, 0.09160241, 0.06457629, 0.05127234, 
    0.06011511,
  9.96372e-09, 1.287421e-05, 5.526486e-05, 0.01119107, 0.002129162, 
    0.00600928, 0.0003305641, 0.04390704, 0.01079673, 0.05156614, 0.09937651, 
    0.1202757, 0.0299959, 0.028477, 0.03073618, 0.09108508, 0.05744313, 
    0.06155042, 0.1236558, 0.1476621, 0.2083166, 0.01654087, 0.00420784, 
    0.0008665925, 0.01578798, 0.04882422, 0.0637857, 0.04127117, -2.063132e-07,
  0.002535698, 2.902852e-06, 1.810992e-08, 2.532637e-06, 6.317229e-06, 
    4.843649e-06, 0.02031583, 0.002595312, 0.01913434, 0.02501524, 0.112888, 
    0.02584006, 0.0002766328, 0.003853971, 0.002199508, 0.0681345, 
    0.01951897, 0.06858283, 0.1110997, 0.05568841, 0.02683167, 0.003375458, 
    0.01052356, 0.00075567, 0.002163067, 0.01373948, 0.03411807, 0.06061464, 
    0.0661187,
  0.05303678, 0.007080167, 0.01813481, 0.009582603, 0.005043467, 0.01354811, 
    0.04583296, 0.01393445, 0.000274627, 0.02672151, 0.05618642, 0.0706341, 
    0.07178563, 0.05505819, 0.08904252, 0.1167204, 0.09716021, 0.03942879, 
    0.07212865, 0.02856147, 0.08400819, 0.09054829, 0.04232766, 0.07187755, 
    0.03885417, 0.0194262, 0.04875476, 0.03095764, 0.06657425,
  0.05555815, 0.0402599, 0.1177679, 0.1327237, 0.2039837, 0.2283434, 
    0.02680373, 0.1232121, 0.07175546, 0.05279854, 0.1022957, 0.1534072, 
    0.1169988, 0.1625565, 0.1338367, 0.1952042, 0.2863796, 0.165032, 
    0.1356906, 0.1630125, 0.06840007, 0.07721927, 0.1152808, 0.1749276, 
    0.1675359, 0.2458377, 0.1124222, 0.09188335, 0.07217789,
  0.18449, 0.1473435, 0.1841913, 0.2568575, 0.1973315, 0.208932, 0.1403881, 
    8.204517e-05, -7.881235e-06, 0.01181728, 0.02120881, 0.009345485, 
    0.06312621, 0.06917353, 0.157043, 0.1628651, 0.2123061, 0.1280934, 
    0.1784532, 0.09325751, 0.08657581, 0.1358969, 0.109772, 0.08359953, 
    0.1432395, 0.2022921, 0.3177753, 0.2817702, 0.1711791,
  0.2472597, 0.1793921, 0.1156424, 0.08053637, 0.1418056, 0.1468212, 
    0.1766936, 0.1528253, 0.0827233, -7.351177e-05, -0.0001394001, 
    -0.0005016651, -0.001207929, 0.003619317, 0.05247934, 0.09813959, 
    0.1395714, 0.1633602, 0.0744573, 0.1098006, 0.154859, 0.1487016, 
    0.07626409, 0.03565054, 0.08723506, 0.09452799, 0.1762702, 0.220575, 
    0.2673147,
  0.07727361, 0.08290108, 0.01302744, 0.005693504, 0.002693068, 0.009015999, 
    0.01503733, -0.0006563548, 0, 0, 0, 0, 0, 0.0009763621, 0.02886432, 
    0.05739374, 0.07277764, 0.08672666, 0.08592068, 0.0614034, 0.01393798, 
    0.006647315, -0.000614159, -0.0009240629, 0.02296757, -6.184303e-05, 
    0.0005689827, 0.09407167, 0.08234781,
  0.02650599, 0.02351273, 0.0037386, -4.957299e-05, 0.004864952, 
    5.544139e-05, 2.117179e-05, 8.740443e-08, 0, 0, 0, 0, -0.0002223016, 
    0.003586723, 0.003955459, 0.003311937, 0.002561591, 0.0003605577, 
    -4.703573e-06, 0, 0, 0, 0, 0, 0, 0, 0, -0.001795128, 0.02258285,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.02577268, 0.09325131, 0.118473, 
    0.1230386, 0.04751639, 0.0003250196, 0, 0, 0, 0.01158996, 0.1477346, 
    0.06821498, 0.0520126, 0.02699513, 0.01255076, 0,
  0.1557086, 0.2474232, 0.1759682, 0.2056953, 0.0001790265, 0.04171313, 
    0.2290922, 0.06324472, -0.00213215, 0.003382862, -0.001166795, 
    -3.689957e-05, 0.001940988, 0.1691511, 0.1415224, 0.1590924, 0.1316346, 
    0.2161572, 0.1578448, 0.2742127, 0.07771336, 0.1156563, 0.1238751, 
    0.2303592, 0.2948733, 0.1919358, 0.2368473, 0.1444126, 0.1134098,
  0.1499088, 0.2840862, 0.2375391, 0.2188682, 0.1367211, 0.1576162, 
    0.1468055, 0.1529262, 0.1701995, 0.1252934, 0.2013345, 0.1908893, 
    0.2195141, 0.2401, 0.171451, 0.1595494, 0.1628246, 0.173039, 0.1872729, 
    0.1717933, 0.2725793, 0.2801972, 0.2896214, 0.2251594, 0.2694817, 
    0.2545009, 0.2148093, 0.1475413, 0.1811412,
  0.1731134, 0.125373, 0.1652698, 0.1971455, 0.185053, 0.1421156, 0.1774441, 
    0.1612898, 0.142828, 0.1370338, 0.1303535, 0.1385924, 0.1725343, 
    0.117381, 0.1907477, 0.152668, 0.1404191, 0.130536, 0.1559536, 0.149604, 
    0.1508434, 0.1585173, 0.1915661, 0.1455952, 0.09490886, 0.1608996, 
    0.1866992, 0.1776352, 0.178514,
  0.0684494, 0.03588338, 0.02647215, 0.08038523, 0.07085802, 0.05669452, 
    0.1060369, 0.1239137, 0.05365697, 0.02131144, 0.02435466, 0.02605382, 
    0.06140568, 0.1258129, 0.1099405, 0.0553579, 0.06678723, 0.07764818, 
    0.06890335, 0.1354211, 0.1346276, 0.1107314, 0.01883932, 0.02283498, 
    0.04544429, 0.05805774, 0.1468594, 0.1197463, 0.09516934,
  0.003499871, -7.227922e-06, 0.07664793, 0.04712221, 0.01852926, 0.09118441, 
    0.1223964, 0.02681156, 2.252013e-07, -0.0003389043, 0.07390315, 
    0.1420478, 0.05115822, 0.07566698, 0.05023678, 0.1158803, 0.1282043, 
    0.2067119, 0.4026459, 0.06046115, 0.08998255, 0.004458591, 0.001664797, 
    0.004612563, 0.05392144, 0.06057179, 0.1244756, 0.04573486, 0.005136657,
  1.217375e-06, 0.07973421, 0.1254085, 0.01152288, 0.03716712, 0.02905564, 
    0.06129212, 0.02195668, -3.190694e-05, 3.110787e-09, 0.0178661, 0.018321, 
    0.02696966, 0.0080269, 0.1073175, 0.03739185, 0.05851325, 0.04542569, 
    0.006441401, 1.344177e-07, 0.0001017154, 7.773414e-08, 6.552397e-06, 
    0.06085303, 0.07088497, 0.1953065, 0.06580891, 3.970219e-06, 6.789124e-07,
  5.457104e-05, 0.02514783, 0.1083506, 0.01376276, 0.1254598, 0.1712148, 
    0.06848362, 0.07615485, 0.009107815, 0.003910275, 0.004417914, 
    0.04749959, 0.01794919, 0.01398567, 0.02559309, 0.03467786, 0.06188932, 
    0.005769869, 4.53768e-05, 0, -8.333317e-11, 1.64972e-07, 0.002470567, 
    0.05337059, 0.2078958, 0.03099036, 0.0003656248, -3.803095e-05, 
    -2.813182e-07,
  0.04200431, 0.009985456, 0.0684211, 0.005574379, 0.02093158, 0.07011482, 
    0.04644365, 0.03191608, 0.01372023, 0.05743343, 0.02162764, 0.02575441, 
    0.02756441, 0.01693771, 0.0170772, 0.003626934, 0.008871597, 
    -8.340922e-07, 1.344175e-06, 2.133256e-07, 0.0003545408, 0.00181055, 
    0.04823187, 0.08012522, 0.1285189, 0.08641359, 0.07543245, 0.06575961, 
    0.07032013,
  -2.996543e-10, 5.67737e-06, -3.659979e-06, 0.01420725, 0.000506143, 
    0.007144209, 6.98037e-05, 0.03084981, 0.005905357, 0.05729418, 0.1056916, 
    0.106828, 0.02770167, 0.02785673, 0.03532613, 0.1160444, 0.06565283, 
    0.06387623, 0.1116339, 0.155306, 0.1976474, 0.02380736, 0.005898983, 
    0.001402711, 0.01565498, 0.03971893, 0.04839341, 0.02582685, -2.593122e-07,
  5.745454e-05, 2.4923e-06, 3.654883e-08, 1.480744e-07, 3.476149e-06, 
    9.053628e-05, 0.0212247, 0.00395608, 0.002223794, 0.0186251, 0.1020928, 
    0.01782555, 0.0004015069, 0.003066231, 0.0008371561, 0.06151024, 
    0.0110661, 0.04911186, 0.1013459, 0.04334953, 0.0275893, 0.0006846263, 
    0.005862365, 0.0004875456, 0.003584462, 0.005221919, 0.02984575, 
    0.02895625, 0.01127447,
  0.03718416, 0.01885438, 0.01899884, 0.01398483, 0.005769007, 0.01450651, 
    0.0600422, 0.01539895, 0.01505738, 0.02892069, 0.05065612, 0.05861731, 
    0.07429781, 0.07173859, 0.0600023, 0.112749, 0.08378405, 0.02948229, 
    0.0481618, 0.0138013, 0.08686338, 0.07110585, 0.03859072, 0.0396304, 
    0.02432577, 0.01268802, 0.04562252, 0.009240398, 0.06437891,
  0.03962832, 0.04349159, 0.1174425, 0.2122779, 0.17373, 0.2138577, 
    0.05259034, 0.1376089, 0.08628848, 0.09587634, 0.1138037, 0.1451292, 
    0.1354537, 0.1694675, 0.1385149, 0.1866421, 0.2744105, 0.1532348, 
    0.1366741, 0.1904704, 0.08185024, 0.07729855, 0.1158747, 0.1801655, 
    0.1595232, 0.220213, 0.09067743, 0.0809406, 0.06876653,
  0.1735437, 0.172922, 0.2440068, 0.318106, 0.2230582, 0.251512, 0.2321475, 
    0.004392991, 0.008734399, 0.03523748, 0.08408079, 0.02181475, 0.1537922, 
    0.1162696, 0.1895282, 0.2010108, 0.2073453, 0.1475563, 0.1840853, 
    0.1029225, 0.1120801, 0.1713132, 0.1532729, 0.1321266, 0.158105, 
    0.2273887, 0.3180811, 0.2544703, 0.1708594,
  0.2974091, 0.232939, 0.1604805, 0.2106326, 0.2005825, 0.1931486, 0.2092122, 
    0.1677838, 0.1785895, 0.1239211, 0.04239294, 0.02029959, 0.01402529, 
    0.04504666, 0.1301317, 0.1334669, 0.2246487, 0.2614295, 0.1299784, 
    0.1547378, 0.2742852, 0.2052026, 0.1339197, 0.1296232, 0.1611516, 
    0.1479605, 0.1929969, 0.276491, 0.3291432,
  0.09661917, 0.1094169, 0.05812174, 0.03525393, 0.05376043, 0.08240119, 
    0.09039867, 0.06000927, 0.01351578, 0.008665603, -6.348713e-05, 
    -0.0002661927, 0.01100382, 0.02250903, 0.1005233, 0.1109354, 0.1327384, 
    0.1410159, 0.1410137, 0.1014201, 0.07080302, 0.0254599, 0.06928553, 
    0.01363148, 0.1052155, 0.0003359075, 0.009270365, 0.1326511, 0.09368513,
  0.06831595, 0.06973208, 0.04987735, 0.0503353, 0.05679012, 0.03000967, 
    0.02267583, 0.005764253, 0.02225209, 0.01883432, 0.006592336, 
    0.006138317, 0.02163496, 0.02289463, 0.01796875, 0.01274699, 0.01209967, 
    0.02130284, 0.01594267, 0.02011872, 0.02059524, 0.01287436, 
    -1.386036e-08, -3.248611e-06, -1.265345e-06, -2.834472e-05, 
    -0.0009322432, 0.005674319, 0.07467768,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  -0.00100424, -1.481948e-08, -6.728155e-07, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6.720695e-07, 0.08724638, 0.09637573, 0.113269, 0.1736306, 0.2941803, 
    0.01652826, 7.302506e-05, -0.00109961, -0.001055301, 0.07566765, 
    0.1251252, 0.06263699, 0.03662993, 0.03721879, 0.0319824, 0.01346025,
  0.1723279, 0.2658516, 0.1822386, 0.2287185, 0.03704973, 0.1168195, 
    0.2768977, 0.1045677, 0.04481994, 0.05982935, 0.01395318, -0.001215307, 
    0.05419282, 0.186499, 0.1558733, 0.1853155, 0.1329785, 0.2289615, 
    0.166159, 0.2673035, 0.08628083, 0.1210782, 0.1787805, 0.3325699, 
    0.347566, 0.1803631, 0.2401782, 0.1349853, 0.1648151,
  0.1489878, 0.2949023, 0.260375, 0.2360091, 0.1612678, 0.161756, 0.1546218, 
    0.1343809, 0.1885312, 0.1261663, 0.2175308, 0.2310983, 0.2354784, 
    0.2549507, 0.1755064, 0.1833564, 0.1610671, 0.1599433, 0.1842114, 
    0.186832, 0.3198597, 0.2850486, 0.2792165, 0.238832, 0.2826177, 
    0.2539454, 0.2011659, 0.1340154, 0.1746824,
  0.1762168, 0.1261979, 0.1579493, 0.179248, 0.1669226, 0.1535704, 0.1913185, 
    0.1869665, 0.1581193, 0.1500058, 0.1257669, 0.164305, 0.1768093, 
    0.119789, 0.1666919, 0.1214157, 0.1129274, 0.1083293, 0.1120399, 
    0.1372831, 0.1471236, 0.1646766, 0.1869593, 0.1517145, 0.082647, 
    0.1535242, 0.1725975, 0.177657, 0.1765449,
  0.06855389, 0.03022257, 0.01947129, 0.08897328, 0.06430813, 0.04013875, 
    0.1077166, 0.1125523, 0.04021671, 0.02204867, 0.02763014, 0.02343484, 
    0.05713847, 0.1143272, 0.08211832, 0.04773724, 0.04407033, 0.06766796, 
    0.05740465, 0.1079149, 0.1455202, 0.09216035, 0.01989941, 0.02201036, 
    0.04401079, 0.06622387, 0.1258728, 0.1147877, 0.09089579,
  0.001294808, -8.284707e-07, 0.06239352, 0.03368484, 0.01784022, 0.09612425, 
    0.1046266, 0.02970227, 9.07069e-06, -0.0001627769, 0.09906369, 0.1320885, 
    0.04629463, 0.07045408, 0.03562522, 0.1074569, 0.0978045, 0.1997316, 
    0.3515893, 0.0630056, 0.09982824, 0.0007784404, 0.001464947, 0.003830132, 
    0.05940888, 0.06466924, 0.1276406, 0.05169651, 0.009230049,
  8.983288e-07, 0.07906463, 0.1156871, 0.01299428, 0.04169128, 0.01885376, 
    0.07384727, 0.02647589, -6.396993e-06, -1.273078e-09, 0.02149612, 
    0.01613701, 0.02017632, 0.007613977, 0.1031361, 0.02191784, 0.07653806, 
    0.02298615, 0.005551831, -5.837317e-06, 0.0001208337, 9.820861e-08, 
    2.98438e-06, 0.04237279, 0.07984438, 0.2055429, 0.05327393, 3.267398e-06, 
    7.610323e-07,
  0.0001577628, 0.02551183, 0.1054493, 0.03781594, 0.1365152, 0.1655721, 
    0.06803911, 0.07367315, 0.00753556, 0.003632202, 0.003858849, 0.0441657, 
    0.01499947, 0.01740024, 0.01965844, 0.03870997, 0.05663956, 0.005826251, 
    9.686965e-05, -3.894765e-13, 6.038067e-11, 1.878028e-08, 0.006715786, 
    0.04960282, 0.2007627, 0.0323486, 0.0001638516, -3.713143e-05, 
    1.649516e-05,
  0.04786363, 0.007501319, 0.0781159, 0.01024144, 0.01066903, 0.05844013, 
    0.03095392, 0.03664009, 0.01337203, 0.06437365, 0.02715009, 0.0208223, 
    0.02201633, 0.01365772, 0.0184342, 0.001175429, 0.00938923, 
    -2.044323e-05, -1.464592e-06, 3.903069e-07, 0.00565967, 0.00478835, 
    0.06452318, 0.08001546, 0.1039102, 0.08043379, 0.07852466, 0.06984382, 
    0.08180195,
  -6.343787e-10, 2.9053e-06, 3.450404e-06, 0.01082899, 0.00034356, 
    0.006097166, 0.000102674, 0.01614195, 0.001282522, 0.05348483, 0.1222022, 
    0.1102037, 0.03181122, 0.02611188, 0.04097829, 0.1147958, 0.0670769, 
    0.07200614, 0.1118305, 0.1584847, 0.178012, 0.02307265, 0.005660074, 
    0.002690393, 0.01920925, 0.02209598, 0.02471716, 0.00148437, -3.368253e-09,
  2.244303e-06, 3.089572e-06, 4.147727e-08, 3.251377e-07, -2.669144e-06, 
    5.140292e-07, 0.01626051, 0.0005476567, 7.217571e-05, 0.02200389, 
    0.1023637, 0.02050684, 0.0003570492, 0.005222414, 0.0006553685, 
    0.05749673, 0.01209383, 0.03985447, 0.09369732, 0.03117579, 0.02841879, 
    0.0002110523, 0.002560581, 0.0002954187, 0.002795391, 0.001123037, 
    0.03087023, 0.01291541, -0.0002011898,
  0.03077185, 0.01593483, 0.02091956, 0.01686845, 0.006732315, 0.0153, 
    0.0645755, 0.01256973, 0.03601013, 0.02675125, 0.04158901, 0.0547439, 
    0.06849765, 0.07015395, 0.0319223, 0.1170317, 0.05753598, 0.02115134, 
    0.03995604, 0.007243441, 0.09173702, 0.05877113, 0.03972052, 0.03437825, 
    0.02406922, 0.008546783, 0.04016613, 0.00377854, 0.05445214,
  0.03431335, 0.04684526, 0.1053474, 0.2523223, 0.1407359, 0.1945502, 
    0.1213793, 0.1172223, 0.09732954, 0.1011928, 0.1056161, 0.1366818, 
    0.1373693, 0.1793182, 0.1205161, 0.1976002, 0.2436615, 0.1395592, 
    0.1256736, 0.1858733, 0.08801877, 0.05970631, 0.1159858, 0.1813763, 
    0.1688746, 0.2070935, 0.06547421, 0.07371282, 0.05351909,
  0.1384905, 0.1859041, 0.2666557, 0.3238182, 0.2525215, 0.2808024, 
    0.2322581, 0.07331341, 0.03898145, 0.08918687, 0.150989, 0.06836699, 
    0.1954479, 0.2013996, 0.2177988, 0.2463987, 0.2583058, 0.1814629, 
    0.205707, 0.1345586, 0.1317189, 0.2100572, 0.1712535, 0.1650143, 
    0.1788492, 0.236117, 0.3412653, 0.2293174, 0.1573903,
  0.3065103, 0.2827128, 0.2339031, 0.2925279, 0.2904887, 0.2506993, 
    0.2394881, 0.203443, 0.2368007, 0.2538515, 0.1063478, 0.02635227, 
    0.01810776, 0.1442093, 0.1746586, 0.1616804, 0.3018843, 0.359779, 
    0.2393795, 0.226092, 0.3178917, 0.2280463, 0.1558415, 0.256749, 
    0.1877159, 0.1804966, 0.2367664, 0.274182, 0.3274885,
  0.1216359, 0.1761232, 0.1952112, 0.1008881, 0.08960634, 0.1657262, 
    0.2044961, 0.1752702, 0.09013837, 0.05575161, 0.003956924, 0.07367479, 
    0.04032594, 0.1419428, 0.1520984, 0.1379427, 0.195283, 0.2442007, 
    0.2591221, 0.1726643, 0.1283495, 0.07246628, 0.1574734, 0.1007638, 
    0.151309, 0.009028251, 0.03254518, 0.2045537, 0.1134835,
  0.1355256, 0.11224, 0.1521348, 0.155859, 0.1362025, 0.05689605, 0.07245199, 
    0.05358708, 0.03929468, 0.01069739, 0.03325517, 0.04660368, 0.04882864, 
    0.04198243, 0.02842082, 0.03636061, 0.0513085, 0.04519325, 0.1083461, 
    0.1309606, 0.09384222, 0.04870487, 0.00546263, -0.001578901, 
    -0.0007403266, 0.000739145, -0.005283376, 0.0622296, 0.1578107,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0.04740304, -0.002822329, -2.281479e-05, -2.842573e-06, 0, -0.001225611, 
    -0.0008349817, -0.0003485702, 0.0002259188, 0.003436735, -0.001008978, 0, 
    0.0001178537, 0.0905522, 0.1024411, 0.09393346, 0.1707575, 0.2937367, 
    0.09440593, 0.01628421, 0.01125539, 0.0224317, 0.1063013, 0.1072049, 
    0.05015572, 0.02598424, 0.02881357, 0.03690198, 0.06519789,
  0.1538557, 0.2415672, 0.1635264, 0.2361991, 0.2204552, 0.2017232, 
    0.3241106, 0.1767958, 0.1188162, 0.1517485, 0.08439428, 0.00216998, 
    0.09343019, 0.1629768, 0.1451872, 0.2023474, 0.1319063, 0.2188872, 
    0.160085, 0.2467187, 0.09205589, 0.1138312, 0.1783332, 0.3376634, 
    0.311296, 0.1587431, 0.234619, 0.1164079, 0.1622057,
  0.149439, 0.2989813, 0.3037284, 0.2508737, 0.1806539, 0.1677155, 0.1629214, 
    0.1254785, 0.1978081, 0.1352681, 0.2447999, 0.2630958, 0.2278226, 
    0.2584469, 0.1847144, 0.2021108, 0.155661, 0.1788554, 0.2040556, 
    0.2132084, 0.3138432, 0.293415, 0.2610591, 0.2464022, 0.2662151, 
    0.2468012, 0.205982, 0.1349917, 0.1794539,
  0.1836815, 0.1256045, 0.1553837, 0.176306, 0.1646588, 0.155556, 0.1920425, 
    0.1902164, 0.1702045, 0.1412559, 0.1319983, 0.1235696, 0.1572897, 
    0.1190706, 0.1562144, 0.08556623, 0.09469428, 0.09717707, 0.105827, 
    0.1351684, 0.1349362, 0.1493921, 0.1806725, 0.1611487, 0.07267433, 
    0.1490612, 0.1666591, 0.175838, 0.1730358,
  0.06333793, 0.02940497, 0.0175374, 0.09883554, 0.05983371, 0.03787135, 
    0.1134761, 0.1015158, 0.03330098, 0.01334704, 0.03397202, 0.02134605, 
    0.05672555, 0.1108883, 0.07184979, 0.03343023, 0.02941912, 0.06094171, 
    0.05045677, 0.1187818, 0.1268592, 0.07296475, 0.01754223, 0.01787445, 
    0.05315156, 0.06323456, 0.113924, 0.1058093, 0.07247803,
  0.004905699, -7.278363e-07, 0.05700291, 0.02922437, 0.02410933, 0.09724091, 
    0.08781293, 0.01891633, 1.959071e-06, 0.0003157629, 0.1045689, 0.1076248, 
    0.04348727, 0.0638238, 0.02614086, 0.1004931, 0.0573768, 0.1849441, 
    0.3137631, 0.05644911, 0.1043679, 0.0002596541, 0.002497688, 0.002931273, 
    0.06412016, 0.06713232, 0.1218684, 0.04765128, 0.01319397,
  1.290092e-06, 0.08674949, 0.1052916, 0.02246626, 0.04835002, 0.01568334, 
    0.06570832, 0.04481974, 1.560103e-06, -3.85788e-06, 0.03332557, 
    0.02044629, 0.0142067, 0.007315034, 0.09997338, 0.01848501, 0.08876658, 
    0.02068112, 0.006616032, -7.883365e-06, 0.001266166, 1.4855e-07, 
    5.778274e-06, 0.03284712, 0.1021842, 0.2326012, 0.04415025, 5.036584e-06, 
    5.770071e-07,
  0.006382731, 0.0413974, 0.1138711, 0.04780073, 0.1506065, 0.1663543, 
    0.07124367, 0.07162818, 0.009332171, 0.004360703, 0.004756288, 
    0.04732301, 0.01939892, 0.02247223, 0.02602549, 0.04209481, 0.05153945, 
    0.009691902, 0.0001952347, 9.408614e-10, 4.194984e-09, 5.787144e-09, 
    0.006190146, 0.05567094, 0.216308, 0.0403681, 0.0007597909, 
    -3.488517e-07, 0.0004090249,
  0.1037723, 0.01114589, 0.08390801, 0.02198828, 0.01122497, 0.04404709, 
    0.02015902, 0.05115426, 0.01964003, 0.08051812, 0.03075611, 0.01343865, 
    0.01433359, 0.0111414, 0.01843016, 0.0004611911, 0.003311215, 
    4.310644e-05, 1.664792e-07, 1.107713e-07, 0.0141824, 0.0002830735, 
    0.07589338, 0.1057602, 0.1030052, 0.07972994, 0.09759905, 0.05486508, 
    0.08303823,
  7.640383e-08, 1.924577e-06, -3.823988e-06, 0.008564014, 0.0002201261, 
    0.004813668, 0.0001257188, 0.009008927, 0.00186081, 0.04111412, 
    0.1533525, 0.1060982, 0.03811724, 0.03060283, 0.04571417, 0.1118887, 
    0.06623631, 0.08057267, 0.1185289, 0.1509517, 0.165004, 0.02423702, 
    0.007454135, 0.003940293, 0.0224867, 0.006144682, 0.007905817, 
    1.543903e-05, 2.700977e-08,
  5.94505e-07, 1.131876e-06, 3.623316e-08, -3.996121e-09, -9.913284e-05, 
    1.666649e-05, 0.01392348, 0.0001334332, -4.406526e-06, 0.02570507, 
    0.1136312, 0.01941884, 0.001336942, 0.01249119, 0.0007825329, 0.04959052, 
    0.01207703, 0.03766913, 0.09193122, 0.02300339, 0.0254219, 0.0003641095, 
    0.001603849, 0.001031823, 0.004009937, 0.002903767, 0.044712, 
    0.009594688, -4.551519e-05,
  0.009685897, 0.01438592, 0.02603701, 0.01509651, 0.008723598, 0.01236251, 
    0.05384422, 0.007594316, 0.09095387, 0.03646836, 0.03600888, 0.05097885, 
    0.06971649, 0.07613856, 0.02773484, 0.108376, 0.03729126, 0.01581029, 
    0.02980983, 0.002682364, 0.09416416, 0.05831453, 0.04308548, 0.03119872, 
    0.01540274, 0.00849963, 0.0405869, 0.003715887, 0.04418315,
  0.03353928, 0.04301113, 0.09028694, 0.2549643, 0.1290287, 0.1845185, 
    0.1623688, 0.1040846, 0.09379499, 0.09057473, 0.1003328, 0.1251363, 
    0.1280912, 0.1815607, 0.1011236, 0.1970177, 0.222357, 0.1241963, 
    0.1045357, 0.1780144, 0.09262791, 0.04221997, 0.1085165, 0.1713491, 
    0.1627009, 0.2105658, 0.05663424, 0.0730252, 0.06107284,
  0.1356554, 0.1755936, 0.2467037, 0.3236273, 0.2633087, 0.3106115, 
    0.2350682, 0.1818258, 0.06391945, 0.1038842, 0.1854939, 0.1255241, 
    0.2437691, 0.2336601, 0.2473742, 0.2533217, 0.2701009, 0.1854887, 
    0.2133705, 0.173287, 0.1332683, 0.2256845, 0.1691143, 0.1754035, 
    0.2037023, 0.2368475, 0.3477106, 0.2075887, 0.1441577,
  0.2982838, 0.2840711, 0.2414363, 0.3293518, 0.334826, 0.2821985, 0.225194, 
    0.2421134, 0.261939, 0.3063246, 0.1699634, 0.03083841, 0.06837933, 
    0.1795946, 0.2230063, 0.2030687, 0.3020497, 0.4269411, 0.3173007, 
    0.2322161, 0.3428298, 0.2298916, 0.1652341, 0.3218419, 0.2107954, 
    0.1985855, 0.2507926, 0.2597414, 0.335195,
  0.1624886, 0.2308644, 0.251337, 0.1452863, 0.1281488, 0.2496635, 0.223866, 
    0.2147788, 0.1497849, 0.1773039, 0.1006156, 0.1378532, 0.1465175, 
    0.2325999, 0.2319755, 0.1777783, 0.2047889, 0.258774, 0.2752391, 
    0.2187165, 0.1594286, 0.09255709, 0.2950537, 0.1749627, 0.1508093, 
    0.01782132, 0.05213339, 0.211016, 0.1132334,
  0.1805883, 0.1611085, 0.2452423, 0.1820764, 0.1725871, 0.0847727, 
    0.1394169, 0.1095899, 0.1120226, 0.07998516, 0.07820693, 0.09624511, 
    0.08876593, 0.07072802, 0.07775316, 0.1380907, 0.1459778, 0.16261, 
    0.2511141, 0.27337, 0.2157432, 0.1119989, 0.02144233, 0.01213858, 
    0.05712833, 0.01332299, 0.004434182, 0.1141403, 0.2582082,
  0.01928804, 0.01793282, 0.01657761, 0.01522239, 0.01386718, 0.01251196, 
    0.01115674, 0.002321166, 0.001937922, 0.001554678, 0.001171434, 
    0.0007881901, 0.0004049462, 2.170235e-05, -0.002446099, -0.001292832, 
    -0.0001395658, 0.001013701, 0.002166967, 0.003320234, 0.0044735, 
    0.01855199, 0.01913718, 0.01972237, 0.02030757, 0.02089276, 0.02147795, 
    0.02206315, 0.02037221,
  0.06665791, 0.01341033, 0.0006143667, 0.006529803, 0.00985131, 0.002609137, 
    0.008764177, 0.01703808, 0.0176223, 0.01544506, 0.00673556, 3.27606e-05, 
    0.0046704, 0.07008307, 0.1181578, 0.0956723, 0.1587864, 0.2576873, 
    0.07296041, 0.09221154, 0.02485522, 0.07255183, 0.1580939, 0.1068382, 
    0.04117099, 0.01638357, 0.02425906, 0.02905518, 0.07286996,
  0.149234, 0.2239173, 0.1475598, 0.2369126, 0.3304378, 0.2820016, 0.3176329, 
    0.2784794, 0.2051122, 0.15958, 0.1379813, 0.01814813, 0.1523078, 
    0.1467232, 0.1442909, 0.1892422, 0.1316383, 0.2140899, 0.1675122, 
    0.238512, 0.09635305, 0.1115006, 0.173251, 0.3403257, 0.291449, 
    0.1581731, 0.2000313, 0.1071609, 0.1476423,
  0.1599663, 0.2847285, 0.3180047, 0.2727061, 0.2005356, 0.1761822, 
    0.1937455, 0.1571976, 0.224812, 0.12657, 0.2724028, 0.2869081, 0.2260433, 
    0.2661991, 0.2019362, 0.218834, 0.1870203, 0.196939, 0.2404217, 
    0.2446619, 0.3208684, 0.3030967, 0.2682761, 0.2613726, 0.2553577, 
    0.2353412, 0.2180107, 0.1475498, 0.1704005,
  0.1902982, 0.1509227, 0.1515179, 0.1696176, 0.170035, 0.1604049, 0.1849004, 
    0.2045271, 0.1423673, 0.1458935, 0.1333423, 0.1468477, 0.1516369, 
    0.1154636, 0.1436765, 0.08491097, 0.08139428, 0.111303, 0.09993502, 
    0.1373815, 0.1270674, 0.1335645, 0.1585493, 0.1523761, 0.0737983, 
    0.1569173, 0.1538127, 0.1831786, 0.1679366,
  0.06704253, 0.03374305, 0.02400263, 0.09227522, 0.05380451, 0.03326032, 
    0.1212787, 0.100747, 0.03850218, 0.01367202, 0.03937043, 0.01796919, 
    0.06023319, 0.1115484, 0.06536071, 0.03231779, 0.02431666, 0.05971044, 
    0.04205886, 0.1133345, 0.1175288, 0.06497192, 0.02033753, 0.01616673, 
    0.0721776, 0.0523246, 0.1049454, 0.09769729, 0.06586463,
  0.009195398, -1.193607e-05, 0.06711525, 0.02832327, 0.03099008, 0.09444743, 
    0.08227074, 0.01917275, 8.198935e-07, 0.003948625, 0.07278176, 
    0.08743812, 0.04507872, 0.05687509, 0.0324509, 0.08470956, 0.04910463, 
    0.2005911, 0.2881392, 0.04790931, 0.1111051, 0.0002522974, 0.002606266, 
    0.003511105, 0.08689147, 0.07238933, 0.1192463, 0.04188038, 0.01243376,
  0.0001728689, 0.1192448, 0.1147203, 0.02669533, 0.05415341, 0.02258914, 
    0.05887296, 0.0473571, 1.142612e-05, 0.000139179, 0.06205472, 0.02895048, 
    0.01798424, 0.008929349, 0.1204177, 0.02450275, 0.09961294, 0.02704121, 
    0.009469006, 0.0002096981, 0.0005848091, 1.934582e-07, 7.576293e-06, 
    0.02857532, 0.1356553, 0.264388, 0.04758959, 1.714328e-05, 2.276645e-06,
  0.008702875, 0.08080884, 0.1491907, 0.07178889, 0.1659382, 0.1893146, 
    0.07158035, 0.0778347, 0.01256292, 0.004388659, 0.006182084, 0.05122594, 
    0.03661684, 0.02199906, 0.03999572, 0.04246121, 0.0467444, 0.01848252, 
    0.0001232609, 9.341042e-09, 1.410409e-08, 5.707567e-08, 0.004558949, 
    0.06985157, 0.2616722, 0.06197523, 0.0006984768, 1.899946e-07, 0.006366336,
  0.1092874, 0.02645036, 0.09763218, 0.02360745, 0.01379493, 0.04512987, 
    0.01963715, 0.08239169, 0.03054531, 0.1042897, 0.03390983, 0.01457618, 
    0.0187019, 0.01266378, 0.01533957, 0.0003414694, 0.002268119, 
    8.533914e-05, 8.412418e-07, 2.665502e-05, 0.01592096, 0.01011933, 
    0.09428525, 0.1375096, 0.1325191, 0.0745935, 0.1054844, 0.05445285, 
    0.09310386,
  3.334534e-07, 1.566384e-06, -4.060549e-07, 0.004597072, 0.0003197463, 
    0.01113355, 0.0007556098, 0.007540744, 0.00980151, 0.04502454, 0.183805, 
    0.1213479, 0.04805436, 0.03359824, 0.05444747, 0.111446, 0.06630587, 
    0.07979769, 0.1188557, 0.1585292, 0.1587511, 0.02680597, 0.01512869, 
    0.005497827, 0.02375231, 0.0153068, 0.01421435, 4.199113e-06, 1.139954e-07,
  2.459798e-06, 3.234764e-07, 3.219098e-08, 4.521099e-05, -0.0003558196, 
    8.749678e-05, 0.0185881, 0.003691063, 3.915083e-07, 0.03869695, 
    0.1372088, 0.02729297, 0.002079674, 0.01439878, 0.0009675255, 0.05044353, 
    0.01534514, 0.04322348, 0.07846623, 0.02176112, 0.02396767, 0.0009230696, 
    0.002646114, 0.001625758, 0.006529254, 0.003441081, 0.03877785, 
    0.00260998, 3.034168e-06,
  0.01803641, 0.01216051, 0.008535129, 0.01220199, 0.01093754, 0.0158693, 
    0.03607017, 0.01452799, 0.1140604, 0.02558855, 0.03806895, 0.04906962, 
    0.06620726, 0.07299429, 0.03186807, 0.0889084, 0.02366417, 0.01145462, 
    0.01805113, 0.007299605, 0.08551672, 0.05599048, 0.06183814, 0.04163675, 
    0.008074922, 0.02163677, 0.04215552, 0.005374672, 0.03597662,
  0.03001823, 0.03772506, 0.08535089, 0.2582347, 0.113126, 0.17678, 
    0.2129794, 0.09121739, 0.07510971, 0.08539785, 0.07834382, 0.09986966, 
    0.1285212, 0.1684124, 0.0982678, 0.197986, 0.1957838, 0.113701, 
    0.08892841, 0.176456, 0.09486851, 0.02695943, 0.1057661, 0.17, 0.1691378, 
    0.198062, 0.05015685, 0.07929284, 0.05864182,
  0.1213115, 0.1972286, 0.2590279, 0.3416868, 0.264216, 0.2895209, 0.228867, 
    0.1805593, 0.07406915, 0.1064088, 0.2132982, 0.1463658, 0.2546114, 
    0.2412176, 0.2308238, 0.2505648, 0.2460697, 0.1875797, 0.2052497, 
    0.1918052, 0.1299895, 0.2285529, 0.1693738, 0.195353, 0.2111194, 
    0.2230052, 0.3449768, 0.1900108, 0.1474132,
  0.2797417, 0.2848665, 0.27742, 0.3097165, 0.3388147, 0.2903242, 0.1864081, 
    0.215087, 0.2758116, 0.3021449, 0.1828714, 0.07132727, 0.0956429, 
    0.1970406, 0.2204049, 0.2165352, 0.3155978, 0.4277409, 0.3687603, 
    0.2258421, 0.3322443, 0.2309344, 0.2005878, 0.3300107, 0.2259041, 
    0.2218382, 0.2413468, 0.2562945, 0.3372914,
  0.1695327, 0.2275007, 0.2485013, 0.1632364, 0.1676055, 0.2831503, 
    0.2772748, 0.28463, 0.166959, 0.2483433, 0.2138098, 0.2126196, 0.1810057, 
    0.2545273, 0.2770835, 0.1884083, 0.2141508, 0.239752, 0.2716466, 
    0.2160352, 0.1726134, 0.1015759, 0.3169096, 0.235405, 0.1561757, 
    0.09501228, 0.06711081, 0.2125359, 0.1216765,
  0.1669265, 0.1477025, 0.2320147, 0.1636776, 0.1489803, 0.09494659, 
    0.1492623, 0.1542965, 0.1778245, 0.1526099, 0.1431664, 0.1841323, 
    0.2134493, 0.1467245, 0.13296, 0.1425091, 0.1706787, 0.2083704, 
    0.2713768, 0.2631064, 0.2275495, 0.1384902, 0.1007189, 0.04250091, 
    0.1613553, 0.06998297, 0.06572665, 0.2456559, 0.262033,
  0.0173764, 0.01779843, 0.01822047, 0.0186425, 0.01906453, 0.01948656, 
    0.01990859, 0.02669377, 0.02653978, 0.02638578, 0.02623179, 0.0260778, 
    0.02592381, 0.02576982, 0.02550416, 0.02594514, 0.02638613, 0.02682712, 
    0.02726811, 0.02770909, 0.02815008, 0.02312566, 0.02241664, 0.02170761, 
    0.02099858, 0.02028955, 0.01958053, 0.0188715, 0.01703878,
  0.08174979, 0.01748203, -0.0005449777, 0.01896414, 0.01420932, 0.005391232, 
    0.03369257, 0.03265461, 0.01679165, 0.02078542, 0.006738094, 0.03289081, 
    0.03361417, 0.05560476, 0.1332364, 0.1213372, 0.1859957, 0.1946669, 
    0.04005292, 0.09039269, 0.05728771, 0.1963674, 0.1480035, 0.1006002, 
    0.0364067, 0.01237392, 0.02063006, 0.02405842, 0.0658957,
  0.1698385, 0.2393535, 0.1499372, 0.2394272, 0.4083303, 0.3475728, 
    0.3207838, 0.2973716, 0.2081368, 0.1548038, 0.1313635, 0.03055222, 
    0.1674082, 0.161349, 0.185005, 0.1872936, 0.1577, 0.2356146, 0.1835394, 
    0.1933331, 0.09445382, 0.1190639, 0.1777382, 0.3328421, 0.3184816, 
    0.1671854, 0.175352, 0.09769707, 0.1367743,
  0.1696935, 0.2605125, 0.3364408, 0.3009357, 0.2649218, 0.1767713, 
    0.2164383, 0.128466, 0.2406073, 0.1672444, 0.300142, 0.2733987, 
    0.2516519, 0.2996896, 0.2307999, 0.2635252, 0.1939434, 0.2055365, 
    0.2558158, 0.2543288, 0.3785514, 0.3063211, 0.2713139, 0.2623332, 
    0.2624598, 0.2498649, 0.2522981, 0.1725298, 0.1659833,
  0.2121465, 0.1624066, 0.1508904, 0.1774631, 0.189872, 0.1935488, 0.1839624, 
    0.2078765, 0.1409682, 0.1758711, 0.1278531, 0.1403477, 0.1484009, 
    0.1071855, 0.1322798, 0.09239024, 0.07764053, 0.09808376, 0.08851738, 
    0.1557906, 0.1428012, 0.170491, 0.1594515, 0.1442027, 0.08406887, 
    0.1785498, 0.13554, 0.1775889, 0.1745825,
  0.05650809, 0.03565011, 0.01079203, 0.0816294, 0.05120836, 0.03420668, 
    0.1195609, 0.1073733, 0.03333578, 0.01400463, 0.03702891, 0.01774649, 
    0.06195881, 0.1146373, 0.05911054, 0.03252878, 0.02979315, 0.04745125, 
    0.03601614, 0.1076338, 0.123652, 0.05864421, 0.0245832, 0.01912885, 
    0.08594767, 0.0499737, 0.1078036, 0.09360662, 0.07054143,
  0.005351748, -1.078993e-06, 0.09067474, 0.03469282, 0.04052053, 0.08810627, 
    0.08103099, 0.005578053, 1.648617e-06, 0.005790634, 0.03554534, 
    0.07474071, 0.05545893, 0.05572879, 0.03694722, 0.07018974, 0.04423486, 
    0.2044212, 0.2815469, 0.04548994, 0.1158347, 3.82647e-06, 0.001764812, 
    0.004335613, 0.1071518, 0.0969402, 0.1232071, 0.0442214, 0.02161636,
  0.002753202, 0.1606559, 0.1398349, 0.03154476, 0.055705, 0.03549987, 
    0.05514704, 0.05440577, 1.258947e-05, 1.131109e-06, 0.06895887, 
    0.02727711, 0.02673933, 0.007747358, 0.1254546, 0.03562893, 0.09750667, 
    0.03796979, 0.01314742, 0.0004264954, 1.595162e-05, 9.436247e-08, 
    2.232995e-06, 0.0261388, 0.1695653, 0.2924613, 0.04842637, 8.077885e-05, 
    9.974319e-06,
  0.001458782, 0.09509122, 0.183245, 0.08989532, 0.1891117, 0.1904602, 
    0.08189661, 0.08902174, 0.01478875, 0.004342925, 0.006639001, 0.05174465, 
    0.04551908, 0.02719688, 0.05406288, 0.04881638, 0.04265105, 0.03914879, 
    0.002941922, 1.403832e-06, 2.015495e-08, 3.366029e-08, 0.00201689, 
    0.1028454, 0.2981203, 0.08584812, 0.0009727892, 2.106792e-07, 0.007242391,
  0.1142622, 0.04303896, 0.1166219, 0.02089932, 0.01955498, 0.04227512, 
    0.03238845, 0.1196129, 0.0456665, 0.125697, 0.03503131, 0.01833072, 
    0.02041968, 0.01883579, 0.01757406, 0.0003356977, -0.0001233335, 
    0.0008868865, 6.56727e-07, 0.0001016883, 0.007058949, 0.005066988, 
    0.1100294, 0.1792725, 0.166565, 0.07486181, 0.1081013, 0.06008714, 
    0.09647978,
  6.143268e-07, 3.991699e-06, 3.365935e-05, 0.0009605096, 0.001114301, 
    0.01689355, 0.002494314, 0.01383208, 0.01216491, 0.05137001, 0.2136296, 
    0.1266086, 0.0533609, 0.03536452, 0.06175369, 0.117828, 0.06730168, 
    0.08747655, 0.1196923, 0.1498662, 0.1673335, 0.03222091, 0.02765977, 
    0.007009376, 0.02501187, 0.01522644, 0.01239215, 1.258446e-06, 
    3.223931e-07,
  1.620014e-06, 2.720747e-07, 8.56444e-08, 0.0007533125, -0.0004970111, 
    5.130896e-05, 0.02322662, 0.008238348, 2.631947e-07, 0.04521514, 
    0.1881579, 0.03242727, 0.004305656, 0.01679288, 0.00150344, 0.05294415, 
    0.02370811, 0.0407021, 0.06834047, 0.01759911, 0.02569994, 0.007499506, 
    0.002856853, 0.00320051, 0.008535963, 0.004635304, 0.03507818, 
    -2.790971e-05, -0.0002372955,
  0.005212637, 0.007337618, -0.0004447381, 0.0139607, 0.009713918, 0.023478, 
    0.02741791, 0.01848583, 0.1280433, 0.03131877, 0.03781525, 0.04357089, 
    0.06278266, 0.08027316, 0.04712788, 0.09240884, 0.02342458, 0.01097172, 
    0.01592284, 0.009451646, 0.06730057, 0.06200153, 0.06698796, 0.03277216, 
    0.009711869, 0.02686661, 0.04720996, 0.01277164, 0.04064132,
  0.02591881, 0.03175033, 0.09201142, 0.271663, 0.1142784, 0.1552012, 
    0.2281938, 0.0805046, 0.05688184, 0.07248205, 0.06275342, 0.08412192, 
    0.1370268, 0.1409076, 0.1032436, 0.1888843, 0.1895332, 0.1029557, 
    0.07582476, 0.1646062, 0.1080501, 0.01958741, 0.1036154, 0.1786962, 
    0.1657787, 0.1965317, 0.05881444, 0.094159, 0.05363869,
  0.1244167, 0.2071563, 0.2577317, 0.3607354, 0.2557805, 0.2705529, 
    0.2349776, 0.1788855, 0.08168499, 0.09777597, 0.2012804, 0.156627, 
    0.2505018, 0.2364737, 0.2248653, 0.2215803, 0.2453576, 0.1788203, 
    0.220202, 0.2136126, 0.1449802, 0.2200813, 0.1708066, 0.2111882, 
    0.209689, 0.230867, 0.3479098, 0.1782151, 0.1429973,
  0.2631557, 0.2808748, 0.2929935, 0.3140116, 0.3018642, 0.2845311, 
    0.1681489, 0.1954434, 0.2517041, 0.3151724, 0.2099926, 0.1003651, 
    0.1094136, 0.1932728, 0.2134679, 0.2431428, 0.2813821, 0.4367213, 
    0.3456942, 0.2388388, 0.3460597, 0.2230785, 0.2476531, 0.337891, 
    0.2524272, 0.212972, 0.2369138, 0.2460871, 0.3026913,
  0.1593298, 0.2117013, 0.2470283, 0.1662869, 0.1699121, 0.3009782, 
    0.3086993, 0.3472073, 0.1975479, 0.3123837, 0.2818557, 0.203957, 
    0.1873424, 0.31625, 0.2936398, 0.1879022, 0.2217835, 0.2404385, 
    0.2699804, 0.1903608, 0.176338, 0.1122314, 0.3127989, 0.2300634, 
    0.1620013, 0.1381, 0.09840803, 0.2133667, 0.1196495,
  0.1496109, 0.1498923, 0.211614, 0.1500647, 0.1274458, 0.09244128, 
    0.1588445, 0.1632123, 0.1800426, 0.178775, 0.1803759, 0.2270039, 
    0.2378862, 0.2002635, 0.1583343, 0.1576095, 0.1563046, 0.2279301, 
    0.3249426, 0.3336618, 0.2342214, 0.1744039, 0.1661346, 0.05443578, 
    0.2185987, 0.1121349, 0.111656, 0.267989, 0.2544203,
  0.01373157, 0.01418531, 0.01463905, 0.0150928, 0.01554654, 0.01600028, 
    0.01645402, 0.01774929, 0.01788789, 0.0180265, 0.0181651, 0.0183037, 
    0.01844231, 0.01858091, 0.01944239, 0.01909094, 0.01873949, 0.01838804, 
    0.0180366, 0.01768515, 0.0173337, 0.01740892, 0.01716802, 0.01692712, 
    0.01668623, 0.01644533, 0.01620443, 0.01596353, 0.01336858,
  0.07081497, 0.05544846, 0.01093174, 0.04698236, 0.04148982, 0.03337805, 
    0.04836712, 0.04515111, 0.03385691, 0.02657039, 0.02381436, 0.07178587, 
    0.03861383, 0.0363613, 0.1459063, 0.1727107, 0.1874013, 0.1577497, 
    0.02566485, 0.06658846, 0.0590037, 0.1943939, 0.1410345, 0.1140101, 
    0.02709185, 0.009555542, 0.01862106, 0.02286922, 0.06209382,
  0.1789121, 0.2596498, 0.1706747, 0.2446678, 0.4384571, 0.3648804, 
    0.3340131, 0.2708064, 0.1865319, 0.1507717, 0.09960307, 0.07031517, 
    0.1713267, 0.1608342, 0.2162165, 0.224767, 0.2247697, 0.238754, 
    0.1991997, 0.2070716, 0.1486217, 0.1292019, 0.1756722, 0.3449117, 
    0.3281823, 0.1876382, 0.1680455, 0.08619668, 0.1086991,
  0.2627272, 0.2880513, 0.2984214, 0.2774767, 0.3056574, 0.2740465, 
    0.2887117, 0.2276992, 0.2209031, 0.1780887, 0.2823861, 0.2984276, 
    0.2612438, 0.3149104, 0.2255138, 0.271205, 0.2016758, 0.1851646, 
    0.2529229, 0.2804425, 0.3852289, 0.2832785, 0.3026642, 0.3000951, 
    0.2895937, 0.2406417, 0.2372172, 0.2003076, 0.2021404,
  0.1824835, 0.1643211, 0.1627494, 0.1914571, 0.1832983, 0.187476, 0.1723883, 
    0.2063244, 0.1568852, 0.144509, 0.1527555, 0.1585836, 0.1489387, 
    0.1159958, 0.1208828, 0.09924003, 0.0875003, 0.09258793, 0.09893408, 
    0.1740219, 0.145516, 0.1611879, 0.1406406, 0.1406517, 0.0944218, 0.17348, 
    0.1227048, 0.1794315, 0.1867068,
  0.06995258, 0.03736642, 0.01574672, 0.07005688, 0.05468042, 0.03410889, 
    0.1214337, 0.1162323, 0.03078921, 0.01635218, 0.02208889, 0.01740456, 
    0.0628351, 0.1267366, 0.06098377, 0.02734462, 0.0338046, 0.0514584, 
    0.04142051, 0.1191251, 0.1221012, 0.06817094, 0.03271125, 0.02473145, 
    0.1032508, 0.04219782, 0.1060126, 0.0946769, 0.07158002,
  0.008639346, -1.760472e-07, 0.1041417, 0.03090906, 0.05038135, 0.0886948, 
    0.07452883, 0.0007332183, 3.567221e-06, 0.007549788, 0.01518908, 
    0.06686419, 0.05897867, 0.05951731, 0.04724385, 0.08067197, 0.04548765, 
    0.2116498, 0.2868899, 0.03777057, 0.1320508, 0.000142867, 0.0001225302, 
    0.004875956, 0.1017617, 0.1028027, 0.1387479, 0.05047331, 0.03428416,
  0.004458109, 0.1836302, 0.1782852, 0.02649953, 0.05461399, 0.03042638, 
    0.05681192, 0.04741098, 9.862222e-06, 2.596341e-07, 0.06563622, 
    0.04645682, 0.01485214, 0.0051363, 0.1221588, 0.02973637, 0.07569171, 
    0.04049531, 0.01202398, 0.006159202, 3.440253e-06, 2.98434e-08, 
    5.138573e-07, 0.00912948, 0.1395994, 0.3439746, 0.03618883, 0.0005297322, 
    2.487553e-05,
  0.0001241664, 0.05108501, 0.232554, 0.1011201, 0.1473592, 0.175669, 
    0.07901311, 0.0718658, 0.01693111, 0.004253315, 0.006829031, 0.03452811, 
    0.0314272, 0.02623049, 0.04572999, 0.05029109, 0.04539817, 0.06018553, 
    0.004646109, -1.894436e-06, 1.689963e-08, 2.91992e-08, 0.00021622, 
    0.09816566, 0.2783901, 0.1073957, 0.004488199, -7.395926e-07, 0.002178126,
  0.1022686, 0.07087249, 0.1399537, 0.03233939, 0.02263983, 0.0352963, 
    0.04041139, 0.1101496, 0.05950793, 0.1450551, 0.03453156, 0.01146217, 
    0.01080344, 0.02235634, 0.01839451, 0.0003786016, -0.0001351598, 
    0.0003743994, 3.703232e-07, 7.770691e-05, 0.00121803, 0.002949315, 
    0.1323232, 0.1825466, 0.1596041, 0.06657162, 0.1002048, 0.06951034, 
    0.09731092,
  4.623898e-07, 1.366208e-06, 1.149711e-05, 0.0007651825, 0.006028443, 
    0.02446629, 0.003372634, 0.006121288, 0.01120244, 0.04467909, 0.2117769, 
    0.1046088, 0.05350955, 0.03568482, 0.06027493, 0.101043, 0.06509327, 
    0.1053861, 0.1242494, 0.1476323, 0.1665797, 0.03504258, 0.04548953, 
    0.00782709, 0.02419298, 0.01141545, 0.004873784, -9.921295e-07, 
    6.847982e-06,
  4.948355e-07, 2.820839e-07, 8.765171e-08, 0.00404812, 0.001108884, 
    0.0002982022, 0.02828635, 0.02561672, 0.0001713051, 0.04386676, 
    0.1925212, 0.03012452, 0.006685576, 0.01437649, 0.003085998, 0.05926796, 
    0.03376634, 0.0343253, 0.07824443, 0.02753313, 0.02713761, 0.01145431, 
    0.00532006, 0.006623505, 0.02424343, 0.01326483, 0.03678349, 0.002125323, 
    -1.567683e-05,
  -1.305333e-05, 0.00690776, -1.321426e-05, 0.01851908, 0.01782126, 
    0.02675978, 0.03445096, 0.02544366, 0.1322832, 0.03527945, 0.04907028, 
    0.03638143, 0.06116523, 0.08476928, 0.06922553, 0.1124528, 0.02945457, 
    0.01158029, 0.01867133, 0.01619735, 0.05867829, 0.07065815, 0.07436681, 
    0.03441011, 0.02784302, 0.02897354, 0.05795381, 0.01594867, 0.02343474,
  0.02457108, 0.0294964, 0.1201457, 0.2867911, 0.1171614, 0.1440123, 
    0.2330834, 0.06130035, 0.04492778, 0.05944901, 0.05274947, 0.07985649, 
    0.1448427, 0.1289544, 0.1049485, 0.1870352, 0.17773, 0.08531692, 
    0.06837358, 0.1690674, 0.1161359, 0.02408572, 0.1143126, 0.1845522, 
    0.1808937, 0.1882045, 0.0780424, 0.08599712, 0.05062072,
  0.1309215, 0.2323657, 0.2761362, 0.3138207, 0.2240541, 0.2666665, 
    0.2381739, 0.1728055, 0.1009859, 0.08756613, 0.183658, 0.1557893, 
    0.2391171, 0.2302415, 0.2375265, 0.2317013, 0.2617202, 0.197567, 
    0.2377189, 0.2100841, 0.1417469, 0.2027419, 0.16868, 0.1943554, 
    0.2164777, 0.2311254, 0.3345222, 0.1758233, 0.1434536,
  0.2882098, 0.3322974, 0.3554989, 0.3179464, 0.3551426, 0.27186, 0.1718298, 
    0.1792093, 0.2197789, 0.3313188, 0.2649076, 0.1100572, 0.1432426, 
    0.1813824, 0.1997504, 0.2475359, 0.2780232, 0.4272366, 0.3305419, 
    0.245991, 0.3407515, 0.2110767, 0.2582952, 0.3235911, 0.230577, 
    0.2119616, 0.2524828, 0.2480185, 0.3114841,
  0.1728835, 0.2383886, 0.2462218, 0.2141553, 0.167765, 0.3325612, 0.3195488, 
    0.3742147, 0.2363784, 0.3136969, 0.3106299, 0.2023875, 0.197928, 
    0.3302615, 0.3198281, 0.1869484, 0.191759, 0.2531424, 0.2526376, 
    0.195848, 0.1753799, 0.118442, 0.3365135, 0.2199643, 0.1641232, 
    0.1595117, 0.1323038, 0.2214652, 0.1393891,
  0.1375715, 0.1527124, 0.1742023, 0.1600761, 0.1372079, 0.1043672, 
    0.1694048, 0.190494, 0.1977179, 0.2090381, 0.2468208, 0.2358637, 
    0.2359584, 0.2324042, 0.207557, 0.1730839, 0.1544222, 0.2178079, 
    0.3224688, 0.3390788, 0.3024254, 0.2661813, 0.1887612, 0.05740255, 
    0.2172642, 0.1340754, 0.1656633, 0.2543055, 0.2334418,
  0.01948795, 0.01999178, 0.0204956, 0.02099943, 0.02150326, 0.02200708, 
    0.02251091, 0.02121833, 0.02115464, 0.02109096, 0.02102728, 0.0209636, 
    0.02089992, 0.02083623, 0.02214329, 0.02199246, 0.02184163, 0.0216908, 
    0.02153997, 0.02138914, 0.02123831, 0.02178883, 0.02149951, 0.0212102, 
    0.02092089, 0.02063157, 0.02034226, 0.02005295, 0.01908489,
  0.06006323, 0.04815568, 0.009812225, 0.04693641, 0.0674551, 0.07058007, 
    0.06797649, 0.04290587, 0.07494526, 0.07582253, 0.04295386, 0.0556556, 
    0.03411328, 0.01612616, 0.07360415, 0.1114655, 0.1377219, 0.1429565, 
    0.01932906, 0.04994477, 0.05891785, 0.1942648, 0.1349849, 0.100089, 
    0.03070481, 0.0122659, 0.01674683, 0.02183134, 0.06208333,
  0.1498075, 0.2378662, 0.193638, 0.2436757, 0.4250152, 0.3866665, 0.3125326, 
    0.2900988, 0.1645001, 0.1126129, 0.07829773, 0.07545809, 0.1784429, 
    0.1627757, 0.2061235, 0.2136167, 0.18536, 0.3039055, 0.2166773, 
    0.2812903, 0.1425502, 0.1683239, 0.1738625, 0.3900398, 0.3299363, 
    0.3408439, 0.1662917, 0.07539722, 0.09231729,
  0.3867838, 0.3806664, 0.4711367, 0.4318385, 0.3575238, 0.3379093, 
    0.3686211, 0.2033549, 0.2717041, 0.223889, 0.3684433, 0.2510142, 
    0.2649046, 0.2929145, 0.2463438, 0.2330945, 0.2171993, 0.2305739, 
    0.3275294, 0.3004706, 0.3378247, 0.284784, 0.3245278, 0.2962834, 
    0.2547039, 0.212008, 0.249094, 0.2233504, 0.2700662,
  0.2068284, 0.192081, 0.1707616, 0.1845437, 0.2112128, 0.1831297, 0.17318, 
    0.2306288, 0.1647563, 0.1678603, 0.1807967, 0.15583, 0.1576457, 
    0.1105188, 0.1259306, 0.1216592, 0.09722733, 0.08277744, 0.1007626, 
    0.1809264, 0.1474272, 0.1587311, 0.1454181, 0.1351069, 0.0875667, 
    0.1649727, 0.1089916, 0.175436, 0.1780649,
  0.08107994, 0.03430621, 0.0184648, 0.05921375, 0.05348497, 0.04286224, 
    0.1304345, 0.1273403, 0.03738252, 0.01709128, 0.01671606, 0.01813672, 
    0.05935643, 0.1568563, 0.06735469, 0.02500194, 0.05001394, 0.06896953, 
    0.04934811, 0.1290736, 0.1193468, 0.08003195, 0.04971467, 0.03353621, 
    0.07435917, 0.04882771, 0.1011484, 0.09469591, 0.09056913,
  0.007173665, 1.550153e-08, 0.1102379, 0.02805991, 0.07890212, 0.09090043, 
    0.06608274, -0.0001793548, 5.198408e-06, 0.002478154, 0.004073878, 
    0.03584837, 0.07270751, 0.06565304, 0.06953185, 0.09320506, 0.05124229, 
    0.23631, 0.2967461, 0.03158962, 0.1481751, 0.001906959, 4.124846e-06, 
    0.003907991, 0.06927349, 0.1111365, 0.1763212, 0.06661871, 0.01824183,
  0.001167986, 0.1312409, 0.1841904, 0.01764293, 0.05539639, 0.03234063, 
    0.05497064, 0.03482069, 3.526436e-06, 1.186073e-07, 0.04401726, 
    0.05150576, 0.00996243, 0.006470676, 0.1334649, 0.02946944, 0.0615619, 
    0.04259056, 0.02353509, 0.01422393, 3.034779e-06, 7.596544e-09, 
    1.060995e-07, 0.0029569, 0.1223404, 0.3530416, 0.01781147, 0.0002466536, 
    2.562445e-05,
  7.797296e-05, 0.01110461, 0.2515158, 0.09623672, 0.1165547, 0.1546423, 
    0.0723749, 0.06567483, 0.01624136, 0.004574748, 0.00777198, 0.02743629, 
    0.02699477, 0.02474041, 0.03935194, 0.05178468, 0.03981283, 0.07014912, 
    0.004680522, 5.771556e-05, 1.406107e-08, 9.892655e-09, 4.85944e-05, 
    0.07043356, 0.1816188, 0.08709621, 0.004552804, -6.617427e-06, 
    -0.0003538612,
  0.07573183, 0.0861784, 0.113264, 0.04474678, 0.02588014, 0.03386982, 
    0.03506492, 0.1066058, 0.07540133, 0.1498351, 0.03201937, 0.008835451, 
    0.00878535, 0.0192466, 0.01639737, 0.0004718071, -5.671527e-05, 
    1.607602e-05, 2.3749e-07, 0.001182027, 0.001012407, 0.0001022002, 
    0.1163633, 0.1482398, 0.1372095, 0.05041967, 0.1086355, 0.06106612, 
    0.09852993,
  3.240002e-07, 3.030666e-05, 0.0002781055, 0.00877671, 0.01269952, 
    0.02363317, 0.0069287, 0.00529831, 0.02067083, 0.04423135, 0.2132792, 
    0.09291708, 0.05229574, 0.03864666, 0.06054597, 0.08703795, 0.06703975, 
    0.1142242, 0.1104571, 0.1302403, 0.149644, 0.03839524, 0.06027221, 
    0.01438154, 0.03952662, 0.007314778, 0.003230215, -5.201602e-06, 
    9.951057e-05,
  2.863036e-07, 3.102786e-07, 5.099705e-08, 0.009306379, 0.00926662, 
    -1.411665e-05, 0.02824264, 0.03765879, 0.008808747, 0.0396166, 0.1866361, 
    0.02998307, 0.008155995, 0.01186927, 0.005893541, 0.0600549, 0.03741642, 
    0.03135844, 0.09359322, 0.03333838, 0.01332536, 0.03426455, 0.00542301, 
    0.01585217, 0.03353387, 0.02050066, 0.02142833, 0.000331036, 6.976729e-06,
  1.70992e-05, 0.009708933, 0.0005123422, 0.02267947, 0.03677471, 0.03482333, 
    0.04087769, 0.04033615, 0.1226544, 0.04767346, 0.04531419, 0.02681681, 
    0.06668941, 0.1004588, 0.1009441, 0.1430968, 0.03774584, 0.01461667, 
    0.03217886, 0.02323029, 0.05179132, 0.08516004, 0.06185156, 0.05056803, 
    0.04246012, 0.03269774, 0.05995753, 0.01613339, 0.007770641,
  0.02578368, 0.03309543, 0.1195092, 0.3074122, 0.1086541, 0.1398721, 
    0.2411717, 0.0500522, 0.03450016, 0.0511772, 0.04054974, 0.08691698, 
    0.1592832, 0.1204166, 0.1172667, 0.1820985, 0.1764782, 0.0870335, 
    0.07355368, 0.1736893, 0.1201483, 0.03359965, 0.1146693, 0.1738272, 
    0.1917219, 0.2046256, 0.09293208, 0.08945365, 0.05096475,
  0.1326513, 0.2479236, 0.2494228, 0.2731403, 0.2523279, 0.2869194, 
    0.2319674, 0.1826928, 0.1036653, 0.08454183, 0.162214, 0.1446349, 
    0.2283365, 0.2328887, 0.2541385, 0.2329691, 0.2631033, 0.2124401, 
    0.2322839, 0.2229724, 0.1794164, 0.1885101, 0.1676697, 0.2363138, 
    0.2371595, 0.2356894, 0.3461286, 0.1779339, 0.1442853,
  0.2596534, 0.3404025, 0.3104829, 0.309601, 0.3567082, 0.2941984, 0.1965254, 
    0.1639358, 0.2199867, 0.3302667, 0.2809783, 0.1155047, 0.1558618, 
    0.1871365, 0.1974415, 0.2340889, 0.2581405, 0.4434469, 0.3204863, 
    0.2215078, 0.3379123, 0.2082468, 0.2964773, 0.3381293, 0.2295616, 
    0.236739, 0.2545466, 0.2471269, 0.3107815,
  0.1745648, 0.2437185, 0.233208, 0.2654443, 0.2184076, 0.4307477, 0.4132003, 
    0.3951569, 0.2788002, 0.3166504, 0.3211245, 0.2178777, 0.2061147, 
    0.3365104, 0.3654704, 0.1918211, 0.1835729, 0.2869803, 0.234323, 
    0.1981672, 0.1877092, 0.1420124, 0.348472, 0.2801143, 0.1698928, 
    0.169394, 0.2115765, 0.2308752, 0.1485511,
  0.1290794, 0.1525822, 0.1956342, 0.2219906, 0.2031874, 0.1462736, 
    0.2153878, 0.2677741, 0.281213, 0.303999, 0.2822263, 0.2723008, 
    0.2979657, 0.2722217, 0.2712581, 0.2482421, 0.1783354, 0.2481438, 
    0.3398486, 0.3273682, 0.2976224, 0.3139067, 0.2224656, 0.06409279, 
    0.1951286, 0.1616117, 0.1736764, 0.2635897, 0.2215142,
  0.02719259, 0.02769588, 0.02819918, 0.02870247, 0.02920576, 0.02970905, 
    0.03021234, 0.02562701, 0.02509082, 0.02455464, 0.02401845, 0.02348226, 
    0.02294608, 0.02240989, 0.02253769, 0.02243512, 0.02233256, 0.02222999, 
    0.02212742, 0.02202485, 0.02192228, 0.0235111, 0.02364657, 0.02378203, 
    0.02391749, 0.02405296, 0.02418842, 0.02432388, 0.02678996,
  0.0475177, 0.04383528, 0.007915915, 0.04667599, 0.1145565, 0.1071266, 
    0.1010349, 0.05631923, 0.1043368, 0.07277079, 0.04120353, 0.05011315, 
    0.02948635, 0.01239933, 0.06792817, 0.08599116, 0.09212975, 0.09871039, 
    0.01134358, 0.03305379, 0.05970234, 0.1790986, 0.1367156, 0.07865607, 
    0.07951884, 0.02753223, 0.01847403, 0.0226054, 0.06097312,
  0.1082174, 0.2737448, 0.1991122, 0.2284859, 0.4091099, 0.4332309, 
    0.3505346, 0.2941485, 0.1474647, 0.08590186, 0.07484142, 0.07086755, 
    0.209057, 0.2029838, 0.2443377, 0.2660426, 0.3082881, 0.3879696, 
    0.3799009, 0.3731348, 0.2449835, 0.3123291, 0.2535588, 0.4269422, 
    0.345449, 0.2695646, 0.1140919, 0.08123728, 0.07542748,
  0.3843673, 0.3414748, 0.4517972, 0.4699566, 0.3753988, 0.3251869, 
    0.3899913, 0.2949378, 0.3180582, 0.2630922, 0.4008064, 0.3230011, 
    0.2830374, 0.314926, 0.2820315, 0.29382, 0.2801078, 0.2993537, 0.3729208, 
    0.3838014, 0.4285014, 0.3024714, 0.270285, 0.3328418, 0.2964988, 
    0.2695709, 0.2521643, 0.2074177, 0.3411389,
  0.2105867, 0.1782358, 0.1730837, 0.203291, 0.2057859, 0.2056039, 0.1752818, 
    0.2217857, 0.1643525, 0.1858955, 0.1962725, 0.1669005, 0.1773539, 
    0.1056467, 0.1305673, 0.1753335, 0.1060002, 0.1027941, 0.1355159, 
    0.1749473, 0.1661825, 0.1432483, 0.1550174, 0.1457586, 0.07618069, 
    0.1479787, 0.1083462, 0.1667173, 0.1942988,
  0.08744366, 0.04159018, 0.02606639, 0.06218204, 0.06782982, 0.0608265, 
    0.1578957, 0.1594945, 0.05548157, 0.0291479, 0.02290969, 0.01901369, 
    0.05907042, 0.1680383, 0.08211965, 0.02568415, 0.0742895, 0.07466073, 
    0.06639785, 0.1340086, 0.1157835, 0.08934634, 0.0588077, 0.03775641, 
    0.04167167, 0.06577469, 0.1000297, 0.099985, 0.09868345,
  0.007440474, -3.112383e-08, 0.09991111, 0.03073412, 0.07100151, 0.08826253, 
    0.07101228, 0.004933831, 3.742499e-05, 0.0002292634, 0.001659793, 
    0.01368738, 0.07849213, 0.07038995, 0.04822981, 0.09594388, 0.05932553, 
    0.2360551, 0.209487, 0.02299855, 0.1530122, 0.004060379, -5.523103e-06, 
    0.002308911, 0.04472301, 0.1218948, 0.1666568, 0.07061411, 0.01443843,
  4.99508e-05, 0.08300485, 0.1442507, 0.01584758, 0.05955156, 0.04100966, 
    0.05908011, 0.03077427, 5.342757e-05, 7.476217e-08, 0.02446435, 
    0.02934457, 0.01374316, 0.007512236, 0.1300682, 0.03147001, 0.05735802, 
    0.04731863, 0.03129772, 0.04748788, 0.0004033518, 3.259088e-08, 
    2.829051e-08, 0.001835892, 0.1098149, 0.3041127, 0.01240162, 
    0.0003044561, 2.988519e-05,
  0.0002194867, 0.005697122, 0.1851938, 0.08846474, 0.1038341, 0.1475254, 
    0.07422569, 0.05637887, 0.01321751, 0.00395202, 0.008279132, 0.02668019, 
    0.02679051, 0.0247663, 0.03417808, 0.05660952, 0.04011589, 0.08330428, 
    0.01054023, 0.001194356, 6.036444e-07, -1.19852e-09, 5.027809e-05, 
    0.06419477, 0.1417686, 0.07944766, 0.005565959, -1.738454e-06, 0.001006133,
  0.06408967, 0.09192268, 0.1102918, 0.06283387, 0.04069723, 0.03113438, 
    0.03429689, 0.09670554, 0.09962226, 0.1494637, 0.03196122, 0.00836704, 
    0.009902476, 0.01932897, 0.02146614, 0.000371454, -3.893434e-05, 
    4.020091e-06, -5.665332e-07, 0.001768075, 0.0006870776, 0.006525662, 
    0.0831036, 0.1232378, 0.1393808, 0.04029889, 0.1256834, 0.05800679, 
    0.1052721,
  1.578957e-07, 0.000479793, 0.02201294, 0.03188179, 0.01512263, 0.02196985, 
    0.008844617, 0.009086759, 0.02355647, 0.05120897, 0.2241858, 0.09084541, 
    0.0604812, 0.04741433, 0.06428377, 0.08337763, 0.06948341, 0.1075663, 
    0.097784, 0.1201509, 0.1267652, 0.05047639, 0.07053501, 0.02159523, 
    0.04618233, 0.007328569, 0.003197133, 1.11309e-06, 5.569684e-08,
  2.088648e-07, 1.83267e-07, 2.627562e-08, 0.02092955, 0.04208797, 
    0.0001175976, 0.02036433, 0.05406651, 0.019145, 0.09225094, 0.1700411, 
    0.0314262, 0.01179154, 0.01477363, 0.01837283, 0.04737368, 0.03353094, 
    0.02864987, 0.08890222, 0.03488618, 0.008726454, 0.07195956, 0.01160161, 
    0.01857084, 0.03838566, 0.02999981, 0.02180339, 1.168162e-05, 1.37432e-06,
  1.122109e-06, 0.01211204, 0.01095706, 0.03028422, 0.05463756, 0.03759388, 
    0.02990456, 0.05589844, 0.1182234, 0.08112989, 0.04583121, 0.03222013, 
    0.09375932, 0.1142576, 0.1192042, 0.1465599, 0.06931111, 0.02224422, 
    0.06133564, 0.03024869, 0.05585499, 0.08695408, 0.06622466, 0.05931726, 
    0.05116323, 0.04491521, 0.0679009, 0.03124614, 0.001025228,
  0.02709093, 0.03701668, 0.1401587, 0.3210714, 0.1302509, 0.133661, 
    0.2259856, 0.03535, 0.02795083, 0.05514023, 0.02609393, 0.09157835, 
    0.1826314, 0.1300665, 0.1251978, 0.1786998, 0.1846738, 0.1086495, 
    0.09031053, 0.1758385, 0.119135, 0.01527385, 0.1204266, 0.1925126, 
    0.212837, 0.2116548, 0.1097235, 0.09536099, 0.0601249,
  0.1509931, 0.2615214, 0.2764787, 0.2797974, 0.2697738, 0.2906846, 
    0.2212451, 0.2054282, 0.08995371, 0.08197397, 0.1503659, 0.1330394, 
    0.235835, 0.3044632, 0.2736657, 0.2445616, 0.2866817, 0.2248809, 
    0.2298045, 0.2420993, 0.1777481, 0.1735207, 0.1976888, 0.2316369, 
    0.2160222, 0.2511196, 0.3616263, 0.1848094, 0.1527626,
  0.2388481, 0.3397505, 0.3459008, 0.3547651, 0.3335983, 0.3016067, 
    0.1615924, 0.1800966, 0.2345507, 0.3303204, 0.2900859, 0.1175534, 
    0.1632527, 0.1972359, 0.2050766, 0.2464897, 0.2614519, 0.4486471, 
    0.3379244, 0.2576278, 0.3215598, 0.2231486, 0.3294739, 0.3586429, 
    0.2273765, 0.2612304, 0.271589, 0.2603697, 0.3174483,
  0.2122021, 0.2421073, 0.2886331, 0.2698119, 0.2350913, 0.4358647, 
    0.3614033, 0.4473533, 0.2919912, 0.3324764, 0.3264072, 0.213564, 
    0.2042997, 0.3329846, 0.3821957, 0.1854441, 0.1641078, 0.2897585, 
    0.2200977, 0.1799179, 0.1863009, 0.1615563, 0.314021, 0.2904959, 
    0.1762543, 0.1696557, 0.272306, 0.2524713, 0.1785694,
  0.1818918, 0.229006, 0.3053963, 0.3413319, 0.2995857, 0.2082758, 0.243059, 
    0.2777717, 0.2968999, 0.3146513, 0.3370989, 0.3275495, 0.3439343, 
    0.2823449, 0.2503112, 0.242052, 0.1752612, 0.223342, 0.3009087, 
    0.3393147, 0.3043247, 0.3263856, 0.2553341, 0.06127012, 0.2051881, 
    0.1600729, 0.2002702, 0.2644047, 0.2354967,
  0.04373394, 0.04407591, 0.04441789, 0.04475986, 0.04510184, 0.04544381, 
    0.04578579, 0.03436336, 0.03302938, 0.0316954, 0.03036141, 0.02902743, 
    0.02769345, 0.02635946, 0.02572964, 0.02571855, 0.02570745, 0.02569636, 
    0.02568526, 0.02567416, 0.02566307, 0.02624969, 0.0272528, 0.0282559, 
    0.029259, 0.0302621, 0.03126521, 0.03226831, 0.04346035,
  0.0341759, 0.03787872, 0.006686267, 0.04597476, 0.1324162, 0.1198371, 
    0.1090954, 0.06497909, 0.1270989, 0.0757581, 0.05335721, 0.04791914, 
    0.03802142, 0.01093417, 0.04839002, 0.06164523, 0.055121, 0.0756312, 
    0.01219914, 0.01758301, 0.05149374, 0.1676967, 0.1424996, 0.1164067, 
    0.05941273, 0.06115376, 0.07315033, 0.02741776, 0.067473,
  0.07649701, 0.1698398, 0.1453969, 0.1813955, 0.4176545, 0.4445339, 
    0.3655692, 0.2660339, 0.1258995, 0.08293875, 0.07277357, 0.0796451, 
    0.2333193, 0.1172909, 0.2365859, 0.2686177, 0.3002087, 0.2931285, 
    0.2489236, 0.3542044, 0.2066582, 0.2261041, 0.3082688, 0.4222854, 
    0.3422476, 0.2649322, 0.1417258, 0.1287166, 0.08294918,
  0.3037953, 0.3362964, 0.3636731, 0.4384484, 0.3996338, 0.349304, 0.4162575, 
    0.2709791, 0.3741219, 0.3032601, 0.3923759, 0.3217348, 0.3182807, 
    0.3295946, 0.294882, 0.2930685, 0.2899547, 0.3403519, 0.3685433, 
    0.3851147, 0.3976034, 0.2832104, 0.282316, 0.2984982, 0.3058462, 
    0.2450278, 0.2553402, 0.2559789, 0.2790545,
  0.2213634, 0.1774854, 0.1981365, 0.181952, 0.1991713, 0.216064, 0.1740365, 
    0.226203, 0.2055178, 0.2049632, 0.2061914, 0.1641939, 0.1877568, 
    0.124318, 0.1572541, 0.1932959, 0.1641423, 0.1291806, 0.1588347, 
    0.1683289, 0.1857032, 0.1516735, 0.1563576, 0.1690338, 0.06958223, 
    0.1231272, 0.08997481, 0.1880403, 0.1873172,
  0.1048156, 0.0524806, 0.03768208, 0.06498263, 0.08097099, 0.07305794, 
    0.1732361, 0.1764927, 0.06050209, 0.04505745, 0.03003255, 0.02918986, 
    0.06103173, 0.1535181, 0.1080991, 0.02700563, 0.09462633, 0.09110992, 
    0.06454165, 0.1210581, 0.1096046, 0.08882938, 0.06114625, 0.03014711, 
    0.02851693, 0.07630458, 0.09851668, 0.09866458, 0.108618,
  0.008038818, -9.322017e-08, 0.07369561, 0.02922774, 0.07400223, 0.07028285, 
    0.07312967, 0.006855865, 0.001478684, 0.0001629091, 0.0009203054, 
    0.004420072, 0.06331626, 0.06683426, 0.05204529, 0.09292745, 0.06023335, 
    0.2415347, 0.1774911, 0.01762127, 0.1507598, 0.002559398, 6.092749e-05, 
    0.001295915, 0.0301874, 0.1401933, 0.1602646, 0.08022191, 0.02204625,
  2.5255e-05, 0.05503001, 0.1447259, 0.01790272, 0.0698397, 0.05294841, 
    0.05860344, 0.02885864, 0.001775736, 4.197412e-08, 0.01734187, 0.0130706, 
    0.01726864, 0.007789669, 0.1223853, 0.03945911, 0.06240968, 0.04548887, 
    0.03014305, 0.06997934, 0.01731332, 7.882632e-06, 8.947286e-09, 
    0.001986892, 0.09553759, 0.2609866, 0.02293121, 0.002789365, -2.423118e-05,
  1.589018e-05, 0.008049, 0.1712797, 0.07807095, 0.09082201, 0.1358251, 
    0.07133123, 0.05196306, 0.01427254, 0.003497358, 0.009692435, 0.02591651, 
    0.02701068, 0.02870323, 0.03101419, 0.05787282, 0.05041953, 0.08042909, 
    0.01272175, 0.004965929, 0.0008827836, 5.889656e-08, 3.599214e-05, 
    0.06105821, 0.116418, 0.06664399, 0.01231815, -1.444916e-05, 0.001393853,
  0.05096665, 0.08729602, 0.1042146, 0.06910789, 0.04787256, 0.02985805, 
    0.03420223, 0.08008742, 0.1434599, 0.152709, 0.03128658, 0.008456359, 
    0.01075107, 0.01713529, 0.02597439, 0.002044824, 2.275543e-05, 
    0.0002382421, 1.285959e-05, 0.001803445, 0.0005858876, 0.006370531, 
    0.07787433, 0.1084816, 0.145254, 0.03382937, 0.1285668, 0.07588255, 
    0.1018552,
  6.817935e-08, 3.3838e-05, 0.002578733, 0.08199063, 0.02122526, 0.02428648, 
    0.01324855, 0.01386811, 0.02766274, 0.06364608, 0.2188375, 0.09092081, 
    0.06553438, 0.05051181, 0.06392464, 0.08261012, 0.06733704, 0.1046479, 
    0.10445, 0.1093677, 0.112968, 0.05383397, 0.1001595, 0.02860072, 
    0.03929364, 0.01029538, 0.003316852, -4.170796e-06, 9.760778e-08,
  1.03076e-07, 7.6307e-08, 1.375013e-08, 0.03127539, 0.01495608, 0.001738119, 
    0.02370092, 0.06177088, 0.02316654, 0.1032148, 0.1744853, 0.03107748, 
    0.02683231, 0.02386979, 0.03768997, 0.0425434, 0.03640817, 0.03374758, 
    0.07881484, 0.03947932, 0.004276368, 0.1105377, 0.017788, 0.02987521, 
    0.04176553, 0.0336244, 0.01966481, 2.098353e-06, 7.999677e-07,
  5.873191e-07, 0.01288801, 0.01783487, 0.05005753, 0.0808633, 0.03721707, 
    0.02362707, 0.06561212, 0.1086765, 0.09654914, 0.04412996, 0.03966222, 
    0.116442, 0.1196055, 0.1309036, 0.1479081, 0.05258898, 0.03795174, 
    0.07098397, 0.02497956, 0.07084617, 0.09474861, 0.07325985, 0.07189405, 
    0.05886963, 0.05829212, 0.07514301, 0.04512346, -1.97577e-05,
  0.02842475, 0.04166617, 0.1351498, 0.348501, 0.1345368, 0.1405547, 
    0.2058922, 0.02599909, 0.01936306, 0.05457237, 0.02199344, 0.1190867, 
    0.2020164, 0.1468013, 0.1498372, 0.1705488, 0.2116759, 0.123868, 
    0.09822999, 0.1767202, 0.1141676, 0.00367632, 0.110911, 0.2009522, 
    0.2265774, 0.232437, 0.1119844, 0.09983789, 0.07826674,
  0.1606607, 0.2737602, 0.2785287, 0.2506298, 0.2370533, 0.2687449, 
    0.2245081, 0.2294183, 0.08256375, 0.07419612, 0.1351555, 0.1295656, 
    0.2807597, 0.3272891, 0.2641748, 0.2647072, 0.2882194, 0.2241682, 
    0.2369925, 0.2425333, 0.2010328, 0.1599869, 0.2084546, 0.191484, 
    0.2066322, 0.2808462, 0.3624012, 0.193012, 0.1638478,
  0.2319235, 0.2784552, 0.344632, 0.3053947, 0.2253238, 0.2808613, 0.1722997, 
    0.1724578, 0.2029801, 0.322486, 0.2992398, 0.1128922, 0.1846343, 
    0.2267608, 0.21311, 0.23995, 0.3039077, 0.4595106, 0.323434, 0.2256401, 
    0.2871894, 0.2191322, 0.3091972, 0.3286626, 0.2756776, 0.2776831, 
    0.2852211, 0.2699506, 0.3316027,
  0.2359735, 0.2355721, 0.2458172, 0.2701419, 0.2546706, 0.4252574, 
    0.3425875, 0.4716192, 0.3324938, 0.3594317, 0.3556469, 0.2138046, 
    0.1895096, 0.3100474, 0.3715638, 0.1743892, 0.1486848, 0.2462928, 
    0.1878708, 0.18806, 0.2205441, 0.1283473, 0.3220551, 0.2415232, 
    0.1671407, 0.1952722, 0.2892277, 0.2454504, 0.1777403,
  0.2776703, 0.2680989, 0.2856461, 0.3590858, 0.2929624, 0.2547771, 
    0.2761294, 0.3314583, 0.3477379, 0.3028431, 0.2965387, 0.305299, 
    0.3052238, 0.2909081, 0.23315, 0.2325732, 0.15821, 0.1996695, 0.2819123, 
    0.34799, 0.2941033, 0.2857482, 0.2547214, 0.06727158, 0.1977558, 
    0.1459933, 0.1900068, 0.252098, 0.2689827,
  0.05982209, 0.06071055, 0.06159902, 0.06248749, 0.06337596, 0.06426442, 
    0.06515289, 0.05561569, 0.05399634, 0.05237698, 0.05075762, 0.04913826, 
    0.04751891, 0.04589955, 0.03093547, 0.03028661, 0.02963774, 0.02898888, 
    0.02834001, 0.02769115, 0.02704229, 0.02585632, 0.02723607, 0.02861582, 
    0.02999558, 0.03137533, 0.03275509, 0.03413484, 0.05911132,
  0.03490298, 0.03459252, 0.005841703, 0.03746973, 0.1280962, 0.1174138, 
    0.11025, 0.08639516, 0.1366841, 0.09413046, 0.07410448, 0.05733232, 
    0.07420786, 0.0152525, 0.06834687, 0.09581799, 0.06541018, 0.06632616, 
    0.01242082, 0.007316295, 0.05824092, 0.1808896, 0.1959056, 0.222991, 
    0.1181815, 0.1182785, 0.07507711, 0.08627898, 0.07502332,
  0.09611301, 0.1156032, 0.1380213, 0.1395052, 0.4180613, 0.4675233, 
    0.3221276, 0.2849309, 0.1182485, 0.08566918, 0.08517404, 0.1037489, 
    0.215391, 0.07261652, 0.2545094, 0.265814, 0.2634886, 0.2488884, 
    0.114128, 0.2748244, 0.1450326, 0.1684076, 0.2078085, 0.3542646, 
    0.3060994, 0.190081, 0.3366863, 0.2239404, 0.08804273,
  0.2303168, 0.2950611, 0.4404598, 0.3198986, 0.3480813, 0.3276164, 0.338841, 
    0.277995, 0.3501528, 0.2785618, 0.3589554, 0.2988696, 0.2772779, 
    0.3449141, 0.2992512, 0.2917076, 0.2590776, 0.3076682, 0.3247501, 
    0.3208722, 0.3767435, 0.3318933, 0.3360853, 0.2516146, 0.2737713, 
    0.2344176, 0.2712241, 0.2762882, 0.2373762,
  0.2227741, 0.1842441, 0.2073002, 0.186617, 0.2107969, 0.2089369, 0.1980047, 
    0.2225514, 0.2149542, 0.2131471, 0.2411101, 0.1985787, 0.2067135, 
    0.1571736, 0.174262, 0.203574, 0.1562823, 0.1400445, 0.1828357, 
    0.1770622, 0.1956297, 0.1637079, 0.1974344, 0.1858699, 0.06478672, 
    0.1165839, 0.08837762, 0.2008921, 0.1938151,
  0.1054139, 0.06129548, 0.05683713, 0.08717366, 0.0982626, 0.08766926, 
    0.1768956, 0.1610182, 0.07048791, 0.05177342, 0.04216142, 0.04086595, 
    0.0696154, 0.1551239, 0.1323348, 0.04402399, 0.09101482, 0.103399, 
    0.08106128, 0.1353119, 0.1081759, 0.1092864, 0.08386665, 0.02876117, 
    0.02048774, 0.07509496, 0.09332781, 0.08660065, 0.1158372,
  0.01556408, 8.428881e-08, 0.06305574, 0.02501635, 0.1071935, 0.04857701, 
    0.0982969, 0.01935275, 0.007540718, 0.001021278, 0.0003168216, 
    0.0006773922, 0.0503037, 0.06455767, 0.05486302, 0.1069848, 0.0619177, 
    0.227646, 0.1720994, 0.02123191, 0.1382046, 0.0189649, 0.003301793, 
    0.0008926186, 0.01589329, 0.148671, 0.1591827, 0.09854707, 0.04619912,
  5.481861e-06, 0.0339181, 0.1325505, 0.01771242, 0.07605471, 0.05245781, 
    0.06432819, 0.0213619, 0.007141889, 2.829263e-08, 0.01489481, 0.01123144, 
    0.0195659, 0.008570007, 0.1182023, 0.03836137, 0.06303588, 0.03668191, 
    0.02883796, 0.05648921, 0.05653867, 0.003104558, 1.782748e-07, 
    0.001132444, 0.08596898, 0.2370481, 0.02607347, 0.02035806, 0.0001528369,
  3.542905e-06, 0.005785901, 0.1589604, 0.06660924, 0.07306737, 0.1330649, 
    0.06444407, 0.04845294, 0.02014276, 0.00569227, 0.0191788, 0.02272017, 
    0.02792001, 0.02774047, 0.0240438, 0.0592793, 0.04763501, 0.06922793, 
    0.02140356, 0.01037092, 0.006854172, 4.783369e-07, 9.993126e-06, 
    0.05838991, 0.08923966, 0.05195364, 0.01737462, 0.0002438601, 0.006893083,
  0.04373249, 0.1017816, 0.1185865, 0.08786385, 0.05194052, 0.02884172, 
    0.03088075, 0.06199045, 0.1626516, 0.1599416, 0.02868193, 0.00858915, 
    0.01160968, 0.0140881, 0.02701805, 0.007497832, 0.001453986, 0.004146713, 
    0.000670961, 0.0002954365, 0.0004441736, 0.01504176, 0.07897145, 
    0.09938753, 0.1179541, 0.03025286, 0.1261068, 0.08973511, 0.09112775,
  2.634512e-08, 1.536325e-06, -2.114284e-05, 0.09774888, 0.04046205, 
    0.03360889, 0.02960833, 0.01773272, 0.03617968, 0.06619924, 0.2061876, 
    0.07780642, 0.05552015, 0.04705731, 0.05947153, 0.08338846, 0.06485082, 
    0.09763069, 0.1181894, 0.1090116, 0.104839, 0.04939802, 0.1138825, 
    0.02779365, 0.03498723, 0.01623027, 0.004421226, -8.608247e-06, 
    5.978004e-08,
  3.745037e-08, 2.336242e-08, 4.267039e-09, 0.04330797, 0.003128562, 
    0.006413518, 0.03867799, 0.06693897, 0.02215669, 0.1073629, 0.1824514, 
    0.06115933, 0.03735018, 0.03132561, 0.03616457, 0.05328225, 0.04332728, 
    0.06329082, 0.06345998, 0.05499729, 0.001529525, 0.1309377, 0.03033532, 
    0.04387473, 0.03978933, 0.02637426, 0.0167471, -2.551942e-07, 5.802835e-07,
  5.52641e-07, 0.02045959, 0.02786004, 0.0506899, 0.09437673, 0.02922369, 
    0.01728194, 0.05945838, 0.09455932, 0.07226393, 0.07326858, 0.08462004, 
    0.1092087, 0.1258815, 0.1331993, 0.1640696, 0.0573579, 0.05446942, 
    0.07202953, 0.02317, 0.07251468, 0.1045131, 0.09116911, 0.06495612, 
    0.07400902, 0.07096536, 0.06665702, 0.06214578, -3.60485e-05,
  0.02854951, 0.05030369, 0.1395133, 0.3693795, 0.1347416, 0.1276403, 
    0.1941262, 0.02368213, 0.01561721, 0.06332847, 0.03335201, 0.1583461, 
    0.2205281, 0.2023444, 0.1984898, 0.1940902, 0.2397859, 0.1841095, 
    0.1395618, 0.1737752, 0.1053211, 0.0008311105, 0.1010361, 0.1974026, 
    0.2556588, 0.2401378, 0.1173725, 0.09097899, 0.07241577,
  0.1531831, 0.2609869, 0.2590238, 0.248507, 0.1715392, 0.2448538, 0.196055, 
    0.2429232, 0.09720846, 0.07178134, 0.1282338, 0.1303215, 0.3630089, 
    0.3426423, 0.2917983, 0.2888816, 0.2878213, 0.2158294, 0.2509214, 
    0.252467, 0.1787015, 0.1548017, 0.1874982, 0.2190858, 0.2403157, 
    0.2992367, 0.3647472, 0.2050447, 0.1699894,
  0.243566, 0.2829763, 0.2935765, 0.3793567, 0.2223341, 0.2694745, 0.1805859, 
    0.1516031, 0.2208924, 0.3470617, 0.3143898, 0.09453799, 0.2094774, 
    0.2380088, 0.2508895, 0.2632251, 0.2956338, 0.4814645, 0.3303701, 
    0.2033661, 0.2317116, 0.1819502, 0.2696016, 0.2967319, 0.3109588, 
    0.2645495, 0.2948496, 0.2901124, 0.340354,
  0.2124367, 0.2433092, 0.2673224, 0.287752, 0.1952809, 0.3867396, 0.3128695, 
    0.4893417, 0.3598304, 0.4026859, 0.3987049, 0.2176234, 0.1895572, 
    0.2999442, 0.4245208, 0.2093395, 0.1515033, 0.2403001, 0.1345235, 
    0.1722032, 0.1977087, 0.1478973, 0.3165177, 0.2111212, 0.1715444, 
    0.1916137, 0.2924268, 0.250267, 0.1986445,
  0.1870318, 0.2198311, 0.3284915, 0.3017207, 0.2169661, 0.1804586, 
    0.2367208, 0.3166785, 0.3164604, 0.3044666, 0.3162396, 0.3021207, 
    0.279029, 0.2935248, 0.2320567, 0.2157777, 0.1608575, 0.2010294, 
    0.2685458, 0.3674201, 0.3055716, 0.3311597, 0.2488162, 0.06372534, 
    0.1738937, 0.1274058, 0.1903661, 0.2266141, 0.3155366,
  0.06886089, 0.07022113, 0.07158138, 0.07294162, 0.07430187, 0.07566211, 
    0.07702236, 0.07005467, 0.06749191, 0.06492915, 0.0623664, 0.05980364, 
    0.05724088, 0.05467813, 0.03693035, 0.03631238, 0.03569441, 0.03507644, 
    0.03445846, 0.03384049, 0.03322252, 0.03091115, 0.03273163, 0.03455211, 
    0.03637259, 0.03819308, 0.04001356, 0.04183405, 0.06777269,
  0.05226711, 0.04197386, 0.004871788, 0.03570026, 0.1188755, 0.1205526, 
    0.1224912, 0.09658534, 0.1662362, 0.1384487, 0.09085359, 0.05739021, 
    0.1149419, 0.02534453, 0.1079403, 0.1691715, 0.119167, 0.05987019, 
    0.01442352, -0.0001507883, 0.136936, 0.2186644, 0.2567966, 0.2846477, 
    0.2415767, 0.1406559, 0.1528327, 0.0802315, 0.1058517,
  0.06995356, 0.1197401, 0.1836292, 0.1068244, 0.3918947, 0.4839183, 
    0.2661793, 0.3018301, 0.09384181, 0.08700721, 0.08904719, 0.1135731, 
    0.1907513, 0.1180739, 0.221559, 0.270911, 0.29586, 0.3051294, 0.1847992, 
    0.2836064, 0.2118447, 0.1688177, 0.2397365, 0.2839669, 0.3567984, 
    0.2542707, 0.1898924, 0.1747265, 0.08386689,
  0.246157, 0.3373723, 0.5065727, 0.3582387, 0.3189594, 0.31837, 0.3699131, 
    0.288828, 0.318063, 0.3054516, 0.3374195, 0.3140885, 0.3429767, 
    0.3751805, 0.3432594, 0.2992716, 0.2452345, 0.2980977, 0.3414099, 
    0.3617262, 0.4126059, 0.3856062, 0.3313135, 0.263558, 0.2777466, 
    0.2340704, 0.3071459, 0.3793578, 0.3158486,
  0.2668502, 0.2199695, 0.239655, 0.2333961, 0.2398449, 0.2357808, 0.2152352, 
    0.2462167, 0.2624475, 0.241723, 0.2785114, 0.2660465, 0.2681269, 
    0.198373, 0.1716327, 0.2232128, 0.1957364, 0.2197073, 0.2180853, 
    0.2102442, 0.1915189, 0.1856245, 0.2397209, 0.1947302, 0.0527438, 
    0.1214542, 0.1110995, 0.232672, 0.2466736,
  0.1280776, 0.08793521, 0.1088468, 0.1273015, 0.1209002, 0.1308785, 
    0.1968306, 0.1665261, 0.08806306, 0.07923702, 0.05598532, 0.06823853, 
    0.09235303, 0.2041496, 0.1707947, 0.04302991, 0.1138033, 0.1359368, 
    0.1091432, 0.1569609, 0.1622735, 0.1542746, 0.116291, 0.03109105, 
    0.01429006, 0.08460338, 0.1311496, 0.09095934, 0.126724,
  0.02141272, 4.090789e-05, 0.05598509, 0.03509303, 0.1110304, 0.04911739, 
    0.1280834, 0.04050404, 0.02662635, 0.005091453, 9.692253e-05, 
    6.825455e-05, 0.04390283, 0.06665652, 0.06166011, 0.131294, 0.06641973, 
    0.2607745, 0.1748988, 0.02443239, 0.1582016, 0.06464288, 0.0209389, 
    0.0004455308, 0.009167918, 0.16126, 0.1444999, 0.1080323, 0.05578969,
  3.871624e-07, 0.0180206, 0.1114072, 0.01704002, 0.08387508, 0.05180575, 
    0.06256703, 0.02369452, 0.03105625, 1.672034e-08, 0.01177029, 0.01095114, 
    0.01968374, 0.00904925, 0.1119257, 0.03147817, 0.05840269, 0.03004367, 
    0.02644536, 0.06298015, 0.1046859, 0.04589025, 4.134683e-06, 
    0.0007983854, 0.0914864, 0.2183874, 0.03011443, 0.06967551, 0.01359242,
  1.782426e-05, 0.002637596, 0.1496329, 0.05640159, 0.05159453, 0.1103868, 
    0.05825979, 0.049609, 0.02943696, 0.008849671, 0.02874514, 0.0214724, 
    0.02709053, 0.02417941, 0.02035052, 0.05717421, 0.04197387, 0.05984623, 
    0.02352542, 0.0129257, 0.009912772, 0.0002594332, 3.654967e-06, 
    0.05421351, 0.07146785, 0.04332867, 0.03504117, 0.007219498, 0.004962938,
  0.02979114, 0.1206291, 0.1286513, 0.09119371, 0.05001941, 0.03161043, 
    0.03036411, 0.04801503, 0.1717538, 0.1836853, 0.0285493, 0.01067155, 
    0.01313978, 0.01385575, 0.03057819, 0.01202363, 0.006501569, 0.007844164, 
    0.003495717, 0.001561165, 0.002040441, 0.02016741, 0.06307368, 
    0.08802924, 0.09185018, 0.03050325, 0.1122876, 0.07223545, 0.07373156,
  6.137491e-09, 1.119628e-07, -7.948846e-06, 0.06832297, 0.07550225, 
    0.04390536, 0.02401862, 0.02706503, 0.04908833, 0.06072854, 0.1903874, 
    0.0590506, 0.04685675, 0.04314257, 0.04984442, 0.08291948, 0.06060098, 
    0.08683254, 0.1205187, 0.106889, 0.1001394, 0.03875545, 0.1386591, 
    0.02860133, 0.03391851, 0.02787699, 0.01023033, -8.765213e-06, 
    1.647148e-08,
  1.745195e-08, 9.323977e-09, -1.551027e-09, 0.06738212, 0.0006036788, 
    0.02176539, 0.04392055, 0.06460018, 0.03622023, 0.1359442, 0.2193796, 
    0.06732401, 0.04729839, 0.04068721, 0.03474914, 0.05911607, 0.06453356, 
    0.08289313, 0.06462541, 0.09155534, 0.0007610366, 0.1703985, 0.03944962, 
    0.04135044, 0.03935364, 0.02701037, 0.02342488, -2.695919e-05, 
    3.384489e-07,
  7.49969e-07, 0.02868979, 0.07715606, 0.06362013, 0.09501165, 0.01339381, 
    0.01233426, 0.04106109, 0.08052552, 0.09771892, 0.1230046, 0.1408461, 
    0.1299824, 0.1710587, 0.1391626, 0.1701126, 0.06180516, 0.07461813, 
    0.116086, 0.0418394, 0.07160345, 0.1572703, 0.1042754, 0.1036211, 
    0.1020255, 0.1145111, 0.07734726, 0.0972762, -3.342829e-05,
  0.02812605, 0.06171845, 0.1343725, 0.3819718, 0.1504765, 0.1311073, 
    0.1806113, 0.01986552, 0.01358191, 0.0713829, 0.04216037, 0.1922158, 
    0.2604114, 0.2760609, 0.2463754, 0.2396641, 0.268722, 0.2093204, 
    0.225485, 0.186122, 0.09748367, 0.004727097, 0.1254543, 0.2098625, 
    0.3095855, 0.258177, 0.1329415, 0.09437802, 0.0784945,
  0.1747872, 0.2796032, 0.340131, 0.2845556, 0.1868138, 0.2586364, 0.181589, 
    0.2591181, 0.08650983, 0.07455494, 0.1459431, 0.1449816, 0.3885034, 
    0.3507388, 0.2952541, 0.2842486, 0.2706262, 0.2326936, 0.2687968, 
    0.3022765, 0.1413221, 0.149692, 0.1930371, 0.2683726, 0.2214884, 
    0.3158512, 0.3552724, 0.2122804, 0.2279569,
  0.2797137, 0.3078154, 0.3236229, 0.3617365, 0.3237996, 0.3089489, 
    0.2390162, 0.1674404, 0.2991553, 0.3524268, 0.3691338, 0.09623471, 
    0.2379084, 0.2545909, 0.3634627, 0.3210374, 0.3099673, 0.4982863, 
    0.3295847, 0.2157209, 0.2054336, 0.1652756, 0.2651708, 0.3152165, 
    0.4168064, 0.2402688, 0.3274701, 0.3061239, 0.3543175,
  0.2474869, 0.2893568, 0.1937191, 0.3437592, 0.2504039, 0.3556945, 
    0.3347101, 0.4685766, 0.3605981, 0.4519267, 0.4305314, 0.2096902, 
    0.2049502, 0.3206769, 0.4721447, 0.1950932, 0.1714839, 0.2511941, 
    0.1120501, 0.2005603, 0.206672, 0.2031664, 0.2961232, 0.1954881, 
    0.1647557, 0.1802781, 0.3015459, 0.3174872, 0.2266253,
  0.2138095, 0.1732007, 0.278414, 0.2320627, 0.2273256, 0.1821997, 0.2361556, 
    0.3184129, 0.3214697, 0.3095103, 0.3178458, 0.292852, 0.2912741, 
    0.3196455, 0.2327283, 0.2023854, 0.1704788, 0.217012, 0.2760557, 
    0.3793214, 0.2960125, 0.3673228, 0.2379613, 0.06352759, 0.1757463, 
    0.116384, 0.1943857, 0.2070502, 0.3045635,
  0.1022699, 0.1038334, 0.105397, 0.1069605, 0.108524, 0.1100875, 0.1116511, 
    0.1057704, 0.100603, 0.09543564, 0.09026825, 0.08510086, 0.07993347, 
    0.07476608, 0.08472119, 0.08671375, 0.0887063, 0.09069885, 0.09269141, 
    0.09468395, 0.09667651, 0.09490447, 0.09651579, 0.0981271, 0.09973842, 
    0.1013497, 0.102961, 0.1045724, 0.1010191,
  0.08949219, 0.05606827, 0.01133147, 0.07043464, 0.1382616, 0.1308978, 
    0.12035, 0.125387, 0.2814066, 0.2677275, 0.1946009, 0.07988255, 
    0.1260357, -0.006029502, 0.1899065, 0.1088956, 0.09922308, 0.05972811, 
    0.04158281, 0.02650859, 0.1596647, 0.2474904, 0.2889661, 0.1743004, 
    0.2328877, 0.1707146, 0.0856318, 0.1400423, 0.1478035,
  0.1343997, 0.1215709, 0.1630117, 0.07261359, 0.3562886, 0.4693286, 
    0.2484251, 0.2946099, 0.08669256, 0.1030834, 0.09637426, 0.1460208, 
    0.1677514, 0.1052205, 0.2711175, 0.3330881, 0.403219, 0.3545833, 
    0.2876696, 0.3813219, 0.2391532, 0.2077316, 0.2217024, 0.3061299, 
    0.3895468, 0.438874, 0.2237659, 0.1592232, 0.101719,
  0.3590917, 0.4103061, 0.5562276, 0.3772637, 0.3826848, 0.4467855, 
    0.4157865, 0.3639678, 0.38592, 0.3771825, 0.4035505, 0.3851316, 0.402794, 
    0.4292526, 0.3546603, 0.3457288, 0.3233424, 0.3423849, 0.3830459, 
    0.407567, 0.4786576, 0.4680917, 0.4283347, 0.3466629, 0.375334, 
    0.3362344, 0.3445784, 0.406565, 0.4831981,
  0.2984175, 0.2538691, 0.2738046, 0.2958838, 0.2958545, 0.2878788, 
    0.2864344, 0.3223675, 0.3011781, 0.2849253, 0.3557208, 0.3191792, 
    0.3147287, 0.2482016, 0.1679077, 0.2531192, 0.2283391, 0.2609372, 
    0.2812206, 0.3075121, 0.2608148, 0.237647, 0.2504613, 0.1955951, 
    0.04714772, 0.122987, 0.162202, 0.3047408, 0.3088531,
  0.2092876, 0.1568264, 0.1553969, 0.167304, 0.1720534, 0.1641144, 0.2681121, 
    0.2874011, 0.1773695, 0.1543119, 0.0895612, 0.09019427, 0.1187411, 
    0.2244213, 0.1814064, 0.1007153, 0.1613452, 0.203373, 0.1926835, 
    0.2087195, 0.2385108, 0.2078882, 0.1659548, 0.03239296, 0.008870999, 
    0.1236399, 0.1693919, 0.152152, 0.1677853,
  0.06716922, 0.01918198, 0.05724051, 0.0456155, 0.1256723, 0.06878192, 
    0.163756, 0.08833326, 0.07491283, 0.02025641, 0.0001894061, 3.997019e-06, 
    0.02407996, 0.07787123, 0.07389968, 0.1552475, 0.07114451, 0.2698354, 
    0.1782345, 0.04158606, 0.1539313, 0.1391188, 0.1231871, 0.0001655438, 
    0.009785384, 0.1823396, 0.1513797, 0.1148133, 0.07854156,
  0.003906294, 0.007926505, 0.08791135, 0.01742625, 0.1069411, 0.04805134, 
    0.07104868, 0.06053765, 0.06848168, -1.021132e-08, 0.004978826, 
    0.009028864, 0.02458786, 0.01310347, 0.1085629, 0.03525016, 0.05082832, 
    0.02619975, 0.03004087, 0.0575774, 0.1088512, 0.1767614, 0.002770019, 
    0.0007012505, 0.08876447, 0.2032978, 0.03970704, 0.08102693, 0.1182081,
  0.00253753, 0.005363438, 0.1444393, 0.04580766, 0.04017982, 0.09775677, 
    0.0508959, 0.05099609, 0.04033577, 0.01844081, 0.02553356, 0.02815302, 
    0.02735405, 0.02388667, 0.02288649, 0.05285512, 0.05150539, 0.05691904, 
    0.02660399, 0.0308537, 0.05051249, 0.01520072, 0.0002824544, 0.05185016, 
    0.05858291, 0.03526736, 0.05400721, 0.03713586, 0.0168062,
  0.03358138, 0.08672514, 0.1111746, 0.09298994, 0.04966635, 0.03067121, 
    0.0334367, 0.03867412, 0.1784178, 0.2082287, 0.03285951, 0.01526656, 
    0.01613794, 0.01765562, 0.03488565, 0.01365076, 0.01015963, 0.009410566, 
    0.0120628, 0.007267088, 0.02837988, 0.01237846, 0.05897298, 0.07072409, 
    0.07818228, 0.03202462, 0.09297226, 0.05247862, 0.07573174,
  1.429091e-09, 1.968689e-08, -3.572369e-07, 0.02402349, 0.1108746, 
    0.03991952, 0.01671579, 0.04820957, 0.09345699, 0.06641503, 0.1750847, 
    0.05004717, 0.03790532, 0.04255486, 0.04457524, 0.07796267, 0.05712937, 
    0.08505395, 0.1127144, 0.09538892, 0.08890516, 0.03941489, 0.1512332, 
    0.02947674, 0.03943747, 0.03552606, 0.02457902, -1.265094e-05, 
    1.729294e-09,
  6.941082e-09, 1.378859e-09, -4.118335e-07, 0.09621997, 0.005260998, 
    0.1199247, 0.02855596, 0.0881726, 0.06673104, 0.3045905, 0.3473787, 
    0.1116474, 0.04350444, 0.07123014, 0.03666025, 0.06812909, 0.1140793, 
    0.09324938, 0.1090473, 0.124258, 0.001848521, 0.2382306, 0.08308054, 
    0.04622941, 0.04087928, 0.03560385, 0.04141337, -0.0003896463, 
    9.200026e-08,
  -5.130307e-07, 0.08138448, 0.10472, 0.08325557, 0.09858643, 0.00305516, 
    0.01092788, 0.02775, 0.06732874, 0.140465, 0.2557758, 0.1865541, 
    0.1539029, 0.1691964, 0.1962633, 0.1909017, 0.110865, 0.1237565, 
    0.2164169, 0.07000574, 0.08258811, 0.2254737, 0.1283246, 0.2724133, 
    0.1610506, 0.2033516, 0.1625181, 0.1415465, -0.0001102835,
  0.02867808, 0.05867701, 0.1549446, 0.4047578, 0.1298327, 0.1541252, 
    0.1575153, 0.01185145, 0.01049336, 0.06949174, 0.06583781, 0.246447, 
    0.308082, 0.3101524, 0.2633673, 0.244958, 0.302267, 0.2310397, 0.2460805, 
    0.2135167, 0.09884019, 0.003060247, 0.1729262, 0.2334059, 0.3097612, 
    0.2418605, 0.1269319, 0.107025, 0.129026,
  0.2050377, 0.3163437, 0.4208856, 0.2851327, 0.2721737, 0.27909, 0.2062493, 
    0.2787462, 0.06482219, 0.08437583, 0.1478818, 0.16365, 0.4024834, 
    0.3348446, 0.2259574, 0.2735112, 0.2536326, 0.2271949, 0.2482195, 
    0.3524451, 0.1364847, 0.1484833, 0.270327, 0.3184766, 0.2731019, 
    0.3123654, 0.3182501, 0.2048994, 0.2414995,
  0.3247637, 0.3044427, 0.3884697, 0.4442898, 0.4088355, 0.3894, 0.3054438, 
    0.2571673, 0.299012, 0.3941918, 0.4579429, 0.1239403, 0.2582146, 
    0.2464072, 0.546374, 0.3539153, 0.3263361, 0.5092377, 0.3667062, 
    0.2376297, 0.2164149, 0.1528421, 0.307031, 0.3345305, 0.600328, 
    0.1989865, 0.3371225, 0.3049196, 0.3707675,
  0.3217043, 0.3300163, 0.196043, 0.3440754, 0.4295298, 0.395132, 0.4473876, 
    0.4556453, 0.3852174, 0.5111424, 0.4299013, 0.2097245, 0.2487956, 
    0.3487692, 0.4918922, 0.1716677, 0.2086426, 0.2511116, 0.1262958, 
    0.2456486, 0.1903667, 0.2422397, 0.3009128, 0.1679876, 0.128668, 
    0.1769919, 0.3045538, 0.3256537, 0.3033587,
  0.2199932, 0.1424439, 0.225676, 0.2298299, 0.2174531, 0.1790204, 0.2164425, 
    0.2813968, 0.2751963, 0.3015937, 0.3042964, 0.2977166, 0.3143456, 
    0.3637653, 0.2506545, 0.2159391, 0.1884149, 0.2407315, 0.3087448, 
    0.3817878, 0.3371037, 0.4136776, 0.2731148, 0.06870703, 0.1707079, 
    0.09478541, 0.2018815, 0.2015494, 0.2884554,
  0.1907186, 0.1937128, 0.1967069, 0.1997011, 0.2026952, 0.2056894, 
    0.2086836, 0.1798706, 0.1718809, 0.1638913, 0.1559017, 0.147912, 
    0.1399224, 0.1319328, 0.1708668, 0.1756445, 0.1804223, 0.1852001, 
    0.1899778, 0.1947556, 0.1995334, 0.1685241, 0.1687418, 0.1689595, 
    0.1691772, 0.1693949, 0.1696126, 0.1698303, 0.1883233,
  0.1125208, 0.07677264, 0.05669436, 0.114416, 0.1847829, 0.1419904, 
    0.1341105, 0.153255, 0.3176842, 0.2740352, 0.2154037, 0.1180738, 
    0.1665134, -0.02264009, 0.1813539, 0.1023893, 0.08953895, 0.05316275, 
    0.09407537, 0.09875597, 0.2734913, 0.2645603, 0.2812727, 0.1673338, 
    0.239706, 0.2193329, 0.1461346, 0.1555828, 0.1254679,
  0.1563843, 0.1916258, 0.122964, 0.05196664, 0.3034921, 0.4579657, 
    0.2143493, 0.2734995, 0.1129242, 0.1209171, 0.1271839, 0.249619, 
    0.122213, 0.129577, 0.2841092, 0.4519945, 0.3812654, 0.3966946, 
    0.3584945, 0.4263472, 0.2465331, 0.2154675, 0.2674464, 0.3150054, 
    0.3588232, 0.478851, 0.3627476, 0.2815069, 0.1294134,
  0.3881263, 0.4275925, 0.6042716, 0.4811969, 0.4933734, 0.4823361, 
    0.4532616, 0.4145314, 0.4182327, 0.3745279, 0.4828523, 0.4136285, 
    0.4594303, 0.4559749, 0.3419255, 0.358913, 0.3825759, 0.3957157, 
    0.4536228, 0.4298479, 0.4927446, 0.4309394, 0.4300148, 0.4228103, 
    0.4993181, 0.4118621, 0.4302538, 0.4119236, 0.4787363,
  0.3964947, 0.3474047, 0.3442301, 0.3316765, 0.3894503, 0.4122261, 0.340692, 
    0.3676062, 0.3201075, 0.3567964, 0.3777212, 0.3190241, 0.3524555, 
    0.2865539, 0.1849459, 0.2317591, 0.2615038, 0.2733768, 0.2916646, 
    0.3278187, 0.3389199, 0.2924545, 0.3141693, 0.1949847, 0.04754227, 
    0.130645, 0.2126129, 0.3864577, 0.358275,
  0.3266493, 0.2441409, 0.2017085, 0.1878582, 0.2613494, 0.1982298, 
    0.3369584, 0.3137175, 0.261538, 0.3373996, 0.1466747, 0.1062465, 
    0.1377935, 0.2823813, 0.2024012, 0.2110266, 0.2489671, 0.2684786, 
    0.3413761, 0.288338, 0.2904162, 0.1962779, 0.2121117, 0.04770418, 
    0.03568812, 0.1667568, 0.2026668, 0.1992717, 0.2179817,
  0.2180479, 0.06184667, 0.04391488, 0.1184542, 0.1764854, 0.1352324, 
    0.1794938, 0.2142904, 0.1953847, 0.07608329, 0.0001121214, 0.001131706, 
    0.00782972, 0.09760663, 0.1320172, 0.1608815, 0.1176836, 0.2702964, 
    0.1825673, 0.1065132, 0.1618823, 0.1619676, 0.2546403, 0.0001237515, 
    0.01090466, 0.2315543, 0.1640663, 0.1740254, 0.2227554,
  0.1263556, 0.008643235, 0.06120611, 0.02718103, 0.1228894, 0.06387512, 
    0.07666732, 0.09080236, 0.1707047, -0.0002250993, 0.002312053, 
    0.004935933, 0.0380096, 0.02811172, 0.10983, 0.063176, 0.07586943, 
    0.02865674, 0.04029263, 0.0580006, 0.09260292, 0.308382, 0.138494, 
    0.0007399457, 0.0692446, 0.1894812, 0.04967628, 0.108425, 0.2008771,
  0.03351199, 0.01127459, 0.1139569, 0.0435656, 0.04453293, 0.09450477, 
    0.05317928, 0.05609766, 0.05011467, 0.03596581, 0.03338479, 0.04805038, 
    0.04147759, 0.0319389, 0.04929175, 0.08320768, 0.04698045, 0.06863831, 
    0.04272266, 0.08629107, 0.09636422, 0.1509177, 0.0069436, 0.03285658, 
    0.04747418, 0.02361217, 0.07476065, 0.095718, 0.05409367,
  0.02809419, 0.04363488, 0.06568665, 0.09108951, 0.04936299, 0.03656816, 
    0.04057418, 0.03776148, 0.1993556, 0.2308554, 0.03753429, 0.02390627, 
    0.02497434, 0.04343391, 0.06217932, 0.04463729, 0.01280107, 0.01093168, 
    0.01099521, 0.01568194, 0.05940659, 0.01837733, 0.0605289, 0.0490278, 
    0.06121435, 0.04170823, 0.08337275, 0.04150195, 0.05395972,
  4.477753e-10, 6.326935e-09, 3.146231e-07, 0.009644927, 0.1309402, 
    0.0987459, 0.004451738, 0.1359244, 0.1823848, 0.08518395, 0.1516396, 
    0.05077543, 0.04821297, 0.05523172, 0.06657898, 0.09427596, 0.06320512, 
    0.08226701, 0.110171, 0.08989823, 0.08412652, 0.05432299, 0.1894264, 
    0.04223218, 0.0546882, 0.0503388, 0.1745935, -0.0004254938, 6.83089e-10,
  1.602568e-09, -1.030597e-05, 7.658835e-05, 0.06506838, 0.004893575, 
    0.1993216, 0.03059294, 0.1410471, 0.03942081, 0.3844402, 0.3597265, 
    0.1530498, 0.06554167, 0.07215837, 0.08059356, 0.1010907, 0.1186061, 
    0.1039615, 0.1772575, 0.1820464, 0.009471771, 0.2498806, 0.1162418, 
    0.05430057, 0.05125758, 0.0441949, 0.09874631, 0.005625774, 2.041427e-08,
  -1.50023e-06, 0.17095, 0.08336189, 0.1376788, 0.09663734, -4.831921e-05, 
    0.006429414, 0.01966454, 0.04549155, 0.1248352, 0.3501013, 0.1074318, 
    0.1382218, 0.1499694, 0.1847055, 0.2046378, 0.1257899, 0.1721993, 
    0.1870051, 0.06436378, 0.1018137, 0.2388774, 0.1513555, 0.259375, 
    0.128935, 0.1663783, 0.1334185, 0.1791047, -0.0001104622,
  0.02537002, 0.09406783, 0.1713138, 0.418975, 0.1177412, 0.1565667, 
    0.1431689, 0.007264753, 0.00736149, 0.08768771, 0.1047833, 0.2243605, 
    0.3056591, 0.2051301, 0.1900255, 0.2094807, 0.3153726, 0.2739615, 
    0.2480707, 0.2768004, 0.1043803, 0.001259746, 0.2145981, 0.2787234, 
    0.2263138, 0.1881579, 0.1111536, 0.1622351, 0.2046297,
  0.2075869, 0.3862319, 0.4372393, 0.3867474, 0.3187567, 0.2961435, 
    0.2172084, 0.3086459, 0.05894036, 0.1116168, 0.1609101, 0.1839929, 
    0.2830817, 0.2717077, 0.1584074, 0.2776145, 0.2576499, 0.2232564, 
    0.2500562, 0.3839018, 0.1449208, 0.1908831, 0.3307205, 0.3921799, 
    0.2784846, 0.2750436, 0.2813783, 0.1975757, 0.2426176,
  0.3090215, 0.2731338, 0.4333636, 0.4513248, 0.4722103, 0.4270453, 
    0.2908859, 0.3067693, 0.3472064, 0.4593835, 0.5163124, 0.1721499, 
    0.2662708, 0.2290583, 0.5971703, 0.3481204, 0.3392087, 0.5107108, 
    0.4444638, 0.2636068, 0.232684, 0.1944766, 0.3233875, 0.3716314, 
    0.4906512, 0.1708975, 0.2859695, 0.3044805, 0.3677712,
  0.3150297, 0.2425535, 0.1676071, 0.2775102, 0.482181, 0.4354731, 0.407069, 
    0.4493653, 0.4297398, 0.5463206, 0.421476, 0.2221672, 0.2918149, 
    0.3574184, 0.5371805, 0.2049223, 0.237319, 0.2695669, 0.1540196, 
    0.2952518, 0.2357804, 0.2509001, 0.3327254, 0.1942476, 0.09138025, 
    0.1834026, 0.3132063, 0.2795519, 0.4399779,
  0.2325686, 0.1737638, 0.23089, 0.2155821, 0.1961242, 0.1353823, 0.2273127, 
    0.2853627, 0.2365313, 0.3043785, 0.3527959, 0.325491, 0.3407149, 
    0.4075687, 0.2698771, 0.2460271, 0.2091206, 0.2857158, 0.3496596, 
    0.4052076, 0.3509648, 0.4350588, 0.2708608, 0.07110754, 0.1583666, 
    0.0800585, 0.1876258, 0.193657, 0.3242571,
  0.2481331, 0.2487615, 0.2493898, 0.2500181, 0.2506465, 0.2512749, 
    0.2519032, 0.3013948, 0.2972936, 0.2931925, 0.2890914, 0.2849903, 
    0.2808892, 0.276788, 0.2765387, 0.2796103, 0.282682, 0.2857536, 
    0.2888253, 0.2918969, 0.2949686, 0.2883337, 0.2887348, 0.2891359, 
    0.289537, 0.2899382, 0.2903393, 0.2907404, 0.2476304,
  0.1134536, 0.1115486, 0.1018203, 0.1252254, 0.2142633, 0.1579452, 
    0.1402985, 0.1857208, 0.3897045, 0.2931544, 0.2294725, 0.249533, 
    0.2127569, -0.01952144, 0.1510114, 0.1601721, 0.1191654, 0.07277025, 
    0.1042932, 0.136532, 0.3934182, 0.3318761, 0.3069722, 0.1294486, 
    0.202544, 0.2075187, 0.1164594, 0.1541787, 0.1591219,
  0.1314711, 0.248922, 0.2402466, 0.06392389, 0.1795245, 0.4725145, 
    0.1664255, 0.1943125, 0.109792, 0.09259234, 0.1639783, 0.2824364, 
    0.1076406, 0.1246506, 0.2655824, 0.4365579, 0.386705, 0.3247626, 
    0.3289339, 0.4228823, 0.2786046, 0.2167637, 0.2648969, 0.2804518, 
    0.3571146, 0.3672396, 0.3523568, 0.3232802, 0.1702173,
  0.4255013, 0.4280103, 0.5849158, 0.4853776, 0.5899796, 0.503409, 0.5136046, 
    0.4459442, 0.4814217, 0.4404179, 0.4760877, 0.4240862, 0.4525614, 
    0.4579715, 0.3433393, 0.3805133, 0.4628997, 0.4721117, 0.4993855, 
    0.41969, 0.4812991, 0.3986189, 0.3907139, 0.4313802, 0.501837, 0.4858237, 
    0.5470374, 0.4027856, 0.4279575,
  0.4373251, 0.4084418, 0.3909135, 0.4063576, 0.4265054, 0.4121214, 
    0.4124689, 0.3951191, 0.3625507, 0.4311847, 0.3628369, 0.2796425, 
    0.2834426, 0.215147, 0.1770969, 0.242017, 0.3138863, 0.3227478, 0.307856, 
    0.3163813, 0.3328394, 0.287482, 0.3213773, 0.197308, 0.03668492, 
    0.1513405, 0.2426268, 0.4532455, 0.3565985,
  0.3198743, 0.2573373, 0.1592109, 0.1745487, 0.2091871, 0.2041246, 
    0.2866944, 0.3084052, 0.3591406, 0.3098442, 0.2704746, 0.08831441, 
    0.1491915, 0.2903308, 0.1776264, 0.2930666, 0.2933619, 0.3673244, 
    0.3420515, 0.2388662, 0.2537726, 0.2071018, 0.1757835, 0.05529882, 
    0.0113802, 0.1373535, 0.2728905, 0.275134, 0.2292127,
  0.3382896, 0.05268391, 0.03747553, 0.1274412, 0.1682557, 0.1653736, 
    0.245135, 0.3120902, 0.3570876, 0.02855258, 0.000168501, 4.052556e-05, 
    0.00305435, 0.1178924, 0.09252604, 0.1823304, 0.1491869, 0.2902447, 
    0.1921041, 0.1082346, 0.1859659, 0.1298459, 0.2638013, 0.0001201154, 
    0.01400771, 0.2821742, 0.1911144, 0.1633291, 0.3297152,
  0.4494172, 0.01352792, 0.04919837, 0.06265149, 0.1169428, 0.08187896, 
    0.09277781, 0.09150964, 0.2248356, 0.003543097, 0.000537152, 0.001491687, 
    0.06344543, 0.1204999, 0.1171388, 0.06659028, 0.08318172, 0.04882442, 
    0.0490443, 0.07069588, 0.038962, 0.2476026, 0.6270872, 0.002820698, 
    0.0444098, 0.1719687, 0.08620547, 0.1446469, 0.3091135,
  0.1174921, 0.03171993, 0.08183338, 0.0443971, 0.07422075, 0.0950555, 
    0.06770409, 0.07376684, 0.09442266, 0.1098963, 0.0307452, 0.04805807, 
    0.07753142, 0.08273415, 0.09530178, 0.07775941, 0.03682798, 0.04758552, 
    0.06774063, 0.08181623, 0.1110022, 0.270637, 0.1925225, 0.01532214, 
    0.03255389, 0.01182943, 0.1152693, 0.124783, 0.1518822,
  0.0183776, 0.01772363, 0.03794529, 0.1027692, 0.07065737, 0.05500273, 
    0.05672695, 0.06386869, 0.2173299, 0.2009696, 0.04693903, 0.1221268, 
    0.1237766, 0.1715193, 0.0859035, 0.09334479, 0.03008638, 0.02205998, 
    0.01436797, 0.07303263, 0.07109465, 0.09714417, 0.07068, 0.02634068, 
    0.04482833, 0.06179297, 0.07161997, 0.03633646, 0.03459102,
  2.175133e-10, 2.830904e-09, -6.209059e-08, -1.258301e-05, 0.1963864, 
    0.1079495, -9.951254e-05, 0.05767962, 0.2035433, 0.09463919, 0.1487564, 
    0.04788577, 0.03842775, 0.05184585, 0.07136878, 0.08495958, 0.06955114, 
    0.089421, 0.1032155, 0.09162324, 0.07789991, 0.08503472, 0.2909839, 
    0.05648157, 0.04183979, 0.02748365, 0.08869242, 0.0002046001, 5.49897e-10,
  3.743663e-10, -1.714109e-05, 0.001678971, 0.02269929, 9.197278e-05, 
    0.04009575, 0.011713, 0.06020866, 0.03319909, 0.3561037, 0.2420234, 
    0.1193906, 0.04061441, 0.04956803, 0.05594671, 0.07816684, 0.06433595, 
    0.06713725, 0.1126065, 0.1976677, 0.06361149, 0.2368667, 0.114102, 
    0.04827602, 0.03031453, 0.03044385, 0.06674445, 0.001443911, 2.623405e-09,
  -2.234778e-05, 0.1351512, 0.1064294, 0.1338564, 0.09477731, -0.0005479809, 
    0.00237222, 0.01223049, 0.03207094, 0.1024741, 0.2178703, 0.07248942, 
    0.1022565, 0.1186474, 0.1528966, 0.1895353, 0.1207213, 0.1787867, 
    0.1468688, 0.2276465, 0.1272125, 0.2642795, 0.1554367, 0.1391593, 
    0.07937946, 0.1005578, 0.08201316, 0.1183931, -0.0001579503,
  0.03461478, 0.1378641, 0.2064184, 0.4250731, 0.06804871, 0.153978, 
    0.1367888, 0.003793468, 0.006700563, 0.1113762, 0.1608463, 0.1515199, 
    0.2037001, 0.1240984, 0.1720004, 0.2177015, 0.3060721, 0.3092665, 
    0.2050395, 0.3271418, 0.1045778, 0.002316917, 0.2199395, 0.2536658, 
    0.1572655, 0.1561467, 0.09983744, 0.1594843, 0.179334,
  0.2587293, 0.4654427, 0.4858966, 0.5044174, 0.3862135, 0.3422588, 
    0.2393726, 0.3023543, 0.05224163, 0.1456579, 0.1635815, 0.218788, 
    0.1455691, 0.1818446, 0.126126, 0.2682586, 0.2690083, 0.2867374, 
    0.2868668, 0.4121109, 0.1446454, 0.2176837, 0.3507029, 0.4495072, 
    0.2693214, 0.2065476, 0.2511462, 0.2162598, 0.3145106,
  0.3100343, 0.2622691, 0.4827771, 0.4700591, 0.5056245, 0.4703466, 
    0.2843115, 0.3058855, 0.4089232, 0.5477802, 0.541981, 0.2202149, 
    0.248565, 0.2068976, 0.5225198, 0.3759326, 0.3577002, 0.5050268, 
    0.4277996, 0.2619909, 0.3030713, 0.2372589, 0.3331318, 0.3862703, 
    0.3003216, 0.09946997, 0.2541865, 0.3061443, 0.3736468,
  0.2706251, 0.1675602, 0.1688424, 0.2235443, 0.4249683, 0.4994788, 
    0.3618862, 0.4360506, 0.436941, 0.5823084, 0.4331875, 0.2497035, 
    0.2776512, 0.4087978, 0.5523405, 0.2281036, 0.2711372, 0.2948934, 
    0.1981111, 0.2972038, 0.2584933, 0.302142, 0.322965, 0.1694743, 
    0.1074132, 0.1971977, 0.3291435, 0.2159022, 0.3743927,
  0.2968457, 0.1592963, 0.1303291, 0.1877926, 0.1369709, 0.1315467, 
    0.2565995, 0.3258966, 0.2728227, 0.3182504, 0.3511278, 0.3440473, 
    0.3872162, 0.4185764, 0.2863661, 0.2830766, 0.2466328, 0.3256166, 
    0.3806581, 0.4269575, 0.3855862, 0.4157773, 0.2791097, 0.0844228, 
    0.1674107, 0.06856687, 0.1791516, 0.2115667, 0.3040419,
  0.2357024, 0.2390266, 0.2423509, 0.2456751, 0.2489993, 0.2523236, 
    0.2556478, 0.2446175, 0.2453152, 0.2460128, 0.2467105, 0.2474081, 
    0.2481057, 0.2488034, 0.2996006, 0.3001851, 0.3007696, 0.3013541, 
    0.3019386, 0.3025231, 0.3031076, 0.2802583, 0.2756519, 0.2710455, 
    0.2664391, 0.2618327, 0.2572263, 0.25262, 0.233043,
  0.1648434, 0.1219504, 0.1029129, 0.123241, 0.2271243, 0.1541512, 0.1572371, 
    0.2067099, 0.3773784, 0.2417344, 0.1990076, 0.273287, 0.2674027, 
    -0.01265156, 0.3006364, 0.2352304, 0.1819521, 0.1087417, 0.07530495, 
    0.1020968, 0.2644539, 0.3045588, 0.3219256, 0.1321141, 0.1308941, 
    0.1969776, 0.1963174, 0.1531812, 0.1016439,
  0.1559519, 0.1666054, 0.1801426, 0.06966891, 0.08076013, 0.4643625, 
    0.139333, 0.1135791, 0.05601573, 0.04730263, 0.1126385, 0.2550423, 
    0.08378287, 0.08227442, 0.2567946, 0.3273629, 0.351964, 0.3119285, 
    0.4328023, 0.4721138, 0.2598677, 0.2646244, 0.2469606, 0.29934, 
    0.3703509, 0.2909791, 0.2895049, 0.2088766, 0.2797695,
  0.406399, 0.4159562, 0.5261307, 0.5379565, 0.5599956, 0.5231296, 0.585991, 
    0.4997454, 0.578661, 0.4789854, 0.484392, 0.3110209, 0.4301361, 
    0.4321508, 0.3136038, 0.3571105, 0.5089779, 0.5509917, 0.4979536, 
    0.3767671, 0.4500972, 0.4162134, 0.3794062, 0.4605983, 0.4492032, 
    0.480757, 0.5728377, 0.35786, 0.4188572,
  0.3894868, 0.3711455, 0.4182866, 0.3740016, 0.383837, 0.3737936, 0.3810329, 
    0.3981941, 0.4127502, 0.4385018, 0.3149661, 0.2428462, 0.2075006, 
    0.1497375, 0.1632075, 0.2863742, 0.3390736, 0.3736913, 0.3209526, 
    0.2672472, 0.3048124, 0.3110057, 0.3358534, 0.1854006, 0.02671058, 
    0.1466685, 0.3174371, 0.447487, 0.3554301,
  0.3377001, 0.2358799, 0.0980961, 0.1895802, 0.1361213, 0.1205944, 
    0.2428552, 0.2626485, 0.4508412, 0.2978485, 0.2779958, 0.04941294, 
    0.164488, 0.2373331, 0.172261, 0.2335424, 0.2450036, 0.3255221, 
    0.3209133, 0.2173425, 0.214129, 0.2219651, 0.1125875, 0.06721703, 
    0.004565633, 0.1164691, 0.1840878, 0.2541234, 0.2781021,
  0.2565965, 0.07694409, 0.02823665, 0.1491413, 0.2310163, 0.1567554, 
    0.2073198, 0.2083022, 0.1892706, 0.04198748, 0.0008044097, -2.074831e-05, 
    -0.0008049574, 0.08415952, 0.07975673, 0.152205, 0.05377272, 0.2717721, 
    0.1948503, 0.1497413, 0.2015874, 0.08821576, 0.2305804, 0.004338091, 
    0.01568815, 0.1971824, 0.2188099, 0.1029131, 0.1687501,
  0.4065779, 0.008760318, 0.03833631, 0.1719539, 0.04712165, 0.06805824, 
    0.05034836, 0.02147028, 0.07139588, 0.06857923, 0.0002128114, 
    0.0004418188, 0.06034313, 0.04211146, 0.08625613, 0.05608095, 0.06137145, 
    0.04013327, 0.02362991, 0.01937227, 0.004874205, 0.09141936, 0.3459889, 
    0.06307068, 0.03258351, 0.164708, 0.04016909, 0.0947151, 0.1609042,
  0.4109699, 0.106504, 0.06130775, 0.07041544, 0.05476732, 0.08782018, 
    0.05333603, 0.03518511, 0.07718635, 0.2115258, 0.03328251, 0.03215122, 
    0.03248189, 0.02779212, 0.0253878, 0.02482881, 0.01479255, 0.01591399, 
    0.0134963, 0.0152219, 0.02598668, 0.09814574, 0.565995, 0.005672439, 
    0.02070124, 0.004160581, 0.04261119, 0.06397073, 0.2151328,
  0.01995557, 0.008785341, 0.02386075, 0.1115152, 0.0554483, 0.1249204, 
    0.1155473, 0.04820148, 0.1394754, 0.1547954, 0.02477879, 0.0400026, 
    0.02656113, 0.02918741, 0.04091183, 0.03109671, 0.01853674, 0.0279489, 
    0.05934047, 0.04554246, 0.1698066, 0.2522876, 0.1100519, 0.01113719, 
    0.02389733, 0.03749778, 0.05997556, 0.0406961, 0.04665439,
  1.291307e-10, 1.598094e-09, -5.298024e-08, -0.001702662, 0.1790202, 
    0.03800024, -0.002447263, 0.01025549, 0.06384332, 0.06920807, 0.1308806, 
    0.02170961, 0.01481331, 0.02603088, 0.03278466, 0.06984974, 0.03838221, 
    0.05734456, 0.08645, 0.1288576, 0.06741417, 0.03825857, 0.4266933, 
    0.1319448, 0.0093699, 0.009200238, 0.02222612, 4.604428e-07, 4.980196e-10,
  4.189953e-10, -5.31985e-05, 0.0009855928, 0.00477819, 7.926932e-06, 
    0.009673417, 0.003909725, 0.03890788, 0.02566879, 0.2954403, 0.1479825, 
    0.05684428, 0.01127252, 0.01514891, 0.02690968, 0.03074705, 0.03472873, 
    0.0339674, 0.05093558, 0.2193043, 0.1136478, 0.2077082, 0.03793662, 
    0.0117849, 0.006840012, 0.01207658, 0.01234503, 0.0006541398, 6.056051e-10,
  -1.966184e-05, 0.06904916, 0.03993452, 0.0793374, 0.1108086, -0.0001065206, 
    0.00124922, 0.007703488, 0.02339466, 0.1113569, 0.1360585, 0.05084498, 
    0.08098508, 0.09464215, 0.1091246, 0.178256, 0.1373326, 0.1147628, 
    0.09659562, 0.1251832, 0.1341783, 0.2495904, 0.132675, 0.1033804, 
    0.06843369, 0.03883656, 0.03565659, 0.05304679, 0.00056782,
  0.04909518, 0.126832, 0.1674084, 0.4351631, 0.04198352, 0.1508991, 
    0.1318208, 0.00117945, 0.009036101, 0.09599962, 0.1740772, 0.1013483, 
    0.1580062, 0.09293979, 0.1278224, 0.1578027, 0.2939756, 0.2408898, 
    0.1340548, 0.3639005, 0.1051227, 0.009007729, 0.1974253, 0.1998122, 
    0.1133492, 0.1367458, 0.08013484, 0.09203001, 0.1362087,
  0.4209184, 0.5037538, 0.4943725, 0.5110463, 0.4349407, 0.3791303, 
    0.2690226, 0.2715505, 0.04066915, 0.1644748, 0.1656922, 0.2537572, 
    0.1015147, 0.1197643, 0.08984464, 0.2422045, 0.2705431, 0.3004163, 
    0.2583064, 0.470822, 0.1698154, 0.2224655, 0.311207, 0.4858243, 
    0.2584118, 0.1637169, 0.2252248, 0.2609727, 0.3765063,
  0.3234305, 0.2837479, 0.5279827, 0.5642357, 0.5849841, 0.5111297, 
    0.2712662, 0.3331305, 0.4507697, 0.6095651, 0.598104, 0.2999081, 
    0.2275201, 0.1744385, 0.4223468, 0.3576399, 0.4157156, 0.4650209, 
    0.3806514, 0.2537139, 0.4448967, 0.2925743, 0.3294191, 0.3828634, 
    0.1887872, 0.07219618, 0.2243483, 0.2752658, 0.3572179,
  0.1903446, 0.11534, 0.1965817, 0.1387794, 0.2912325, 0.4825369, 0.3707538, 
    0.4645779, 0.4662157, 0.563244, 0.4676673, 0.2893655, 0.2960496, 
    0.4723757, 0.5736545, 0.2617324, 0.2999143, 0.3103002, 0.2170164, 
    0.2911415, 0.2455486, 0.303546, 0.3448008, 0.189277, 0.1247102, 
    0.2108462, 0.3298088, 0.1796183, 0.365763,
  0.3077671, 0.1783935, 0.1205114, 0.1603961, 0.1223473, 0.1722191, 0.289811, 
    0.3326885, 0.324582, 0.3194, 0.3983615, 0.3993734, 0.4354773, 0.4571131, 
    0.3457136, 0.3307915, 0.3162585, 0.3530212, 0.4193451, 0.4604628, 
    0.4468934, 0.4094989, 0.267834, 0.1270015, 0.1603161, 0.06270023, 
    0.167216, 0.2141689, 0.3119896,
  0.1903012, 0.1965569, 0.2028125, 0.2090682, 0.2153239, 0.2215795, 
    0.2278352, 0.2152054, 0.213451, 0.2116967, 0.2099424, 0.2081881, 
    0.2064338, 0.2046794, 0.2641436, 0.2624334, 0.2607231, 0.2590128, 
    0.2573026, 0.2555923, 0.2538821, 0.2088978, 0.2061067, 0.2033156, 
    0.2005246, 0.1977335, 0.1949424, 0.1921513, 0.1852966,
  0.1320664, 0.0900026, 0.07794213, 0.09837383, 0.2040183, 0.1118662, 
    0.1670179, 0.2636123, 0.2761762, 0.1674013, 0.1267473, 0.1855603, 
    0.2006753, -0.004582988, 0.2648108, 0.221719, 0.1820576, 0.145103, 
    0.03983897, 0.06502005, 0.1383861, 0.2146715, 0.2265415, 0.1170027, 
    0.05933221, 0.1263973, 0.1545605, 0.130785, 0.07510684,
  0.1444859, 0.1405237, 0.1591387, 0.06815469, 0.02865046, 0.3955939, 
    0.1367085, 0.07300501, 0.02297674, 0.02058499, 0.0697649, 0.1840939, 
    0.05270705, 0.102651, 0.2438895, 0.3134431, 0.3344204, 0.2938473, 
    0.4208861, 0.5003445, 0.2707315, 0.2989939, 0.2174167, 0.2998548, 
    0.4069708, 0.2992607, 0.2021713, 0.1306587, 0.3131533,
  0.3563053, 0.4094126, 0.4949823, 0.5031103, 0.5564598, 0.505654, 0.5870373, 
    0.5046088, 0.6238772, 0.4900934, 0.4249386, 0.2404831, 0.4291714, 
    0.3865235, 0.3238971, 0.3789445, 0.4994461, 0.5598795, 0.4982394, 
    0.3435138, 0.4311578, 0.3938048, 0.36468, 0.4082732, 0.3859471, 
    0.4400792, 0.4950811, 0.3253442, 0.4067885,
  0.4094135, 0.3675027, 0.4050218, 0.3427086, 0.3554105, 0.3636856, 
    0.3506764, 0.3382053, 0.4263396, 0.3883933, 0.2716442, 0.2037319, 
    0.1719125, 0.1133757, 0.1995665, 0.3082902, 0.3100548, 0.3538624, 
    0.2815748, 0.2464364, 0.2587911, 0.2985668, 0.3475394, 0.1619271, 
    0.0212389, 0.1505242, 0.3499899, 0.4372562, 0.3741655,
  0.3080156, 0.1669973, 0.06772593, 0.1664673, 0.1245206, 0.07429502, 
    0.2334362, 0.3090254, 0.3130972, 0.2903478, 0.1502402, 0.05863096, 
    0.1357429, 0.2244855, 0.180599, 0.1759396, 0.1710572, 0.19989, 0.2853529, 
    0.1918773, 0.2121236, 0.2154863, 0.08859407, 0.07955826, 0.007689935, 
    0.1100068, 0.1664507, 0.1764554, 0.2618177,
  0.1498173, 0.05126091, 0.02051807, 0.1338011, 0.185906, 0.06279419, 
    0.2054246, 0.08626503, 0.06856448, 0.01169937, 0.003089317, 
    -4.259509e-05, -0.001622661, 0.05365376, 0.03555783, 0.12165, 0.01751418, 
    0.2437671, 0.199242, 0.1387831, 0.0840111, 0.03309689, 0.1021675, 
    0.04146747, 0.01693379, 0.1529805, 0.1971204, 0.0618476, 0.1164466,
  0.1415965, 0.03646755, 0.03003123, 0.08602184, 0.01497972, 0.02537095, 
    0.01491473, 0.005607277, 0.02462062, 0.01942531, 0.000116887, 
    -6.03656e-05, 0.01220366, 0.004723257, 0.05577042, 0.02853931, 
    0.03687218, 0.01504825, 0.002723395, 0.003057972, 0.0005341308, 
    0.02897947, 0.1355964, 0.214386, 0.02313684, 0.1645255, 0.005951341, 
    0.02663094, 0.04291974,
  0.1535214, 0.1140783, 0.05129695, 0.09158, 0.01247528, 0.05263254, 
    0.01820133, 0.01295722, 0.01913767, 0.04179822, 0.01324949, 0.007244034, 
    0.01000017, 0.004260183, 0.004087606, 0.01299825, 0.005412147, 
    0.004603987, 0.001831961, 0.002721575, 0.005254121, 0.02558363, 
    0.2247777, 0.00179692, 0.01445564, 0.00117424, 0.002480781, 0.01086034, 
    0.07772487,
  0.01255313, 0.006885449, 0.01632641, 0.1008459, 0.03985341, 0.03127766, 
    0.02262023, 0.01607191, 0.08744103, 0.1166656, 0.006155486, 0.006670073, 
    0.003572546, 0.006178392, 0.009757323, 0.005092692, 0.004583355, 
    0.01676149, 0.01936869, 0.02153865, 0.07955852, 0.282477, 0.3552932, 
    0.006260211, 0.0108726, 0.01221649, 0.04891676, 0.02537134, 0.02223189,
  1.00971e-10, 1.236189e-09, 1.254769e-09, -0.001431172, 0.118596, 
    0.01451071, -0.003485313, 0.002525402, 0.01615048, 0.0230136, 0.07677023, 
    0.005892654, 0.005729231, 0.01021303, 0.0116503, 0.04482474, 0.02265297, 
    0.03463304, 0.04684721, 0.1115834, 0.037943, 0.009812432, 0.4474281, 
    0.125789, 0.0006538617, 0.0006310605, 0.006090642, -5.548205e-07, 
    4.802505e-10,
  6.64497e-10, -7.821928e-05, 0.00022818, 0.0007901537, 2.035417e-06, 
    0.004199077, 0.01348932, 0.02618158, 0.01974713, 0.1870752, 0.1000409, 
    0.02013231, 0.001161574, 0.003148002, 0.01010094, 0.01505961, 0.01553583, 
    0.016522, 0.03223829, 0.1473803, 0.05426696, 0.1479975, 0.007615954, 
    -0.002538116, 0.0003074181, 0.004048958, 0.002877278, 0.000123316, 
    7.385009e-10,
  -5.96038e-06, 0.03772084, 0.02055301, 0.03869886, 0.1068813, -8.645804e-05, 
    0.001190907, 0.006659572, 0.01728393, 0.09876718, 0.09831192, 0.02770307, 
    0.06296511, 0.06900971, 0.08860253, 0.1954659, 0.1056313, 0.05997172, 
    0.04920437, 0.06691046, 0.1378245, 0.2221742, 0.1208789, 0.08900593, 
    0.04187047, 0.02096353, 0.01701009, 0.0183771, 0.002529805,
  0.03389379, 0.07410868, 0.1043644, 0.4253387, 0.02964535, 0.1466383, 
    0.1315699, -0.0004507907, 0.003905378, 0.07914133, 0.1595572, 0.07589408, 
    0.1186343, 0.06888387, 0.1087586, 0.1235451, 0.2806861, 0.1813609, 
    0.09261184, 0.3777911, 0.08630447, 0.01175991, 0.1804195, 0.168682, 
    0.08580936, 0.1046639, 0.07068592, 0.05691228, 0.1245433,
  0.4668487, 0.4923871, 0.5463312, 0.4940201, 0.429111, 0.3900013, 0.2136657, 
    0.2355088, 0.04134766, 0.1711631, 0.1806963, 0.2692814, 0.07281779, 
    0.0831432, 0.0667342, 0.2178602, 0.2724214, 0.2585639, 0.1959124, 
    0.500052, 0.1446706, 0.2008479, 0.2758764, 0.5271576, 0.2163951, 
    0.1359759, 0.1929038, 0.2450827, 0.3786159,
  0.2829481, 0.2965336, 0.5213385, 0.6109088, 0.6221293, 0.5735077, 0.334315, 
    0.3773642, 0.5020351, 0.6605061, 0.6191524, 0.4145475, 0.2151828, 
    0.1578109, 0.3498576, 0.3530774, 0.4570613, 0.4129936, 0.3583366, 
    0.2682284, 0.56033, 0.3271059, 0.366419, 0.3552275, 0.1247905, 
    0.04686426, 0.1938579, 0.235509, 0.2894918,
  0.1186053, 0.08141823, 0.2235049, 0.08161423, 0.1819405, 0.4659405, 
    0.4206369, 0.468733, 0.4959527, 0.5468978, 0.5179468, 0.3237544, 
    0.3179217, 0.5208973, 0.5913343, 0.3084962, 0.3476793, 0.3186279, 
    0.2392547, 0.3086245, 0.2664546, 0.3172017, 0.3949581, 0.2201203, 
    0.1397363, 0.2253011, 0.3378604, 0.1705697, 0.2807625,
  0.4030319, 0.3247904, 0.1453629, 0.1435747, 0.1705275, 0.2264897, 
    0.3134388, 0.3191935, 0.3474837, 0.3853073, 0.4645678, 0.4466444, 
    0.4962237, 0.4999811, 0.3972284, 0.385056, 0.3607944, 0.3691777, 
    0.4870635, 0.4872243, 0.5184139, 0.4007506, 0.290815, 0.1654666, 
    0.1468018, 0.06107107, 0.1595194, 0.2091016, 0.3980175,
  0.2090821, 0.2139375, 0.218793, 0.2236484, 0.2285038, 0.2333593, 0.2382147, 
    0.2179647, 0.216782, 0.2155992, 0.2144165, 0.2132337, 0.212051, 
    0.2108682, 0.2587067, 0.254143, 0.2495793, 0.2450156, 0.2404519, 
    0.2358882, 0.2313244, 0.1935677, 0.1944587, 0.1953497, 0.1962408, 
    0.1971318, 0.1980228, 0.1989138, 0.2051977,
  0.09585206, 0.06167449, 0.04555555, 0.07078583, 0.1500295, 0.07776929, 
    0.1474255, 0.2253804, 0.1971819, 0.09847434, 0.0765809, 0.08698364, 
    0.1045569, -0.001112507, 0.1520436, 0.2056284, 0.2069074, 0.1124609, 
    0.02782727, 0.04208105, 0.07927141, 0.13425, 0.1605057, 0.08526153, 
    0.02392342, 0.05949777, 0.1023121, 0.07990179, 0.07181192,
  0.1803779, 0.1047407, 0.127685, 0.06321162, 0.01024345, 0.3292333, 
    0.128256, 0.0432619, 0.01206429, 0.009207364, 0.04171303, 0.1201949, 
    0.03180987, 0.1145459, 0.2259716, 0.2790599, 0.3008286, 0.2896452, 
    0.3445945, 0.483408, 0.2589578, 0.3117469, 0.2281171, 0.2298008, 
    0.3844062, 0.3475287, 0.1411257, 0.1029426, 0.2255813,
  0.2990599, 0.385847, 0.4370481, 0.4033361, 0.50581, 0.4907935, 0.5722699, 
    0.4159671, 0.6051789, 0.471091, 0.3718185, 0.2081555, 0.3960995, 
    0.3491316, 0.3029755, 0.3888727, 0.477088, 0.5384392, 0.4772811, 
    0.2848112, 0.3863865, 0.3535004, 0.3313226, 0.3356918, 0.348791, 
    0.4115535, 0.4227993, 0.2707032, 0.3474117,
  0.3782046, 0.3237096, 0.3658938, 0.2981907, 0.3363045, 0.3279309, 
    0.3311664, 0.299326, 0.4104592, 0.3264856, 0.2350403, 0.1639945, 
    0.1262441, 0.09716024, 0.2160845, 0.3254489, 0.2854612, 0.3068025, 
    0.2453396, 0.2275966, 0.2214283, 0.2472239, 0.303104, 0.1294321, 
    0.01875131, 0.1643531, 0.3425035, 0.4102414, 0.3896089,
  0.2522383, 0.1289453, 0.04955751, 0.1306427, 0.103679, 0.05407769, 
    0.2234727, 0.2573098, 0.1859615, 0.1605576, 0.06694544, 0.05352028, 
    0.1178625, 0.21584, 0.1817886, 0.1328934, 0.1008371, 0.1337676, 
    0.2417573, 0.1746703, 0.199054, 0.1915259, 0.07981707, 0.09011615, 
    0.01433977, 0.07685474, 0.1513447, 0.1453113, 0.2336916,
  0.08067978, 0.02306624, 0.01711907, 0.0691789, 0.1200976, 0.03169224, 
    0.1392292, 0.05169421, 0.0320644, 0.005327191, 0.003426533, 
    -1.955301e-06, -0.0008633499, 0.03365882, 0.02158465, 0.07388131, 
    0.005898164, 0.2103061, 0.204593, 0.100381, 0.03976782, 0.0134171, 
    0.03939096, 0.04734097, 0.01057114, 0.1230486, 0.1577816, 0.03671937, 
    0.07840361,
  0.05162588, 0.04494081, 0.01813493, 0.02389415, 0.004036176, 0.004853729, 
    0.005499008, 0.002299024, 0.0108358, 0.00844488, 5.264609e-05, 
    -0.0001546944, 0.002941353, 0.001200701, 0.02548172, 0.00728246, 
    0.009671347, 0.001671362, 0.0001257506, 0.0006548645, 0.0002035275, 
    0.01119335, 0.05268998, 0.1001933, 0.01718432, 0.1586882, 0.001439983, 
    0.00967752, 0.01365457,
  0.05300855, 0.03027048, 0.04583924, 0.08724241, 0.003796842, 0.02566838, 
    0.006659964, 0.005856014, 0.003463301, 0.009770731, 0.006072818, 
    0.002412734, 0.001692425, 0.0004324895, 0.001122165, 0.006489135, 
    0.002451526, 0.00203189, 0.000732158, 0.001217524, 0.002200742, 
    0.008923302, 0.08497386, 0.000562163, 0.01669842, 0.0002772278, 
    -0.0001753136, 0.003119042, 0.02147185,
  0.00194585, 0.006220055, 0.0170639, 0.092767, 0.005972906, 0.005510802, 
    0.002746762, 0.00245564, 0.05937471, 0.0922789, 0.0006359273, 
    0.002620238, 0.0008694908, 0.00246859, 0.005324512, 0.001584827, 
    0.0003046777, 0.001983804, 0.003481918, 0.003621442, 0.01880707, 
    0.1128719, 0.1322352, 0.006234325, 0.005927943, 0.005456628, 0.0328706, 
    0.006756959, 0.004225254,
  9.189651e-11, 1.143152e-09, 7.828148e-09, 0.007224286, 0.05628905, 
    0.003211391, -0.003619448, 0.001154026, 0.006592467, 0.005255654, 
    0.03550898, 0.001339084, 0.00209415, 0.001493839, 0.003230386, 
    0.02263064, 0.01342442, 0.0128128, 0.01398664, 0.03405039, 0.01902715, 
    0.001214353, 0.3748036, 0.09422476, 7.303851e-05, 2.040714e-05, 
    0.002794274, -3.115175e-07, 4.688535e-10,
  7.896935e-10, -6.265638e-05, 8.296193e-05, 0.0001961336, 1.029739e-06, 
    0.002426598, 0.02561593, 0.01171101, 0.01691188, 0.1013694, 0.05532619, 
    0.003761334, 0.0002459328, 0.0008736569, 0.001929363, 0.006633524, 
    0.01011236, 0.008387705, 0.02456329, 0.1055097, 0.0203152, 0.1127217, 
    0.00263907, -0.003084338, 6.938061e-05, 0.0006444256, 0.001349194, 
    5.389434e-05, 9.351423e-10,
  -1.49433e-06, 0.02866599, 0.0123299, 0.02405198, 0.0958932, -0.0001551627, 
    0.0006949875, 0.008150911, 0.01886349, 0.07445014, 0.07958737, 
    0.01613833, 0.04404871, 0.04740669, 0.09654504, 0.174535, 0.05521344, 
    0.02580903, 0.02568632, 0.03428579, 0.130203, 0.216042, 0.1086963, 
    0.07455536, 0.02094334, 0.01040416, 0.008170487, 0.008594679, 0.002818948,
  0.02149134, 0.03265591, 0.06098941, 0.4056603, 0.01682598, 0.107098, 
    0.1320574, -0.0007348417, 0.002652344, 0.05633151, 0.1500133, 0.06094096, 
    0.08939587, 0.05238418, 0.09636007, 0.09737276, 0.2503115, 0.1435611, 
    0.06306513, 0.362299, 0.07170358, 0.009563308, 0.1716369, 0.1508787, 
    0.06696935, 0.06855338, 0.04634141, 0.02972561, 0.0795678,
  0.4099824, 0.470645, 0.5029877, 0.4497997, 0.3986843, 0.3861403, 0.1445505, 
    0.193042, 0.04775376, 0.1530464, 0.1765294, 0.2909183, 0.04710052, 
    0.06321957, 0.05040576, 0.1902578, 0.2569465, 0.2108231, 0.1423837, 
    0.5095259, 0.1079913, 0.1691542, 0.2377444, 0.5607316, 0.1538691, 
    0.1132859, 0.1526286, 0.2002286, 0.3214834,
  0.2256773, 0.305198, 0.4836008, 0.6575007, 0.6846742, 0.5916176, 0.4520655, 
    0.4048085, 0.5495583, 0.6585657, 0.6272128, 0.4949407, 0.222502, 
    0.1722566, 0.2897134, 0.3591655, 0.5006548, 0.3613667, 0.3659748, 
    0.2685604, 0.6291867, 0.3951563, 0.3650512, 0.3291257, 0.08042882, 
    0.03585571, 0.1624296, 0.183263, 0.2101547,
  0.08304726, 0.06021231, 0.2395733, 0.04356528, 0.1210473, 0.4503981, 
    0.4533544, 0.5017774, 0.4532369, 0.5514369, 0.5749816, 0.4054948, 
    0.3753639, 0.6373606, 0.6059282, 0.3685859, 0.3721385, 0.3222696, 
    0.2868666, 0.2840458, 0.3580351, 0.3677397, 0.4813559, 0.2470737, 
    0.2590857, 0.2028446, 0.3338538, 0.133571, 0.2197638,
  0.4537773, 0.3444995, 0.1791432, 0.1869328, 0.2183654, 0.2681484, 
    0.3380666, 0.388248, 0.4017891, 0.4723528, 0.5364762, 0.532111, 
    0.6002731, 0.5594719, 0.5289934, 0.5517714, 0.4498632, 0.4825875, 
    0.5714704, 0.5389305, 0.5799705, 0.3780885, 0.3465115, 0.2680779, 
    0.1255253, 0.07498697, 0.126315, 0.1783788, 0.4589868,
  0.1642161, 0.1686779, 0.1731397, 0.1776015, 0.1820634, 0.1865252, 0.190987, 
    0.1623627, 0.1627142, 0.1630657, 0.1634172, 0.1637687, 0.1641202, 
    0.1644717, 0.218619, 0.2127485, 0.2068779, 0.2010074, 0.1951368, 
    0.1892662, 0.1833957, 0.1492897, 0.150347, 0.1514042, 0.1524615, 
    0.1535187, 0.154576, 0.1556332, 0.1606466,
  0.06492731, 0.03827018, 0.02688468, 0.05722777, 0.1062443, 0.05397099, 
    0.1210872, 0.163138, 0.130038, 0.0613963, 0.04394806, 0.04048589, 
    0.04176216, 0.0005468159, 0.09604938, 0.1786542, 0.2086231, 0.08404554, 
    0.02070507, 0.04120919, 0.04199581, 0.09049868, 0.1032026, 0.05753045, 
    0.01514287, 0.03761579, 0.07598186, 0.05633309, 0.04725083,
  0.1791029, 0.074373, 0.08827729, 0.0628745, 0.004812399, 0.2615159, 
    0.1200179, 0.02398988, 0.008234579, 0.003709233, 0.0275887, 0.07826835, 
    0.01806504, 0.09958175, 0.227079, 0.2251385, 0.278032, 0.2487542, 
    0.288781, 0.4190741, 0.2438186, 0.2989539, 0.2153075, 0.1635474, 
    0.3341343, 0.3387835, 0.1055078, 0.07884175, 0.1545708,
  0.2447205, 0.3172745, 0.3327086, 0.3283063, 0.4186716, 0.4220924, 
    0.5140024, 0.3280781, 0.5211112, 0.4029836, 0.2856138, 0.1751001, 
    0.3331009, 0.3061601, 0.2540138, 0.3512084, 0.4240106, 0.4874631, 
    0.4012326, 0.2339996, 0.342185, 0.269083, 0.2607769, 0.2534159, 
    0.3126865, 0.3783009, 0.3534557, 0.2103323, 0.2688632,
  0.3044979, 0.2568625, 0.2858907, 0.2300495, 0.2792455, 0.2760365, 
    0.2756243, 0.2579858, 0.37045, 0.2640546, 0.1779139, 0.1129833, 
    0.08738786, 0.06368944, 0.1970356, 0.2878915, 0.252221, 0.2222212, 
    0.1896486, 0.1871573, 0.1636434, 0.1851273, 0.209797, 0.1009836, 
    0.01784547, 0.1378721, 0.2812498, 0.350944, 0.3230821,
  0.2089854, 0.1028231, 0.03777815, 0.1008058, 0.08213571, 0.03978652, 
    0.1911561, 0.1866862, 0.1220103, 0.09120525, 0.04893592, 0.03804788, 
    0.08858157, 0.1877083, 0.1558742, 0.1017411, 0.07146835, 0.103169, 
    0.2036461, 0.1609892, 0.1658648, 0.1383279, 0.05625163, 0.09356361, 
    0.01060909, 0.0553381, 0.1116052, 0.1107172, 0.1940157,
  0.05345103, 0.01321814, 0.01108329, 0.035094, 0.06671689, 0.0181354, 
    0.09624067, 0.0377023, 0.01925654, 0.00314105, 0.001778862, 2.065599e-05, 
    9.681798e-05, 0.01096299, 0.02009019, 0.03931336, 0.00269605, 0.1822609, 
    0.1802849, 0.06411749, 0.01855449, 0.005992041, 0.019781, 0.02610234, 
    0.00634676, 0.08243249, 0.1272433, 0.02261534, 0.05241719,
  0.02494507, 0.05119039, 0.01122877, 0.01123201, -0.0001293736, 
    0.0009883982, 0.002168351, 0.001315075, 0.006141258, 0.004702847, 
    1.448441e-05, -8.989229e-05, 0.001230723, 0.0006157676, 0.00818449, 
    0.002843594, 0.002760017, 0.0002497355, 2.049877e-05, 0.000196491, 
    0.0001095066, 0.00573609, 0.02542149, 0.05168032, 0.01460111, 0.1351169, 
    0.0007754313, 0.005187618, 0.00645904,
  0.02663174, 0.01297475, 0.04774478, 0.07186574, 0.001362563, 0.01160186, 
    0.002494958, 0.002399307, 0.001458275, 0.004875012, 0.00312334, 
    0.001411672, 0.0003341569, 0.0001150108, 0.0006837968, 0.002109526, 
    0.0009510643, 0.0008129624, 0.0004193601, 0.0007028335, 0.001265189, 
    0.004529226, 0.04507372, 0.0003098717, 0.02186305, -1.909682e-05, 
    0.0002151589, 0.001557347, 0.008933919,
  0.001116688, 0.003358401, 0.02285338, 0.07831162, 0.001409616, 0.002050075, 
    0.0005781017, 0.001113369, 0.04513285, 0.07459076, 0.0001923858, 
    0.001509327, 0.0004228411, 0.00135709, 0.002891453, 0.0008081527, 
    0.0001076709, 0.0005941499, 0.001488323, 0.001499469, 0.007517784, 
    0.03359724, 0.058654, 0.007003799, 0.004127893, 0.001922785, 0.01499779, 
    0.002337019, 0.001538008,
  9.258939e-11, 1.122597e-09, 7.505355e-09, 0.006208784, 0.02740415, 
    0.001225359, -0.003614697, 0.0007300325, 0.00357108, 0.002220568, 
    0.01638753, 0.0003815958, 0.0007290164, 0.0002074767, 0.0007796842, 
    0.0176662, 0.008517751, 0.004636841, 0.003740732, 0.01345408, 0.01182553, 
    0.0003346369, 0.2952569, 0.06694016, 3.018505e-05, 5.457913e-06, 
    0.001636069, -3.217748e-07, 4.674671e-10,
  9.290253e-10, -2.819563e-05, 4.327076e-05, 0.0001658606, 6.298557e-07, 
    0.001639332, 0.02598526, 0.005357937, 0.02043504, 0.05471805, 0.02259793, 
    0.000848634, 0.0001342101, 0.0004219302, 0.0009939428, 0.002774774, 
    0.005245504, 0.003734532, 0.02241674, 0.0655046, 0.009190053, 0.08707148, 
    0.001456404, -0.00260274, 2.16482e-05, 0.0002282193, 0.0008042498, 
    3.038092e-05, 1.084506e-09,
  -5.530512e-06, 0.02629256, 0.0086984, 0.01623086, 0.08429903, 
    -0.0001395621, 0.001313228, 0.008490286, 0.01988295, 0.05438516, 
    0.06631174, 0.009558347, 0.02549913, 0.03090131, 0.04608789, 0.1128156, 
    0.02436872, 0.01385576, 0.01161533, 0.02280914, 0.1148068, 0.2071743, 
    0.09369431, 0.04976897, 0.007724358, 0.005203755, 0.004070391, 
    0.004673663, 0.0009064176,
  0.01333649, 0.01834888, 0.03719751, 0.3853842, 0.008357371, 0.07596666, 
    0.1162928, -0.0004871471, 0.001259492, 0.05023451, 0.1424843, 0.0501306, 
    0.07165516, 0.03736065, 0.0772615, 0.07459916, 0.2136167, 0.1005061, 
    0.04226446, 0.3359427, 0.05783534, 0.007624197, 0.145081, 0.1322315, 
    0.04842648, 0.04247219, 0.02141162, 0.01393306, 0.05858394,
  0.3371131, 0.4238721, 0.4420171, 0.3826278, 0.320744, 0.3363609, 
    0.09443133, 0.1480732, 0.05888997, 0.1442124, 0.1679311, 0.305186, 
    0.02666852, 0.04958802, 0.03657785, 0.1535302, 0.2219053, 0.1634847, 
    0.09811848, 0.4744482, 0.08105853, 0.1208775, 0.2150165, 0.5514444, 
    0.116845, 0.09458103, 0.1137481, 0.1460527, 0.2391076,
  0.156837, 0.3007386, 0.4175221, 0.6753238, 0.7037835, 0.5670294, 0.5055485, 
    0.4544719, 0.5884855, 0.6391428, 0.6120564, 0.535303, 0.2240573, 
    0.2184657, 0.2418003, 0.3347883, 0.5638, 0.3123324, 0.3392063, 0.2944776, 
    0.6570975, 0.3635535, 0.3335256, 0.3368236, 0.05397316, 0.02876557, 
    0.1424485, 0.1316296, 0.1442542,
  0.06519327, 0.04538013, 0.2921245, 0.01924635, 0.08975494, 0.4164144, 
    0.4489317, 0.4577147, 0.4409648, 0.5510119, 0.6985769, 0.5135553, 
    0.6035851, 0.6159799, 0.593008, 0.4055298, 0.3699377, 0.2895006, 
    0.3368246, 0.25722, 0.4508716, 0.5141127, 0.5505475, 0.3161283, 
    0.3347593, 0.1794109, 0.3131558, 0.112578, 0.1858138,
  0.5044605, 0.3020464, 0.2405319, 0.2804871, 0.2739854, 0.328561, 0.4058727, 
    0.422971, 0.4361253, 0.5173734, 0.5059446, 0.6178747, 0.6750445, 
    0.7087557, 0.638221, 0.6334982, 0.6059582, 0.5822061, 0.631201, 
    0.6321325, 0.5981994, 0.3264024, 0.3849686, 0.3463102, 0.1049299, 
    0.08750113, 0.1108238, 0.1484899, 0.521639,
  0.1151061, 0.1179393, 0.1207726, 0.1236059, 0.1264391, 0.1292724, 
    0.1321056, 0.1000621, 0.1004082, 0.1007542, 0.1011003, 0.1014463, 
    0.1017924, 0.1021384, 0.1452283, 0.1407921, 0.1363559, 0.1319197, 
    0.1274835, 0.1230474, 0.1186112, 0.09534474, 0.09660161, 0.09785847, 
    0.09911534, 0.1003722, 0.1016291, 0.1028859, 0.1128395,
  0.05076362, 0.02477964, 0.01767227, 0.05597783, 0.07882905, 0.03401319, 
    0.09197623, 0.1101169, 0.08527919, 0.0419936, 0.02809788, 0.0191326, 
    0.02527875, 0.001322989, 0.07081317, 0.1551077, 0.1996531, 0.07548731, 
    0.01562707, 0.03249228, 0.02228332, 0.06327636, 0.06946661, 0.03848766, 
    0.011771, 0.02916158, 0.05128432, 0.04316786, 0.03467957,
  0.1616633, 0.06194706, 0.07210921, 0.05443026, 0.002524082, 0.2096765, 
    0.1223884, 0.01497591, 0.005357874, 0.001761827, 0.01827725, 0.05272607, 
    0.01086938, 0.09052669, 0.1858235, 0.164039, 0.2087389, 0.1888487, 
    0.2091968, 0.3173639, 0.1978373, 0.2474571, 0.1745576, 0.1181966, 
    0.2824923, 0.2774074, 0.07926586, 0.05881497, 0.1256859,
  0.1729656, 0.2054494, 0.2226687, 0.2288669, 0.3011385, 0.3074422, 0.40777, 
    0.2441507, 0.4253055, 0.3004519, 0.2008216, 0.1307116, 0.2622441, 
    0.2497328, 0.1891798, 0.2706662, 0.3389492, 0.3992725, 0.3138673, 
    0.1772763, 0.2583214, 0.1700367, 0.1731683, 0.1717062, 0.2559272, 
    0.323915, 0.2627189, 0.1548496, 0.1988398,
  0.2276984, 0.201166, 0.2277823, 0.1692919, 0.2073907, 0.2267737, 0.2021853, 
    0.1856075, 0.2855124, 0.1914339, 0.1124586, 0.06976434, 0.0517581, 
    0.0380284, 0.1856415, 0.2113062, 0.1808069, 0.1435319, 0.1274087, 
    0.1263249, 0.1078607, 0.1272884, 0.1475069, 0.07803259, 0.01227413, 
    0.1033612, 0.2060361, 0.2713562, 0.246826,
  0.158148, 0.06473104, 0.0297485, 0.06982581, 0.04497765, 0.02786314, 
    0.1367671, 0.1327364, 0.08273386, 0.05628503, 0.03597272, 0.02759582, 
    0.06257749, 0.1474169, 0.1264095, 0.0657887, 0.0505867, 0.07928594, 
    0.1450714, 0.1199871, 0.117309, 0.09139834, 0.03434638, 0.09851114, 
    0.007176225, 0.03556276, 0.07383825, 0.07002668, 0.1356356,
  0.03536739, 0.008317951, 0.006151367, 0.02015975, 0.03944676, 0.01229939, 
    0.06269419, 0.0303409, 0.01357405, 0.002097809, 0.0009154725, 
    3.378881e-06, 0.0003540572, 0.004230223, 0.0128662, 0.0179655, 
    0.001771406, 0.1496459, 0.1257601, 0.03620238, 0.007858748, 0.003648777, 
    0.01277833, 0.0158235, 0.003808086, 0.04446591, 0.08803464, 0.009589458, 
    0.02598318,
  0.01496532, 0.03693257, 0.00546913, 0.006747913, -0.00107918, 0.0005196505, 
    0.0007687421, 0.0008866232, 0.004083758, 0.003096495, 3.994046e-06, 
    9.060313e-06, 0.0007428705, 0.0004062961, 0.002661939, 0.001632036, 
    0.00127313, 0.0001303891, 8.139836e-06, 9.67491e-05, 7.112398e-05, 
    0.003567128, 0.01525368, 0.03328909, 0.0121475, 0.1091549, 0.0005208406, 
    0.003424844, 0.003913484,
  0.01702296, 0.006353971, 0.05032036, 0.05589083, 0.0006551782, 0.004528074, 
    0.0006588429, 0.0008677, 0.000886469, 0.003497661, 0.001109634, 
    0.0006955462, 0.000253558, 7.076254e-05, 0.0004602673, 0.0007040959, 
    0.0003945282, 0.000384353, 0.0002785445, 0.0004722529, 0.0008538324, 
    0.002841328, 0.0295141, 0.0004829609, 0.02090976, 4.604963e-05, 
    0.0003008892, 0.0009802368, 0.005333701,
  0.0008496873, 0.004408826, 0.02317574, 0.06340091, 0.0009454404, 
    0.001012241, 0.0003176347, 0.0005629131, 0.04197353, 0.06901493, 
    0.0001041684, 0.001017061, 0.0002563027, 0.0008773382, 0.001296543, 
    0.0005073564, 6.316308e-05, 0.0002876183, 0.0008941285, 0.0008884257, 
    0.004663145, 0.01797048, 0.03117159, 0.00511173, 0.002551897, 
    0.0007733771, 0.005697859, 0.0009881972, 0.0006676094,
  9.372772e-11, 1.119006e-09, 7.04095e-09, 0.006093263, 0.01380116, 
    0.0007771453, -0.00288052, 0.0005229383, 0.002370513, 0.001371427, 
    0.007314412, 0.000161975, 0.000335175, 9.71192e-06, 0.0003297934, 
    0.01078511, 0.004207537, 0.001817827, 0.001098932, 0.006480446, 
    0.005332631, 0.0001858238, 0.2441365, 0.0498141, 1.72699e-05, 
    2.785905e-06, 0.001103872, -5.264576e-07, 4.695122e-10,
  1.063262e-09, -1.607817e-05, 2.7852e-05, 0.0001770518, 4.363744e-07, 
    0.001226661, 0.0150857, 0.003003154, 0.0165688, 0.03113156, 0.009284479, 
    0.0004195933, 8.738972e-05, 0.0002792985, 0.0006595221, 0.001366871, 
    0.002462148, 0.001644763, 0.01244056, 0.03165253, 0.005611572, 
    0.06562524, 0.0009839397, -0.002290497, 1.198635e-05, 0.000143742, 
    0.000551054, 1.99538e-05, 1.135801e-09,
  -1.438943e-05, 0.01953645, 0.006601011, 0.01148488, 0.06985746, 
    -0.000145032, 0.002272714, 0.01188159, 0.02408339, 0.03524135, 
    0.05315689, 0.005498905, 0.01116327, 0.01609367, 0.02206567, 0.07124726, 
    0.01137659, 0.007788105, 0.006524181, 0.01623323, 0.09860947, 0.1794953, 
    0.07809366, 0.02918732, 0.003446226, 0.002941743, 0.0024625, 0.003149903, 
    0.0001858385,
  0.01078896, 0.01056757, 0.02551041, 0.3614002, 0.004737844, 0.0551121, 
    0.09606594, -0.0003048316, 0.0003878341, 0.04104252, 0.1296628, 
    0.03821028, 0.05467498, 0.02544877, 0.05719035, 0.05466388, 0.1601875, 
    0.07350268, 0.02542128, 0.3085908, 0.04735585, 0.006568988, 0.1230697, 
    0.1049602, 0.03405308, 0.02342748, 0.01054592, 0.007797356, 0.0363339,
  0.2489521, 0.3532161, 0.3667173, 0.3095582, 0.2479555, 0.2780144, 
    0.06960747, 0.1266559, 0.08739352, 0.1240693, 0.1567934, 0.300035, 
    0.01564304, 0.03960761, 0.02633992, 0.1222497, 0.1683649, 0.1221453, 
    0.06419352, 0.43145, 0.06511867, 0.08505616, 0.1753901, 0.5125409, 
    0.09824315, 0.07525022, 0.07729632, 0.09826883, 0.1621671,
  0.1048451, 0.2946263, 0.3536707, 0.6071925, 0.6526579, 0.4870683, 
    0.4868994, 0.4319427, 0.5791979, 0.5931771, 0.5899677, 0.5796738, 
    0.2502266, 0.2492462, 0.2086563, 0.3124035, 0.6079752, 0.2691328, 
    0.3163463, 0.3112128, 0.6500012, 0.3081977, 0.2547634, 0.4055002, 
    0.04050185, 0.02255853, 0.1095793, 0.08576547, 0.09906875,
  0.0519469, 0.03561386, 0.3600209, 0.01080605, 0.07291837, 0.3260708, 
    0.4479049, 0.4622376, 0.4506387, 0.5966457, 0.6835464, 0.4957522, 
    0.7603397, 0.5017387, 0.4838501, 0.3500813, 0.3605011, 0.2008279, 
    0.3137334, 0.2382029, 0.5240028, 0.6154947, 0.4943681, 0.4343159, 
    0.3848487, 0.1460417, 0.2831443, 0.09135678, 0.1535375,
  0.4851466, 0.2659999, 0.2640692, 0.2815238, 0.3406365, 0.3774038, 0.412447, 
    0.4551378, 0.5023334, 0.4694507, 0.5054253, 0.5418931, 0.6076173, 
    0.6983948, 0.6598243, 0.5814155, 0.5889478, 0.5568643, 0.5592581, 
    0.4789572, 0.5095509, 0.2993264, 0.3842137, 0.4246954, 0.09773063, 
    0.07913936, 0.09716619, 0.1337001, 0.526122,
  0.08991197, 0.09149998, 0.093088, 0.09467603, 0.09626404, 0.09785206, 
    0.09944008, 0.07241698, 0.07138316, 0.07034933, 0.0693155, 0.06828167, 
    0.06724785, 0.06621402, 0.08737243, 0.08529633, 0.08322024, 0.08114414, 
    0.07906805, 0.07699195, 0.07491586, 0.0696598, 0.07118171, 0.07270361, 
    0.07422552, 0.07574742, 0.07726932, 0.07879123, 0.08864155,
  0.04553084, 0.01698917, 0.01751745, 0.0641911, 0.05457126, 0.02339314, 
    0.06819545, 0.08166731, 0.04964029, 0.02452592, 0.01786528, 0.01606631, 
    0.0179825, 0.001294372, 0.0593107, 0.1329544, 0.1948243, 0.06522014, 
    0.01330429, 0.02860216, 0.01420909, 0.04587627, 0.05016017, 0.02875976, 
    0.009593111, 0.02469371, 0.04083534, 0.03537486, 0.0256342,
  0.151239, 0.05356894, 0.06712376, 0.05202996, 0.001765398, 0.1690702, 
    0.1094837, 0.01213132, 0.002978312, 0.001231826, 0.01259122, 0.04078354, 
    0.007544668, 0.08131397, 0.1554494, 0.1205259, 0.1551265, 0.1488286, 
    0.1577237, 0.2385043, 0.1737752, 0.1943839, 0.1466102, 0.08724956, 
    0.2253254, 0.2347349, 0.05927429, 0.04774744, 0.1095456,
  0.1296602, 0.1441261, 0.1614666, 0.1719946, 0.2291196, 0.233978, 0.318364, 
    0.1936783, 0.3339452, 0.2388216, 0.1566578, 0.106424, 0.2023161, 
    0.2078187, 0.1506721, 0.2196727, 0.2796192, 0.3272802, 0.2501717, 
    0.1378717, 0.1928638, 0.1161582, 0.1264195, 0.1204086, 0.2030977, 
    0.2514119, 0.1869272, 0.1205169, 0.156993,
  0.1813188, 0.1649219, 0.186434, 0.1328488, 0.1657216, 0.1960325, 0.1571267, 
    0.1341762, 0.2228365, 0.1475548, 0.0780085, 0.04547504, 0.03280077, 
    0.02805121, 0.1446196, 0.1539391, 0.126699, 0.09387901, 0.08444165, 
    0.08779021, 0.07405511, 0.09018011, 0.1115893, 0.06596122, 0.005560888, 
    0.08334257, 0.156112, 0.2245096, 0.1982976,
  0.1086279, 0.03948366, 0.02250623, 0.04410352, 0.02479951, 0.01781073, 
    0.09044878, 0.08572128, 0.05954871, 0.04078578, 0.0278785, 0.02126568, 
    0.04259226, 0.1065416, 0.1038142, 0.0396307, 0.03513759, 0.05883997, 
    0.1003005, 0.07934967, 0.07135528, 0.0608228, 0.02174623, 0.09738135, 
    0.00472545, 0.02030981, 0.04689519, 0.04631728, 0.09485111,
  0.02343774, 0.006013076, 0.003238069, 0.01281658, 0.02383855, 0.009073872, 
    0.04037399, 0.01718707, 0.01058996, 0.001606062, 0.0005396485, 
    -7.691734e-07, 0.0009217809, 0.002265991, 0.00423987, 0.009511154, 
    0.001360044, 0.1107493, 0.08040565, 0.01842112, 0.004160285, 0.002680184, 
    0.009514503, 0.01177584, 0.00274804, 0.02457061, 0.05365101, 0.004397512, 
    0.01343977,
  0.01050283, 0.02554296, 0.00310052, 0.004587207, -0.0009408311, 
    0.0003595818, 0.0004905082, 0.0006717751, 0.003076787, 0.002289666, 
    5.529028e-07, -3.239673e-06, 0.0005281765, 0.0003033447, 0.0009562859, 
    0.001072088, 0.0007666451, 8.698317e-05, 5.24949e-06, 7.936673e-05, 
    5.268507e-05, 0.002555492, 0.01074486, 0.02487078, 0.01001554, 0.0859957, 
    0.0003905525, 0.002551085, 0.002738043,
  0.01255543, 0.004187624, 0.0495426, 0.05319721, 0.0004372943, 0.00227646, 
    0.000269925, 0.0003783798, 0.0006292178, 0.00267717, 0.0004779547, 
    0.0004008944, 0.0002506632, 5.61664e-05, 0.0003173569, 0.0003455839, 
    0.0002215954, 0.0002094766, 0.0002075266, 0.0003566327, 0.0006468801, 
    0.002055018, 0.02195383, 0.003931255, 0.0161204, 0.0007757882, 
    0.0002641557, 0.000707506, 0.003764235,
  0.0004243424, 0.01006524, 0.0187868, 0.05549134, 0.0007303649, 0.000615869, 
    0.000264467, 0.0002898806, 0.04925774, 0.07535307, 7.38873e-05, 
    0.0007655635, 0.0001795034, 0.0006373976, 0.0007803931, 0.0003663424, 
    4.385752e-05, 0.0001735668, 0.0006286668, 0.0006155411, 0.003413462, 
    0.01216568, 0.02059302, 0.00626645, 0.001742223, 0.0003783993, 
    0.002254618, 0.0004355051, 0.0003594834,
  9.627309e-11, 1.126639e-09, 6.714541e-09, 0.009269476, 0.009255267, 
    0.0005704314, -0.002048844, 0.0004114051, 0.001742459, 0.001021032, 
    0.00394535, 9.765943e-05, 0.0001964843, 2.35211e-05, 0.0001905666, 
    0.00526507, 0.001920175, 0.0009403018, 0.0005008744, 0.003530732, 
    0.002501688, 0.0001285086, 0.1967751, 0.03648688, 1.201497e-05, 
    1.958743e-06, 0.0008287172, -4.990299e-07, 4.714109e-10,
  1.134448e-09, -9.681668e-06, 2.04269e-05, 0.000170612, 3.308704e-07, 
    0.000989847, 0.009847481, 0.002111774, 0.01248717, 0.01936048, 
    0.004914129, 0.0002869146, 6.461018e-05, 0.000211248, 0.0004993171, 
    0.0008484377, 0.00122548, 0.0008000358, 0.005490785, 0.01790129, 
    0.004105524, 0.05234401, 0.0007483267, -0.001934976, 8.560516e-06, 
    0.0001049149, 0.0004225597, 1.480996e-05, 1.046372e-09,
  -1.800573e-05, 0.0135229, 0.004610434, 0.009020716, 0.05994889, 
    -0.000131759, 0.00638968, 0.0221836, 0.03086398, 0.02366435, 0.03805421, 
    0.003389357, 0.005374381, 0.006850703, 0.01281309, 0.04627812, 
    0.006382768, 0.004877867, 0.004022058, 0.01254146, 0.08643527, 0.1504758, 
    0.067935, 0.0192761, 0.00219408, 0.002008076, 0.001727797, 0.002413644, 
    0.0001362356,
  0.01008602, 0.007716683, 0.02016021, 0.3383305, 0.003205344, 0.0407435, 
    0.07860807, -0.0001539324, 0.0002781446, 0.03636006, 0.1205376, 
    0.02779897, 0.0439181, 0.01732528, 0.0461142, 0.04332393, 0.121728, 
    0.05241059, 0.01527911, 0.2848966, 0.04275177, 0.006984604, 0.1130697, 
    0.08440418, 0.02347319, 0.01344051, 0.005660873, 0.005197087, 0.02257635,
  0.1935746, 0.307058, 0.3210377, 0.2589208, 0.2005992, 0.2358512, 
    0.05909649, 0.1265153, 0.169488, 0.109844, 0.1475611, 0.3032736, 
    0.01145124, 0.03317484, 0.02108031, 0.1003833, 0.1319139, 0.09167466, 
    0.0449984, 0.4051325, 0.05623282, 0.06841572, 0.1555374, 0.4954681, 
    0.08647477, 0.06118865, 0.05481967, 0.06506194, 0.1129098,
  0.07741226, 0.3162304, 0.3282377, 0.5502677, 0.5867256, 0.4085928, 
    0.4053965, 0.3763753, 0.5035368, 0.4939177, 0.5450363, 0.6179402, 
    0.2986202, 0.2828367, 0.184741, 0.2896915, 0.5784833, 0.2465549, 
    0.2923063, 0.3378868, 0.5988058, 0.2788765, 0.2011309, 0.3967923, 
    0.03376036, 0.02085683, 0.08485505, 0.05878696, 0.0704961,
  0.04215575, 0.03016517, 0.3785455, 0.007454432, 0.06318226, 0.2722388, 
    0.4888021, 0.4440668, 0.4777471, 0.6237121, 0.6823139, 0.4517018, 
    0.7515838, 0.3737204, 0.373899, 0.2640376, 0.3779507, 0.1538198, 
    0.2630268, 0.1978518, 0.4821765, 0.5692836, 0.505957, 0.4840134, 
    0.386788, 0.09985206, 0.3716778, 0.07457685, 0.1307938,
  0.498836, 0.2427349, 0.2515836, 0.2705835, 0.30288, 0.3652399, 0.368722, 
    0.3568502, 0.3586487, 0.3382948, 0.3881122, 0.3867258, 0.4363232, 
    0.509382, 0.4411786, 0.436958, 0.476602, 0.3936258, 0.3995194, 0.3427987, 
    0.3891856, 0.2725961, 0.3857348, 0.5142663, 0.1031421, 0.04940819, 
    0.0983767, 0.1461025, 0.4888394,
  0.0681904, 0.06946099, 0.07073158, 0.07200217, 0.07327276, 0.07454335, 
    0.07581393, 0.05947545, 0.05850072, 0.057526, 0.05655127, 0.05557655, 
    0.05460182, 0.0536271, 0.06627633, 0.06478909, 0.06330187, 0.06181464, 
    0.06032741, 0.05884018, 0.05735295, 0.05712727, 0.05831863, 0.05951, 
    0.06070136, 0.06189273, 0.06308409, 0.06427545, 0.06717393,
  0.04449594, 0.01249589, 0.02495449, 0.07469007, 0.0515782, 0.01993208, 
    0.05671283, 0.08003597, 0.03524838, 0.01759019, 0.013679, 0.01439018, 
    0.01641501, 0.001212219, 0.05505277, 0.1197302, 0.1943943, 0.06081341, 
    0.01196413, 0.04280983, 0.01128733, 0.03577934, 0.03676278, 0.02558552, 
    0.008511445, 0.02208818, 0.03631662, 0.03098612, 0.02148177,
  0.1466166, 0.0488786, 0.0686131, 0.04954228, 0.001385547, 0.1499191, 
    0.09911247, 0.01074658, 0.00195412, 0.001063276, 0.01050626, 0.03453818, 
    0.005220238, 0.07914399, 0.1424491, 0.1014707, 0.1310848, 0.1307242, 
    0.1318098, 0.2031968, 0.1506822, 0.1619422, 0.1251881, 0.07116061, 
    0.1942487, 0.1945823, 0.05120405, 0.04199645, 0.1035223,
  0.1105572, 0.1236469, 0.1288993, 0.147409, 0.19914, 0.2022745, 0.2695021, 
    0.1669803, 0.2778286, 0.2069198, 0.1301895, 0.08526731, 0.1681832, 
    0.1711164, 0.1258011, 0.179434, 0.2383967, 0.2800377, 0.2117257, 
    0.1145912, 0.1509792, 0.0895411, 0.09794223, 0.09297861, 0.1676041, 
    0.2056397, 0.1554552, 0.1042711, 0.1351454,
  0.1538809, 0.1410625, 0.1594734, 0.1131542, 0.1389065, 0.1699532, 
    0.1270263, 0.1051217, 0.1819714, 0.1245328, 0.06196808, 0.03415915, 
    0.02501904, 0.02333953, 0.1081334, 0.117221, 0.0961586, 0.06887525, 
    0.06232235, 0.06371106, 0.05643113, 0.07057868, 0.08830341, 0.06668268, 
    0.003886728, 0.06766569, 0.1254014, 0.1885269, 0.1678814,
  0.07789616, 0.02646124, 0.01531102, 0.03024344, 0.01591874, 0.01253682, 
    0.06713894, 0.05547425, 0.04053865, 0.03308672, 0.02322916, 0.01789468, 
    0.02495338, 0.07567003, 0.09701727, 0.02687671, 0.02388098, 0.04226187, 
    0.07370929, 0.05353675, 0.0466829, 0.04514814, 0.01537899, 0.09789384, 
    0.00291377, 0.01415391, 0.03320216, 0.03488744, 0.07056683,
  0.01573507, 0.00491686, 0.003178427, 0.008733136, 0.01447214, 0.006945534, 
    0.0272452, 0.01124147, 0.009056865, 0.001397104, 0.0003545922, 
    2.109262e-07, 0.009427571, 0.001627874, 0.00290074, 0.006578248, 
    0.001171324, 0.07048407, 0.05252897, 0.01041659, 0.003102262, 
    0.002210116, 0.007930147, 0.009581226, 0.003197528, 0.01454178, 
    0.03026306, 0.002698643, 0.009234073,
  0.008464177, 0.01992713, 0.001617166, 0.003623041, -0.0009887055, 
    0.0002705395, 0.0003887649, 0.000567149, 0.002595913, 0.001893492, 
    3.339626e-07, -1.921992e-06, 0.0004309185, 0.0002334023, 0.0006097413, 
    0.0008039462, 0.0005779748, 7.885916e-05, 4.744383e-06, 7.118364e-05, 
    4.395853e-05, 0.002100772, 0.008711615, 0.02058457, 0.02567862, 
    0.1829003, 0.0003240728, 0.002105378, 0.002201402,
  0.01029154, 0.003096028, 0.09763747, 0.1005486, 0.0003295537, 0.001509037, 
    0.0001789977, 0.0002377244, 0.0004993852, 0.001909316, 0.0003223875, 
    0.0002975368, 0.0002093849, 4.747797e-05, 0.0002503661, 0.0002463803, 
    0.000160052, 0.0001512838, 0.0001711222, 0.0003008989, 0.000545534, 
    0.001685258, 0.01815228, 0.1076565, 0.02809585, 0.01110071, 0.0002328132, 
    0.0005839441, 0.003029332,
  0.0002962709, 0.01428851, 0.02090368, 0.06136626, 0.0003411664, 
    0.000467035, 0.0002196708, 0.0002103908, 0.09172846, 0.1308774, 
    6.023696e-05, 0.0006354308, 0.0001421324, 0.0005140156, 0.0005801179, 
    0.0003018242, 3.863198e-05, 0.0001345699, 0.0005064718, 0.0004945003, 
    0.002801458, 0.009588917, 0.01623017, 0.08008671, 0.03767638, 
    0.0002578151, 0.001353806, 0.0002778235, 0.0002638823,
  1.011051e-10, 1.141035e-09, 6.480306e-09, 0.01898565, 0.007426438, 
    0.000472561, -0.001553836, 0.0003557951, 0.001394163, 0.0008650331, 
    0.002677558, 7.307057e-05, 0.0001453153, 3.530856e-05, 0.000150198, 
    0.002862612, 0.001123649, 0.0006181039, 0.000363062, 0.002394651, 
    0.001524208, 0.000108836, 0.2395078, 0.03402475, 9.078555e-06, 
    1.615817e-06, 0.0007054411, -1.127036e-07, 4.765515e-10,
  1.175756e-09, -6.317314e-06, 1.580881e-05, 0.0001624844, 2.689743e-07, 
    0.0008622612, 0.01126942, 0.001536034, 0.01309887, 0.01457085, 
    0.003460836, 0.0002366742, 5.428238e-05, 0.0001802323, 0.0004208573, 
    0.0006656112, 0.0008167944, 0.0004969526, 0.003116768, 0.01181905, 
    0.003355252, 0.0445169, 0.000636147, -0.001888307, 7.108727e-06, 
    8.624768e-05, 0.0003643539, 1.25399e-05, 1.029653e-09,
  -1.883265e-05, 0.01074788, 0.003584746, 0.008543084, 0.05804619, 
    -0.0001037785, 0.02098962, 0.06838282, 0.05660981, 0.02028961, 
    0.02877971, 0.002515235, 0.003324989, 0.003764248, 0.008789016, 
    0.0307719, 0.00476282, 0.003702952, 0.003004387, 0.01038029, 0.07677367, 
    0.1379504, 0.07722636, 0.0143404, 0.001755822, 0.001629838, 0.001431646, 
    0.002056024, 0.0008590496,
  0.01158944, 0.006041253, 0.01744494, 0.3341247, 0.002562793, 0.03409123, 
    0.07405473, 0.001274466, 0.0001964586, 0.0355934, 0.1253457, 0.02101247, 
    0.03907713, 0.01352284, 0.04123325, 0.03568596, 0.0964584, 0.0404217, 
    0.01110085, 0.2788795, 0.04501203, 0.007748815, 0.1104421, 0.06740201, 
    0.01858312, 0.008895209, 0.003866645, 0.004164998, 0.01908637,
  0.1656031, 0.3048982, 0.3076151, 0.2395717, 0.1819955, 0.2105428, 
    0.05548809, 0.2028879, 0.314116, 0.1124241, 0.1660308, 0.3374614, 
    0.009632409, 0.02827278, 0.01899217, 0.08456688, 0.1110279, 0.07436247, 
    0.03527153, 0.4240413, 0.0530068, 0.06734706, 0.1711764, 0.50741, 
    0.08767484, 0.05321095, 0.04194361, 0.04958961, 0.08617133,
  0.06356259, 0.3962265, 0.3285971, 0.5225387, 0.5433562, 0.431522, 
    0.4132012, 0.4104361, 0.5116165, 0.4963837, 0.5226175, 0.5312907, 
    0.3899905, 0.3556534, 0.1747681, 0.281387, 0.6099328, 0.2454823, 
    0.3134317, 0.4487432, 0.580955, 0.3122602, 0.175255, 0.4093128, 
    0.03097797, 0.02159883, 0.07343128, 0.04698035, 0.05605431,
  0.03703619, 0.02749078, 0.4343421, 0.005130751, 0.05869493, 0.2200496, 
    0.4670256, 0.4517674, 0.525245, 0.5983763, 0.6768637, 0.5145379, 
    0.6218007, 0.320293, 0.3308969, 0.2147725, 0.3928711, 0.1588796, 
    0.2571781, 0.1637147, 0.4618435, 0.5248522, 0.5354455, 0.5136203, 
    0.3679169, 0.09430744, 0.4486911, 0.07435939, 0.1197387,
  0.4954482, 0.2312361, 0.2315703, 0.2353521, 0.2474896, 0.3342416, 0.323862, 
    0.2981175, 0.2953403, 0.2618829, 0.305004, 0.2763806, 0.3318098, 
    0.419189, 0.3564775, 0.334916, 0.3684416, 0.3047583, 0.293665, 0.2686014, 
    0.2916448, 0.2590469, 0.4030436, 0.5787988, 0.1111051, 0.02722937, 
    0.1072609, 0.210192, 0.4583623 ;

 lat = -89.5, -79.5, -69.5, -59.5, -49.5, -39.5, -29.5, -19.5, -9.5, 0.5, 
    10.5, 20.5, 30.5, 40.5, 50.5, 60.5, 70.5, 80.5 ;

 lat_bnds =
  -90, -89,
  -80, -79,
  -70, -69,
  -60, -59,
  -50, -49,
  -40, -39,
  -30, -29,
  -20, -19,
  -10, -9,
  0, 1,
  10, 11,
  20, 21,
  30, 31,
  40, 41,
  50, 51,
  60, 61,
  70, 71,
  80, 81 ;

 lon = 0.625, 13.125, 25.625, 38.125, 50.625, 63.125, 75.625, 88.125, 
    100.625, 113.125, 125.625, 138.125, 150.625, 163.125, 175.625, 188.125, 
    200.625, 213.125, 225.625, 238.125, 250.625, 263.125, 275.625, 288.125, 
    300.625, 313.125, 325.625, 338.125, 350.625 ;

 lon_bnds =
  0, 1.25,
  12.5, 13.75,
  25, 26.25,
  37.5, 38.75,
  50, 51.25,
  62.5, 63.75,
  75, 76.25,
  87.5, 88.75,
  100, 101.25,
  112.5, 113.75,
  125, 126.25,
  137.5, 138.75,
  150, 151.25,
  162.5, 163.75,
  175, 176.25,
  187.5, 188.75,
  200, 201.25,
  212.5, 213.75,
  225, 226.25,
  237.5, 238.75,
  250, 251.25,
  262.5, 263.75,
  275, 276.25,
  287.5, 288.75,
  300, 301.25,
  312.5, 313.75,
  325, 326.25,
  337.5, 338.75,
  350, 351.25 ;

 pfull = 0.0252729048206747, 0.0885404738757409, 0.213072411383256, 
    0.41190537807884, 0.671080828691593, 0.987471468515016, 1.36790961365676, 
    1.82562112064242, 2.38097588033244, 3.06218961364243, 3.90121721567151, 
    4.9296281825995, 6.18008131929323, 7.68875807563375, 9.49537809361575, 
    11.643153995098, 14.1786857151188, 17.1517875598959, 20.6152476986609, 
    24.6245259348741, 29.237386591333, 34.5134757786445, 40.5138467378254, 
    47.3004421634272, 54.9355325495126, 63.4811392623337, 72.9984371159701, 
    83.5471442618119, 95.1849171805989, 107.966767294215, 121.944503506415, 
    137.166169497631, 153.675572970355, 171.511834307961, 190.708985325578, 
    211.295632932361, 233.294677858721, 256.723099608772, 281.591803639405, 
    307.905555737256, 335.66293113824, 364.856338389786, 395.47216160598, 
    427.490864234311, 460.887168786725, 495.630391513078, 531.761718445649, 
    569.289185351388, 607.768705103107, 646.445374671436, 684.792067788697, 
    722.468679913451, 759.124006783627, 794.401045766566, 827.769968639223, 
    858.597822486016, 886.389109609622, 910.841030891388, 931.860653469283, 
    949.549679924174, 964.159924710431, 976.012345333387, 985.470174132691, 
    992.77226220014, 997.948601287575 ;

 time = 746.5, 776, 805.5, 836, 866.5, 897, 927.5, 958.5, 989, 1019.5, 1050, 
    1080.5 ;

 time_bnds =
  731, 762,
  762, 790,
  790, 821,
  821, 851,
  851, 882,
  882, 912,
  912, 943,
  943, 974,
  974, 1004,
  1004, 1035,
  1035, 1065,
  1065, 1096 ;
}
