netcdf atmos.1980-1981.aliq.10 {
dimensions:
	time = UNLIMITED ; // (1 currently)
	pfull = 65 ;
	lat = 18 ;
	lon = 29 ;
	bnds = 2 ;
variables:
	float aliq(time, pfull, lat, lon) ;
		aliq:long_name = "Cloud fraction for large-scale liquid clouds" ;
		aliq:units = "dimensionless" ;
		aliq:_FillValue = -999.f ;
		aliq:missing_value = -999.f ;
		aliq:interp_method = "conserve_order2" ;
		aliq:cell_methods = "time: mean within months time: mean over years" ;
		aliq:time_avg_info = "average_T1,average_T2,average_DT" ;
	double average_DT(time) ;
		average_DT:long_name = "Length of average period" ;
		average_DT:units = "days" ;
	double average_T1(time) ;
		average_T1:long_name = "Start time for average period" ;
		average_T1:units = "days since 1979-01-01 00:00:00" ;
	double average_T2(time) ;
		average_T2:long_name = "End time for average period" ;
		average_T2:units = "days since 1979-01-01 00:00:00" ;
	double climatology_bounds(time, bnds) ;
	double lat(lat) ;
		lat:standard_name = "latitude" ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_N" ;
		lat:axis = "Y" ;
		lat:bounds = "lat_bnds" ;
	double lat_bnds(lat, bnds) ;
	double lon(lon) ;
		lon:standard_name = "longitude" ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_E" ;
		lon:axis = "X" ;
		lon:bounds = "lon_bnds" ;
	double lon_bnds(lon, bnds) ;
	double pfull(pfull) ;
		pfull:standard_name = "air_pressure" ;
		pfull:long_name = "ref full pressure level" ;
		pfull:units = "mb" ;
		pfull:positive = "down" ;
		pfull:axis = "Z" ;
	double time(time) ;
		time:standard_name = "time" ;
		time:long_name = "time" ;
		time:climatology = "climatology_bounds" ;
		time:units = "days since 1979-01-01 00:00:00" ;
		time:calendar = "standard" ;
		time:axis = "T" ;

// global attributes:
		:CDI = "Climate Data Interface version 2.4.4 (https://mpimet.mpg.de/cdi)" ;
		:Conventions = "CF-1.6" ;
		:title = "c96L65_am5f9d8r0_amip" ;
		:associated_files = "area: 19800101.grid_spec.nc" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
		:code_release_version = "2024.05" ;
		:git_hash = "5d306c05d9fe755cab04eedc8fd3de0d3c8355a0" ;
		:creationtime = "Mon Aug 25 14:09:46 2025" ;
		:hostname = "pp050" ;
		:history = "Mon Aug 25 13:32:22 2025: ncks -d lat,,,10 -d lon,,,10 atmos.1980-1981.aliq.10.nc reduced/atmos.1980-1981.aliq.10.nc\n",
			"Mon Aug 25 14:40:53 2025: cdo -O -s -select,month=10 merged_output.nc monthly_nc_files/all_years.10.nc\n",
			"Mon Aug 25 14:40:11 2025: cdo -O -s -mergetime /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/shards/ts/regrid-xy/180_288.conserve_order2/atmos_month/P1M/P1Y/atmos_month.198001-198012.aliq.nc /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/shards/ts/regrid-xy/180_288.conserve_order2/atmos_month/P1M/P1Y/atmos_month.198101-198112.aliq.nc merged_output.nc\n",
			"Mon Aug 25 14:12:17 2025: cdo --history splitname 19800101.atmos_month.nc /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/cycle/19800101T0000Z/split/regrid-xy/180_288.conserve_order2/19800101.atmos_month.\n",
			"fregrid --debug --standard_dimension --input_mosaic C96_mosaic.nc --input_dir /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/cycle/19800101T0000Z/history/native --input_file 19800101.atmos_month --associated_file_dir /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/cycle/19800101T0000Z/history/native --interp_method conserve_order2 --remap_file fregrid_remap_file_288_by_180.nc --nlon 288 --nlat 180 --scalar_field (**please see the field list in this file**) --output_file 19800101.atmos_month.nc" ;
		:CDO = "Climate Data Operators version 2.4.4 (https://mpimet.mpg.de/cdo)" ;
		:comment = "FMS time averaging, version 3.0, precision=double" ;
		:NCO = "netCDF Operators version 5.2.4 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco, Citation = 10.1016/j.envsoft.2008.03.004)" ;
data:

 aliq =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.28785e-05, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 3.077326e-05, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.115413e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.797668e-10, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, -4.062229e-06, 0, 0, 0, 0, 0, -3.024428e-06, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, -3.252877e-06, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -3.663882e-05, -3.653159e-05, 0.001046124, 
    0, 0, -1.395827e-05, -7.369554e-06, 0, -2.079772e-06, 0, -3.61489e-06, 0, 
    0, 0.0006390217, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2.148844e-06, 0.0002884606, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, -2.041112e-06, 0, 0, 0, 0, 0, 0, 0, -1.873014e-05, 
    -9.305526e-06, 0, 0, 0, 0, 0, 0, 0, 0, -1.237905e-05, 0, 0, 0, 0, 0,
  0, 0.001059221, 0.0001529191, 0, 0, -2.402918e-11, 0, -1.624891e-05, 0, 0, 
    0, 0, 0, -1.311901e-05, -1.03397e-05, 0, 0, 0, 0, 0, 0, 0, 0, 
    -1.938506e-05, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, -8.424199e-06, 7.393283e-05, 0, -1.931313e-05, 
    -2.662121e-06, -0.000127653, 0.0002536455, 0.002572609, -4.553735e-06, 0, 
    0.0008326187, 0.0003682523, 0, -2.470914e-05, 0.001273177, 0.0004535588, 
    0, -1.134796e-05, 0.001662399, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0.003356201, 0, 0, -4.750814e-05, -2.077235e-06, 
    0.0003937452, -1.542263e-05, 8.064011e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -3.081815e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -6.024458e-06, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -1.315432e-05, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.034311e-05, 0, 0, 0, 0, 
    0, 0, 0, -1.484354e-05, 0, 0, 0, 0,
  0, -4.027626e-06, 0, 0, 0, -3.578624e-05, -5.703768e-05, -1.455136e-05, 0, 
    0, 0, 0, 0, 0.001425016, 0.0001806177, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0003562564, 0, 0, 0, 0, 0,
  0, 0.001941762, 0.001263625, 0, 0, 5.086427e-05, 0, -1.994182e-05, 
    -3.160451e-06, -7.625165e-06, 0, 0, -7.352927e-06, -2.039783e-05, 
    -4.652865e-05, 0, 0, 0, 0, 0, 0, 0, 0, -1.483315e-05, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, -0.0001112963, 0.003031405, 6.2297e-05, -4.025013e-05, 
    -1.183893e-05, 0.0005136461, 0.005291705, 0.005503579, -1.42257e-05, 
    0.000118295, 0.003989509, 0.003235482, 0.0006351958, -0.0001030804, 
    0.002864096, 0.002230146, -1.46434e-05, -7.676573e-06, 0.003135742, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0.005149684, -2.308925e-07, 0, 0.0002739539, 0.000461184, 
    0.0006935676, -0.0001123836, 0.002156049, 0, 0, 0, 0, 0, 0, 0, 
    -4.444045e-05, 0, 0, 0, 0.0004774467, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -6.189666e-06, 4.456319e-05, 0.0002477206, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4.269586e-05, 1.853502e-05, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -5.848921e-05, -2.305696e-05, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.79334e-05, 0.0002558373, 
    -4.774202e-06, 0, 0, 0, 0, 0, 0, -3.66011e-05, 0, 0, 0, 0,
  0, -1.6232e-05, 0, 0, -2.63732e-06, -1.308557e-05, -0.000133448, 
    0.0001094686, -8.304218e-06, 0, 0, 0, -2.578045e-05, 0.001390122, 
    0.000126255, 0, 0, 0, 0, 0, 0, 0, 0, 0.001050768, 0, 0, 0, 0, 0,
  0, 0.006632048, 0.00256126, 0, 0, 0.002074997, 0, -8.80576e-06, 
    -3.124835e-05, -2.049057e-05, 0, 0.0002220524, 7.384006e-07, 0.00140285, 
    -7.487946e-05, 0, 0, 0, 0, 0, 0, 0, 0, -3.139429e-05, 0, 0, 0.001043531, 
    0, 0,
  0, 0, 0, -2.366881e-06, 0, 0, 0.0006650235, 0.0040339, 0.002785584, 
    -0.0001702421, 0.0003194789, 0.003423012, 0.01875453, 0.01307655, 
    0.0007198729, 0.003485608, 0.009489866, 0.008825472, 0.001707932, 
    0.001099773, 0.006031923, 0.005126227, -0.000107527, -4.375159e-05, 
    0.004567691, -3.723307e-06, -3.037505e-05, 0, 0,
  0, 0, 0, 0, 0, 1.731677e-05, 0.007099652, -9.263047e-06, -5.067242e-06, 
    0.001454038, 0.002784122, 0.006383769, 0.002041088, 0.008408375, 0, 
    -1.745905e-05, 0, -1.741993e-05, 0, 0, 4.46659e-06, 0.0005317475, 0, 0, 
    0, 0.001536643, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 3.301136e-08, 0, 6.108866e-05, 3.625737e-05, 
    0.003521742, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0003840811, 0.0008247863, 0, 
    0.0002198956, 0, 0, 0, 0, 0, 0, 8.93206e-05, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3.89958e-05, 0, 0, 0, 0,
  0, 0, 0, 0.0006374982, -5.765111e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 3.990459e-05, 0, 0, 0, 0, 0.0003597101, 0.00248824, -9.791864e-07, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0008064749, 0.001571481, 
    0.001301457, -4.366572e-06, 0, 0, 0, 0, 0, 0.0001480721, 4.628861e-05, 0, 
    0, 0,
  0, -4.161074e-05, 0, 0, -4.008505e-06, 0.001542222, -0.0002015589, 
    0.001794502, -2.491265e-05, 0, 0, -7.559283e-06, -5.790951e-05, 
    0.002324492, 0.0002638703, -9.206056e-05, -3.485262e-05, 0, 0, 0, 0, 0, 
    0, 0.003403035, 0.0008017299, 0, 0, 0, 0,
  -7.333028e-06, 0.01357435, 0.004448621, 0, 0, 0.005706009, 0, 1.06491e-05, 
    -7.136603e-05, -4.380026e-05, 0, 0.0002252169, 3.401968e-05, 0.002837801, 
    6.865236e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0.0002635268, 0, -1.103626e-05, 
    0.002552448, -3.769771e-07, 0,
  0, 0, 0, -3.617557e-05, 0, 0, 0.002407311, 0.006209858, 0.008200975, 
    0.0007588283, 0.0006323833, 0.007046622, 0.03788309, 0.02755925, 
    0.002624498, 0.006916852, 0.01578655, 0.01802102, 0.006713922, 
    0.002924616, 0.009355471, 0.009531936, -0.000328245, 3.662261e-05, 
    0.00556512, 0.0001163516, 6.889757e-05, -5.161919e-06, 0.0004190384,
  0, 0, 0, 0, 0, -2.688698e-05, 0.009022744, 0.0001469711, -1.654935e-05, 
    0.002781069, 0.007327762, 0.01467185, 0.004705405, 0.01444933, 0, 
    -3.649016e-05, 0, 6.388692e-05, 0, 0, -1.097538e-06, 0.001082059, 0, 0, 
    0, 0.002905174, -8.595768e-06, 0, 0,
  0, 0, 0, 0, 0, 0, 0, -4.290794e-05, 0.001623574, 0, 0.001007176, 
    0.0007864958, 0.006652952, 0.0001405725, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -3.512358e-07, -3.477467e-06, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.025024e-07, 0.002262249, 0.005249035, 
    0.001588889, 0.0002685614, 0, -1.536195e-05, 0, 0, 0, 0, 0.001420722, 
    -4.174891e-06, -3.539717e-06, -1.905825e-05, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -9.023758e-06, 4.210187e-05, 
    -1.773413e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.276144e-05, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, -1.981034e-06, 0.0002848532, 0, 0, 0, 0, 0, 0, 0, 0, 
    -3.080433e-06, 0, 0.0004834802, 0, 0, -9.616551e-08, 0, 0, 0, 0, 
    0.001371593, -5.342526e-07, -2.571774e-06, 6.980449e-05, 0,
  0, 0, 0, 0.004646912, -1.075796e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -3.990848e-07, -5.68633e-06, 0, 0.0002360761, 0.002511682, 0, 0, 0, 0, 
    0.000969247, 0.008016023, 0.001240153, 0, 0,
  0, 0, 0, 0, -4.53698e-06, 0, 0, 0.000198077, 0, 0, 0, 0, 0, 0, 0, 
    0.001267529, 0.00251913, 0.004404634, -5.678923e-05, 0, 0, 0, 0, 0, 
    0.0006660407, 0.002584069, 0, 0, 0,
  0, -0.0001108521, -9.202968e-07, 0, 8.117838e-05, 0.006008772, 
    0.0004918993, 0.007593518, -6.958735e-05, 0, -8.976993e-07, 
    -1.943803e-05, 0.0006964155, 0.00545556, 0.001176016, -0.0001818687, 
    0.0008141837, 0, 0, 0, 0, 0, 0, 0.004596694, 0.001611255, 1.641177e-05, 
    0, 0, 0,
  -5.119125e-06, 0.0240855, 0.005798586, 0, 0, 0.01024693, -1.60788e-05, 
    0.0002766397, 0.0002089987, -0.0001063381, 0, 0.0005242861, 0.000388427, 
    0.004178373, 0.00063246, 0, -3.537565e-05, 0, 0, 0, 0, 0, 0, 0.001786649, 
    -1.015061e-06, -9.978489e-06, 0.004515488, -1.507909e-06, 0,
  0, 0, 0, 0.0005302939, 0, 0, 0.008437887, 0.009752105, 0.01751581, 
    0.004234714, 0.002591935, 0.01942775, 0.06430872, 0.05612, 0.007625886, 
    0.008468428, 0.02273119, 0.03401391, 0.01454132, 0.006208321, 0.01600738, 
    0.01463801, 0.001209811, 0.000650329, 0.006906384, 0.001452212, 
    0.001364351, 4.081492e-05, 0.002006393,
  0, 0, 0, 0, 0, 1.08716e-05, 0.01233813, 0.0003289037, -3.45666e-05, 
    0.005052859, 0.01495426, 0.02980518, 0.009528455, 0.02330769, 0, 
    -4.997339e-05, 0, 7.182395e-05, 0, 0, 0.0005095084, 0.001931808, 0, 
    0.0001527694, 0, 0.004255008, 0.0001000865, 0, 0,
  0, 0, 0, 0, 0, 0, 0, -0.0002167471, 0.003327544, 0, 0.002368589, 
    0.004862923, 0.009208082, 0.002890151, 0.0002449585, -4.59985e-06, 0, 0, 
    0, 0, 0, -1.194425e-06, 0, 0, 0.00136589, 3.084973e-06, 0.001059231, 0, 0,
  0.0001058739, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.306883e-06, 0.003454495, 
    0.00588933, 0.01337337, 0.002547282, 0.000496939, 0.0007296542, 
    0.0001289612, 0, 0, 0, 0.0004228526, 0.005039683, 0.0008355949, 
    -2.500323e-05, 0.0001829056, -4.068969e-05, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.857227e-05, 0, 0.003192562, 
    0.00238959, 0.0007976823, 9.984543e-06, 0, 0, 0, -9.9248e-06, 
    -5.090783e-06, 0, -2.972127e-06, -8.103326e-06, 0.001419961, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, -8.61434e-06, 0, 0, 0, 0, 0, 0, 0, 0, -4.141867e-08, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, -1.296756e-06, 0.000547438, 0.001498457, 0.00135915, 0, 0, 0, 0, 
    -3.885448e-06, -2.418611e-05, 3.454646e-05, 2.948909e-05, 0, 0.001385612, 
    0, 0.0002989728, 0.000105068, 0.0006583105, 0, 0, 0, 0.003235025, 
    -3.066088e-05, 0.0002782597, 0.0006325928, 0,
  0, 0, 0, 0.01151548, 0.0005706546, -4.906753e-05, 0, 0, 0, 0, 
    -2.856871e-05, 4.574067e-08, 0, -3.344112e-05, 5.774659e-05, 
    0.0007489754, -3.764578e-05, 4.417718e-05, 0.002277331, 0.005474825, 
    0.000155449, 0, 0, 0, 0.004489202, 0.0201983, 0.007416252, -1.796123e-05, 0,
  0, 9.214806e-05, -8.47202e-06, 0, 0.0002571923, 0, 0, 0.0008587749, 
    -8.898009e-08, 0, 0, 0, 0, -9.059823e-06, 5.847249e-07, 0.002878784, 
    0.006520079, 0.009412055, 0.000463487, -2.271182e-06, 0, 0, 0, 0, 
    0.001205347, 0.004465169, -8.639247e-05, 0, 0,
  0, 0.0005214239, 0.0008377909, 0, -1.258282e-06, 0.01690168, 0.003033165, 
    0.01785562, -0.0001217457, 0, 0.0004448731, 0.0004103672, 0.004248262, 
    0.01442961, 0.003965044, -0.0001019793, 0.004004078, -6.720505e-07, 0, 0, 
    0, 0, 0, 0.0130328, 0.002468754, 0.0001789731, 0, 0, 0,
  -1.111027e-05, 0.03596353, 0.007216333, 0, 0, 0.01491758, 7.388792e-05, 
    0.004191917, 0.002153224, -0.0001204584, -2.567001e-05, 0.00220778, 
    0.001762606, 0.01163611, 0.00170589, -1.112259e-06, 7.083252e-06, 
    8.451607e-06, 0, 0, 0, 0, -6.55112e-09, 0.005016148, 2.9258e-05, 
    2.066319e-05, 0.005878299, -4.736759e-06, 0,
  -1.461258e-06, -3.493718e-05, 0, 0.001782416, 0, -1.399607e-05, 0.01518265, 
    0.01735037, 0.0261745, 0.01221976, 0.007250727, 0.04331057, 0.09647869, 
    0.08444796, 0.01770988, 0.01525446, 0.03323794, 0.05366716, 0.02360424, 
    0.01163353, 0.02757421, 0.02094669, 0.003667056, 0.001925226, 
    0.007783308, 0.003015754, 0.002822277, 0.0006680971, 0.0034272,
  0, 0, 0, 0, 0, 0.0002806428, 0.01545118, 0.002108894, 0.0005182825, 
    0.007756261, 0.02500063, 0.05129719, 0.01595096, 0.03660657, 
    -2.643391e-05, -4.530916e-05, 0.0002443253, 0.001757209, -3.551041e-05, 
    -7.237638e-07, 0.001920307, 0.00512128, 2.635438e-05, 0.0006039792, 
    -1.125983e-05, 0.006954027, 0.003231812, 0, 0,
  0, 0, 0, 8.533251e-05, -1.640547e-06, 0, 0, 0.0002762738, 0.00659998, 
    6.226647e-05, 0.004407303, 0.01054796, 0.0136777, 0.003690894, 
    0.001898967, -7.886778e-05, -1.484419e-05, -9.775897e-07, 0.001190348, 
    0.0005449605, 0, -2.018768e-05, 0.0004375114, 3.510684e-05, 0.005987346, 
    0.0008815242, 0.002100316, 0, 0,
  0.001466497, -1.06293e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0.0004456508, 
    0.008281459, 0.01352587, 0.02098844, 0.007804762, 0.004053503, 
    0.004693407, 0.001105661, -2.117159e-06, 0, 0, 0.003804746, 0.008277635, 
    0.004214363, 0.001479564, 0.003635754, 0.0003264397, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -7.927955e-07, 0.0007931758, 3.389298e-05, 
    0.005438733, 0.00390309, 0.003666888, 0.0007169087, -1.721268e-05, 0, 0, 
    5.56156e-05, -1.27638e-05, 0, 6.673764e-05, 0.00137928, 0.00334593, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -6.310076e-07, 0, 0, 0, 0, -2.309739e-05, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, -4.982909e-06, 0.000939405, -1.145077e-05, -3.012554e-05, 
    0.0001146126, 0, 0, 0, 0, 0, 0.001126218, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.0001356898, 0.0002137787, 0, 0,
  0.0002415625, 0, 3.797648e-05, 0.001634267, 0.004671654, 0.005688151, 
    0.0027549, 0, 0, 0, 0, 0.0004810058, 8.06363e-05, 0.0007234528, 
    0.0003956744, 0.0004054221, 0.00178894, -3.602404e-06, 0.0007084981, 
    0.002030656, 0.002654695, -5.740973e-05, 0, 0, 0.006236841, 0.001479704, 
    0.002446641, 0.001506553, -3.942997e-05,
  0, -4.338489e-06, 0, 0.02136971, 0.005339745, -0.0001413105, 0, 0, 0, 
    -1.488725e-09, 1.10657e-05, 5.897101e-06, 7.409937e-05, 0.001302813, 
    0.004802687, 0.005263952, 0.0002274878, 0.002668686, 0.005539084, 
    0.0132531, 0.002805427, -3.810698e-10, 0, 0, 0.008191941, 0.0406689, 
    0.01780226, 0.001237124, -3.730005e-05,
  -1.032658e-08, 0.0002713861, 3.480645e-05, -3.261593e-06, 0.0010466, 
    -6.038834e-06, 0, 0.001767852, 0.0009683497, 0, 1.013923e-07, 
    -2.019299e-06, 1.015124e-07, 9.71891e-05, 0.007072125, 0.008371626, 
    0.01962347, 0.02185111, 0.005260561, -2.181803e-05, 1.623404e-07, 0, 0, 
    6.674461e-06, 0.003425034, 0.007494143, 0.002754862, 0.0001334896, 0,
  -3.904189e-11, 0.002388397, 0.002510497, 2.044839e-07, 0.001000088, 
    0.03780982, 0.01045736, 0.02780404, 0.001183696, 0, 0.002844774, 
    0.005674385, 0.009905696, 0.02885458, 0.01687292, 0.003794104, 
    0.01135432, -5.158739e-06, 7.325273e-07, 0, 0, 0, 5.492373e-07, 
    0.04261415, 0.02162564, 0.000387608, 4.602673e-13, 1.880337e-05, 0,
  0.001159097, 0.06225094, 0.01712954, 5.95109e-07, 0, 0.02451341, 
    9.899485e-05, 0.01550752, 0.02117976, 0.00332303, 8.293393e-05, 
    0.01672117, 0.01105918, 0.03771041, 0.004877229, 1.638892e-05, 
    0.0004638935, 1.325794e-05, -1.132694e-09, 0.0003941518, 0, 1.729358e-08, 
    4.128664e-05, 0.04056787, 0.001173764, 0.0001206355, 0.007235864, 
    0.0001068794, 0,
  0.0002724251, -5.614145e-05, -1.150917e-05, 0.002878198, -8.389142e-06, 
    -2.327439e-05, 0.02520677, 0.03218761, 0.04781428, 0.03377368, 
    0.02378289, 0.0942868, 0.1605808, 0.1244561, 0.05401061, 0.03644822, 
    0.05711188, 0.08532466, 0.03720949, 0.02156082, 0.04033446, 0.03968918, 
    0.02070099, 0.01239555, 0.01106277, 0.009378763, 0.009595795, 
    0.003568435, 0.00734954,
  0, 0, 0, -7.368951e-07, 0, 0.00119152, 0.0172108, 0.007417595, 0.005710243, 
    0.01243921, 0.03807184, 0.07655324, 0.03486228, 0.04727864, 0.0001294293, 
    0.001748514, 0.0009856474, 0.01140495, 0.0003528854, -6.99424e-06, 
    0.003929737, 0.01049121, 0.0007354467, 0.001146635, 0.0001269505, 
    0.009764207, 0.0115591, 0, -2.800677e-07,
  0, 0, 0, 0.0006621133, -2.300242e-05, 0, 0, 0.0006679646, 0.009509729, 
    0.0016052, 0.009850761, 0.02242317, 0.02628558, 0.008097241, 0.008442152, 
    0.001332602, 0.001567172, 0.000615218, 0.004922932, 0.003365697, 
    0.0002402432, -0.0001383201, 0.001504145, 0.0009647716, 0.009842714, 
    0.002877816, 0.002744392, 0, 0,
  0.001804088, 0.0002065775, 0, 0, 0, 0, 0, 0, 0, 0, 0.00444233, 0.02359646, 
    0.03464611, 0.03619978, 0.02188713, 0.01497416, 0.01093121, 0.00516451, 
    -8.478695e-06, 0, 0, 0.005437229, 0.0136684, 0.01089977, 0.01102048, 
    0.01229994, 0.004416073, 0.002636069, 0,
  0.0006087179, 0.0003906134, -7.156894e-06, 0, 0, 0, 0, 0, 0, 0, 0, 
    -5.224713e-05, 0.003892024, 0.001110256, 0.00716092, 0.005150896, 
    0.01401454, 0.006971464, 0.002598192, -7.704663e-06, 0, 0.001002752, 
    -3.708743e-05, 0.0001832454, 0.002615478, 0.007953199, 0.01271774, 
    0.0002164594, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -3.126918e-06, 0, 0, 0, 
    -6.351674e-06, 0, -7.328557e-07, -1.240572e-05, 8.17028e-05, 
    -6.420041e-05, -1.243259e-05, 7.352456e-05,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  -3.989801e-05, 5.811437e-05, 4.360227e-05, 0.001606526, 0.001176498, 
    0.001116884, 0.00195457, 0.001228629, 0, 0, 0, 0, 0, 0.002835206, 0, 
    9.050935e-05, 2.709315e-05, 0, 0, 0.0001612176, 0, -9.480197e-07, 0, 0, 
    -5.615699e-07, 0.001441743, 0.002291511, -4.35471e-05, -7.202078e-06,
  0.003356155, 8.269308e-05, 0.001470822, 0.00629814, 0.01463579, 0.01177058, 
    0.004449083, -2.487664e-05, 0, 0, -1.230246e-15, 0.002324874, 
    0.004456689, 0.003220654, 0.00578516, 0.00194951, 0.004985509, 
    0.000444025, 0.003437433, 0.006098731, 0.004755009, 0.00200355, 0, 0, 
    0.01147146, 0.007619384, 0.008262599, 0.004988932, 0.001979945,
  -2.621971e-05, 0.002563008, -3.089339e-06, 0.03332051, 0.01391094, 
    0.001114864, 2.180279e-07, -7.229089e-08, -1.021048e-06, 1.730502e-05, 
    0.0009753486, 0.001092684, 0.0009600545, 0.002526685, 0.01373425, 
    0.01391367, 0.002894808, 0.0179247, 0.02768136, 0.03196002, 0.01016914, 
    0.000442899, 4.648263e-05, 0.0002080069, 0.01391038, 0.05959002, 
    0.03698164, 0.005631525, 0.0003456732,
  -1.529378e-07, 0.0008215687, 0.0001530648, 0.000183354, 0.002915262, 
    0.001013679, -5.705839e-05, 0.00390479, 0.005155385, -1.145868e-06, 
    2.061708e-05, -7.752325e-05, 0.002719153, 0.001005555, 0.01127263, 
    0.02094536, 0.0434719, 0.06463644, 0.01630232, 0.00124526, -3.874032e-06, 
    1.745196e-05, 0, 0.0002097196, 0.02006719, 0.01706612, 0.006850811, 
    0.0002827607, 2.369233e-05,
  6.278515e-07, 0.01591953, 0.007573706, 2.463802e-05, 0.002724591, 
    0.06184022, 0.02354475, 0.04794965, 0.01153884, 5.293382e-06, 
    0.008823534, 0.1053376, 0.06530705, 0.1001125, 0.118016, 0.0433066, 
    0.0233527, -1.462011e-05, 0.0003107634, 4.307121e-05, -7.836223e-11, 
    -3.445518e-07, 6.62649e-05, 0.1831019, 0.1464317, 0.005827029, 
    4.484472e-05, 0.0003819416, -6.013792e-08,
  0.001230956, 0.1211842, 0.06146486, 3.027567e-06, 1.965188e-05, 0.03801517, 
    0.001626778, 0.04293095, 0.08316033, 0.04150372, 0.01642272, 0.1435352, 
    0.1275716, 0.1633474, 0.04253066, 3.702967e-05, 0.001466079, 0.002194194, 
    -2.134434e-06, 0.003280119, 5.578944e-07, 3.132491e-05, 0.01466086, 
    0.1954238, 0.06444042, 0.004880091, 0.01034648, 0.001882012, -3.595506e-07,
  0.0006832267, 0.0005975274, 6.643196e-05, 0.005397429, 4.945528e-05, 
    9.37244e-05, 0.08250237, 0.1191896, 0.1619188, 0.1609967, 0.2140395, 
    0.2977297, 0.383536, 0.2893524, 0.2757449, 0.166429, 0.1425185, 
    0.1430862, 0.06273236, 0.06080307, 0.08691424, 0.1727715, 0.07252096, 
    0.0561573, 0.0247305, 0.02763109, 0.02831746, 0.01607505, 0.01187167,
  -3.398117e-06, -9.703623e-06, 0, 5.721472e-06, 1.156787e-05, 0.007331815, 
    0.03201385, 0.08476921, 0.02328992, 0.02027872, 0.07808596, 0.1337405, 
    0.104621, 0.08707678, 0.01651257, 0.006890617, 0.005785037, 0.03299888, 
    0.001599621, 0.00292872, 0.02688673, 0.0366501, 0.01295084, 0.0229665, 
    0.002526987, 0.01418539, 0.01874851, 0.0002000005, 0.0003325279,
  0, 2.133791e-05, -9.698734e-08, 0.001854889, 0.000387057, -5.899165e-06, 
    0.0001427918, 0.001576292, 0.01721112, 0.008986615, 0.0248005, 
    0.08756746, 0.06531031, 0.04171665, 0.03399604, 0.01276729, 0.005008708, 
    0.007098398, 0.01435112, 0.008042224, 0.003393605, 0.004404433, 
    0.008733448, 0.007420665, 0.02001116, 0.009443667, 0.006003642, 
    4.231702e-05, -7.614487e-09,
  0.006207169, 0.001205486, 0.0002404599, 0, -2.320012e-07, -1.699976e-09, 
    -1.462265e-10, 0, 0.0005587736, -7.062526e-06, 0.01013832, 0.05050517, 
    0.07107279, 0.08179131, 0.04537491, 0.04238484, 0.02769979, 0.02036673, 
    0.0005553722, -1.89128e-06, 0, 0.008371777, 0.01920612, 0.01665305, 
    0.02872313, 0.02751098, 0.01391923, 0.01056322, 0,
  0.001703194, 0.003538995, 1.411632e-05, 0.002391091, -2.423564e-05, 0, 
    -3.339028e-06, -1.095567e-05, 0, 0, 0, 0.003753743, 0.006273335, 
    0.005937079, 0.009636239, 0.008393339, 0.03317282, 0.02621272, 
    0.007937129, 0.0008640235, 0, 0.00197381, -9.714344e-05, 0.0007592402, 
    0.01006394, 0.02478284, 0.03741867, 0.006644859, 0.0002109177,
  0, -6.295982e-06, -1.010369e-05, -1.485599e-07, 0, -2.507141e-06, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, -4.01067e-05, 0.002443784, -1.51924e-06, 0.00554278, 
    -0.0001786413, -1.276993e-05, 0, 0.0009620053, -6.908282e-05, 
    0.002873757, 0.001297285, 0.0002847409, 0.002090659,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.186584e-05, 0, 0, 
    0.0002240103, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, -4.063961e-06, 0.000899803, 0, 0, 0, 0, 0, 0, 0, 
    0.0001032211, 0, 0, 0.0003976665, -2.402176e-06, -6.004021e-06, 0, 
    0.0003649367, 0, 0, 0, 0, 0, -3.028524e-05, 0,
  5.030815e-05, 0.001072877, 0.002304796, 0.00258256, 0.002412308, 
    0.004437753, 0.004101212, 0.005566693, 0.00155887, 0.0008596544, 0, 
    6.08687e-05, 0.0001687393, 0.004630296, -3.370001e-06, 0.0002907941, 
    0.001173348, -4.450117e-06, 0.000127136, 0.002838771, 0.0003712312, 
    -1.152684e-05, -2.419015e-05, -1.353771e-05, -1.708681e-05, 0.003573741, 
    0.004922308, 0.0007744752, 0.0008811677,
  0.01550535, 0.008009721, 0.00256367, 0.0114455, 0.02773922, 0.02300726, 
    0.008659371, 0.002467849, -1.630677e-05, 1.497341e-06, 0.0004381074, 
    0.003080457, 0.008644378, 0.009611437, 0.01701839, 0.007907673, 
    0.01948379, 0.002521483, 0.009361254, 0.02188001, 0.01549687, 0.00512048, 
    0.001109163, 0, 0.02228745, 0.01366329, 0.01961276, 0.01651723, 0.01040747,
  0.003936629, 0.01297056, 3.509758e-05, 0.06727348, 0.04034963, 0.003043, 
    0.0009789353, 0.0008034023, 0.001210499, 1.979653e-05, 0.01000384, 
    0.0112928, 0.002850895, 0.009335741, 0.02786676, 0.04080887, 0.02194435, 
    0.03701503, 0.07017451, 0.05502018, 0.02543319, 0.001328532, 0.000941517, 
    0.01017734, 0.02942114, 0.1062345, 0.1244766, 0.04344334, 0.0154666,
  0.0006412278, 0.03246412, 0.01609506, 0.02738946, 0.02145217, 0.04090898, 
    0.0006164839, 0.007946991, 0.01348657, -7.901629e-06, 6.236263e-05, 
    0.006642725, 0.002676864, 0.003931147, 0.02147423, 0.0702255, 0.1360946, 
    0.1883863, 0.1113223, 0.03819045, 0.009892965, 0.00354091, 2.304458e-06, 
    0.02339033, 0.1127404, 0.1243696, 0.08680934, 0.03594026, 0.01662488,
  -2.833896e-07, 0.03899279, 0.1331218, 0.01113741, 0.03492968, 0.1187537, 
    0.06576166, 0.0804287, 0.01275674, 0.0003284197, 0.01148751, 0.1102456, 
    0.05236468, 0.09170263, 0.1234926, 0.07272901, 0.07987982, 0.001505722, 
    0.0008815327, 2.540614e-05, 2.247488e-06, 1.912114e-05, 0.007307671, 
    0.4030812, 0.2728469, 0.05589889, 0.03739516, 0.003686606, 2.179771e-05,
  0.01392166, 0.3472348, 0.4251684, 0.0008253397, 0.0007176332, 0.06049721, 
    0.02282243, 0.07756808, 0.3586562, 0.2694866, 0.03129803, 0.1254774, 
    0.1334307, 0.1540626, 0.02791353, 8.064191e-05, 0.001072499, 0.005614454, 
    0.0001487909, 0.01056633, 6.644249e-05, 0.02379265, 0.0857641, 0.3491651, 
    0.09329665, 0.005899624, 0.02793767, 0.01867752, 0.0004524396,
  0.1093255, 0.04827451, 0.01005244, 0.009474053, -2.633766e-05, 0.000829668, 
    0.1785216, 0.1453187, 0.1757416, 0.1385816, 0.1890789, 0.2453545, 
    0.3358228, 0.2523044, 0.26619, 0.1946685, 0.1866772, 0.176442, 0.121828, 
    0.07917584, 0.1026245, 0.1779354, 0.2866401, 0.1790542, 0.09749845, 
    0.1651774, 0.2296865, 0.17367, 0.06941082,
  0.01416359, 0.004669729, 9.083949e-05, 0.0200898, 0.0007541479, 0.02087273, 
    0.07542109, 0.09222442, 0.05380331, 0.016067, 0.0606368, 0.1052517, 
    0.08238579, 0.08349612, 0.03318175, 0.07121591, 0.07213135, 0.1196525, 
    0.0370916, 0.02090907, 0.1118875, 0.04661491, 0.06583171, 0.06896348, 
    0.1007614, 0.06778247, 0.08652478, 0.1914741, 0.05883055,
  -2.410994e-05, 0.0007688774, -1.632934e-05, 0.002535636, 0.001223102, 
    -1.528113e-05, 0.0005516037, 0.0049357, 0.0239062, 0.03952305, 0.0372447, 
    0.1179101, 0.09283224, 0.05793754, 0.06626004, 0.1030192, 0.07930338, 
    0.04786014, 0.028682, 0.0223855, 0.005066718, 0.04487474, 0.0265445, 
    0.1096222, 0.186437, 0.09134842, 0.02642979, 0.00251875, 0.0002340828,
  0.01294792, 0.005643702, 0.000912227, -2.004221e-06, 4.654864e-05, 
    0.0003155943, -1.523725e-05, 0, 0.000732267, -3.259e-05, 0.02099226, 
    0.08733545, 0.1265114, 0.156065, 0.1042273, 0.09637229, 0.08390769, 
    0.04914806, 0.01058913, 4.389524e-05, 2.936121e-07, 0.01261108, 
    0.02723951, 0.03319366, 0.1049438, 0.07215626, 0.02852938, 0.02086652, 
    0.001100221,
  0.00428455, 0.007284196, 2.460332e-06, 0.004680074, 0.0001786902, 
    0.0008648061, 0.0009472526, -5.754639e-05, -8.345797e-06, 0, 
    -2.409515e-06, 0.008131159, 0.0184576, 0.02874054, 0.01325321, 
    0.02054501, 0.05580305, 0.07190052, 0.01996825, 0.004275694, 
    -5.071379e-07, 0.007362557, 0.001843741, 0.007427091, 0.01806769, 
    0.05313422, 0.08417606, 0.01891158, 0.0103422,
  2.207265e-05, 4.662869e-05, 0.0001144195, -2.160657e-05, 0, 6.876948e-05, 
    8.258887e-05, 0, 0, 0, 0, 0, 0, 0, 0, -3.04422e-06, 0.0003568678, 
    0.01833929, 0.002696841, 0.009653419, 0.0005936695, 2.831532e-05, 
    -3.95343e-11, 0.003833153, 0.002150017, 0.01417591, 0.01154439, 
    0.006170629, 0.004631697,
  -1.284153e-06, 0, 0, -1.551768e-05, -4.410357e-06, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 3.602067e-06, 0.000126858, -1.480907e-05, -5.672806e-06, 
    0.0007107056, 0.0002160901, -3.90655e-08, 0, 0, 0, -5.549738e-07, 
    0.0007170304, -5.003146e-05,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.000364002, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 9.200961e-06, 0, 0, 0, 0,
  5.633891e-05, 0, 0, 0, 0, -1.60194e-05, 0.001877462, 0, -7.045816e-09, 0, 
    0, 0, -2.458845e-05, 1.27619e-06, 0.001475836, 7.429726e-05, 
    0.0002964593, 0.00208132, -1.333375e-05, -3.996321e-05, 0, 0.0007393469, 
    0, 0, 0, 0, -6.443126e-06, 0.0006514578, 7.120292e-07,
  0.002237518, 0.004693265, 0.005063551, 0.01227282, 0.007516158, 0.01326849, 
    0.01247687, 0.01917442, 0.01132426, 0.009126987, 0.004189424, 
    0.001898415, 0.0001893476, 0.01120888, 0.00112159, 0.00201621, 
    0.007069443, 0.004312919, 0.001552759, 0.007707221, 0.0066078, 
    0.001832688, 0.002917895, 0.001619688, 0.001670695, 0.007272591, 
    0.014235, 0.01034546, 0.0090123,
  0.03309784, 0.02182792, 0.03124558, 0.03327956, 0.06408882, 0.08899359, 
    0.03128717, 0.01686015, 0.008230306, 0.001283836, 0.006435565, 
    0.005562998, 0.01500355, 0.0173048, 0.04178567, 0.01953418, 0.03801515, 
    0.01752369, 0.02324824, 0.04093188, 0.02651289, 0.02343047, 0.002898566, 
    0.0002200715, 0.036855, 0.04738665, 0.05725595, 0.03120688, 0.02779029,
  0.09048157, 0.06389881, 0.01569997, 0.114943, 0.1043376, 0.07584538, 
    0.01604614, 0.02099757, 0.01454185, 0.01105138, 0.01804132, 0.02915784, 
    0.01229196, 0.04364606, 0.05162429, 0.07836543, 0.05749456, 0.09071964, 
    0.2170498, 0.169252, 0.1264632, 0.06646497, 0.03831585, 0.05859362, 
    0.04593851, 0.125458, 0.1660029, 0.1333198, 0.09162037,
  0.001544292, 0.03309895, 0.08929218, 0.02214035, 0.05356929, 0.02773688, 
    0.003245483, 0.001821392, 0.01494701, 1.135507e-05, 0.003285636, 
    0.008731426, 0.0004139068, 0.006896495, 0.03485508, 0.07392445, 
    0.1489817, 0.1928009, 0.1230459, 0.05518744, 0.02501395, 0.008884481, 
    5.446584e-07, 0.01999173, 0.07861809, 0.1547039, 0.07779819, 0.0296032, 
    0.01482487,
  -2.887023e-08, 0.02450342, 0.07594776, 0.006396041, 0.02795165, 0.0859483, 
    0.04431394, 0.06790708, 0.01186191, 0.0002092923, 0.005440117, 
    0.08625993, 0.04740297, 0.06735224, 0.0966579, 0.05330025, 0.05987779, 
    0.002241629, 0.0007416455, 1.942832e-06, 3.72013e-07, 5.049798e-07, 
    0.0006072991, 0.3317638, 0.2335369, 0.04308468, 0.03482671, 0.0009215974, 
    2.666564e-06,
  0.003649265, 0.299793, 0.3587213, 0.0001901065, 0.0002287152, 0.05178465, 
    0.009413807, 0.05593866, 0.2687556, 0.1889361, 0.01947453, 0.1007451, 
    0.085466, 0.1196598, 0.01751532, 0.000485325, 6.139101e-05, 0.002616051, 
    0.001837331, 0.003350534, 7.824984e-06, 0.00324053, 0.03999268, 
    0.3241906, 0.05897148, 0.0006342274, 0.0241949, 0.008226883, 1.564541e-05,
  0.06616317, 0.02208504, 0.00361193, 0.05294767, 0.0001730552, 6.576194e-05, 
    0.1235702, 0.1046903, 0.154945, 0.1051721, 0.1512032, 0.2130136, 
    0.288219, 0.2296462, 0.2136073, 0.1442649, 0.1526583, 0.1473414, 
    0.08764294, 0.06970096, 0.07678059, 0.1169258, 0.2209334, 0.1451389, 
    0.06083731, 0.1337615, 0.1643275, 0.1234867, 0.05496965,
  0.04105131, 0.005744276, 0.0005006809, 0.02346216, 0.002360587, 0.01065401, 
    0.06968486, 0.07439488, 0.05486221, 0.01706825, 0.0520368, 0.09784693, 
    0.06792079, 0.06627429, 0.01388331, 0.04259555, 0.06620186, 0.1029862, 
    0.03713115, 0.01965649, 0.09684603, 0.03588059, 0.04844017, 0.04119535, 
    0.06031039, 0.05875932, 0.07952167, 0.2281883, 0.1193749,
  0.0531614, 0.03695349, 0.02492085, 0.01599828, 0.01502021, 0.0121204, 
    0.02299235, 0.009284348, 0.03456596, 0.0616952, 0.04115288, 0.09481727, 
    0.08862618, 0.03643868, 0.04902861, 0.1021161, 0.1045697, 0.08477923, 
    0.07513522, 0.05148679, 0.0271264, 0.08332199, 0.07117557, 0.1307447, 
    0.1764518, 0.1068432, 0.06931734, 0.05508028, 0.05807689,
  0.05103247, 0.02342503, 0.01459945, -5.831602e-06, 0.004195211, 0.00263124, 
    0.0004187462, 2.267251e-05, 0.007703282, 0.004734347, 0.05972418, 
    0.1384773, 0.1897233, 0.1984012, 0.1629985, 0.1551089, 0.1327937, 
    0.1739428, 0.08916169, 0.006496173, 0.0003872624, 0.01871832, 0.03823446, 
    0.05820377, 0.1653342, 0.1987192, 0.1146556, 0.04564642, 0.02412944,
  0.03821596, 0.02143144, 0.001675434, 0.00757539, 0.001140029, 0.001715425, 
    0.002070244, 0.0008540981, -2.469779e-05, 0, -5.053047e-05, 0.0190391, 
    0.02461045, 0.03284949, 0.0414915, 0.05389024, 0.1108698, 0.2091547, 
    0.1436293, 0.01128204, 0.0005920288, 0.01186083, 0.01492423, 0.02443153, 
    0.03866365, 0.1296461, 0.1719823, 0.0998301, 0.06437265,
  0.009201044, 0.002789212, 0.006599235, 0.0008482831, 0, 9.508431e-05, 
    0.001027302, 0, 0, 0, 0, 0, 0, -3.057831e-08, -9.08458e-05, 0.005571076, 
    0.00344522, 0.07200141, 0.01048152, 0.02356016, 0.009054961, 0.005309372, 
    -2.124024e-05, 0.007025933, 0.01293589, 0.03857755, 0.0395714, 
    0.03946466, 0.02818361,
  0.001716723, 1.674191e-05, -2.946844e-05, 8.288303e-06, 0.0004818568, 
    -1.314618e-07, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0001231476, 0.002102316, 
    0.007377657, 0.005597366, 0.005255106, 0.003365029, 0.000136974, 
    0.0008499136, -6.464757e-06, -2.153822e-06, 5.145704e-07, 0.003088419, 
    0.002084573,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -9.743156e-06, 0, 0, 0.001001579, 0, 0, 0, 
    0, 0, -6.817824e-06, 0, 0, 0, 0.0001795695, 3.472001e-05, 0, 0, 0,
  0.002409837, -2.47343e-05, -6.39478e-07, 8.189474e-07, 0, 6.724709e-06, 
    0.004047994, 0.0009384911, 0.00115549, 0.0007261638, 0.0001542831, 
    0.001203743, 0.0005890511, 0.0007986546, 0.00381758, 0.001760517, 
    0.003000717, 0.005827031, -4.478046e-05, 0.001288969, 0.0002035977, 
    0.001627184, -3.851815e-05, 1.456501e-05, -2.064935e-06, 0, 
    -2.909965e-05, 0.003485499, 0.005571091,
  0.02979923, 0.02965134, 0.02636275, 0.03829634, 0.04521342, 0.05284122, 
    0.06168917, 0.1063662, 0.08764149, 0.06861433, 0.02565547, 0.0187523, 
    0.01804993, 0.04266204, 0.02610852, 0.01673717, 0.03204195, 0.04589244, 
    0.03643732, 0.03485925, 0.02293788, 0.006390108, 0.01400221, 0.007879547, 
    0.002857307, 0.01848669, 0.04814336, 0.05717997, 0.03395903,
  0.07763636, 0.08358098, 0.0851552, 0.0960573, 0.1188778, 0.1349907, 
    0.1045499, 0.1174054, 0.07636917, 0.04946974, 0.04455872, 0.03523196, 
    0.04127382, 0.06178769, 0.07248679, 0.116261, 0.127996, 0.08796805, 
    0.1323873, 0.1075495, 0.100504, 0.08831014, 0.03541618, 0.004973587, 
    0.07883294, 0.07745832, 0.1028921, 0.09421359, 0.06716291,
  0.1010932, 0.04525216, 0.09875518, 0.102081, 0.1044906, 0.06891751, 
    0.006632704, 0.01698722, 0.01841987, 0.01299533, 0.02968075, 0.05497143, 
    0.05612318, 0.09537838, 0.1092935, 0.1143432, 0.09309776, 0.1145761, 
    0.2303744, 0.1873977, 0.1381528, 0.08451434, 0.03571624, 0.04810404, 
    0.04348208, 0.1046204, 0.1604467, 0.1386318, 0.1252933,
  -2.819933e-05, 0.02024586, 0.07495268, 0.007140109, 0.03582766, 0.02468036, 
    -0.0001949797, 0.000366825, 0.01994104, 0.0009957789, 0.004481136, 
    0.009135087, 0.001722763, 0.01574707, 0.04816189, 0.09231979, 0.1611368, 
    0.1707689, 0.06325523, 0.0381263, 0.007402705, 0.002802787, 
    -8.838763e-08, 0.01854662, 0.05992924, 0.1476044, 0.06462942, 0.02499079, 
    0.01724954,
  -4.395143e-06, 0.01976515, 0.04570639, 0.003611638, 0.02341863, 0.06742768, 
    0.03503321, 0.06070086, 0.01592279, 0.0007025989, 0.006003645, 
    0.06772205, 0.04988299, 0.06382641, 0.0827827, 0.04818111, 0.05447699, 
    0.002173363, 0.000299267, 3.034139e-07, 1.209635e-07, 2.132556e-07, 
    2.324619e-05, 0.2785556, 0.226523, 0.04280861, 0.0162974, 0.0002349016, 
    8.946158e-07,
  0.002573145, 0.2728358, 0.2954874, 9.522375e-05, 6.413017e-05, 0.05210233, 
    0.008722451, 0.05581237, 0.2107554, 0.1419976, 0.01095992, 0.07590418, 
    0.06852559, 0.1071356, 0.01683355, 0.0001992146, 1.703015e-05, 
    7.144007e-05, 3.421725e-05, 3.085147e-05, 1.305044e-06, 4.972743e-05, 
    0.01780099, 0.2865924, 0.04278096, -1.70126e-05, 0.02150702, 0.008116825, 
    2.200132e-06,
  0.04928783, 0.01470244, 0.004468389, 0.04150973, 9.868767e-05, 
    0.0003734801, 0.1064958, 0.09490965, 0.1403031, 0.0915748, 0.1091369, 
    0.1928499, 0.2503469, 0.2308624, 0.184002, 0.1141048, 0.1441108, 
    0.1401245, 0.07952822, 0.06608456, 0.07063085, 0.09627756, 0.1788857, 
    0.1269782, 0.04505386, 0.1129129, 0.1269478, 0.08803269, 0.04841799,
  0.0362216, 0.007545142, 5.635138e-06, 0.0262376, 0.001287699, 0.008605252, 
    0.06488702, 0.06711389, 0.04964345, 0.01631971, 0.05058723, 0.08997676, 
    0.0676418, 0.0575329, 0.01143483, 0.03860242, 0.05270751, 0.06972077, 
    0.02330972, 0.02108246, 0.08655638, 0.03230614, 0.0378885, 0.03139865, 
    0.03929128, 0.04925377, 0.06300785, 0.1782807, 0.08648872,
  0.0808717, 0.04921416, 0.02318764, 0.02632419, 0.03608396, 0.02462489, 
    0.02390363, 0.01447139, 0.05777756, 0.07962463, 0.04250328, 0.08109162, 
    0.08556825, 0.02037128, 0.04496285, 0.08674532, 0.08233485, 0.08324189, 
    0.07080778, 0.04860266, 0.05377916, 0.0671332, 0.05871623, 0.1118972, 
    0.1423101, 0.08630008, 0.0534261, 0.04360019, 0.08612752,
  0.1339253, 0.09310883, 0.06421888, 0.006312137, 0.03050211, 0.04063024, 
    0.001541246, 0.0007187467, 0.02249826, 0.03414302, 0.1057427, 0.163203, 
    0.215321, 0.1982157, 0.1723445, 0.1845492, 0.16847, 0.2535031, 
    0.08838177, 0.02760636, 0.001865539, 0.07276872, 0.08735485, 0.08431563, 
    0.1699789, 0.1903476, 0.107519, 0.06603436, 0.08114626,
  0.1063808, 0.076161, 0.03364468, 0.05713664, 0.04990489, 0.01957841, 
    0.004983781, 0.002569522, 5.373098e-05, -1.429436e-05, 0.006475342, 
    0.03856074, 0.04805294, 0.05361561, 0.05893889, 0.1150361, 0.1424064, 
    0.3053067, 0.2260851, 0.04391451, 0.03494763, 0.06734157, 0.04794155, 
    0.05193968, 0.09349209, 0.1853329, 0.2245691, 0.1631879, 0.1064866,
  0.05670385, 0.02458332, 0.02449545, 0.01541206, 0.001330037, 0.007500576, 
    0.007846167, 0.001842491, -4.66755e-06, -1.962829e-05, -2.10624e-05, 0, 
    -0.0002354006, -5.907584e-05, 0.004579232, 0.02916476, 0.02366293, 
    0.1642881, 0.05535606, 0.04829983, 0.03390352, 0.04615765, 0.01037214, 
    0.01744589, 0.03433712, 0.06248378, 0.07503862, 0.05773107, 0.07782175,
  0.005618167, 0.005690969, 0.001550258, 0.001994347, 0.0008473312, 
    6.058964e-06, 0, -1.954302e-05, 0, 0, 0, 0, 0, 0, 0, -1.025827e-06, 
    0.003959908, 0.0193619, 0.04583798, 0.07421339, 0.0494587, 0.01843406, 
    0.006692438, 0.003092613, 0.001097805, -2.348266e-05, -3.518498e-07, 
    0.01600343, 0.01074474,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -3.085137e-07, 
    4.568968e-05, -3.533238e-07, 0, 1.284779e-07, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0.0004851418, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.709254e-06, -1.948631e-05, 0, 
    0.0003687477, 0.002077334, 0, -1.087221e-05, -0.0001041136, 4.270171e-06, 
    0, 0.001035867, 1.83007e-05, 1.247701e-06, 0.0003943875, 0.004847368, 
    7.496507e-05, -1.938019e-06, 9.985472e-06, 0.000444833,
  0.04399145, 0.01592107, 0.007917561, 0.0001064303, -1.790403e-05, 
    0.004691415, 0.008007935, 0.008444128, 0.01106714, 0.0104595, 0.01588958, 
    0.01738505, 0.01175292, 0.01609535, 0.03073845, 0.02017303, 0.02840153, 
    0.04839205, 0.04891899, 0.04505339, 0.01855123, 0.02337328, 0.02049667, 
    0.01017138, 0.006088872, 0.009352544, 0.01114811, 0.03783197, 0.05120116,
  0.08070243, 0.08032085, 0.09435864, 0.1276989, 0.1118745, 0.1207033, 
    0.1166185, 0.1764893, 0.1644748, 0.124661, 0.09533124, 0.09131712, 
    0.07472373, 0.1069772, 0.08347633, 0.1523659, 0.1444616, 0.1192278, 
    0.1069593, 0.120694, 0.09242044, 0.0785906, 0.05658136, 0.01880573, 
    0.03737152, 0.101992, 0.1514218, 0.1528969, 0.1070459,
  0.1439798, 0.1129593, 0.09557906, 0.1054654, 0.1123342, 0.1187479, 
    0.1087863, 0.1309965, 0.09321143, 0.08856881, 0.08233681, 0.05375268, 
    0.09360939, 0.123021, 0.1305484, 0.135887, 0.1726098, 0.1556118, 
    0.1445194, 0.112084, 0.1061783, 0.1163907, 0.07842462, 0.02501382, 
    0.1218028, 0.115667, 0.1505126, 0.1120241, 0.1002919,
  0.0819348, 0.03274909, 0.07906559, 0.09187286, 0.08612038, 0.04993722, 
    0.008486639, 0.009554821, 0.01593455, 0.02235781, 0.02571018, 0.0516852, 
    0.07285358, 0.08875876, 0.1119787, 0.07552611, 0.07875787, 0.0919714, 
    0.2165014, 0.1707964, 0.132726, 0.06078143, 0.03764364, 0.01942259, 
    0.03487583, 0.08703633, 0.1391841, 0.1122655, 0.1301221,
  7.475532e-05, 0.008842049, 0.05374099, 0.001386596, 0.01533247, 0.02276512, 
    -7.765141e-05, -0.0006977628, 0.01992421, 0.0067963, 0.00270597, 
    0.007883623, 0.007107515, 0.01252656, 0.05926374, 0.08926924, 0.1588838, 
    0.1418834, 0.04499558, 0.0291359, 0.002056989, 0.001637561, 
    -4.703423e-09, 0.00829391, 0.04897447, 0.144873, 0.06408116, 0.02535863, 
    0.02263454,
  0.001207618, 0.01969173, 0.03560213, 0.002008084, 0.02624123, 0.05190317, 
    0.03825157, 0.0546174, 0.02127262, 0.0006915246, 0.00920191, 0.05773562, 
    0.05208281, 0.06506444, 0.06492948, 0.05109401, 0.04833087, 0.0005198442, 
    0.0009700835, 5.685667e-08, 6.54373e-09, 9.480976e-08, 6.562695e-06, 
    0.2107561, 0.185316, 0.04533163, 0.001238452, 0.0001255932, 1.365552e-07,
  0.007433592, 0.2385451, 0.2018438, 0.0001123884, 5.135576e-05, 0.05080659, 
    0.01159003, 0.05721066, 0.1504656, 0.08862876, 0.01018958, 0.05629439, 
    0.05856994, 0.08541023, 0.01901178, 5.46547e-05, -3.695541e-05, 
    -4.973438e-05, 4.276738e-06, -3.866091e-06, 1.043974e-06, 7.752282e-06, 
    0.006594693, 0.2200305, 0.02703574, -6.171624e-07, 0.02526194, 0.0138834, 
    -7.844326e-06,
  0.03739507, 0.01350083, 0.005948562, 0.02783543, 0.0002510039, 0.000876171, 
    0.08998476, 0.08677982, 0.1257502, 0.0787297, 0.08544753, 0.1769278, 
    0.2158998, 0.2191619, 0.1479733, 0.08564592, 0.1525096, 0.1519585, 
    0.07207341, 0.05816989, 0.0611283, 0.07307909, 0.1391578, 0.09057765, 
    0.03853823, 0.1104395, 0.09830783, 0.05627447, 0.04408786,
  0.02943446, 0.005321456, 9.875619e-06, 0.02600264, 0.0007141524, 
    0.007797293, 0.05600659, 0.05989166, 0.05505966, 0.01691874, 0.05008891, 
    0.08226786, 0.05768353, 0.04891231, 0.009148113, 0.03061827, 0.03564208, 
    0.03942065, 0.01592808, 0.01903268, 0.07167883, 0.0299273, 0.03068411, 
    0.02627804, 0.027143, 0.04556566, 0.06034391, 0.1408807, 0.05131878,
  0.07894991, 0.04945254, 0.02612846, 0.02756258, 0.0283737, 0.01875334, 
    0.01912886, 0.01752359, 0.08670384, 0.1041691, 0.04534846, 0.07925394, 
    0.07128701, 0.01935976, 0.02727706, 0.08184202, 0.07068987, 0.06791022, 
    0.04747729, 0.04586696, 0.05127317, 0.0475599, 0.04733147, 0.09193801, 
    0.1183274, 0.06414917, 0.0446022, 0.03248938, 0.05666658,
  0.1843401, 0.1038606, 0.06236068, 0.02976742, 0.07318806, 0.07569297, 
    0.005816364, 0.0638012, 0.0821889, 0.07215781, 0.1230104, 0.1602345, 
    0.2264044, 0.1937914, 0.1744538, 0.1801606, 0.1906075, 0.2441113, 
    0.07619052, 0.03419926, 0.04261102, 0.09703781, 0.1189504, 0.08944325, 
    0.1627678, 0.1625181, 0.09884425, 0.06661423, 0.1012052,
  0.1377053, 0.1432005, 0.07225762, 0.1020314, 0.1288815, 0.09309236, 
    0.04930274, 0.004991812, 0.0004202401, 0.0008431406, 0.02141088, 
    0.06453815, 0.08485276, 0.06743915, 0.1035935, 0.1639402, 0.1565599, 
    0.3272327, 0.2446479, 0.0973822, 0.07302056, 0.1329317, 0.09188311, 
    0.130169, 0.1300421, 0.1835757, 0.2207499, 0.1457772, 0.1121646,
  0.1318286, 0.1016102, 0.1043638, 0.1118825, 0.08116701, 0.06378441, 
    0.07494362, 0.03506009, 0.007304186, 0.003503991, -2.312523e-05, 0, 
    0.00240084, 0.01232001, 0.02023258, 0.0793514, 0.06543529, 0.214415, 
    0.1213524, 0.08989433, 0.08689168, 0.09115344, 0.0302353, 0.04522933, 
    0.09918, 0.1319334, 0.1416719, 0.1066892, 0.1263573,
  0.04853741, 0.05318019, 0.01958566, 0.03679504, 0.02260027, 0.006953363, 
    0.006454898, 8.732014e-05, -8.176411e-08, 2.676562e-05, 5.305963e-08, 0, 
    0, 0, 7.035013e-08, 0.004249482, 0.04156528, 0.09313289, 0.1190911, 
    0.1270988, 0.08757336, 0.06817846, 0.0322901, 0.008454245, 0.02111886, 
    0.0001810816, -0.0001700235, 0.07071649, 0.04121074,
  -9.78004e-06, 0, -4.415453e-05, 0.0001256374, 0.0002579094, -1.585798e-05, 
    6.355207e-07, 0, -7.350799e-07, 4.630098e-07, 0, 0, 0, 2.848698e-06, 
    -7.283379e-05, 0.006449352, 0.0226203, 0.02332761, 0.009804692, 
    0.002558922, 0.0001636027, 0.0008741086, 7.423724e-05, -1.106498e-05, 
    -3.925865e-09, 0, 0, -2.500277e-05, 5.80745e-06,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2.20213e-05, 
    0.0001182304, 0, 0, 0, 0, 9.540206e-05, 0.001868639, -8.439854e-05, 
    8.365813e-05, 0, 0,
  0.03176903, 0.01196651, 0, 0, 0, 0, 0, 0, 0, 0, -1.709254e-06, 
    4.859055e-05, -5.672664e-06, 0.0009777094, 0.004406703, -0.0003873311, 
    0.006671892, 0.005355752, 0.0001172356, 0.0001713806, 0.007784367, 
    0.0201517, 0.01769936, 0.01194923, 0.02394841, 0.006408927, 0.003069827, 
    0.01480012, 0.01780829,
  0.113218, 0.1036023, 0.0862269, 0.0396386, 0.01685612, 0.02890099, 
    0.05134975, 0.04988277, 0.06825958, 0.07291826, 0.06818961, 0.06770791, 
    0.06603053, 0.07721733, 0.08518723, 0.0810913, 0.07714127, 0.1707425, 
    0.1451787, 0.1290621, 0.09072602, 0.08466761, 0.0537687, 0.06620716, 
    0.05229725, 0.04817162, 0.07680984, 0.1041815, 0.1184487,
  0.1305068, 0.1222558, 0.1334887, 0.166778, 0.1554572, 0.1549972, 0.1517904, 
    0.1884398, 0.2022911, 0.1605172, 0.1325763, 0.0998469, 0.1101977, 
    0.1263307, 0.1258137, 0.1903114, 0.1678893, 0.1403187, 0.1433031, 
    0.1756559, 0.1607161, 0.1424813, 0.1369597, 0.06080198, 0.09325497, 
    0.2063993, 0.2422206, 0.203439, 0.1510727,
  0.1376372, 0.1104102, 0.09057535, 0.1031312, 0.10627, 0.105533, 0.1056681, 
    0.1094808, 0.09181202, 0.08771136, 0.07393047, 0.05321626, 0.09921204, 
    0.1220864, 0.1439079, 0.1262522, 0.1564688, 0.1350212, 0.1315939, 
    0.10058, 0.0932088, 0.1103985, 0.08820062, 0.04383709, 0.1179197, 
    0.1120828, 0.1490417, 0.1024158, 0.1015248,
  0.07014412, 0.02745476, 0.05448239, 0.08581751, 0.07364552, 0.0428878, 
    0.0061802, 0.002429807, 0.01124373, 0.00516721, 0.02120289, 0.04804469, 
    0.08584425, 0.08489692, 0.09179833, 0.06315535, 0.07207779, 0.08403251, 
    0.212493, 0.1526876, 0.1079802, 0.04129016, 0.02499085, 0.007903145, 
    0.03615748, 0.07982349, 0.1158498, 0.08928191, 0.1373211,
  0.001522377, 0.004961534, 0.03056856, 0.0005432811, 0.008761775, 0.0167695, 
    0.0006811984, -0.0005564437, 0.02953574, 0.004852, 0.004125427, 
    0.006200265, 0.01100239, 0.007613712, 0.058685, 0.09508246, 0.1597228, 
    0.1278723, 0.03557088, 0.01916289, 0.001671238, 0.0001019273, 
    -1.248388e-09, 0.003937393, 0.03796501, 0.1286941, 0.06136604, 
    0.02434488, 0.0169176,
  0.002790274, 0.02266653, 0.02445537, 0.002699045, 0.02363614, 0.04811995, 
    0.04371073, 0.04741279, 0.01897988, 0.0004471635, 0.01246331, 0.04438407, 
    0.05226718, 0.06110599, 0.04541238, 0.06072564, 0.04165003, 0.0008127395, 
    0.0001441937, 2.56888e-08, 2.577978e-09, 6.220499e-08, 1.33536e-05, 
    0.1499162, 0.1386797, 0.03783925, 0.0003445968, 8.036946e-06, 2.57204e-08,
  0.01563828, 0.2303278, 0.1354863, 0.0007692671, 0.0002347239, 0.04978622, 
    0.0148658, 0.0611529, 0.1072297, 0.06558749, 0.008029627, 0.03427335, 
    0.04256614, 0.06240477, 0.01241458, 0.0001599849, 0.0005869925, 
    0.0001107688, 9.488333e-06, 1.069892e-06, 2.978608e-07, 3.708743e-06, 
    0.000361906, 0.1545624, 0.0186641, 0.0001311485, 0.02389356, 0.009354866, 
    -2.445154e-06,
  0.03112901, 0.01402098, 0.007544869, 0.023501, 0.0003813084, 0.001217574, 
    0.06582411, 0.06948857, 0.11106, 0.06702951, 0.06353845, 0.1554637, 
    0.1799821, 0.2206222, 0.1244794, 0.06545127, 0.1531875, 0.1511237, 
    0.06592861, 0.05279509, 0.05808702, 0.05853025, 0.1162156, 0.05763008, 
    0.04123875, 0.1058214, 0.08314043, 0.0331107, 0.03782573,
  0.01945182, 0.002494817, -1.710231e-05, 0.02002862, 0.0002767967, 
    0.009762138, 0.0449047, 0.05122381, 0.04616383, 0.0169608, 0.04605927, 
    0.07513436, 0.05295989, 0.04032128, 0.008109052, 0.01997572, 0.02141391, 
    0.03377607, 0.01995499, 0.01845109, 0.05327774, 0.02637986, 0.02032125, 
    0.01743509, 0.0166121, 0.0372017, 0.05967295, 0.1139897, 0.03224518,
  0.07488328, 0.04300811, 0.01961602, 0.01428562, 0.02101569, 0.0143567, 
    0.01379203, 0.02218501, 0.1323628, 0.09707999, 0.04951, 0.07014555, 
    0.07067423, 0.01982942, 0.02273423, 0.06717482, 0.05846973, 0.05642818, 
    0.03540993, 0.03259953, 0.04392186, 0.03744579, 0.04703561, 0.07620743, 
    0.09872124, 0.06302632, 0.04247891, 0.02511288, 0.03986344,
  0.1686151, 0.09929121, 0.0490386, 0.03950902, 0.05931704, 0.06566299, 
    0.01359073, 0.09227419, 0.1052879, 0.1004366, 0.113415, 0.1482116, 
    0.21726, 0.1896461, 0.1854081, 0.1766601, 0.1759051, 0.2215541, 
    0.06431414, 0.03060922, 0.06950906, 0.0964777, 0.122232, 0.08701743, 
    0.1462026, 0.1443517, 0.1047865, 0.05866623, 0.08098798,
  0.1253848, 0.1606252, 0.1297868, 0.1064076, 0.1327034, 0.1227555, 0.121682, 
    0.0173942, 0.009337173, 0.02568262, 0.1145042, 0.102673, 0.1269088, 
    0.09225328, 0.1628096, 0.2222821, 0.1580547, 0.3205216, 0.2341891, 
    0.1076117, 0.1058121, 0.1389416, 0.1350768, 0.1833537, 0.142, 0.160775, 
    0.2227354, 0.14995, 0.1130708,
  0.1955068, 0.1949681, 0.1708477, 0.2192926, 0.1894635, 0.1640296, 
    0.1898096, 0.1262814, 0.08497065, 0.03361988, 0.02379381, -1.606415e-06, 
    0.006869257, 0.03544988, 0.0384858, 0.1374882, 0.1261084, 0.2527974, 
    0.1697521, 0.09688029, 0.1272543, 0.09415627, 0.07654122, 0.09981903, 
    0.1437661, 0.1810966, 0.161909, 0.1160307, 0.1856491,
  0.1595506, 0.1545401, 0.1043021, 0.1147239, 0.126082, 0.09254099, 
    0.05695505, 0.03983413, 0.01298799, 0.004963906, 0.005420957, 
    0.002023453, 0.004733123, 0.00500326, 0.02090656, 0.08778632, 0.1281708, 
    0.1547426, 0.1604611, 0.1623012, 0.1111104, 0.0943986, 0.09909413, 
    0.04358386, 0.0802412, 0.005351164, 0.0004116567, 0.1771769, 0.1427775,
  0.004003334, 0.004512526, 0.003705736, 0.0124477, 0.01452174, 0.01919238, 
    0.01750515, 0.01236522, 0.009722157, 0.02257449, -0.0006842143, 
    8.500915e-05, 0.002446698, 0.006544804, 0.01984045, 0.05435082, 
    0.07389166, 0.06471477, 0.04530787, 0.02233136, 0.01586363, 0.01399171, 
    0.004747127, -0.0004476751, 8.922879e-05, -6.947112e-06, 0, 0.000229381, 
    0.001179287,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.000189998, -7.024922e-05, 
    0.001441283, -6.350787e-06, 0, 0, 5.275572e-05, 0.0008657373, 0.00350654, 
    0.001868157, 0.01846574, 0.01283306, 0,
  0.06455927, 0.02411174, 0.005057172, 0.0003189824, -2.246036e-05, 
    -1.012712e-05, -0.000206296, -1.905034e-05, -5.906798e-05, 0, 
    0.0001323459, 0.0001170469, -0.0004815694, 0.01055534, 0.01508964, 
    0.01437925, 0.03538349, 0.03461446, 0.0216519, 0.01661908, 0.02700522, 
    0.0448494, 0.05369063, 0.05339889, 0.05094628, 0.08316499, 0.1056567, 
    0.08389779, 0.07642811,
  0.2215076, 0.1755783, 0.186765, 0.134241, 0.09603125, 0.1071195, 0.1077911, 
    0.1066406, 0.1316457, 0.1267747, 0.1221404, 0.1402985, 0.1198401, 
    0.1463286, 0.1325171, 0.1238088, 0.1395855, 0.2258581, 0.1933549, 
    0.1912253, 0.1646114, 0.1539432, 0.1358597, 0.179639, 0.1752053, 
    0.1593915, 0.1618134, 0.2047225, 0.2207821,
  0.1294937, 0.108522, 0.1515977, 0.1850603, 0.1608402, 0.1520339, 0.1685844, 
    0.1910627, 0.2136211, 0.1683187, 0.1631219, 0.1143486, 0.1245196, 
    0.1543427, 0.1388513, 0.1667489, 0.1506685, 0.1347132, 0.1475566, 
    0.1832772, 0.1729303, 0.1546178, 0.1656235, 0.1110597, 0.1325019, 
    0.2052358, 0.2353838, 0.2057003, 0.1642095,
  0.130915, 0.1134986, 0.08149856, 0.101257, 0.1076325, 0.1021162, 0.1044547, 
    0.09902441, 0.07875814, 0.07568087, 0.04564175, 0.05059116, 0.09448158, 
    0.1156094, 0.1387441, 0.1166964, 0.1426017, 0.1247994, 0.1235086, 
    0.08666242, 0.07994971, 0.09993237, 0.0933209, 0.05637548, 0.1094085, 
    0.105227, 0.1440273, 0.1022424, 0.0951338,
  0.05651741, 0.01655113, 0.05779904, 0.08670916, 0.06505962, 0.04984232, 
    0.008883875, 0.005807833, 0.007863711, 4.263681e-05, 0.01372915, 
    0.0547361, 0.08944093, 0.07951866, 0.09881167, 0.05773523, 0.08140527, 
    0.08217829, 0.2126892, 0.1341864, 0.08893049, 0.02390347, 0.009582639, 
    0.004330509, 0.0393443, 0.07301112, 0.1086516, 0.07756012, 0.1188417,
  0.0006721928, 0.004453761, 0.02468812, 0.0004996384, 0.0117584, 0.01380411, 
    0.0001217754, -0.0004230459, 0.01591145, 0.007495579, 0.002470825, 
    0.005566051, 0.02029666, 0.01353118, 0.05323248, 0.09457058, 0.1673776, 
    0.1091433, 0.04038101, 0.02350518, 0.001223438, 0.000183442, 
    2.907142e-10, 0.002965097, 0.03510039, 0.1225919, 0.06290451, 0.02084379, 
    0.006563256,
  0.006127856, 0.02447541, 0.02329073, 0.00223007, 0.0282672, 0.05102627, 
    0.05114669, 0.04462456, 0.01336747, 0.0007974569, 0.01450062, 0.03782585, 
    0.06001034, 0.05932779, 0.03896101, 0.06675906, 0.04139701, 0.0004767241, 
    2.489545e-06, 2.158068e-08, 2.041151e-09, 3.244091e-08, 5.440403e-06, 
    0.127645, 0.09882165, 0.0334712, -3.193918e-05, 2.650205e-06, 
    -1.582303e-07,
  0.0199532, 0.2224303, 0.0961314, 0.001070621, 0.00115282, 0.05600279, 
    0.02528853, 0.0699539, 0.08193888, 0.06727113, 0.006978131, 0.02644252, 
    0.03415417, 0.04420442, 0.008412592, 0.001024533, 0.005008355, 
    -5.777653e-05, 0.0002505257, 1.087851e-06, 2.000479e-07, 1.474737e-06, 
    0.001354773, 0.1095312, 0.01321831, 0.0001623685, 0.01818887, 0.01558494, 
    1.087779e-05,
  0.02227577, 0.01719508, 0.007168768, 0.02102025, 0.0003547241, 0.001759039, 
    0.05818481, 0.06465808, 0.09614192, 0.06137796, 0.05093129, 0.1300263, 
    0.1560077, 0.2161497, 0.1127881, 0.06450228, 0.1465345, 0.1463532, 
    0.06537268, 0.05420461, 0.07663666, 0.05016413, 0.09683362, 0.03529354, 
    0.04291325, 0.1022873, 0.07551906, 0.01995089, 0.02560462,
  0.009859895, 0.0009508392, 6.502128e-06, 0.01317659, 0.0001838672, 
    0.008817414, 0.03355137, 0.04510057, 0.03891359, 0.02399737, 0.04635123, 
    0.07193904, 0.05423671, 0.03378686, 0.007066016, 0.01087487, 0.01882869, 
    0.02994706, 0.01741669, 0.0218909, 0.04188355, 0.02770893, 0.0126576, 
    0.01638824, 0.01104213, 0.03028014, 0.04901436, 0.09328432, 0.02453904,
  0.04863662, 0.03985649, 0.01798606, 0.01351111, 0.01710543, 0.01012127, 
    0.01069624, 0.03410911, 0.1785315, 0.09429158, 0.04726703, 0.06729515, 
    0.07313496, 0.01582329, 0.01786135, 0.05151867, 0.04871977, 0.04473768, 
    0.02730632, 0.02551386, 0.03737105, 0.02944715, 0.0514598, 0.05960852, 
    0.07719618, 0.05467969, 0.03363769, 0.02111855, 0.04421945,
  0.1584048, 0.1045149, 0.0423192, 0.03481473, 0.04618611, 0.0558312, 
    0.03843777, 0.08454669, 0.1044563, 0.10317, 0.1038896, 0.1367544, 
    0.2092478, 0.1757152, 0.1775314, 0.1723805, 0.1750787, 0.2114116, 
    0.0598447, 0.0263352, 0.07797177, 0.09533785, 0.117803, 0.07855802, 
    0.1440834, 0.1215075, 0.1030948, 0.04842923, 0.08210538,
  0.1413224, 0.1757013, 0.1265273, 0.1216471, 0.1322786, 0.1247705, 
    0.1366757, 0.06486739, 0.04700712, 0.101872, 0.1894392, 0.1364768, 
    0.1412314, 0.118383, 0.1733869, 0.2471147, 0.1763871, 0.3215128, 
    0.2099365, 0.102346, 0.1047795, 0.1485571, 0.1546657, 0.1971664, 
    0.1480618, 0.1450435, 0.217066, 0.1408855, 0.1251654,
  0.2179954, 0.2145944, 0.181407, 0.2341759, 0.2340052, 0.201842, 0.2225953, 
    0.1932912, 0.1505859, 0.09447828, 0.04108987, 0.03553203, 0.03051233, 
    0.1024209, 0.1038617, 0.2130381, 0.1817402, 0.298563, 0.1792897, 
    0.1260509, 0.1397801, 0.1009551, 0.1178949, 0.131292, 0.2158226, 
    0.2226406, 0.194885, 0.1804084, 0.2179969,
  0.2457449, 0.2075715, 0.1627915, 0.2170589, 0.2145327, 0.167066, 0.1700014, 
    0.1019611, 0.03102195, 0.02170116, 0.04783724, 0.09229799, 0.06052261, 
    0.05694307, 0.07151192, 0.2086195, 0.2149397, 0.2222396, 0.2377725, 
    0.2009885, 0.1351261, 0.1238233, 0.1202297, 0.09141938, 0.1609996, 
    0.03168073, 0.006431776, 0.2507855, 0.2261106,
  0.03843921, 0.04569184, 0.05750678, 0.07428385, 0.05875646, 0.03603887, 
    0.04385599, 0.04993374, 0.03674383, 0.02719938, 0.01960875, 0.02995115, 
    0.0613649, 0.1023056, 0.144856, 0.190831, 0.1232063, 0.0976, 0.06008267, 
    0.05219586, 0.07747938, 0.08713166, 0.04448445, 0.01485019, 0.008813294, 
    2.336939e-05, -0.001666629, 0.01339098, 0.07503182,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  -0.0001300029, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.931398e-06, 
    0.000158045, 0.004063245, 0.01048547, -0.0005039963, 0.002237868, 
    -9.70122e-06, 0, 0, 0.0008921532, 0.02276804, 0.02484782, 0.02489877, 
    0.05942499, 0.03601896, 0.003454213,
  0.1853989, 0.08145081, 0.029088, 0.01095535, -0.0002821996, 6.125482e-05, 
    0.02066509, -7.977146e-05, 1.938148e-05, -0.0002198692, 0.001612919, 
    0.001593039, 0.004446974, 0.03924319, 0.05346386, 0.07659946, 0.08717823, 
    0.0989176, 0.09959763, 0.07317011, 0.06934599, 0.07680089, 0.09374832, 
    0.1153464, 0.1859562, 0.1943287, 0.2107122, 0.1942873, 0.2154776,
  0.2407947, 0.1943687, 0.2308619, 0.1994791, 0.1601207, 0.1726327, 
    0.1559686, 0.1550877, 0.1767673, 0.1803811, 0.1645613, 0.1892676, 
    0.2070517, 0.2053142, 0.1627185, 0.1693689, 0.1711137, 0.2631218, 
    0.2282464, 0.2206537, 0.2025093, 0.2122465, 0.1735266, 0.2336116, 
    0.2121534, 0.1865038, 0.191881, 0.2063011, 0.2359038,
  0.1284446, 0.1005094, 0.1226307, 0.1913363, 0.1752158, 0.1495235, 
    0.1587014, 0.1979232, 0.2112793, 0.1760467, 0.1707231, 0.1328304, 
    0.1252143, 0.1598865, 0.1359919, 0.1473254, 0.1425638, 0.1352757, 
    0.140629, 0.1729246, 0.1608794, 0.155522, 0.1692443, 0.1241994, 
    0.1273949, 0.1922144, 0.2051937, 0.2030668, 0.1530909,
  0.1229988, 0.1027106, 0.07849954, 0.0947412, 0.1070355, 0.0950516, 
    0.1083771, 0.08718696, 0.08546265, 0.04824013, 0.03424012, 0.0508631, 
    0.09161965, 0.1056601, 0.1407579, 0.1171563, 0.1333392, 0.1092632, 
    0.1106275, 0.07164516, 0.08306226, 0.08888474, 0.07215974, 0.06391291, 
    0.1086849, 0.1040574, 0.138448, 0.09281018, 0.09878002,
  0.04702361, 0.01531235, 0.06691317, 0.09103541, 0.05863852, 0.03994802, 
    0.003876154, 0.001048302, 0.00113868, 2.998195e-05, 0.01832669, 
    0.06400644, 0.08878094, 0.07548918, 0.09383112, 0.0546556, 0.08012482, 
    0.07232893, 0.1974306, 0.1310582, 0.08494969, 0.0152679, 0.00157573, 
    0.0006194311, 0.04349119, 0.06633365, 0.1053694, 0.06593326, 0.09977549,
  -1.112926e-05, 0.00517463, 0.02130046, 0.0006392214, 0.01295182, 
    0.005127931, 0.0001139044, -0.0003385279, 0.007844345, 0.007253175, 
    0.002818037, 0.002545816, 0.02278141, 0.0228144, 0.04644765, 0.09688313, 
    0.1500767, 0.09335481, 0.03683206, 0.02841595, 6.542374e-05, 
    1.498214e-06, 2.196512e-09, 0.001077568, 0.03129984, 0.1153062, 
    0.05438668, 0.01882033, 0.001486676,
  0.008215035, 0.03119162, 0.01875304, 0.001504347, 0.02578789, 0.05732447, 
    0.06425148, 0.04107079, 0.00834544, 0.00127446, 0.01595555, 0.03269643, 
    0.06412585, 0.0663728, 0.04125022, 0.07321798, 0.03894714, 0.0005067147, 
    0.0004137179, 2.052514e-08, -1.286047e-10, 5.594443e-10, 8.756171e-06, 
    0.1118601, 0.07034115, 0.01511796, -1.386016e-05, 6.599111e-07, 
    -2.900311e-05,
  0.02957307, 0.230081, 0.07902579, 0.002644471, 0.009707545, 0.06613466, 
    0.03193992, 0.07815246, 0.06715699, 0.05328856, 0.008011756, 0.01623361, 
    0.02781087, 0.03243277, 0.006768906, 0.001147337, 0.003813337, 
    5.430393e-05, 7.09386e-05, 9.369573e-06, 1.179746e-07, 7.957798e-07, 
    0.0008674503, 0.08631386, 0.01051643, 0.0006133857, 0.009694209, 
    0.0247938, 0.0003876112,
  0.01819274, 0.02034961, 0.008352442, 0.03400411, 0.00101326, 0.001813703, 
    0.05547234, 0.05577819, 0.100818, 0.05160937, 0.04948316, 0.1172473, 
    0.1441773, 0.2146624, 0.1029598, 0.06824318, 0.1365883, 0.1535881, 
    0.06876304, 0.06322214, 0.08571604, 0.04503966, 0.09001152, 0.02358895, 
    0.04132098, 0.09442791, 0.06622826, 0.01325847, 0.02254433,
  0.004210277, 1.944052e-05, -4.312819e-05, 0.005328692, 7.517847e-05, 
    0.008863343, 0.0292986, 0.04910326, 0.03444063, 0.02154686, 0.04925569, 
    0.06962291, 0.05572864, 0.03332011, 0.008541992, 0.007520996, 0.01878911, 
    0.02639738, 0.01622698, 0.02423471, 0.02896717, 0.03338663, 0.00929301, 
    0.01563177, 0.007996871, 0.02273203, 0.02829875, 0.07997945, 0.004561284,
  0.03419896, 0.03304199, 0.01822077, 0.0149941, 0.01787006, 0.007307392, 
    0.009988088, 0.04538125, 0.2037346, 0.09198283, 0.0419126, 0.05641147, 
    0.07865396, 0.02143325, 0.02325651, 0.05045373, 0.03409264, 0.04380051, 
    0.02426768, 0.02308792, 0.02327986, 0.02854734, 0.04891569, 0.04562455, 
    0.06663266, 0.04528299, 0.02649925, 0.01227043, 0.04645242,
  0.1362044, 0.1038347, 0.04140755, 0.02926858, 0.04167804, 0.0521281, 
    0.04940629, 0.07728662, 0.09903868, 0.1017613, 0.09070516, 0.1238199, 
    0.1995799, 0.1848691, 0.1674082, 0.1642773, 0.1686617, 0.1840008, 
    0.04085962, 0.02536324, 0.06986114, 0.09781763, 0.1210162, 0.07857177, 
    0.1328843, 0.1023011, 0.07876504, 0.05669028, 0.08688181,
  0.1350875, 0.1800514, 0.1292253, 0.136465, 0.1231132, 0.1210059, 0.1312278, 
    0.1369151, 0.1193788, 0.1628128, 0.2140661, 0.1592138, 0.1485162, 
    0.1175412, 0.1760602, 0.2353857, 0.1726746, 0.2952785, 0.1953503, 
    0.09509803, 0.121864, 0.1598994, 0.1805324, 0.2054851, 0.1604754, 
    0.15682, 0.2055384, 0.1299309, 0.1194666,
  0.2437616, 0.2240564, 0.1817808, 0.2696844, 0.2463919, 0.1937595, 
    0.2009538, 0.2279358, 0.2060881, 0.1757531, 0.09851597, 0.09419757, 
    0.1630075, 0.181907, 0.1644271, 0.2731426, 0.2215881, 0.3135111, 
    0.2118353, 0.1356432, 0.1498679, 0.1657912, 0.1731721, 0.2240814, 
    0.2828014, 0.2568431, 0.2162079, 0.1852057, 0.2453176,
  0.2902755, 0.2312196, 0.2296269, 0.2590517, 0.2832031, 0.2143209, 
    0.2778763, 0.2449035, 0.1153798, 0.1144347, 0.08767484, 0.2022502, 
    0.132156, 0.09871908, 0.1386367, 0.2229399, 0.2682634, 0.2607269, 
    0.2747387, 0.2660055, 0.1912791, 0.1343159, 0.169942, 0.1475537, 
    0.1906781, 0.07088709, 0.03746942, 0.2833335, 0.2397905,
  0.1279229, 0.1087899, 0.1156353, 0.1630919, 0.1841233, 0.140129, 0.1010828, 
    0.1010239, 0.06641705, 0.06840076, 0.113536, 0.1650758, 0.1986755, 
    0.2155911, 0.2305766, 0.2388548, 0.151967, 0.1137418, 0.09565745, 
    0.07975157, 0.1000028, 0.145844, 0.1356446, 0.09174129, 0.09071361, 
    0.01035875, -0.005598078, 0.1091642, 0.1758973,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  -0.0005295048, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.003311346, 0.02085501, 
    0.02361818, 0.03337649, 0.02532579, 0.01167429, 5.475237e-05, 
    -1.90677e-06, 0, 0.003538149, 0.2042885, 0.1993337, 0.1128997, 0.135168, 
    0.06028283, 0.01548919,
  0.2534801, 0.1317954, 0.06443103, 0.041519, -0.0007251399, 0.001010084, 
    0.05371426, 0.001500609, 0.0018648, -0.0013581, 0.004640884, 0.005087816, 
    0.0101822, 0.120311, 0.1261073, 0.1366124, 0.1793672, 0.1562152, 
    0.1645369, 0.1472826, 0.1240895, 0.1450732, 0.2104297, 0.2287358, 
    0.2526411, 0.2625553, 0.2544838, 0.2476045, 0.3103879,
  0.2377503, 0.2106211, 0.2611725, 0.2288219, 0.1908633, 0.1961421, 
    0.1823105, 0.1738092, 0.1919322, 0.2210869, 0.2013331, 0.2345928, 
    0.2400087, 0.253085, 0.2079085, 0.2138053, 0.171436, 0.2735208, 
    0.2459754, 0.2469559, 0.2502569, 0.2400193, 0.241762, 0.2856961, 
    0.2516944, 0.1923745, 0.2085019, 0.2031705, 0.2081157,
  0.1292031, 0.09418563, 0.1101803, 0.1790106, 0.1757448, 0.1459967, 
    0.1478696, 0.1964025, 0.2026508, 0.1658663, 0.1683647, 0.1316884, 
    0.1298804, 0.1627349, 0.1309762, 0.1454268, 0.1268417, 0.1280775, 
    0.1331088, 0.1683642, 0.162196, 0.1574952, 0.173351, 0.1187219, 
    0.1165771, 0.1866506, 0.189557, 0.1885553, 0.1477496,
  0.1121978, 0.09878306, 0.06896076, 0.07723629, 0.1016436, 0.09996985, 
    0.0979364, 0.09944853, 0.07928573, 0.03395939, 0.03141324, 0.05592474, 
    0.08672922, 0.1013335, 0.1467319, 0.1149715, 0.1284578, 0.09496611, 
    0.1034542, 0.05848712, 0.08911677, 0.08664429, 0.07834835, 0.06391375, 
    0.1050335, 0.1069244, 0.1212209, 0.08605194, 0.08979326,
  0.0387585, 0.01792685, 0.06393293, 0.09920081, 0.04873934, 0.03436305, 
    0.007555652, 0.003927376, 0.0005206452, 0.00215482, 0.02479883, 
    0.07983682, 0.08890027, 0.07222021, 0.07781135, 0.04832026, 0.07703343, 
    0.06375206, 0.1918893, 0.1237179, 0.07412158, 0.01083335, 0.0001865064, 
    -4.234083e-05, 0.04707473, 0.07066774, 0.1060567, 0.05728171, 0.1147046,
  0.0005565129, 0.01925687, 0.01797089, 0.0004863655, 0.0163775, 
    0.0006635752, 0.0001310955, -0.0001102499, 0.001830876, 0.003286652, 
    0.009466164, 0.006588284, 0.02698695, 0.03539988, 0.04079347, 0.08638497, 
    0.1293952, 0.0857875, 0.03771963, 0.03600784, 7.893344e-05, 3.774724e-05, 
    1.507155e-09, 8.757872e-05, 0.03093349, 0.1139462, 0.05944692, 
    0.005377513, 0.0007618815,
  0.00199489, 0.0453316, 0.01374955, 0.0017139, 0.02698337, 0.05507089, 
    0.07633594, 0.03801262, 0.008949898, 0.001583318, 0.01616456, 0.03260076, 
    0.07384612, 0.07176931, 0.05393639, 0.07311833, 0.02770643, 0.0009720173, 
    0.0001682565, -2.527495e-09, 4.208335e-11, 3.782948e-09, 9.756422e-06, 
    0.1025016, 0.05411109, 0.01105276, 8.313435e-06, 3.057363e-07, 0.004569193,
  0.0394272, 0.2386266, 0.07881799, 0.005736664, 0.0150098, 0.05479871, 
    0.03471293, 0.08409902, 0.05355917, 0.03898931, 0.01575595, 0.01074828, 
    0.01602289, 0.02780826, 0.006793094, 0.001808797, 0.002671166, 
    5.472229e-05, 6.485972e-06, 1.075783e-05, 1.834079e-07, 1.284322e-07, 
    0.005246619, 0.06834771, 0.008136341, 0.001184304, 0.005257443, 
    0.03459512, 0.003943755,
  0.01512755, 0.01500021, 0.007969442, 0.04536624, 0.001095384, 0.00163204, 
    0.0488449, 0.04986709, 0.1045745, 0.04433008, 0.05142083, 0.1083729, 
    0.1381524, 0.2183567, 0.09271942, 0.07825036, 0.1275108, 0.1471035, 
    0.08073154, 0.06410615, 0.1034201, 0.05004372, 0.09579189, 0.01935309, 
    0.04388542, 0.09457691, 0.06693283, 0.009846251, 0.02274665,
  0.001586853, 1.918228e-06, 4.692317e-07, 0.00491225, 4.548423e-05, 
    0.008423816, 0.0309083, 0.0519562, 0.02671179, 0.01850595, 0.04908185, 
    0.07302029, 0.05996131, 0.03654886, 0.01441862, 0.006231398, 0.0184959, 
    0.01489206, 0.01321706, 0.02263331, 0.02083666, 0.04090998, 0.00846302, 
    0.0163187, 0.007143977, 0.02104956, 0.01886332, 0.05744094, 0.001589473,
  0.03118924, 0.0381243, 0.01833614, 0.01632963, 0.01855058, 0.00433727, 
    0.009686899, 0.0811407, 0.2214933, 0.1019668, 0.04199231, 0.05396722, 
    0.08419047, 0.01471639, 0.02218772, 0.05490529, 0.02691261, 0.03898358, 
    0.02033219, 0.01425079, 0.0157878, 0.02759858, 0.05182272, 0.03973481, 
    0.06263582, 0.03947169, 0.02402108, 0.009552714, 0.04127883,
  0.1225346, 0.1000527, 0.04451303, 0.02890156, 0.04144625, 0.04922801, 
    0.05343574, 0.06662173, 0.09351927, 0.1030445, 0.07104625, 0.09625491, 
    0.1811395, 0.1850538, 0.1605844, 0.1620191, 0.1658589, 0.1756478, 
    0.03031501, 0.02455043, 0.0688829, 0.103525, 0.1286257, 0.07848598, 
    0.1328131, 0.08448582, 0.06721746, 0.06551684, 0.0800932,
  0.1290499, 0.1757562, 0.1192408, 0.1353538, 0.1092583, 0.1005256, 
    0.1190372, 0.1940965, 0.1885505, 0.173806, 0.2051286, 0.1821036, 
    0.1576212, 0.1300376, 0.1822523, 0.2571585, 0.1882069, 0.2841379, 
    0.1900685, 0.1026137, 0.1252549, 0.166867, 0.2192133, 0.220486, 
    0.1820124, 0.1619676, 0.1948751, 0.1296523, 0.1175326,
  0.2453549, 0.2298404, 0.1783579, 0.2860687, 0.2642207, 0.1874399, 0.200853, 
    0.227358, 0.2514651, 0.2110079, 0.1631466, 0.1521246, 0.2307913, 
    0.1755714, 0.1865369, 0.2910152, 0.2328691, 0.3169923, 0.2529067, 
    0.1295736, 0.1648778, 0.1816792, 0.2269267, 0.276133, 0.2998002, 
    0.2749833, 0.2047237, 0.1907491, 0.2237441,
  0.2722788, 0.2376608, 0.2567895, 0.2978975, 0.3137997, 0.2383354, 
    0.3223071, 0.3188455, 0.2039127, 0.2103166, 0.1381346, 0.3062255, 
    0.1537288, 0.133761, 0.1428613, 0.1969698, 0.2760327, 0.255733, 
    0.2806175, 0.2811466, 0.2256015, 0.1513238, 0.2003062, 0.1889746, 
    0.222567, 0.1123017, 0.09386043, 0.2762929, 0.2722837,
  0.1609389, 0.1343212, 0.1755194, 0.2277415, 0.2363834, 0.1987417, 
    0.1863558, 0.1746869, 0.1515511, 0.1375341, 0.1564041, 0.2336833, 
    0.2596396, 0.2599745, 0.2699398, 0.2726347, 0.1743152, 0.1263642, 
    0.1148231, 0.09684162, 0.1057265, 0.1648776, 0.1707258, 0.1306021, 
    0.1774816, 0.05499224, 0.0754405, 0.1303258, 0.22181,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0.0124918, -3.309479e-06, -1.070779e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0002195299, 0.04458348, 0.05590422, 0.04651151, 0.09534875, 0.06459048, 
    0.03343213, 0.001380666, 0.002117227, 0.001264363, 0.03811188, 0.2982576, 
    0.2589813, 0.2385101, 0.2493174, 0.1088905, 0.02253532,
  0.26618, 0.1585084, 0.1032272, 0.09715675, 0.002353139, 0.006289893, 
    0.116561, 0.002387718, 0.002303367, 0.003902867, 0.009486387, 0.01079228, 
    0.07201549, 0.2235488, 0.2022801, 0.2329704, 0.2512805, 0.2480974, 
    0.2445833, 0.2482676, 0.2221503, 0.2304706, 0.2976531, 0.3113299, 
    0.272322, 0.2658607, 0.2480998, 0.256545, 0.3441784,
  0.2393076, 0.2162228, 0.2655471, 0.2447739, 0.2361561, 0.2158092, 
    0.1971412, 0.1986202, 0.2272003, 0.2535506, 0.2465752, 0.2511838, 
    0.2510986, 0.2721006, 0.2391356, 0.2208949, 0.175211, 0.2636334, 
    0.2473522, 0.2563583, 0.2520525, 0.2548649, 0.2757467, 0.300302, 
    0.2478226, 0.1924254, 0.2083463, 0.1974438, 0.2091673,
  0.1276789, 0.09437238, 0.1053777, 0.16969, 0.1692987, 0.1378635, 0.1389914, 
    0.1957168, 0.2002299, 0.1763192, 0.1494249, 0.1246719, 0.1200419, 
    0.1624379, 0.1251825, 0.1264583, 0.1164559, 0.121047, 0.1177096, 
    0.1610139, 0.1592728, 0.1571469, 0.1612723, 0.1174052, 0.11035, 
    0.1902804, 0.176205, 0.1739183, 0.1378231,
  0.1006939, 0.1008957, 0.05852947, 0.07522373, 0.1016376, 0.1012025, 
    0.1070108, 0.0964637, 0.08162036, 0.0267499, 0.03202788, 0.06100075, 
    0.08579412, 0.0990444, 0.1451795, 0.1061423, 0.1159034, 0.09621507, 
    0.08974349, 0.04898033, 0.08759019, 0.07882156, 0.07659863, 0.07209033, 
    0.09145302, 0.09764145, 0.1070717, 0.08003388, 0.07528028,
  0.03490726, 0.02003111, 0.06379157, 0.1023001, 0.04437478, 0.02994153, 
    0.008229956, 0.0009553119, 0.001817819, 0.007692468, 0.03717336, 
    0.07921633, 0.09040296, 0.06814624, 0.06808871, 0.0378748, 0.06491877, 
    0.05906585, 0.1830878, 0.1168318, 0.05746236, 0.0207581, 0.000273187, 
    -1.083601e-05, 0.056693, 0.06734825, 0.1106202, 0.05044322, 0.1301471,
  0.003823226, 0.0338807, 0.02202028, 0.001247605, 0.02266429, 0.0001783188, 
    0.0002851896, -0.0002647422, 0.0009177321, 0.003404193, 0.02490539, 
    0.01730212, 0.02760718, 0.04037043, 0.04243448, 0.07967267, 0.106394, 
    0.07939643, 0.04173613, 0.04170405, 3.554e-06, 0.003646107, 1.070922e-08, 
    3.994277e-05, 0.03640722, 0.1154755, 0.07009953, 0.002954279, 0.003776314,
  0.001550411, 0.05656676, 0.02148763, 0.005351578, 0.02457584, 0.06163342, 
    0.08718835, 0.03353622, 0.01487793, 0.001496009, 0.01711623, 0.04029937, 
    0.08049215, 0.07008851, 0.07361731, 0.07083695, 0.02757623, 0.00559849, 
    5.649424e-05, 7.18762e-09, 1.196176e-08, 6.696634e-08, 0.0008929649, 
    0.1141647, 0.05480878, 0.01103777, 1.225559e-05, 1.95129e-07, 0.0002655007,
  0.08051215, 0.2683992, 0.1030148, 0.008561631, 0.01275226, 0.04479917, 
    0.03309602, 0.08628265, 0.05356695, 0.02922493, 0.01248153, 0.008452212, 
    0.01248552, 0.02889456, 0.006815271, 0.002243802, 0.005274738, 
    0.001283664, 0.0009925371, -1.124171e-05, 3.680412e-07, -5.32629e-06, 
    0.02483669, 0.06709345, 0.007367638, 0.0009377906, 0.006192577, 
    0.03347417, 0.01071835,
  0.0143981, 0.0144956, 0.01038297, 0.05054007, 0.001214348, 0.002627665, 
    0.05911686, 0.04342004, 0.1232911, 0.0441277, 0.06462076, 0.1115367, 
    0.1434852, 0.2262885, 0.09659734, 0.0817136, 0.1459506, 0.1428134, 
    0.09108607, 0.07036225, 0.1141207, 0.05694837, 0.09646322, 0.02151714, 
    0.0481078, 0.1021439, 0.06195037, 0.01175919, 0.0169626,
  0.003449076, -1.58987e-06, 0.0002595372, 0.01000537, 2.659855e-05, 
    0.009836815, 0.02876562, 0.05648995, 0.02000413, 0.01902369, 0.05091786, 
    0.09274532, 0.07228045, 0.03595894, 0.01722181, 0.005785275, 0.01243826, 
    0.01036484, 0.01059881, 0.03777729, 0.01663908, 0.05192457, 0.008369578, 
    0.02477818, 0.008711101, 0.02039832, 0.01878227, 0.0359997, 0.0006557618,
  0.03257094, 0.03872349, 0.02320537, 0.01826083, 0.0222344, 0.002894298, 
    0.009013634, 0.1052778, 0.233951, 0.1017194, 0.0483185, 0.07189766, 
    0.07885248, 0.01612362, 0.02516584, 0.06334057, 0.01662103, 0.03771244, 
    0.02264599, 0.01121402, 0.01668684, 0.02790826, 0.05708105, 0.03831297, 
    0.06327565, 0.03161088, 0.02403536, 0.01052978, 0.04221691,
  0.1204818, 0.08495376, 0.05466238, 0.02941854, 0.04312739, 0.04290209, 
    0.05440282, 0.05706621, 0.08364147, 0.104436, 0.06447901, 0.09178817, 
    0.1767816, 0.1651181, 0.1636569, 0.1654118, 0.152321, 0.1586605, 
    0.02797435, 0.023257, 0.06823738, 0.1045934, 0.1200031, 0.07782193, 
    0.1224181, 0.07779309, 0.0681024, 0.05347528, 0.08206381,
  0.134614, 0.1703232, 0.1372488, 0.1371199, 0.1023989, 0.09231322, 
    0.1171221, 0.2039491, 0.2018652, 0.1571636, 0.186764, 0.1812816, 
    0.1526039, 0.1436137, 0.1767899, 0.2472937, 0.1850654, 0.2713175, 
    0.1713621, 0.1063795, 0.1221151, 0.1705903, 0.2401359, 0.2549555, 
    0.1743473, 0.152321, 0.1770104, 0.1266305, 0.1214863,
  0.242708, 0.2417294, 0.1804024, 0.2832986, 0.2534252, 0.1870555, 0.1914271, 
    0.222726, 0.2655154, 0.2430076, 0.1957368, 0.1830865, 0.2728351, 
    0.1691406, 0.1890474, 0.2824206, 0.2243586, 0.3195572, 0.2639307, 
    0.1195924, 0.1694219, 0.1943182, 0.2277664, 0.2883944, 0.3062941, 
    0.2847856, 0.2136002, 0.1944429, 0.2498657,
  0.2439185, 0.2495198, 0.2663762, 0.2890288, 0.3097119, 0.2419749, 
    0.3403261, 0.3164373, 0.2836565, 0.2679076, 0.2166766, 0.3327928, 
    0.146343, 0.1389867, 0.1478814, 0.1796513, 0.2753932, 0.2560544, 
    0.2801148, 0.2832821, 0.2501833, 0.1603364, 0.2090345, 0.2464419, 
    0.2193142, 0.1904067, 0.1894696, 0.2710629, 0.2481014,
  0.159965, 0.1595245, 0.1930566, 0.2584009, 0.2779674, 0.2180127, 0.1992663, 
    0.1938228, 0.1675106, 0.1496614, 0.1590362, 0.2147883, 0.2288924, 
    0.2345583, 0.2575269, 0.2390586, 0.1647416, 0.1041614, 0.1035441, 
    0.121185, 0.1348534, 0.1948767, 0.1913135, 0.1669032, 0.2014483, 
    0.1092033, 0.1170347, 0.1389082, 0.2360923,
  0.0003970285, 0.0002160506, 3.507261e-05, -0.0001459053, -0.0003268833, 
    -0.0005078612, -0.0006888392, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -0.00088936, -0.0007083821, -0.0005274042, -0.0003464262, -0.0001654483, 
    1.552965e-05, 0.0001965076, 0.0005418108,
  0.01380973, 0.02004084, 0.0006848198, 0, 0, 0, 0, 0, 0, 0, 0, 0.0002574608, 
    0.001538536, 0.1176415, 0.05954433, 0.07019792, 0.1180465, 0.130093, 
    0.07167362, 0.01493035, 0.005029887, 0.003712631, 0.09711372, 0.2983712, 
    0.267404, 0.2543125, 0.2592764, 0.2060817, 0.04142476,
  0.2640466, 0.1626594, 0.1146857, 0.1667693, 0.009619977, 0.03025736, 
    0.1777752, 0.01099142, 0.002814665, 0.02277957, 0.02458159, 0.02699174, 
    0.1609921, 0.297618, 0.2585971, 0.2504315, 0.2849894, 0.2684091, 
    0.2695885, 0.2773899, 0.2509678, 0.2517824, 0.3137431, 0.3525414, 
    0.2843771, 0.2409259, 0.2498908, 0.2569993, 0.3327237,
  0.2300435, 0.2218723, 0.2569225, 0.2525598, 0.2641601, 0.2281579, 
    0.2190664, 0.2125608, 0.2389386, 0.2597928, 0.2681571, 0.2612891, 
    0.2661298, 0.2702495, 0.2536566, 0.2341125, 0.1885464, 0.2669405, 
    0.2488954, 0.2706651, 0.2430232, 0.2510489, 0.2678905, 0.287365, 
    0.2466347, 0.1925308, 0.1976402, 0.1913481, 0.1808318,
  0.1383727, 0.1161734, 0.09565648, 0.1647311, 0.172389, 0.1286191, 
    0.1484109, 0.1941302, 0.1996777, 0.1754586, 0.1484925, 0.1450492, 
    0.1170553, 0.1600521, 0.1294927, 0.124696, 0.1189265, 0.1235591, 
    0.1242375, 0.1622673, 0.1683108, 0.1610632, 0.1525989, 0.1144551, 
    0.1027771, 0.2008031, 0.1771357, 0.1575143, 0.1233504,
  0.09863167, 0.1053492, 0.05175992, 0.07474249, 0.1045609, 0.104922, 
    0.1087611, 0.1085445, 0.0808726, 0.02392964, 0.03014198, 0.06469817, 
    0.08762461, 0.1176905, 0.1478105, 0.0979872, 0.1051538, 0.08855048, 
    0.08939226, 0.05535445, 0.08560219, 0.0821657, 0.08199055, 0.08560621, 
    0.08023832, 0.1145242, 0.1072238, 0.08051214, 0.08073984,
  0.01747854, 0.01032586, 0.0620443, 0.1045921, 0.04983472, 0.02780634, 
    0.01096873, 0.001638785, 0.006065671, 0.007528965, 0.02657847, 
    0.07755651, 0.08980526, 0.06282248, 0.06169126, 0.03126885, 0.05013416, 
    0.0530016, 0.1746936, 0.1131327, 0.05759846, 0.03101283, 6.333807e-05, 
    -3.386722e-06, 0.06553294, 0.0686494, 0.1183865, 0.04835404, 0.1339218,
  0.002941725, 0.02351359, 0.04533368, 0.006488793, 0.02556943, 0.0004469775, 
    0.0002707719, -0.0001644549, 0.001051282, 0.001586652, 0.08455137, 
    0.0603778, 0.02568879, 0.04565673, 0.04100888, 0.07258989, 0.0905949, 
    0.07005036, 0.04257067, 0.04405509, 6.574921e-06, 0.006731412, 
    2.597596e-07, 4.788004e-05, 0.04824077, 0.1174863, 0.07935185, 
    0.004590072, 0.00596782,
  0.004718277, 0.06857461, 0.04746494, 0.01034636, 0.0214477, 0.07845399, 
    0.1119397, 0.03462313, 0.01860233, 0.002076841, 0.01715375, 0.05988077, 
    0.1011411, 0.0877383, 0.09435497, 0.0756415, 0.02977322, 0.009424478, 
    0.000233877, 2.439876e-07, 8.568594e-08, 1.32699e-06, 0.005732897, 
    0.133074, 0.06858131, 0.03134286, 2.343427e-05, 8.450868e-07, 
    -9.146817e-05,
  0.09646401, 0.2961387, 0.1594248, 0.008827121, 0.007455851, 0.04740427, 
    0.0300003, 0.09482552, 0.06684613, 0.03720224, 0.01168072, 0.009573121, 
    0.02187157, 0.03923624, 0.008532731, 0.001862565, 0.003200537, 
    0.001351417, 0.003127764, 0.0004639964, 1.501906e-06, 0.000565088, 
    0.0356932, 0.08061145, 0.00614239, 0.0009583778, 0.006688811, 0.02377487, 
    0.03984676,
  0.01804932, 0.01653234, 0.01518636, 0.06375194, 0.001085415, 0.002677378, 
    0.06890628, 0.04705331, 0.1448326, 0.05106227, 0.09390438, 0.1416227, 
    0.1613357, 0.2489904, 0.116131, 0.1010621, 0.165338, 0.1586296, 
    0.1144664, 0.08715914, 0.1242344, 0.07257025, 0.1102812, 0.03210592, 
    0.05748036, 0.1137777, 0.06130272, 0.02018777, 0.01690875,
  0.01244251, 3.357372e-05, 3.794669e-05, 0.01423708, 2.740142e-05, 
    0.01140776, 0.02808535, 0.06970415, 0.01864255, 0.01938999, 0.06120387, 
    0.1144879, 0.08334921, 0.04258095, 0.02537029, 0.01029774, 0.01007048, 
    0.008062609, 0.006096432, 0.03615501, 0.02736579, 0.07482783, 0.01195881, 
    0.03591457, 0.01296557, 0.02312128, 0.03393278, 0.02711109, 0.001867675,
  0.02791052, 0.02092832, 0.02054989, 0.01910971, 0.02178851, 0.002938133, 
    0.01426292, 0.1155426, 0.2445905, 0.09440053, 0.05347556, 0.0941851, 
    0.08107257, 0.01631261, 0.02692866, 0.07372626, 0.01806248, 0.04195429, 
    0.01985926, 0.01095792, 0.02220689, 0.03838908, 0.06817009, 0.04582738, 
    0.06917648, 0.02951922, 0.02701754, 0.0114551, 0.04312044,
  0.1106475, 0.07523908, 0.05696441, 0.03588013, 0.05168095, 0.03820882, 
    0.056095, 0.05010526, 0.07246158, 0.100414, 0.05977227, 0.08934699, 
    0.1558754, 0.157047, 0.1706528, 0.1609838, 0.1506657, 0.1528676, 
    0.02764799, 0.01963685, 0.06327184, 0.1105864, 0.1094992, 0.07108435, 
    0.1199419, 0.0748743, 0.06467102, 0.05278403, 0.06419301,
  0.1275187, 0.189339, 0.1291164, 0.1299855, 0.09178264, 0.09431793, 
    0.1105924, 0.208538, 0.2031994, 0.14382, 0.1713681, 0.182241, 0.1419518, 
    0.1463352, 0.1603645, 0.2739808, 0.1897132, 0.255131, 0.1550992, 
    0.104439, 0.1124371, 0.1698153, 0.2479209, 0.2833653, 0.1914096, 
    0.1505944, 0.1667691, 0.1191682, 0.1168736,
  0.2412872, 0.2622305, 0.1923994, 0.2794356, 0.2548864, 0.1837406, 0.183849, 
    0.2165605, 0.2649983, 0.2824373, 0.229266, 0.1896114, 0.2705802, 
    0.1563898, 0.1988031, 0.2939075, 0.2401357, 0.33851, 0.2615928, 
    0.1149972, 0.1789453, 0.2012555, 0.2416762, 0.2723542, 0.3283868, 
    0.305981, 0.2261296, 0.1874206, 0.2327761,
  0.2336699, 0.2415387, 0.2607049, 0.3110956, 0.3189259, 0.237583, 0.3419508, 
    0.3344782, 0.3109983, 0.2577161, 0.2071252, 0.3297433, 0.1342678, 
    0.1357831, 0.1463965, 0.1799145, 0.2724344, 0.2497791, 0.290038, 
    0.2898027, 0.2398858, 0.2082682, 0.1881729, 0.266962, 0.2158835, 
    0.2454062, 0.2810191, 0.289946, 0.2307528,
  0.1351204, 0.1684278, 0.196611, 0.2609126, 0.291121, 0.2216027, 0.1994293, 
    0.197988, 0.1742602, 0.1409453, 0.1374456, 0.178532, 0.1833756, 0.195866, 
    0.2169656, 0.1781946, 0.1421051, 0.08665637, 0.0894489, 0.1237111, 
    0.1459856, 0.2331157, 0.1932357, 0.1650422, 0.1829564, 0.142169, 
    0.1483082, 0.137541, 0.2279409,
  0.01043131, 0.009305734, 0.008180157, 0.007054581, 0.005929005, 
    0.004803428, 0.003677852, 0.005199137, 0.004737262, 0.004275388, 
    0.003813513, 0.003351638, 0.002889764, 0.002427889, -0.0003887502, 
    -6.000604e-05, 0.0002687381, 0.0005974823, 0.0009262264, 0.001254971, 
    0.001583715, 0.002937179, 0.004195886, 0.005454592, 0.0067133, 
    0.007972006, 0.009230713, 0.01048942, 0.01133177,
  0.02775702, 0.0250874, 0.02047222, 0.006650193, -0.0001081852, 0, 0, 0, 0, 
    0, 0.001315886, 0.02354884, 0.005751247, 0.1551722, 0.0581453, 
    0.06604121, 0.1191122, 0.1457637, 0.1419946, 0.07131425, 0.05532978, 
    0.04485558, 0.1821555, 0.2924344, 0.2529213, 0.2447653, 0.2510258, 
    0.263411, 0.08635058,
  0.2673642, 0.1665087, 0.1134437, 0.1781729, 0.03002411, 0.077347, 
    0.1911128, 0.03611447, 0.02887758, 0.04475974, 0.06495435, 0.03230251, 
    0.229747, 0.297938, 0.2714621, 0.2474712, 0.2857641, 0.2780128, 
    0.2850099, 0.266265, 0.2683491, 0.2647719, 0.3247151, 0.3727976, 
    0.2813905, 0.2237229, 0.2551978, 0.2588447, 0.3311757,
  0.2250781, 0.2200211, 0.2750393, 0.2602848, 0.2600283, 0.2283572, 
    0.2149806, 0.2211965, 0.251781, 0.2654355, 0.2788625, 0.2645939, 
    0.2632918, 0.2610105, 0.2587726, 0.2503849, 0.1906517, 0.2665241, 
    0.2584721, 0.2800605, 0.2352825, 0.2345669, 0.2660605, 0.2899952, 
    0.2375787, 0.1912559, 0.1766956, 0.1926413, 0.1721186,
  0.1454181, 0.09601731, 0.1047089, 0.1762262, 0.1757923, 0.1315955, 
    0.147149, 0.1847508, 0.1877997, 0.1818476, 0.1495537, 0.1348137, 
    0.1118285, 0.1642873, 0.1298059, 0.121034, 0.1254465, 0.1231315, 
    0.1167408, 0.1604548, 0.1743818, 0.1701079, 0.1642988, 0.1198518, 
    0.09530389, 0.1839941, 0.1701581, 0.1454794, 0.1171473,
  0.09744372, 0.1063617, 0.05162507, 0.07646713, 0.09705257, 0.1125217, 
    0.1096655, 0.107899, 0.07870045, 0.02258179, 0.03005327, 0.0620564, 
    0.09128534, 0.1179357, 0.153081, 0.09616921, 0.1041911, 0.08068591, 
    0.09793919, 0.05464554, 0.09513989, 0.0808219, 0.07475158, 0.1015962, 
    0.07467178, 0.1126957, 0.1126487, 0.07270217, 0.08772378,
  0.007644347, 0.001252602, 0.06431036, 0.117151, 0.06205385, 0.03260787, 
    0.01132911, 0.002262215, 0.0108107, 0.004757032, 0.01531812, 0.06193694, 
    0.09121247, 0.06616585, 0.05885792, 0.03691837, 0.04363655, 0.04817531, 
    0.1716846, 0.1208616, 0.06992534, 0.02853242, -1.533486e-06, 
    -5.877733e-07, 0.0733825, 0.07189193, 0.1177376, 0.04932526, 0.106417,
  0.004571222, 0.01692793, 0.07448512, 0.007236064, 0.02511782, 0.001620908, 
    0.0006571842, 0.0006358224, 0.001010223, 0.0004356512, 0.1078379, 
    0.06252094, 0.02176576, 0.04427671, 0.04218511, 0.07709761, 0.08162773, 
    0.07568529, 0.04965359, 0.04622898, -6.497357e-05, 0.0002157132, 
    2.49386e-07, 2.276421e-06, 0.06954704, 0.1391924, 0.07555851, 0.01000338, 
    0.002504803,
  0.009493224, 0.08436465, 0.1328233, 0.01037603, 0.02389619, 0.09807651, 
    0.1341352, 0.04594353, 0.02109741, 0.002027913, 0.01998393, 0.07520145, 
    0.1052417, 0.09957525, 0.1175922, 0.07631008, 0.03454298, 0.01480192, 
    0.0001375742, 5.813808e-07, 2.623372e-07, 0.0001444027, 0.003381753, 
    0.1599848, 0.09666827, 0.1319567, 3.472736e-05, 1.549045e-05, -3.99233e-05,
  0.107829, 0.3469385, 0.208272, 0.007067425, 0.001853746, 0.04636439, 
    0.03534907, 0.1021746, 0.09205026, 0.06509785, 0.01247982, 0.01137262, 
    0.02909099, 0.05235199, 0.0117352, 0.003222221, 0.0009956263, 0.01033864, 
    0.001157489, 0.001183723, 0.01036962, 0.009616728, 0.07571697, 0.1039725, 
    0.007974923, 0.000903812, 0.007117369, 0.02072773, 0.02575545,
  0.02149173, 0.02136968, 0.01887113, 0.07993317, 0.001289878, 0.002595079, 
    0.07852279, 0.0537659, 0.1615951, 0.06225431, 0.109623, 0.1496935, 
    0.1762194, 0.2551112, 0.1343831, 0.1182862, 0.1796788, 0.1820827, 
    0.1304568, 0.09614792, 0.1411207, 0.09002042, 0.1248321, 0.03691363, 
    0.06607991, 0.1307416, 0.06369347, 0.04083222, 0.02017003,
  0.01071019, 1.196405e-05, -5.112957e-05, 0.009746335, 0.0007593938, 
    0.01465022, 0.0345746, 0.06609585, 0.02322261, 0.02525888, 0.06319133, 
    0.1271675, 0.08368507, 0.05016738, 0.03326511, 0.01886039, 0.0129004, 
    0.009002418, 0.004223685, 0.05658532, 0.04006064, 0.09847482, 0.0142546, 
    0.04118078, 0.01410976, 0.02793968, 0.02505256, 0.03641339, 0.0005194704,
  0.01161393, 0.01019883, 0.02055415, 0.01457722, 0.022593, 0.003332997, 
    0.01520206, 0.116635, 0.2504932, 0.07617678, 0.05769752, 0.1077656, 
    0.08031789, 0.01798431, 0.03011932, 0.07607421, 0.02215962, 0.04858998, 
    0.0211685, 0.0117397, 0.03861046, 0.05316659, 0.06879406, 0.05301663, 
    0.09082963, 0.03306745, 0.03344572, 0.008928209, 0.04415689,
  0.1026499, 0.06870449, 0.06484614, 0.0484925, 0.06640117, 0.02666753, 
    0.05679219, 0.04678727, 0.06004894, 0.09214044, 0.06265303, 0.07908175, 
    0.1403734, 0.1598814, 0.1725119, 0.1638102, 0.1544848, 0.1548995, 
    0.02799607, 0.01773468, 0.06146464, 0.1265085, 0.1093189, 0.06734535, 
    0.12333, 0.09237382, 0.06808674, 0.0527192, 0.06839168,
  0.132731, 0.1874719, 0.1500632, 0.1303696, 0.0891002, 0.1004758, 0.1270261, 
    0.2116698, 0.1962038, 0.1326585, 0.164077, 0.1804786, 0.1452401, 
    0.157622, 0.1809815, 0.2672719, 0.1933127, 0.245272, 0.1348216, 
    0.1009106, 0.1121903, 0.1785263, 0.2449231, 0.2905434, 0.1945335, 
    0.1440131, 0.169783, 0.1150141, 0.1147056,
  0.22774, 0.2537722, 0.1864931, 0.2547272, 0.251737, 0.1639977, 0.1822957, 
    0.2158371, 0.254429, 0.3031481, 0.2497502, 0.1834348, 0.2862229, 
    0.1521147, 0.2034615, 0.2806118, 0.2515905, 0.3517351, 0.2462216, 
    0.1227396, 0.1975528, 0.1876141, 0.2384163, 0.2965195, 0.3601539, 
    0.3203942, 0.2092844, 0.2062485, 0.2700176,
  0.2632734, 0.2591019, 0.2466625, 0.3179441, 0.3353756, 0.2821416, 
    0.3201256, 0.3579395, 0.299004, 0.2538448, 0.207439, 0.3022941, 
    0.1329836, 0.1291959, 0.1356574, 0.1781654, 0.2906001, 0.2467729, 
    0.2910002, 0.307564, 0.2625664, 0.2141155, 0.1866264, 0.251714, 
    0.2279116, 0.3042069, 0.3400433, 0.2792616, 0.2395938,
  0.1186111, 0.1779616, 0.1990753, 0.2267094, 0.2773218, 0.2249287, 
    0.2158085, 0.207268, 0.1614851, 0.1244402, 0.1126668, 0.1498184, 
    0.1506172, 0.1754228, 0.1803115, 0.1368683, 0.1322019, 0.08108748, 
    0.09626766, 0.1407214, 0.1848583, 0.270611, 0.2030002, 0.1587778, 
    0.1616788, 0.1520572, 0.1681957, 0.1222015, 0.2135593,
  0.02662281, 0.02587743, 0.02513206, 0.02438669, 0.02364131, 0.02289594, 
    0.02215057, 0.01980616, 0.0185438, 0.01728144, 0.01601907, 0.01475671, 
    0.01349435, 0.01223199, 0.01147202, 0.01231596, 0.0131599, 0.01400384, 
    0.01484777, 0.01569171, 0.01653565, 0.01727252, 0.01843632, 0.01960012, 
    0.02076391, 0.02192771, 0.02309151, 0.02425531, 0.0272191,
  0.05691364, 0.02939671, 0.02437822, 0.02201968, 0.01105898, 0.001883519, 0, 
    0, 0, 0.0003140963, 0.02630493, 0.02761178, 0.02395334, 0.1574417, 
    0.05694401, 0.06090103, 0.1062685, 0.1577805, 0.1510363, 0.1416979, 
    0.1861547, 0.1708339, 0.2296596, 0.2988175, 0.2529364, 0.2197592, 
    0.2406965, 0.2632499, 0.1604843,
  0.2696794, 0.1773062, 0.120656, 0.1759443, 0.09067498, 0.1266176, 
    0.2020315, 0.09137741, 0.05671065, 0.07440399, 0.09664775, 0.07955103, 
    0.259866, 0.3097741, 0.2634089, 0.2419354, 0.2802796, 0.2915989, 
    0.2940168, 0.2650285, 0.2759855, 0.2655919, 0.3359758, 0.3886256, 
    0.2771142, 0.2168437, 0.2503915, 0.2625049, 0.3166988,
  0.2242534, 0.2337496, 0.2810304, 0.270449, 0.278568, 0.2414937, 0.2243876, 
    0.2339286, 0.2673118, 0.2706294, 0.2811736, 0.2786627, 0.2707689, 
    0.2596493, 0.2696185, 0.2385048, 0.1943103, 0.2599734, 0.2617558, 
    0.2823728, 0.232125, 0.2340069, 0.2838837, 0.2816786, 0.2173103, 
    0.1970801, 0.1647272, 0.2128638, 0.1690089,
  0.1412596, 0.1185796, 0.1166164, 0.1646336, 0.1739992, 0.1524376, 
    0.1439969, 0.1861998, 0.1899951, 0.1782987, 0.1603898, 0.163713, 
    0.1186448, 0.1583585, 0.1130943, 0.1195715, 0.1234707, 0.1199511, 
    0.1171879, 0.1441742, 0.1707809, 0.1841357, 0.1654254, 0.126283, 
    0.09108461, 0.1700934, 0.1603785, 0.1325379, 0.1312615,
  0.1107, 0.1051221, 0.05327356, 0.07436049, 0.08708251, 0.1039981, 
    0.1039737, 0.1136866, 0.08187201, 0.03135858, 0.03398484, 0.05994717, 
    0.08992712, 0.1111485, 0.1545156, 0.09300168, 0.1012414, 0.08288464, 
    0.0944899, 0.06064328, 0.09740344, 0.08433893, 0.0855825, 0.1175457, 
    0.0799392, 0.1011747, 0.115147, 0.08061387, 0.09203619,
  0.002334802, 6.018736e-05, 0.0661162, 0.1243909, 0.06212705, 0.04346328, 
    0.01550531, 0.006557033, 0.01327179, 0.001402423, 0.009688749, 
    0.03085935, 0.08736083, 0.06054818, 0.0535031, 0.03610821, 0.04671571, 
    0.05042669, 0.1696606, 0.1319234, 0.08313143, 0.03430997, 0.0002241704, 
    -3.569339e-07, 0.08593865, 0.07101049, 0.1151581, 0.05265613, 0.09464704,
  9.42077e-05, 0.02215987, 0.09654839, 0.008952991, 0.0233627, 0.0006215677, 
    0.001521256, 0.0006779379, 0.0003488745, 0.0001045774, 0.07374223, 
    0.0391744, 0.01202347, 0.03972966, 0.02458566, 0.07795035, 0.08000334, 
    0.0756033, 0.05973146, 0.04488969, -0.0001087919, 3.41727e-06, 
    1.672248e-07, -1.261815e-05, 0.07437764, 0.1663303, 0.07379465, 
    0.003548105, 2.47735e-05,
  0.008878508, 0.06336727, 0.2006263, 0.01703917, 0.03269146, 0.1073401, 
    0.1347475, 0.04755854, 0.0200986, 0.002302161, 0.02296271, 0.04231344, 
    0.08995728, 0.08064032, 0.1028668, 0.07323818, 0.04174558, 0.01371719, 
    0.0004344775, 3.41127e-07, 7.105148e-08, 5.823708e-05, 0.0003369594, 
    0.1518669, 0.08600046, 0.2761516, 0.0002065909, 2.827616e-05, 
    -1.187119e-05,
  0.07456613, 0.4153667, 0.2148957, 0.009252699, 0.001659652, 0.04771002, 
    0.04124714, 0.08807275, 0.1168662, 0.08293594, 0.01338207, 0.007026484, 
    0.02272346, 0.03606543, 0.01147334, 0.00304857, 9.410667e-05, 
    0.008550672, 0.003919498, 0.0002141367, 0.001092258, 0.006925603, 
    0.07042071, 0.1009993, 0.03346027, 0.0004884272, 0.01409987, 0.01812638, 
    0.01757983,
  0.01516637, 0.01995734, 0.01656558, 0.1016146, 0.004898401, 0.003746084, 
    0.08383869, 0.04325049, 0.1501878, 0.05270292, 0.09531727, 0.1198779, 
    0.1367734, 0.2218084, 0.1085748, 0.1157263, 0.1686536, 0.1776927, 
    0.1295111, 0.1044057, 0.1421356, 0.08042455, 0.138006, 0.04057357, 
    0.06074446, 0.1308783, 0.06478927, 0.03258007, 0.0186173,
  0.001328486, 2.700602e-07, -1.602245e-07, 0.006588283, 0.001532083, 
    0.0139278, 0.04459552, 0.06505991, 0.03292227, 0.02800969, 0.05946767, 
    0.1231317, 0.08004043, 0.05087832, 0.04034689, 0.02611657, 0.01484019, 
    0.01325552, 0.00519129, 0.05830332, 0.03468146, 0.1188584, 0.01299673, 
    0.03773259, 0.0140436, 0.03582624, 0.02483164, 0.05851155, 0.0001060016,
  0.001401915, 0.007338674, 0.02493186, 0.020418, 0.01808683, 0.003869852, 
    0.02172409, 0.1095118, 0.2629444, 0.04760084, 0.05437665, 0.1020575, 
    0.0789748, 0.01839971, 0.03409424, 0.07356001, 0.03267499, 0.05343025, 
    0.02063823, 0.01093614, 0.04157151, 0.0647888, 0.06811963, 0.0591016, 
    0.1052291, 0.03417078, 0.03478833, 0.007139947, 0.03934473,
  0.08595271, 0.0647644, 0.07660121, 0.0681738, 0.06332684, 0.01820033, 
    0.06204309, 0.04565667, 0.04420922, 0.08509297, 0.06505644, 0.06753229, 
    0.1269256, 0.1620239, 0.1737267, 0.1646938, 0.158063, 0.1710496, 
    0.03115599, 0.01858177, 0.06376179, 0.1230958, 0.1130162, 0.06702067, 
    0.1294191, 0.09140858, 0.07404976, 0.0546645, 0.06842131,
  0.1250678, 0.1784445, 0.1558175, 0.121705, 0.09341151, 0.1014809, 
    0.1269678, 0.2194915, 0.1871976, 0.1243716, 0.1692291, 0.184147, 
    0.1471501, 0.1668687, 0.1845549, 0.2887735, 0.2082011, 0.2451331, 
    0.124869, 0.1071807, 0.1083746, 0.1783429, 0.2755053, 0.2895852, 
    0.2031253, 0.140542, 0.1710827, 0.1143211, 0.1126451,
  0.2230682, 0.2462847, 0.1912598, 0.2556165, 0.2610232, 0.1614422, 
    0.1955004, 0.1938041, 0.2531681, 0.330138, 0.2468711, 0.196672, 
    0.2899727, 0.1711573, 0.213298, 0.296302, 0.2653627, 0.3685501, 0.241834, 
    0.1229128, 0.1913619, 0.1795714, 0.2422865, 0.2931936, 0.3223045, 
    0.3488269, 0.2047653, 0.2214902, 0.2542475,
  0.2497387, 0.2587794, 0.2455181, 0.3234162, 0.3100592, 0.3104751, 
    0.2905921, 0.3526253, 0.3001773, 0.234137, 0.2099916, 0.2683822, 
    0.1457957, 0.137384, 0.133396, 0.1954653, 0.2852102, 0.2584275, 
    0.2866146, 0.3235304, 0.2553214, 0.2140809, 0.1934955, 0.24021, 
    0.2684223, 0.3293992, 0.3711613, 0.2894126, 0.2350265,
  0.1275953, 0.2037445, 0.2275995, 0.2128407, 0.2613758, 0.23614, 0.2485579, 
    0.2219317, 0.1695602, 0.1046719, 0.09936847, 0.1233973, 0.1244068, 
    0.1388548, 0.1436228, 0.1068067, 0.09471075, 0.06498419, 0.09170512, 
    0.1782372, 0.230135, 0.3010184, 0.1962781, 0.1471707, 0.1505199, 
    0.1519913, 0.1554536, 0.1130863, 0.2088451,
  0.03044799, 0.02970061, 0.02895324, 0.02820586, 0.02745848, 0.02671111, 
    0.02596373, 0.02681958, 0.02582505, 0.02483052, 0.02383598, 0.02284145, 
    0.02184692, 0.02085239, 0.01866151, 0.01971105, 0.02076058, 0.02181012, 
    0.02285965, 0.02390919, 0.02495872, 0.02410449, 0.02479687, 0.02548924, 
    0.02618161, 0.02687399, 0.02756636, 0.02825873, 0.03104589,
  0.1341597, 0.03341874, 0.02632235, 0.02614591, 0.01304228, 0.003596886, 
    4.722085e-05, 0.001586924, 0.001987875, 0.026063, 0.03899927, 0.04148019, 
    0.07629806, 0.1498, 0.05248011, 0.05834666, 0.1016213, 0.1596131, 
    0.1537493, 0.1536962, 0.2647123, 0.3294888, 0.2437688, 0.3097261, 
    0.2768917, 0.229849, 0.2594435, 0.2529578, 0.2248121,
  0.2797284, 0.1871302, 0.1248515, 0.1790754, 0.1540332, 0.1701526, 0.221586, 
    0.1691577, 0.1188369, 0.1224188, 0.1585731, 0.1605041, 0.2499455, 
    0.3231669, 0.2946442, 0.2305386, 0.3045278, 0.3178524, 0.2874245, 
    0.2809967, 0.2932026, 0.2800971, 0.3608797, 0.4117731, 0.2831379, 
    0.230826, 0.25521, 0.2649965, 0.313352,
  0.2386549, 0.2249544, 0.2894261, 0.2861814, 0.2935372, 0.2529231, 
    0.2368306, 0.259833, 0.3071579, 0.2993774, 0.3075431, 0.2928223, 
    0.2866814, 0.2705083, 0.2739434, 0.2392541, 0.1944236, 0.2445961, 
    0.2509746, 0.2795199, 0.2614287, 0.2623294, 0.2969899, 0.26594, 
    0.2059103, 0.1678949, 0.1812846, 0.2211026, 0.1626697,
  0.1463087, 0.1182177, 0.1248653, 0.1826217, 0.187122, 0.1605729, 0.1576446, 
    0.1907896, 0.1777474, 0.1931459, 0.181649, 0.1645452, 0.1276409, 
    0.1518145, 0.1032517, 0.1056753, 0.1391925, 0.115743, 0.1296359, 
    0.1451684, 0.1767152, 0.1765577, 0.1636647, 0.1346551, 0.09541354, 
    0.1785842, 0.1724417, 0.1283334, 0.1403898,
  0.115422, 0.115495, 0.06083184, 0.07421651, 0.09747723, 0.1179115, 
    0.1019762, 0.114813, 0.08082831, 0.02899906, 0.03614812, 0.06154965, 
    0.09420606, 0.1177407, 0.1644682, 0.1028999, 0.1099021, 0.08278714, 
    0.1030498, 0.06401759, 0.09352887, 0.09174356, 0.08909318, 0.1322736, 
    0.075399, 0.102984, 0.1186619, 0.09878077, 0.09539434,
  0.001756363, -4.225993e-06, 0.06444012, 0.1180023, 0.06589332, 0.07016278, 
    0.02326306, 0.009714359, 0.01423051, 8.958556e-05, 0.005887602, 
    0.01378535, 0.08165537, 0.06358875, 0.04805892, 0.03363579, 0.05189553, 
    0.0539851, 0.1837462, 0.1327828, 0.09278055, 0.04258634, 0.0008305914, 
    -5.368496e-07, 0.08490308, 0.06955772, 0.1293108, 0.05239359, 0.1004842,
  5.762309e-06, 0.01323131, 0.07639781, 0.0124048, 0.02298879, 0.004418636, 
    0.002554539, -0.0001410877, 1.306855e-05, 2.733939e-05, 0.02370579, 
    0.02006154, 0.004439653, 0.04114883, 0.005763887, 0.0652947, 0.06931514, 
    0.06919663, 0.06563011, 0.04783133, 0.0006789017, 3.877464e-07, 
    7.394882e-08, -1.013858e-05, 0.07220128, 0.1785478, 0.04731205, 
    0.0002439848, 3.291347e-06,
  0.002218829, 0.03492371, 0.1672582, 0.03187821, 0.04552905, 0.1115761, 
    0.1301634, 0.04699118, 0.02356665, 0.003592204, 0.02252374, 0.0233147, 
    0.08322271, 0.06757328, 0.08209035, 0.07519005, 0.04675249, 0.01934626, 
    0.001497092, -1.057691e-07, 1.090613e-05, 2.518187e-07, 2.174285e-05, 
    0.1006716, 0.0415133, 0.1933512, 8.477211e-05, 1.585988e-07, 0.0001315433,
  0.04362011, 0.3714777, 0.1296183, 0.01256029, 0.001994581, 0.04524476, 
    0.05040628, 0.06824587, 0.1190839, 0.08134836, 0.01229572, 0.005047658, 
    0.0198188, 0.03024218, 0.01195103, 0.002059885, 0.0002441268, 
    0.002131721, 0.001556575, 0.006782134, 0.02041418, 0.01961448, 
    0.05806956, 0.06200957, 0.1532325, 0.0004749173, 0.01646134, 0.008856846, 
    0.007461349,
  0.005968236, 0.0108513, 0.008840308, 0.192835, 0.01331623, 0.007451488, 
    0.09067781, 0.03998635, 0.1409121, 0.04909251, 0.09726233, 0.1019048, 
    0.09715514, 0.1796521, 0.09319417, 0.1095773, 0.1522974, 0.1699519, 
    0.1314939, 0.1169727, 0.1393016, 0.07923272, 0.1388755, 0.03753575, 
    0.0519771, 0.1092801, 0.05568835, 0.01504315, 0.009236101,
  5.572994e-05, 8.252677e-07, 2.401215e-07, 0.001754227, 0.0003062374, 
    0.01082454, 0.0448978, 0.05376037, 0.04262824, 0.03004584, 0.05903864, 
    0.1212685, 0.07020284, 0.04608578, 0.04528775, 0.0293163, 0.01302888, 
    0.02181234, 0.008758616, 0.04571097, 0.02539768, 0.1289707, 0.0130684, 
    0.03313623, 0.01470165, 0.03450367, 0.005237434, 0.03431303, 6.404477e-05,
  0.0002939467, 0.01104615, 0.01833907, 0.02382581, 0.01239465, 0.005131895, 
    0.01603334, 0.1136032, 0.2810488, 0.02608632, 0.05566576, 0.09120855, 
    0.0816227, 0.02636933, 0.04033135, 0.07495359, 0.04002513, 0.05917843, 
    0.0235864, 0.01137862, 0.04095761, 0.05826598, 0.04887468, 0.05883662, 
    0.08747004, 0.02777661, 0.03062702, 0.01174005, 0.0297714,
  0.0754674, 0.06154039, 0.08667681, 0.09605473, 0.06590045, 0.005853401, 
    0.07113937, 0.04394655, 0.03212728, 0.07834445, 0.07669139, 0.06509374, 
    0.1331178, 0.1623344, 0.1700692, 0.1755238, 0.1611132, 0.1847586, 
    0.03356949, 0.01745437, 0.07376711, 0.1209975, 0.1092688, 0.06529827, 
    0.1414512, 0.09584387, 0.0915691, 0.06017832, 0.0715244,
  0.1305013, 0.1837509, 0.1548054, 0.1306849, 0.09756744, 0.09385853, 
    0.1240803, 0.2497752, 0.1745605, 0.1247171, 0.1784574, 0.1896094, 
    0.1498583, 0.1659698, 0.1808131, 0.2904534, 0.210686, 0.2478821, 
    0.1273983, 0.120377, 0.1142462, 0.1814095, 0.2647435, 0.2878283, 
    0.2099142, 0.1440253, 0.1723163, 0.1284395, 0.1132851,
  0.2060215, 0.2429245, 0.1947022, 0.2473064, 0.2370075, 0.188524, 0.173978, 
    0.2192184, 0.2851303, 0.3490764, 0.2914732, 0.2273445, 0.3075153, 
    0.2012857, 0.2000703, 0.3138251, 0.307084, 0.3827658, 0.2751025, 
    0.1086759, 0.1919459, 0.1797075, 0.2341831, 0.2855602, 0.3402632, 
    0.3530627, 0.1966442, 0.2091801, 0.2629513,
  0.2976465, 0.2633268, 0.254539, 0.3299341, 0.3459954, 0.3213486, 0.2693637, 
    0.3595423, 0.2950901, 0.2573544, 0.2145163, 0.2569142, 0.1611256, 
    0.1814941, 0.1593355, 0.1851973, 0.283573, 0.258719, 0.2703974, 
    0.3224109, 0.2917809, 0.2584123, 0.2090908, 0.2499916, 0.2409517, 
    0.3573927, 0.3696073, 0.2779076, 0.2624302,
  0.1806695, 0.2752109, 0.3064542, 0.2777711, 0.3102747, 0.307804, 0.2976355, 
    0.2619152, 0.1840834, 0.09585059, 0.1089228, 0.1182722, 0.1249679, 
    0.1405039, 0.1467412, 0.1036927, 0.08186023, 0.09231712, 0.1342382, 
    0.2335026, 0.2829134, 0.3223563, 0.2350266, 0.1603689, 0.1558421, 
    0.1310186, 0.1295223, 0.1260198, 0.2133751,
  0.05484225, 0.05051054, 0.04617883, 0.04184712, 0.03751541, 0.0331837, 
    0.02885199, 0.03361201, 0.03281273, 0.03201343, 0.03121414, 0.03041485, 
    0.02961556, 0.02881627, 0.01757674, 0.02247109, 0.02736544, 0.0322598, 
    0.03715415, 0.0420485, 0.04694286, 0.04999004, 0.05022668, 0.05046333, 
    0.05069997, 0.05093662, 0.05117326, 0.05140991, 0.05830761,
  0.2266804, 0.06645939, 0.04013835, 0.02802701, 0.01269293, 0.002834104, 
    0.0002297506, 0.00428468, 0.006281967, 0.03776615, 0.03884367, 
    0.07544271, 0.1235266, 0.1351142, 0.06206707, 0.05884288, 0.09710661, 
    0.1496264, 0.1567122, 0.1511071, 0.2856261, 0.4147843, 0.2716084, 
    0.2975717, 0.2759164, 0.2314434, 0.2670234, 0.2454872, 0.241751,
  0.2914391, 0.1685584, 0.1306732, 0.1852872, 0.2057456, 0.1979804, 
    0.2416539, 0.2309752, 0.1776692, 0.1675932, 0.2120173, 0.1638343, 
    0.2485176, 0.3086646, 0.284407, 0.236543, 0.2993072, 0.2904775, 
    0.2710146, 0.2927961, 0.2939881, 0.2616173, 0.3459541, 0.4503797, 
    0.3097848, 0.2370738, 0.2627436, 0.2696295, 0.307355,
  0.2413631, 0.2530217, 0.3271592, 0.3126372, 0.3232632, 0.2585931, 
    0.2641759, 0.2703223, 0.3182334, 0.3366723, 0.3258078, 0.3155358, 
    0.2818165, 0.293549, 0.2948862, 0.2611026, 0.2288123, 0.2536044, 
    0.260336, 0.3068138, 0.2832995, 0.2759631, 0.2861886, 0.2762075, 
    0.2281749, 0.1937005, 0.1842207, 0.2383591, 0.2153224,
  0.1665878, 0.1326306, 0.1426616, 0.1775742, 0.1911549, 0.1718711, 
    0.1635832, 0.1982734, 0.1808505, 0.1835572, 0.2020442, 0.2016096, 
    0.1415566, 0.1526219, 0.1059147, 0.1102605, 0.1536596, 0.1431145, 
    0.1424641, 0.1721401, 0.1948682, 0.1733945, 0.1710676, 0.1487181, 
    0.1197919, 0.1961799, 0.1973765, 0.131151, 0.1402012,
  0.1422153, 0.1261512, 0.07456425, 0.08921459, 0.1081323, 0.1293602, 
    0.1092072, 0.1242514, 0.09931526, 0.03947297, 0.05613173, 0.06013418, 
    0.1021705, 0.1223063, 0.1773075, 0.1230705, 0.1274295, 0.09625106, 
    0.1354226, 0.07894762, 0.1056694, 0.1013852, 0.1116894, 0.1480553, 
    0.07970954, 0.107978, 0.1292883, 0.1184938, 0.09841488,
  0.002618727, 2.735207e-05, 0.0459208, 0.09743606, 0.06886873, 0.09137139, 
    0.03988499, 0.008707792, 0.02298272, 4.051608e-05, 0.002528062, 
    0.006682768, 0.06702343, 0.05825673, 0.04959926, 0.03609806, 0.07703081, 
    0.05490913, 0.1958318, 0.161122, 0.09721406, 0.04938352, 0.004387467, 
    2.11539e-07, 0.06260434, 0.07469256, 0.1450131, 0.06163181, 0.1291352,
  8.90575e-07, 0.006104763, 0.02130976, 0.009878114, 0.02957589, 0.009804804, 
    0.005516765, 0.0008389937, 0.0002486843, 4.250577e-06, 0.004505255, 
    0.005077467, 0.001803252, 0.03994899, 0.003415843, 0.05905872, 
    0.05411715, 0.05758192, 0.0810298, 0.05831979, 0.003315205, 
    -1.214939e-07, 2.92449e-08, -2.768477e-06, 0.07737527, 0.1571694, 
    0.03755258, 0.0003897492, 1.577248e-06,
  0.000288377, 0.01837207, 0.09769677, 0.06094122, 0.05474872, 0.1210268, 
    0.1242536, 0.05063118, 0.02084336, 0.003908021, 0.01814101, 0.01704098, 
    0.09105855, 0.06405271, 0.07260045, 0.07526506, 0.05177116, 0.02831119, 
    0.003900719, 0.0002382432, 5.019804e-08, 1.121988e-07, 5.903689e-06, 
    0.09871445, 0.03000295, 0.08535595, 0.0001922662, 7.706209e-08, 
    1.074104e-06,
  0.03478672, 0.3272852, 0.08461855, 0.02422619, 0.003286375, 0.0410997, 
    0.04882924, 0.05844709, 0.1204242, 0.07939111, 0.01052681, 0.005472621, 
    0.01818359, 0.03042509, 0.01372281, 0.002092418, 0.003292701, 
    0.0002124617, 0.0001584167, 0.003232527, 0.007372275, 0.02058117, 
    0.04899385, 0.05575488, 0.1992292, 0.0001713071, 0.01887513, 0.008851847, 
    0.003830684,
  0.002132419, 0.004540041, 0.006020586, 0.2289605, 0.009086533, 0.01418089, 
    0.1026743, 0.04158007, 0.1409562, 0.05037329, 0.0987741, 0.09456479, 
    0.08133458, 0.1502923, 0.09039624, 0.1110409, 0.1387974, 0.1662218, 
    0.1425501, 0.124414, 0.1435525, 0.08252879, 0.1473439, 0.03505739, 
    0.04186965, 0.08287263, 0.05382755, 0.01045031, 0.004244782,
  1.21199e-05, 2.200221e-07, -3.639105e-08, 0.0009217666, 0.0005386564, 
    0.01010907, 0.04779322, 0.04858794, 0.05713458, 0.03514587, 0.06307238, 
    0.1179882, 0.06807789, 0.04206994, 0.04997259, 0.03670359, 0.01572423, 
    0.03261586, 0.01130659, 0.03945932, 0.0212808, 0.1377947, 0.01737412, 
    0.03622398, 0.01932634, 0.0359132, 0.009334518, 0.004621813, 3.026752e-05,
  -9.035915e-05, 0.01511818, 0.01730854, 0.01320346, 0.008478404, 
    0.003370318, 0.0109618, 0.1148236, 0.2920746, 0.01815238, 0.06091164, 
    0.09133138, 0.08279794, 0.03762266, 0.0483641, 0.07755768, 0.04786626, 
    0.05716303, 0.02455469, 0.01282617, 0.04141879, 0.0493898, 0.04153027, 
    0.05424678, 0.07904822, 0.02739921, 0.03327802, 0.01814924, 0.0275903,
  0.06753423, 0.06087122, 0.08907704, 0.1003522, 0.05735201, 0.003935428, 
    0.0810254, 0.03828757, 0.02213463, 0.0779666, 0.08574549, 0.06804815, 
    0.1378379, 0.1639337, 0.1698009, 0.1914385, 0.1643253, 0.1969397, 
    0.03192898, 0.02301212, 0.07836232, 0.08939391, 0.1188688, 0.06944475, 
    0.1300223, 0.08523133, 0.1051796, 0.06626388, 0.0811093,
  0.1413418, 0.1874994, 0.1513522, 0.1137386, 0.09685843, 0.1065712, 
    0.1571363, 0.2692877, 0.1666672, 0.1201514, 0.1769946, 0.1994525, 
    0.1889462, 0.1863506, 0.1996011, 0.2913501, 0.2003069, 0.2534887, 
    0.1346919, 0.1290136, 0.1094988, 0.1829303, 0.2961985, 0.294089, 
    0.2149599, 0.1458904, 0.1677396, 0.1460473, 0.1310722,
  0.2202852, 0.23616, 0.2120602, 0.2970381, 0.258872, 0.1941349, 0.2129977, 
    0.2277802, 0.2841617, 0.3498427, 0.3277242, 0.2350517, 0.3036622, 
    0.2017223, 0.2314554, 0.3399085, 0.3526256, 0.40901, 0.2887162, 
    0.09822121, 0.184972, 0.1606149, 0.25376, 0.2803008, 0.3664114, 
    0.3564106, 0.190572, 0.2318866, 0.2782326,
  0.3176714, 0.2419584, 0.2687275, 0.3396376, 0.3456683, 0.330091, 0.3358116, 
    0.3908763, 0.317784, 0.2784402, 0.2273595, 0.2650729, 0.1301176, 
    0.1512132, 0.1919959, 0.2327302, 0.292856, 0.2796914, 0.3044011, 
    0.4199337, 0.3078533, 0.2732486, 0.2499272, 0.2556835, 0.262989, 
    0.3834196, 0.356966, 0.3032047, 0.2590234,
  0.166254, 0.2646776, 0.3010565, 0.2918076, 0.3284443, 0.3185062, 0.2763699, 
    0.3237362, 0.1665632, 0.1551233, 0.1337709, 0.1383542, 0.1375999, 
    0.1332932, 0.1449443, 0.1413008, 0.135698, 0.1913898, 0.226613, 
    0.2520545, 0.3056498, 0.3869614, 0.2476742, 0.1744376, 0.1659603, 
    0.1164796, 0.1174214, 0.1496746, 0.221692,
  0.1199358, 0.114148, 0.1083601, 0.1025722, 0.09678437, 0.09099649, 
    0.08520862, 0.087462, 0.08921725, 0.09097251, 0.09272775, 0.094483, 
    0.09623826, 0.09799351, 0.09241223, 0.1011973, 0.1099824, 0.1187675, 
    0.1275526, 0.1363377, 0.1451228, 0.1439716, 0.1392191, 0.1344666, 
    0.1297142, 0.1249617, 0.1202092, 0.1154567, 0.1245661,
  0.2813914, 0.1341276, 0.0653999, 0.02771819, 0.01220063, 0.001318829, 
    0.0004175689, 0.003967458, 0.01956261, 0.04192056, 0.05065569, 0.1277758, 
    0.1764945, 0.116146, 0.05887406, 0.05844056, 0.09540616, 0.1410298, 
    0.1425396, 0.1516796, 0.3111903, 0.4495772, 0.3079218, 0.2861356, 
    0.2557662, 0.2171632, 0.2873626, 0.2504769, 0.2426558,
  0.2908956, 0.147245, 0.1206644, 0.1789511, 0.2295506, 0.2035456, 0.2713706, 
    0.2655854, 0.2192698, 0.1960593, 0.2351684, 0.1613197, 0.2507009, 
    0.2915277, 0.2825661, 0.2248311, 0.2837124, 0.2943116, 0.2734246, 
    0.2736979, 0.2740865, 0.2593616, 0.3204702, 0.4283953, 0.3081936, 
    0.2228296, 0.2636138, 0.2841889, 0.3237437,
  0.2335482, 0.2240236, 0.2953969, 0.330763, 0.3282996, 0.2651679, 0.2513632, 
    0.2596713, 0.3234045, 0.3297299, 0.3273753, 0.3036664, 0.2716172, 
    0.3209043, 0.2992586, 0.2724366, 0.2385221, 0.2575544, 0.277327, 
    0.3328407, 0.3033119, 0.2895073, 0.3095355, 0.293598, 0.2444001, 
    0.2066097, 0.1921092, 0.238464, 0.1999819,
  0.1767457, 0.1491414, 0.1455721, 0.1915311, 0.2150365, 0.2047457, 
    0.1779491, 0.2082091, 0.1862881, 0.1817412, 0.2284354, 0.230939, 
    0.1752966, 0.1764326, 0.1122958, 0.1231805, 0.2103654, 0.1576673, 
    0.1558215, 0.1991247, 0.2260008, 0.2027024, 0.1915326, 0.173652, 
    0.1268028, 0.2018647, 0.2094613, 0.1321726, 0.1561173,
  0.1586984, 0.1392051, 0.1022121, 0.1165325, 0.1294548, 0.1421091, 
    0.1240874, 0.1411804, 0.1223117, 0.0411054, 0.06072142, 0.08158698, 
    0.1081809, 0.1383487, 0.206242, 0.1484874, 0.1424834, 0.09861016, 
    0.1431017, 0.08578512, 0.1175725, 0.1147948, 0.1318092, 0.1597514, 
    0.07342265, 0.1173211, 0.1375283, 0.1550294, 0.1237171,
  0.0105804, 0.0009034738, 0.02981391, 0.07940435, 0.07591876, 0.1207371, 
    0.0473754, 0.01586269, 0.02789146, 0.0005992765, 0.0003246345, 
    0.001571407, 0.05517706, 0.05401489, 0.06002833, 0.03828698, 0.09287873, 
    0.06601803, 0.1863868, 0.1595394, 0.09642947, 0.06767658, 0.007023712, 
    1.070235e-06, 0.03942317, 0.0768529, 0.1549633, 0.05649827, 0.142319,
  3.745941e-07, 0.002671666, 0.01060929, 0.008443125, 0.04257894, 0.02116361, 
    0.01238751, 0.002931198, 0.002294879, 9.191635e-07, 0.0006915852, 
    0.001257069, 0.001134431, 0.03636934, 0.005361302, 0.05653155, 
    0.04688849, 0.0588916, 0.09971827, 0.06987031, 0.02197251, 0.00085483, 
    9.089009e-07, 1.751343e-06, 0.07582151, 0.1082611, 0.06415067, 
    0.003551306, 1.890154e-05,
  0.0001894399, 0.01405469, 0.03162726, 0.07674643, 0.05681324, 0.1334114, 
    0.1275607, 0.05415702, 0.01817639, 0.004672639, 0.01746511, 0.01202569, 
    0.1033676, 0.06276292, 0.06431001, 0.07434659, 0.05845307, 0.04022978, 
    0.01357197, 0.003054666, 4.258933e-08, 7.09592e-08, 2.525405e-06, 
    0.1025767, 0.0220136, 0.03604788, 0.002611687, 7.680902e-08, 3.337898e-07,
  0.03230971, 0.3048887, 0.06340118, 0.04734372, 0.005985683, 0.0417197, 
    0.04674586, 0.05145321, 0.1232658, 0.08612206, 0.01048512, 0.006407705, 
    0.01816742, 0.02947765, 0.01601344, 0.005075896, 0.004971249, 
    0.0006393763, 0.000645688, 0.0009772187, 0.00548673, 0.008759944, 
    0.03427474, 0.05519367, 0.1100885, 0.0002185207, 0.023602, 0.0100773, 
    0.001525551,
  0.001252054, 0.001754457, 0.00473048, 0.1710761, 0.005087866, 0.02336024, 
    0.1072647, 0.04202588, 0.1349497, 0.05270986, 0.1099117, 0.09268077, 
    0.0716646, 0.1316828, 0.08236106, 0.1053132, 0.1279873, 0.162631, 
    0.1515883, 0.1342348, 0.1415207, 0.09153308, 0.1476668, 0.03583797, 
    0.0354786, 0.06445698, 0.04991941, 0.007894012, 0.00226356,
  4.71945e-06, 6.469854e-08, -0.000103188, 0.0004950925, 0.0002692228, 
    0.008968464, 0.05099078, 0.04702064, 0.0707178, 0.04330586, 0.07062346, 
    0.1178176, 0.06562936, 0.05185895, 0.05343639, 0.04017636, 0.03045804, 
    0.03970732, 0.009751356, 0.03168585, 0.01430224, 0.1600582, 0.02077446, 
    0.03643396, 0.02257492, 0.04276274, 0.02204986, 0.000341921, 9.967699e-06,
  -9.0673e-05, 0.01573396, 0.02804364, 0.01079337, 0.007911051, 0.000484778, 
    0.008003948, 0.08519301, 0.2933621, 0.0177753, 0.07159755, 0.1009198, 
    0.08812404, 0.04917576, 0.05187424, 0.08739802, 0.05860777, 0.05353247, 
    0.02626118, 0.01205499, 0.04048591, 0.04910464, 0.03354733, 0.06430811, 
    0.07292687, 0.0358448, 0.04754197, 0.01945987, 0.02568111,
  0.0573488, 0.05580329, 0.09489795, 0.1100183, 0.05237564, 0.005572702, 
    0.08315935, 0.0327145, 0.01523608, 0.07976188, 0.08671519, 0.07295921, 
    0.1454057, 0.1625542, 0.1785015, 0.2130594, 0.1722686, 0.2036363, 
    0.03711333, 0.01417521, 0.08603258, 0.06518589, 0.1261635, 0.07966463, 
    0.1243606, 0.08715022, 0.1098116, 0.07792783, 0.09069394,
  0.1537079, 0.2035599, 0.1549721, 0.1343331, 0.1117697, 0.1030336, 0.162096, 
    0.282462, 0.1704462, 0.116304, 0.1663356, 0.211392, 0.2407035, 0.200239, 
    0.226034, 0.3112624, 0.2164302, 0.2582315, 0.1411741, 0.1329265, 
    0.1016929, 0.1804207, 0.3168287, 0.3266649, 0.219576, 0.144474, 
    0.1648561, 0.174865, 0.1486889,
  0.2314941, 0.2512129, 0.2450263, 0.3192267, 0.2825741, 0.1884198, 
    0.2086974, 0.2489752, 0.2391085, 0.3464223, 0.307915, 0.229229, 
    0.2813066, 0.1886662, 0.2403329, 0.3579845, 0.3590758, 0.4368761, 
    0.2889151, 0.1008562, 0.180049, 0.1216241, 0.2800559, 0.2709408, 
    0.3529814, 0.356537, 0.2224083, 0.2491401, 0.3073962,
  0.3438199, 0.2430975, 0.2758436, 0.3620847, 0.3605562, 0.3458405, 
    0.3426962, 0.4061994, 0.3030264, 0.2666058, 0.2315056, 0.2643071, 
    0.1269904, 0.152035, 0.1910262, 0.2875528, 0.2975478, 0.2742049, 
    0.2908737, 0.3771179, 0.2773963, 0.26827, 0.2080053, 0.2927716, 
    0.3192546, 0.4045568, 0.3561782, 0.3434351, 0.2874065,
  0.174115, 0.2460888, 0.3293005, 0.318312, 0.3403419, 0.3289856, 0.3000994, 
    0.311723, 0.1531555, 0.1162038, 0.1576266, 0.1601102, 0.1785109, 
    0.1706709, 0.180312, 0.1512942, 0.1689791, 0.1408297, 0.1958259, 
    0.214391, 0.2824864, 0.3555492, 0.2372026, 0.2097011, 0.1927235, 0.12064, 
    0.1044307, 0.1527127, 0.201336,
  0.152014, 0.1452512, 0.1384884, 0.1317255, 0.1249627, 0.1181998, 0.111437, 
    0.137973, 0.1439384, 0.1499039, 0.1558693, 0.1618348, 0.1678002, 
    0.1737657, 0.1747755, 0.1836733, 0.1925711, 0.2014689, 0.2103667, 
    0.2192645, 0.2281623, 0.2151678, 0.2070674, 0.198967, 0.1908666, 
    0.1827662, 0.1746658, 0.1665654, 0.1574243,
  0.2935669, 0.2261348, 0.09144711, 0.04123563, 0.01286655, 0.0001363856, 
    3.531025e-05, 0.00482683, 0.02667877, 0.04211257, 0.1024812, 0.1750972, 
    0.1938072, 0.08799838, 0.03828922, 0.07253923, 0.07764848, 0.1177817, 
    0.123648, 0.1311073, 0.3296509, 0.4742281, 0.353297, 0.2829602, 
    0.2622301, 0.2274929, 0.2938843, 0.2654543, 0.2471173,
  0.3028524, 0.1348536, 0.1200729, 0.1746483, 0.2489071, 0.196805, 0.2874388, 
    0.2966624, 0.2518677, 0.2119192, 0.2366474, 0.1572747, 0.245062, 
    0.2693368, 0.2545894, 0.2262751, 0.2616155, 0.2999547, 0.259914, 
    0.2662593, 0.2810911, 0.2715422, 0.3046315, 0.3941828, 0.2977858, 
    0.2335592, 0.2682846, 0.3027737, 0.3454306,
  0.2025416, 0.2395563, 0.3212078, 0.3361659, 0.3352004, 0.2780904, 
    0.2314859, 0.2453997, 0.3195662, 0.335998, 0.3537228, 0.2884867, 
    0.271413, 0.3212233, 0.2886214, 0.278371, 0.2356247, 0.2493816, 
    0.2771687, 0.3458983, 0.3052567, 0.3163803, 0.3237093, 0.2871225, 
    0.2214962, 0.1583833, 0.1538258, 0.2242798, 0.1746396,
  0.159759, 0.1553636, 0.1426172, 0.2125493, 0.2473405, 0.1952683, 0.1804788, 
    0.2219755, 0.2119256, 0.2216594, 0.2615921, 0.2466369, 0.205028, 
    0.1927028, 0.1176199, 0.1454977, 0.2133003, 0.1675738, 0.1882201, 
    0.217571, 0.2488976, 0.2428853, 0.2345995, 0.1799733, 0.08858764, 
    0.1656312, 0.2056834, 0.127235, 0.1773685,
  0.1843668, 0.1719762, 0.1232521, 0.1441032, 0.1559431, 0.1586816, 
    0.1435567, 0.1530925, 0.1389795, 0.05818627, 0.08041752, 0.1181749, 
    0.1320279, 0.1638362, 0.2575388, 0.1832705, 0.1534022, 0.1150999, 
    0.1449066, 0.09489255, 0.1314575, 0.1609108, 0.1568208, 0.1741924, 
    0.06132302, 0.1419989, 0.1510223, 0.1759784, 0.1457759,
  0.02298016, 0.005847836, 0.01647758, 0.06446089, 0.07457562, 0.1279351, 
    0.06837779, 0.03405816, 0.03411144, 0.002053221, -5.014507e-05, 
    0.0002316418, 0.04491203, 0.05921005, 0.06626739, 0.04478205, 0.08804605, 
    0.07417978, 0.1890987, 0.1565973, 0.1095912, 0.08247505, 0.01429854, 
    1.097127e-05, 0.02741672, 0.08222701, 0.1564898, 0.06567143, 0.1654522,
  5.165738e-07, 0.001132028, 0.005750478, 0.01139139, 0.05455355, 0.04553292, 
    0.02666416, 0.0164545, 0.009508071, 4.406259e-07, 0.000167749, 
    0.0002567225, 0.003891347, 0.045146, 0.004337352, 0.05443776, 0.0506867, 
    0.05933569, 0.09849048, 0.08038473, 0.05385669, 0.01302949, 0.000449103, 
    1.110981e-06, 0.06206059, 0.09611329, 0.08790121, 0.01269639, 0.001555528,
  4.814483e-06, 0.01118619, 0.01352845, 0.06531665, 0.07627962, 0.1463849, 
    0.1246281, 0.06045619, 0.02124957, 0.007089796, 0.019479, 0.009453829, 
    0.114986, 0.05545918, 0.05427426, 0.06339671, 0.05092964, 0.0404312, 
    0.01521504, 0.01046714, -3.775163e-06, 9.128654e-08, 2.162386e-06, 
    0.09710172, 0.01861654, 0.01388694, 0.01179226, 8.527067e-07, 5.355024e-07,
  0.03045269, 0.2727975, 0.05188231, 0.04809883, 0.008826517, 0.04297493, 
    0.04338337, 0.03933026, 0.1087974, 0.09264909, 0.01309251, 0.008715851, 
    0.01742863, 0.02755268, 0.01834742, 0.008805374, 0.007528744, 
    0.001483922, 0.002446054, 0.0006014938, 0.004091497, 0.006009123, 
    0.02799549, 0.05645119, 0.05012596, 0.0003848077, 0.02593271, 0.01338067, 
    0.001153171,
  0.001002233, 0.0009773602, 0.002624937, 0.1168984, 0.009010181, 0.02484795, 
    0.1082139, 0.03720588, 0.1228164, 0.05104337, 0.1066872, 0.07859733, 
    0.0598641, 0.1102943, 0.06969494, 0.09207501, 0.1154314, 0.1511021, 
    0.149298, 0.1236838, 0.1367624, 0.09649304, 0.1605012, 0.0429803, 
    0.02894433, 0.0516106, 0.04465424, 0.006078907, 0.001309655,
  2.014571e-06, 1.845321e-08, 4.850431e-05, 0.0004624833, 5.448611e-05, 
    0.006057365, 0.05077971, 0.04324165, 0.06478621, 0.04998107, 0.08680825, 
    0.1145976, 0.06280009, 0.05043684, 0.05043257, 0.03721736, 0.04002676, 
    0.05114452, 0.01167801, 0.02636505, 0.00829333, 0.1836326, 0.02149004, 
    0.03395323, 0.02145912, 0.03901595, 0.02543664, 1.143819e-05, 3.257764e-06,
  -1.965207e-05, 0.02184856, 0.04369967, 0.006158223, 0.005303572, 
    -4.070303e-05, 0.003640244, 0.06504122, 0.2688076, 0.02707379, 
    0.08983702, 0.1248595, 0.09432665, 0.06578156, 0.05624007, 0.09833823, 
    0.0675392, 0.06069772, 0.0199539, 0.01200225, 0.02225927, 0.05063776, 
    0.02701315, 0.07330535, 0.06350973, 0.0388746, 0.08319273, 0.03340022, 
    0.01651258,
  0.04644558, 0.06056906, 0.09668139, 0.1085056, 0.0350932, 0.001340211, 
    0.07633403, 0.0271466, 0.01346425, 0.08269177, 0.07346816, 0.08762924, 
    0.1560192, 0.1853826, 0.2023228, 0.2281509, 0.1945331, 0.204604, 
    0.04815545, 0.01214225, 0.1012421, 0.06405611, 0.1268786, 0.1026891, 
    0.1322514, 0.08986293, 0.1133552, 0.09153755, 0.0987986,
  0.1563894, 0.2259736, 0.1694805, 0.1433336, 0.1118134, 0.08825736, 
    0.1630999, 0.2833518, 0.1784032, 0.1144859, 0.1503238, 0.2217203, 
    0.2466232, 0.2282203, 0.2592776, 0.3397956, 0.2379657, 0.2696041, 
    0.1370384, 0.1472047, 0.1183698, 0.1900076, 0.3030757, 0.3670051, 
    0.2223414, 0.156977, 0.1826049, 0.2100848, 0.1468579,
  0.2471467, 0.2406175, 0.2351233, 0.2951327, 0.2891828, 0.1835173, 
    0.1921549, 0.2447517, 0.2445956, 0.340459, 0.3334631, 0.2346988, 
    0.2823597, 0.1848613, 0.2364893, 0.3417916, 0.4075972, 0.4446943, 
    0.2988487, 0.1106968, 0.1666928, 0.1272256, 0.2909258, 0.2584865, 
    0.3456505, 0.3683941, 0.2658088, 0.2797894, 0.3132878,
  0.3492636, 0.2553483, 0.2475747, 0.3756006, 0.3543778, 0.3565079, 
    0.3241055, 0.3707323, 0.3172596, 0.3449246, 0.2541507, 0.2282955, 
    0.1315618, 0.1923867, 0.2251506, 0.2796377, 0.2721447, 0.244289, 
    0.2826528, 0.3700902, 0.2610708, 0.255484, 0.1864891, 0.3189958, 
    0.2989625, 0.4139313, 0.3643723, 0.3615524, 0.3164264,
  0.151115, 0.218057, 0.3023131, 0.2765206, 0.2999553, 0.2912052, 0.2734705, 
    0.2609816, 0.1877038, 0.1017624, 0.1852458, 0.1299702, 0.1391363, 
    0.142822, 0.153578, 0.1365835, 0.1578681, 0.1355479, 0.1646283, 
    0.2426671, 0.2754118, 0.3282974, 0.2544057, 0.1942728, 0.184465, 
    0.1265624, 0.09698161, 0.166063, 0.1927736,
  0.2005169, 0.1936221, 0.1867273, 0.1798325, 0.1729377, 0.1660429, 0.159148, 
    0.1797582, 0.1894086, 0.1990589, 0.2087093, 0.2183597, 0.2280101, 
    0.2376605, 0.2578852, 0.2651201, 0.272355, 0.2795899, 0.2868248, 
    0.2940597, 0.3012946, 0.2723601, 0.2623696, 0.2523791, 0.2423886, 
    0.2323981, 0.2224077, 0.2124172, 0.2060328,
  0.305252, 0.3026243, 0.1184775, 0.06581964, 0.01916397, 0.00578456, 
    0.0006016368, 0.00529471, 0.03032487, 0.07609277, 0.1783132, 0.1835605, 
    0.2087909, 0.0612445, 0.04370777, 0.07213864, 0.07951802, 0.1107439, 
    0.1106431, 0.1177876, 0.3406247, 0.4796298, 0.3977962, 0.296964, 
    0.2633279, 0.2182235, 0.2939448, 0.2725799, 0.2677636,
  0.3188269, 0.1269699, 0.1182667, 0.1608812, 0.2621384, 0.2010881, 
    0.2703693, 0.3169652, 0.251853, 0.2323164, 0.2252342, 0.148614, 
    0.2499115, 0.2476294, 0.2503504, 0.2356255, 0.2801316, 0.3058265, 
    0.2946721, 0.3011576, 0.3186197, 0.2987772, 0.3288508, 0.3969119, 
    0.3023434, 0.2137655, 0.2668839, 0.3383652, 0.352557,
  0.2157589, 0.2524785, 0.32809, 0.344934, 0.3640857, 0.3067285, 0.2854262, 
    0.2870028, 0.3436964, 0.3892317, 0.3801413, 0.3080058, 0.2827831, 
    0.3285809, 0.2928259, 0.2607099, 0.2523027, 0.3037252, 0.3456085, 
    0.3828577, 0.3420503, 0.3452985, 0.3408279, 0.2745329, 0.2231831, 
    0.1823628, 0.1459316, 0.2201731, 0.1736821,
  0.1947576, 0.1879149, 0.2099007, 0.2972322, 0.2995171, 0.2208828, 0.205186, 
    0.2799196, 0.2675309, 0.2519847, 0.3147817, 0.2870423, 0.2234035, 
    0.1967856, 0.1422352, 0.1905366, 0.2277685, 0.2067262, 0.2348716, 
    0.2625112, 0.2770792, 0.259878, 0.2542138, 0.1755646, 0.07015471, 
    0.1736128, 0.236108, 0.1482865, 0.2130272,
  0.2239953, 0.206569, 0.1509962, 0.1960833, 0.2061631, 0.2122968, 0.1802108, 
    0.1954834, 0.1677413, 0.117268, 0.1427423, 0.1447436, 0.1391595, 
    0.1764262, 0.2731593, 0.1946985, 0.1729662, 0.1488257, 0.218587, 
    0.1551232, 0.1800857, 0.2155287, 0.1999961, 0.1953295, 0.06523962, 
    0.1642575, 0.1863585, 0.1892795, 0.1709298,
  0.04309552, 0.03286267, 0.01423368, 0.07451728, 0.08316393, 0.1482686, 
    0.09250938, 0.07317449, 0.03964059, 0.006599244, -0.0002676869, 
    2.823485e-05, 0.03787311, 0.06789859, 0.08466128, 0.06589621, 0.09449654, 
    0.08095924, 0.2062341, 0.1839402, 0.1207383, 0.09659231, 0.03989989, 
    7.133349e-05, 0.02306295, 0.1017178, 0.1700882, 0.08134411, 0.1817085,
  1.614845e-06, 0.0002800566, 0.002997244, 0.01337114, 0.06010216, 
    0.05655861, 0.04583577, 0.05064878, 0.02704578, -3.369569e-06, 
    4.83676e-05, 7.851465e-05, 0.006302377, 0.04160524, 0.007785854, 
    0.06507716, 0.05190522, 0.05458878, 0.08713446, 0.05860525, 0.05117508, 
    0.07095335, 0.004016125, 5.54016e-07, 0.04872201, 0.0876516, 0.1024785, 
    0.04386561, 0.005721002,
  2.521379e-06, 0.00794551, 0.008321594, 0.05081794, 0.07938585, 0.1415757, 
    0.1067695, 0.06395967, 0.02263576, 0.009415443, 0.01873269, 0.01012598, 
    0.1162881, 0.04855459, 0.04260215, 0.05284115, 0.04279065, 0.03594954, 
    0.017715, 0.01678563, 0.001238619, 1.322534e-06, 9.001784e-07, 
    0.08951035, 0.01825862, 0.006555597, 0.03009382, 0.0002430383, 
    2.220915e-06,
  0.03271963, 0.2358351, 0.04572335, 0.03838721, 0.009098727, 0.04243728, 
    0.03713077, 0.03162583, 0.09649852, 0.1104798, 0.01823122, 0.01101222, 
    0.0183659, 0.02473869, 0.02102144, 0.01113609, 0.01001276, 0.005487246, 
    0.008493762, 0.001073006, 0.002543378, 0.02154505, 0.02660551, 
    0.05444108, 0.02216126, 0.001096806, 0.02587745, 0.02161224, 0.002759523,
  0.0009474558, 0.0007144855, 0.00144639, 0.07525951, 0.009063717, 
    0.02336152, 0.1097238, 0.03130032, 0.1090928, 0.04502983, 0.09046765, 
    0.05681219, 0.04721909, 0.09139262, 0.05811341, 0.0734251, 0.09892805, 
    0.1337784, 0.1373911, 0.1036287, 0.1211373, 0.08624464, 0.168025, 
    0.05449754, 0.02473612, 0.04222643, 0.03867017, 0.006146, 0.00125707,
  1.114243e-06, 1.28596e-08, 5.486603e-05, 0.0004201136, 1.876536e-05, 
    0.0132555, 0.04678784, 0.03981668, 0.07566925, 0.07435492, 0.1140237, 
    0.1075574, 0.05665198, 0.04568676, 0.05424453, 0.03985786, 0.04374468, 
    0.08691357, 0.01738184, 0.02410612, 0.005693595, 0.2103922, 0.02379543, 
    0.03089449, 0.02271118, 0.03435893, 0.02539087, 2.427679e-05, 1.438964e-06,
  -2.986632e-06, 0.02571895, 0.02557257, 0.002101938, 0.003455278, 
    -5.203202e-06, 0.00240031, 0.04806309, 0.2664476, 0.03985944, 0.1448631, 
    0.1385545, 0.1088409, 0.08296515, 0.07296152, 0.1168203, 0.1000916, 
    0.08159607, 0.02988262, 0.01357505, 0.01553758, 0.05286998, 0.02487686, 
    0.08821016, 0.05319205, 0.04080125, 0.09606196, 0.06137385, 0.01208507,
  0.03982822, 0.0689454, 0.08620866, 0.1125788, 0.02735083, 2.698011e-05, 
    0.07594687, 0.01932924, 0.01272799, 0.0814224, 0.08185999, 0.09032749, 
    0.1830863, 0.2119871, 0.2731981, 0.270597, 0.2215603, 0.2393173, 
    0.06835187, 0.01365042, 0.07643748, 0.06856685, 0.1475677, 0.1054484, 
    0.149557, 0.09237111, 0.1337912, 0.1301343, 0.09093586,
  0.1772837, 0.2456223, 0.2017513, 0.1474603, 0.111414, 0.1117472, 0.1624108, 
    0.3040906, 0.1662675, 0.09585436, 0.141666, 0.2670959, 0.2729792, 
    0.2716349, 0.3298921, 0.3830773, 0.2710168, 0.2745423, 0.1445177, 
    0.1428614, 0.1566255, 0.2123572, 0.3372858, 0.3983217, 0.2304797, 
    0.1918193, 0.230441, 0.2435208, 0.1450665,
  0.2814516, 0.2427159, 0.2234702, 0.292496, 0.2987567, 0.1704075, 0.2036377, 
    0.2874649, 0.2649594, 0.3717245, 0.3685553, 0.2777434, 0.2721814, 
    0.1945293, 0.3297809, 0.4115731, 0.4236003, 0.4455048, 0.2987971, 
    0.1069577, 0.1856252, 0.1712238, 0.3285944, 0.2829851, 0.3813545, 
    0.3684842, 0.3120255, 0.3100939, 0.3423772,
  0.410001, 0.2929151, 0.2648141, 0.4011476, 0.3770952, 0.385125, 0.3272976, 
    0.4179972, 0.3171367, 0.3673086, 0.2801495, 0.2491689, 0.1713275, 
    0.1900432, 0.2517457, 0.2626051, 0.2821473, 0.2322179, 0.2691927, 
    0.4046848, 0.3083041, 0.296221, 0.2600642, 0.327372, 0.3626303, 
    0.4097548, 0.3433783, 0.3687976, 0.3906822,
  0.1442124, 0.243961, 0.2920505, 0.2507484, 0.2519805, 0.2839966, 0.2882394, 
    0.2588791, 0.1904433, 0.1730796, 0.201732, 0.1296007, 0.1395112, 
    0.1349761, 0.1276052, 0.1311032, 0.150336, 0.1589087, 0.1471403, 
    0.2209188, 0.2770724, 0.2882971, 0.2732385, 0.2030504, 0.1803, 0.1256072, 
    0.1074178, 0.1526966, 0.2559916,
  0.2399209, 0.2333734, 0.226826, 0.2202785, 0.213731, 0.2071835, 0.2006361, 
    0.2051182, 0.2160514, 0.2269846, 0.2379179, 0.2488511, 0.2597843, 
    0.2707175, 0.2988887, 0.3041481, 0.3094076, 0.3146671, 0.3199266, 
    0.325186, 0.3304455, 0.2930267, 0.2833815, 0.2737363, 0.264091, 
    0.2544459, 0.2448006, 0.2351554, 0.2451589,
  0.3164906, 0.3318967, 0.1849849, 0.07362615, 0.02949325, 0.02188493, 
    0.002936545, 0.004451871, 0.03049537, 0.09606802, 0.2240884, 0.1984405, 
    0.2262934, 0.0349236, 0.03143766, 0.05124947, 0.07402883, 0.1061602, 
    0.09732994, 0.1180755, 0.3586735, 0.5133092, 0.4352368, 0.3369598, 
    0.2854707, 0.2333666, 0.2843023, 0.2787767, 0.2923693,
  0.3192303, 0.1212382, 0.1251347, 0.1391483, 0.2504593, 0.2184903, 
    0.2233062, 0.3216357, 0.2515084, 0.2449536, 0.2162457, 0.1511189, 
    0.2465185, 0.2239274, 0.2564261, 0.2173175, 0.3172953, 0.3255314, 
    0.3098285, 0.3562795, 0.3292074, 0.3089769, 0.3157701, 0.4187132, 
    0.2814203, 0.2093514, 0.2832164, 0.3522913, 0.3915428,
  0.2773067, 0.2987067, 0.3577875, 0.4158783, 0.4232746, 0.3511286, 
    0.3383297, 0.330945, 0.3850189, 0.4510474, 0.3545471, 0.3234711, 
    0.3077454, 0.3327571, 0.277043, 0.2830994, 0.3170195, 0.3707003, 
    0.3649867, 0.3675218, 0.3296671, 0.2930072, 0.3174075, 0.2933916, 
    0.2622096, 0.2389148, 0.1776555, 0.2604195, 0.2332079,
  0.2764334, 0.3077758, 0.2924291, 0.3135372, 0.2996957, 0.2270189, 
    0.2431944, 0.2957395, 0.2919232, 0.3202276, 0.3678217, 0.3368814, 
    0.2623425, 0.2188658, 0.1722078, 0.2344629, 0.2594916, 0.2357559, 
    0.2820942, 0.2864407, 0.2979049, 0.2749596, 0.2667076, 0.1787272, 
    0.06151971, 0.2076307, 0.2615511, 0.1833094, 0.2696422,
  0.2720483, 0.2641838, 0.1904134, 0.2467793, 0.2478383, 0.2459845, 
    0.2531392, 0.2523443, 0.2407694, 0.1971776, 0.2324992, 0.1810686, 
    0.1545149, 0.2075328, 0.2772391, 0.2264723, 0.2611209, 0.2126886, 
    0.2641992, 0.2105225, 0.2543101, 0.2367338, 0.2155932, 0.2117006, 
    0.06713501, 0.184785, 0.2039132, 0.1886528, 0.2452459,
  0.1282949, 0.05338919, 0.01327888, 0.1019347, 0.122141, 0.197134, 
    0.1139397, 0.1226495, 0.1040648, 0.03233894, 0.0001952734, 9.153812e-06, 
    0.02452584, 0.09997773, 0.1061458, 0.08345201, 0.1131314, 0.1106492, 
    0.2189853, 0.1910192, 0.1774422, 0.1222455, 0.1301829, 8.238855e-05, 
    0.02795513, 0.1753698, 0.2264274, 0.1449932, 0.2283555,
  0.0007943575, 0.0001475484, 0.001839271, 0.0270123, 0.06560427, 0.06803861, 
    0.1074113, 0.1215358, 0.1339447, -6.407791e-05, 1.434992e-05, 
    2.59632e-05, 0.02532993, 0.03819712, 0.01777984, 0.06903079, 0.05595903, 
    0.05426092, 0.08058568, 0.0503501, 0.1135391, 0.1807183, 0.05606648, 
    2.563635e-06, 0.04486861, 0.08943978, 0.117905, 0.09327804, 0.03085601,
  3.237063e-05, 0.006923334, 0.006146593, 0.03718185, 0.0749313, 0.1191001, 
    0.09260806, 0.06113514, 0.03048369, 0.01345666, 0.01741333, 0.0155543, 
    0.1095091, 0.04294528, 0.03742906, 0.04907062, 0.03966031, 0.03346046, 
    0.02269072, 0.02974811, 0.01922948, 0.001925296, 2.627199e-06, 
    0.07976075, 0.01769625, 0.002971387, 0.07002583, 0.01021002, 9.995481e-05,
  0.04146778, 0.2194353, 0.04442324, 0.03304457, 0.01412183, 0.04317395, 
    0.03522839, 0.02724086, 0.09115739, 0.1545717, 0.02530093, 0.01273911, 
    0.02090946, 0.03136534, 0.02704683, 0.01577336, 0.009667041, 0.01362144, 
    0.02290827, 0.01396755, 0.002408764, 0.007722778, 0.02317129, 0.05261393, 
    0.008817713, 0.006870358, 0.03286217, 0.02961059, 0.009711453,
  0.0006213587, 0.0004202589, 0.0006359809, 0.04715391, 0.01163779, 
    0.0288557, 0.10107, 0.0320456, 0.1085402, 0.05721303, 0.07294515, 
    0.05234618, 0.03810912, 0.08030345, 0.04809458, 0.06177018, 0.08318932, 
    0.1171348, 0.1195039, 0.09121531, 0.105653, 0.07315614, 0.1671942, 
    0.05454373, 0.02562989, 0.04101411, 0.03649983, 0.008743105, 0.0006666891,
  7.262133e-07, 1.037156e-08, 2.347383e-06, 0.0004040775, 7.158625e-06, 
    0.006062469, 0.038996, 0.03913555, 0.08778591, 0.1381591, 0.1208768, 
    0.09581035, 0.05268783, 0.05502845, 0.05719619, 0.04367767, 0.05192716, 
    0.0864419, 0.07071131, 0.03214985, 0.005940436, 0.2181779, 0.04749765, 
    0.03161111, 0.02915523, 0.04354548, 0.03596203, 0.0003513957, 8.217404e-07,
  -1.007217e-05, 0.01412552, 0.02129598, 0.0001689609, 0.002555252, 
    2.622785e-07, 0.001397236, 0.03897181, 0.2888274, 0.04216327, 0.2616541, 
    0.2018301, 0.1419471, 0.1119286, 0.133559, 0.1732729, 0.1182678, 
    0.09816386, 0.08425407, 0.00838236, 0.01547498, 0.05236557, 0.03781971, 
    0.1240507, 0.05235652, 0.04486763, 0.1018907, 0.09152057, 0.01680594,
  0.04337682, 0.06782605, 0.08385226, 0.1314509, 0.04600871, -8.695322e-05, 
    0.07642687, 0.01461363, 0.01472586, 0.06709313, 0.09681419, 0.1091063, 
    0.2322446, 0.2586699, 0.322974, 0.2776209, 0.2540019, 0.2736405, 
    0.1116719, 0.01501135, 0.05339186, 0.07984305, 0.1667542, 0.1320595, 
    0.2033638, 0.1259327, 0.1811516, 0.1473598, 0.08805263,
  0.1980797, 0.2437756, 0.2118253, 0.1620203, 0.1127958, 0.154431, 0.1678893, 
    0.3369095, 0.1755385, 0.1031196, 0.1122256, 0.2727898, 0.3332209, 
    0.3473511, 0.3644612, 0.3932316, 0.296654, 0.2849855, 0.169013, 
    0.1314459, 0.1481353, 0.2174711, 0.3457491, 0.4114047, 0.2436363, 
    0.2496316, 0.2809226, 0.2348864, 0.1765858,
  0.3429563, 0.2429894, 0.2627807, 0.3260236, 0.3184462, 0.1769617, 
    0.2711441, 0.3463124, 0.3175645, 0.4400984, 0.395781, 0.312437, 
    0.2517537, 0.2545946, 0.5537028, 0.5276484, 0.4442926, 0.4505209, 
    0.305867, 0.1187862, 0.2223684, 0.2167223, 0.3373829, 0.342341, 
    0.4051017, 0.3707473, 0.3326109, 0.3716135, 0.3635818,
  0.4138181, 0.3267271, 0.3208319, 0.3963338, 0.4282748, 0.4466802, 0.324362, 
    0.4263393, 0.3270751, 0.4138341, 0.2938532, 0.2786912, 0.1621442, 
    0.2275528, 0.280954, 0.2673294, 0.3050863, 0.2717803, 0.3218333, 
    0.4277281, 0.3220085, 0.3846263, 0.3584373, 0.352951, 0.4045353, 
    0.4236981, 0.3330566, 0.3303242, 0.4594228,
  0.2501894, 0.3115036, 0.3274509, 0.2576383, 0.3405846, 0.3627864, 
    0.4040068, 0.2965854, 0.1981211, 0.1539707, 0.206619, 0.1373273, 
    0.1435264, 0.1383724, 0.1539109, 0.1351224, 0.1535986, 0.1967005, 
    0.1951655, 0.2746237, 0.2713985, 0.2993572, 0.2605862, 0.2184618, 
    0.2066323, 0.1384289, 0.1191881, 0.1729655, 0.2773002,
  0.2506851, 0.2451252, 0.2395654, 0.2340055, 0.2284457, 0.2228858, 0.217326, 
    0.2317873, 0.2420588, 0.2523303, 0.2626018, 0.2728733, 0.2831448, 
    0.2934163, 0.3127954, 0.3164187, 0.320042, 0.3236652, 0.3272885, 
    0.3309118, 0.3345351, 0.300548, 0.2922131, 0.2838781, 0.2755432, 
    0.2672083, 0.2588733, 0.2505384, 0.2551329,
  0.337118, 0.3509603, 0.2098309, 0.08823716, 0.03998611, 0.03764493, 
    0.01175278, 0.005218487, 0.04323441, 0.1173501, 0.2404606, 0.211035, 
    0.2258744, 0.01305033, 0.02875636, 0.04095762, 0.07897975, 0.0883279, 
    0.09059519, 0.1164542, 0.3882014, 0.5187119, 0.4596978, 0.3347841, 
    0.3288368, 0.2399096, 0.2787049, 0.2869242, 0.3161576,
  0.345573, 0.1156609, 0.125945, 0.09613618, 0.221415, 0.2335847, 0.1607412, 
    0.3183474, 0.2399513, 0.2507634, 0.2225972, 0.1551596, 0.2303734, 
    0.1953436, 0.2574037, 0.2285995, 0.3098671, 0.3544539, 0.3168648, 
    0.3763688, 0.3636883, 0.3372894, 0.3298401, 0.4338702, 0.2633157, 
    0.2474236, 0.3180768, 0.3757965, 0.4470068,
  0.3678652, 0.3700978, 0.4173804, 0.5120046, 0.4684259, 0.400389, 0.3426268, 
    0.3821442, 0.3934234, 0.4313172, 0.3378726, 0.3060997, 0.3292111, 
    0.3220628, 0.2876579, 0.3007669, 0.3453177, 0.3865812, 0.3617122, 
    0.3533096, 0.2910962, 0.2394835, 0.3113497, 0.3143736, 0.3107635, 
    0.273711, 0.2815195, 0.3339813, 0.3199734,
  0.3683469, 0.397507, 0.3526446, 0.3225936, 0.3208673, 0.261225, 0.2816751, 
    0.3181453, 0.3450978, 0.3535859, 0.3404039, 0.279543, 0.2556499, 
    0.2413849, 0.2112557, 0.2669894, 0.2996905, 0.3235348, 0.3310451, 
    0.3427002, 0.3053826, 0.3102471, 0.2772271, 0.1947941, 0.06160069, 
    0.2404744, 0.3253413, 0.2371754, 0.3448887,
  0.3321133, 0.2721713, 0.1525981, 0.2342473, 0.2512321, 0.2302106, 
    0.2887957, 0.311614, 0.387197, 0.2407618, 0.2113699, 0.1680095, 
    0.1435988, 0.2029623, 0.2598462, 0.2679732, 0.2814383, 0.2266534, 
    0.3014158, 0.2748431, 0.3496787, 0.2449146, 0.2476379, 0.2231466, 
    0.04864021, 0.1677922, 0.2136567, 0.1945428, 0.2910902,
  0.2350305, 0.05480134, 0.0129414, 0.1300988, 0.1533391, 0.222458, 
    0.1917956, 0.2160044, 0.2002721, 0.06853412, 0.001610997, 2.37583e-05, 
    0.01925999, 0.1146007, 0.1337388, 0.1419549, 0.2076983, 0.1454464, 
    0.2248033, 0.1752237, 0.1993687, 0.1694668, 0.1797536, 0.0008107986, 
    0.03245431, 0.2096249, 0.1982715, 0.1351476, 0.2507463,
  0.1243779, 0.0001003754, 0.0005645494, 0.02402988, 0.06637289, 0.07719627, 
    0.1271929, 0.1945909, 0.2611626, 0.02154303, 5.082942e-06, 6.591103e-06, 
    0.06816199, 0.07939772, 0.05185435, 0.1044524, 0.07299557, 0.07213326, 
    0.08212524, 0.07380524, 0.1362504, 0.337755, 0.1891461, -2.854734e-06, 
    0.06555977, 0.1007606, 0.119465, 0.1544806, 0.1994977,
  0.00365385, 0.004925401, 0.004584228, 0.03036644, 0.06920776, 0.1037983, 
    0.09234199, 0.1033477, 0.05246773, 0.03278613, 0.01943893, 0.02130296, 
    0.125495, 0.04900797, 0.0377344, 0.05777451, 0.05923489, 0.06090305, 
    0.04939815, 0.0581791, 0.09222663, 0.05567051, 0.0001514213, 0.067379, 
    0.01371432, 0.0007556489, 0.1043644, 0.07429573, 0.009965003,
  0.06283806, 0.2052012, 0.03254807, 0.02441436, 0.02825825, 0.04974599, 
    0.03887224, 0.03005049, 0.07881712, 0.1732524, 0.06407852, 0.01728213, 
    0.03238503, 0.04847039, 0.07432081, 0.04617561, 0.01751582, 0.01578384, 
    0.028673, 0.0443987, 0.01943372, 0.003392833, 0.007926694, 0.03711822, 
    0.004375461, 0.02235049, 0.04977784, 0.04339239, 0.02323229,
  0.0002428814, 0.0002246168, 0.0002514147, 0.0335724, 0.01099285, 
    0.06088658, 0.09096077, 0.04144798, 0.1137035, 0.06703476, 0.05745802, 
    0.06220429, 0.04129216, 0.07715598, 0.04401776, 0.05594836, 0.0737966, 
    0.1032292, 0.1090439, 0.07997425, 0.09654476, 0.06537735, 0.1570655, 
    0.05924039, 0.03734924, 0.05182557, 0.04114798, 0.02308121, 0.0001514593,
  4.979409e-07, 1.013007e-08, 5.193911e-09, 0.001242303, 1.347058e-06, 
    0.008618313, 0.02822225, 0.04105591, 0.08622564, 0.1769294, 0.1108316, 
    0.08696306, 0.05734276, 0.05617106, 0.07286733, 0.06173677, 0.06843559, 
    0.1143639, 0.1156421, 0.0538979, 0.02096983, 0.2375185, 0.06992277, 
    0.03900357, 0.04573605, 0.05701324, 0.06592901, 0.03937487, 5.048743e-07,
  -5.344195e-06, 0.006220228, 0.01686278, 5.177111e-06, 0.001728232, 
    3.578511e-07, 0.001180596, 0.03363513, 0.2951917, 0.02731076, 0.2191768, 
    0.2019759, 0.1579443, 0.1430686, 0.2124583, 0.1920397, 0.1092376, 
    0.1257826, 0.2030994, 0.02344728, 0.01771823, 0.06029505, 0.06352217, 
    0.1168139, 0.06261799, 0.06714007, 0.09719092, 0.08334277, 0.02138377,
  0.05230784, 0.03330898, 0.07243765, 0.1503755, 0.03076906, 0.0002416479, 
    0.07367382, 0.01124869, 0.01416592, 0.05808668, 0.09671082, 0.112997, 
    0.3032801, 0.3175198, 0.2962078, 0.2506802, 0.2486557, 0.262464, 
    0.1555665, 0.0125013, 0.0358928, 0.06787539, 0.1801791, 0.1101135, 
    0.2093823, 0.1769114, 0.2280531, 0.189266, 0.09201726,
  0.2409825, 0.252136, 0.2012023, 0.1464971, 0.1129432, 0.1493476, 0.1711763, 
    0.3342708, 0.1750117, 0.09975396, 0.1008256, 0.2672911, 0.3494159, 
    0.3359369, 0.3345363, 0.3881226, 0.3017438, 0.291203, 0.1901802, 
    0.1360559, 0.1348744, 0.2183136, 0.3611009, 0.3963917, 0.2567213, 
    0.3173951, 0.3293299, 0.2847241, 0.2163585,
  0.3293851, 0.2503936, 0.3120827, 0.3587545, 0.3376909, 0.2318994, 
    0.3574619, 0.3923478, 0.3880028, 0.4751232, 0.4277855, 0.3293822, 
    0.2458093, 0.3066514, 0.5837532, 0.4849907, 0.4609903, 0.4504128, 
    0.3531057, 0.1381643, 0.2118708, 0.3026047, 0.2896613, 0.3610413, 
    0.4358974, 0.3515658, 0.3608638, 0.3559353, 0.3406582,
  0.3790149, 0.3116719, 0.3487888, 0.3846569, 0.4328486, 0.4432966, 
    0.4070988, 0.4786221, 0.3585302, 0.3956066, 0.3134646, 0.3351788, 
    0.2252475, 0.2918478, 0.3017637, 0.348406, 0.3756711, 0.3357514, 
    0.3903483, 0.470217, 0.4426901, 0.4094008, 0.3580352, 0.3766854, 
    0.3316808, 0.441985, 0.3066863, 0.3083385, 0.4330147,
  0.3498905, 0.3237614, 0.3438855, 0.3136606, 0.4346947, 0.4337391, 
    0.4395994, 0.3400949, 0.2728628, 0.2622697, 0.2307851, 0.1867587, 
    0.1726984, 0.1563885, 0.2027832, 0.1905487, 0.1930971, 0.1998361, 
    0.2325605, 0.3104913, 0.3390559, 0.3231383, 0.2960791, 0.2942419, 
    0.211143, 0.1475099, 0.1268761, 0.2066571, 0.3281284,
  0.2550113, 0.2492436, 0.2434759, 0.2377082, 0.2319406, 0.2261729, 
    0.2204052, 0.237675, 0.2480085, 0.2583421, 0.2686756, 0.2790091, 
    0.2893426, 0.2996761, 0.3162931, 0.3186414, 0.3209896, 0.3233379, 
    0.3256861, 0.3280344, 0.3303826, 0.2987873, 0.2918732, 0.2849591, 
    0.278045, 0.2711309, 0.2642168, 0.2573028, 0.2596254,
  0.3548526, 0.367483, 0.2382637, 0.1071295, 0.04600915, 0.04944498, 
    0.02217541, 0.004999165, 0.05557267, 0.1327683, 0.2395567, 0.2353063, 
    0.2174888, 0.001485066, 0.02484645, 0.02688924, 0.0687141, 0.08524317, 
    0.09545041, 0.111464, 0.419804, 0.5283629, 0.4660915, 0.3080375, 
    0.3197865, 0.2615722, 0.2476605, 0.2649483, 0.3452103,
  0.3476333, 0.09794509, 0.1176335, 0.0635179, 0.1836693, 0.2227916, 
    0.09467532, 0.3021919, 0.2282269, 0.2476004, 0.224117, 0.1528811, 
    0.193824, 0.1725896, 0.2629701, 0.2641801, 0.317052, 0.3830347, 0.358238, 
    0.3710354, 0.3782203, 0.3416635, 0.3337848, 0.4430256, 0.2476078, 
    0.2894412, 0.3942746, 0.4173739, 0.4959991,
  0.4307025, 0.4457672, 0.5008392, 0.5348998, 0.4211092, 0.4057971, 
    0.3549195, 0.395768, 0.4271825, 0.3932005, 0.3053786, 0.2761855, 
    0.3416548, 0.3223792, 0.2764243, 0.2932139, 0.3765143, 0.3695827, 
    0.3990188, 0.3362319, 0.2501087, 0.2251454, 0.2807112, 0.3315913, 
    0.3156233, 0.3093393, 0.3760338, 0.4190921, 0.4194459,
  0.4777466, 0.4231772, 0.3850145, 0.3336097, 0.3429174, 0.3270432, 
    0.3258103, 0.3153285, 0.3426992, 0.3635164, 0.3107147, 0.2809595, 
    0.2190591, 0.2169157, 0.1874115, 0.2671019, 0.3291145, 0.361659, 
    0.396138, 0.4002813, 0.3585765, 0.3155352, 0.2695953, 0.2156574, 
    0.06692249, 0.2661303, 0.4185902, 0.3228185, 0.4355616,
  0.3089113, 0.2034098, 0.1479308, 0.1929417, 0.1987717, 0.1727941, 
    0.2378148, 0.3138502, 0.329397, 0.2606291, 0.1726345, 0.1347693, 
    0.09287757, 0.1952255, 0.267854, 0.3142872, 0.2761511, 0.2783455, 
    0.3124355, 0.3038541, 0.2481928, 0.2199118, 0.2457717, 0.2477269, 
    0.03888328, 0.1447739, 0.197885, 0.1972816, 0.2233678,
  0.2353572, 0.06797633, 0.01210972, 0.1309808, 0.1448631, 0.22339, 
    0.2396703, 0.3471195, 0.3092004, 0.04704798, 0.005687776, 2.273858e-05, 
    0.01400824, 0.1214533, 0.1595144, 0.1814861, 0.1857896, 0.1972961, 
    0.2181273, 0.1366193, 0.178863, 0.1641637, 0.2037746, 0.00112965, 
    0.02754762, 0.2265794, 0.1699871, 0.079676, 0.2024392,
  0.3020367, -0.0001610778, 0.0001110319, 0.05426969, 0.1170445, 0.0599215, 
    0.07764401, 0.1230306, 0.1563617, 0.02833991, 2.579468e-06, 9.788388e-07, 
    0.09719467, 0.1458519, 0.0791349, 0.160131, 0.07201421, 0.08128385, 
    0.09240544, 0.05590923, 0.1007229, 0.2935074, 0.468748, -5.741258e-05, 
    0.06305218, 0.09954491, 0.1385246, 0.1523311, 0.2883421,
  0.04519745, 0.01986405, 0.002344205, 0.02725051, 0.07873827, 0.1104355, 
    0.1044318, 0.08954494, 0.1160136, 0.1287293, 0.01973977, 0.05056895, 
    0.1336072, 0.05525441, 0.05487556, 0.06332801, 0.0946589, 0.07406431, 
    0.09923702, 0.07625235, 0.2306162, 0.4893852, 0.02714452, 0.04436458, 
    0.0069911, 0.0002373504, 0.1639756, 0.314334, 0.2316723,
  0.08379969, 0.1758841, 0.01743089, 0.02784025, 0.07031312, 0.1500548, 
    0.05255524, 0.06227887, 0.06833683, 0.1103429, 0.1037687, 0.1141284, 
    0.1238965, 0.03758427, 0.08834441, 0.09021665, 0.0337995, 0.03047062, 
    0.03560557, 0.06577708, 0.0967259, 0.02337002, 0.02414228, 0.02154682, 
    0.002037394, 0.1034649, 0.08205814, 0.101953, 0.05385899,
  0.0001002472, 0.0001080783, 0.0001130482, 0.02457404, 0.01387348, 
    0.1382399, 0.09327148, 0.06707148, 0.09686141, 0.06506566, 0.04737495, 
    0.05891021, 0.06032121, 0.07551391, 0.05326378, 0.05856989, 0.08854149, 
    0.1153975, 0.1215697, 0.1138818, 0.134955, 0.06435691, 0.1905099, 
    0.06563696, 0.08903364, 0.06145805, 0.0698857, 0.08660921, -1.572278e-05,
  3.826672e-07, 1.005512e-08, -1.484726e-08, 0.002556925, 8.842483e-08, 
    0.01646272, 0.02011648, 0.1089777, 0.06214803, 0.1307834, 0.08933818, 
    0.07365955, 0.07048309, 0.05274663, 0.06150139, 0.06806368, 0.07771484, 
    0.09666098, 0.1451818, 0.1987784, 0.04331346, 0.2375846, 0.08306158, 
    0.04564244, 0.05946986, 0.07115741, 0.09491415, 0.06876611, 3.752709e-07,
  -4.570823e-06, 0.006774869, 0.006387153, -2.664103e-05, 0.001829526, 
    1.491297e-07, 0.0008722798, 0.03125052, 0.2844987, 0.01363644, 0.1784641, 
    0.1827089, 0.1516287, 0.1341427, 0.1498973, 0.1454649, 0.08313341, 
    0.1434481, 0.2757863, 0.03035429, 0.02055242, 0.04652503, 0.06317328, 
    0.09437963, 0.05073038, 0.08908001, 0.08333005, 0.0907411, 0.02875784,
  0.06766391, 0.03253505, 0.07324706, 0.1601616, 0.01833838, 0.002156584, 
    0.07411894, 0.01002685, 0.01152302, 0.05092386, 0.1066476, 0.09089413, 
    0.2561663, 0.3015321, 0.2379037, 0.2293056, 0.2309903, 0.3224792, 
    0.2096073, 0.009696689, 0.03066609, 0.05458383, 0.1756, 0.08832766, 
    0.1942959, 0.1664368, 0.1871188, 0.1469815, 0.08744834,
  0.2584845, 0.2383174, 0.2410072, 0.1579249, 0.1421931, 0.1374681, 
    0.1808425, 0.3308586, 0.1689361, 0.1029231, 0.1060907, 0.2888034, 
    0.3529179, 0.2596769, 0.2888668, 0.3640218, 0.3052892, 0.3093295, 
    0.2272564, 0.1465392, 0.1321135, 0.2110493, 0.3715695, 0.4105272, 
    0.2602379, 0.3338091, 0.3504639, 0.2835617, 0.2419557,
  0.2542199, 0.2811289, 0.3653705, 0.4212137, 0.3817081, 0.2724715, 
    0.4354475, 0.4134392, 0.4606488, 0.4972454, 0.4244719, 0.4154173, 
    0.3002125, 0.347724, 0.4301483, 0.4263363, 0.4960183, 0.4598999, 
    0.3569371, 0.1439091, 0.2593015, 0.3365758, 0.2455648, 0.404341, 
    0.4451721, 0.3276881, 0.3239098, 0.3231297, 0.3371631,
  0.325397, 0.2326571, 0.314471, 0.3792965, 0.4481281, 0.430686, 0.4588261, 
    0.4961444, 0.3845047, 0.4206972, 0.3464804, 0.3710448, 0.3231052, 
    0.2837822, 0.3259777, 0.501792, 0.4096753, 0.3536897, 0.4312859, 
    0.4372558, 0.431279, 0.4241862, 0.3348492, 0.4237364, 0.2615819, 
    0.4688677, 0.3052601, 0.2800092, 0.4103134,
  0.3551283, 0.4025397, 0.3543845, 0.3291673, 0.4431822, 0.4402452, 
    0.4206495, 0.3965707, 0.2476829, 0.3755213, 0.3110207, 0.3168963, 
    0.2753261, 0.2147863, 0.2487374, 0.2254904, 0.2396106, 0.198948, 
    0.2724668, 0.3518654, 0.3931744, 0.3179788, 0.3233609, 0.3461114, 
    0.2418926, 0.1742473, 0.1571305, 0.3015946, 0.3177737,
  0.2571882, 0.2510844, 0.2449806, 0.2388767, 0.2327729, 0.2266691, 
    0.2205653, 0.2222541, 0.2317687, 0.2412833, 0.2507978, 0.2603124, 
    0.269827, 0.2793416, 0.2951939, 0.2967471, 0.2983002, 0.2998533, 
    0.3014064, 0.3029596, 0.3045127, 0.2936336, 0.2886696, 0.2837058, 
    0.2787419, 0.273778, 0.2688141, 0.2638502, 0.2620712,
  0.3730161, 0.3904701, 0.2437951, 0.1127155, 0.0493355, 0.05764352, 
    0.03314583, 0.002661346, 0.04959793, 0.1142429, 0.2252786, 0.273932, 
    0.2453802, -0.01021692, 0.02801658, 0.02485047, 0.06294961, 0.09905942, 
    0.1064056, 0.1434044, 0.437304, 0.5150235, 0.4642889, 0.2879903, 
    0.3203114, 0.294896, 0.2091837, 0.2311265, 0.3628449,
  0.3644099, 0.08196083, 0.1026952, 0.03857266, 0.1390138, 0.1974774, 
    0.04969588, 0.2575823, 0.2232249, 0.2254642, 0.2061939, 0.148936, 
    0.1467026, 0.1461933, 0.2748904, 0.2977194, 0.34985, 0.4194561, 0.384558, 
    0.3699968, 0.3844511, 0.3747689, 0.3359781, 0.454072, 0.2341933, 
    0.3412875, 0.4551027, 0.4883132, 0.5122565,
  0.5320949, 0.5156695, 0.5523955, 0.4445137, 0.3519958, 0.3880621, 
    0.3507805, 0.4003071, 0.4299968, 0.3419899, 0.2612588, 0.2415878, 
    0.3211089, 0.298158, 0.2442363, 0.2987819, 0.3753607, 0.4002776, 
    0.4127687, 0.3220672, 0.2282505, 0.2063564, 0.2562589, 0.3064274, 
    0.3141424, 0.3520871, 0.4190144, 0.4716537, 0.511781,
  0.4529587, 0.3882408, 0.3976503, 0.3378909, 0.3301699, 0.3327642, 
    0.3131611, 0.292337, 0.3159932, 0.338514, 0.3080807, 0.237431, 0.1806336, 
    0.1816708, 0.1788327, 0.2651291, 0.3630632, 0.3635671, 0.4282505, 
    0.4135459, 0.3490743, 0.3050098, 0.2470027, 0.2061848, 0.05506612, 
    0.2789619, 0.4855219, 0.3829552, 0.4841738,
  0.2661264, 0.1660725, 0.1162728, 0.1588078, 0.1675253, 0.1522934, 
    0.2065998, 0.2655915, 0.25598, 0.2024902, 0.1080688, 0.06148284, 
    0.06116103, 0.1814561, 0.2645939, 0.2943859, 0.293944, 0.2664353, 
    0.2636531, 0.2153432, 0.2255155, 0.226986, 0.1912524, 0.2557949, 
    0.03997649, 0.1421913, 0.1645876, 0.1421498, 0.2051726,
  0.1423545, 0.08265427, 0.01167091, 0.091663, 0.1345323, 0.1970862, 
    0.1578689, 0.2101739, 0.2340883, 0.01672232, 0.007120677, -1.214643e-05, 
    0.01154342, 0.05579085, 0.1449383, 0.1120107, 0.1497942, 0.1142842, 
    0.2154312, 0.1145965, 0.1361293, 0.08273797, 0.1436459, 0.004678502, 
    0.03189319, 0.1773457, 0.1371611, 0.04397185, 0.1505164,
  0.2762853, -0.0001950883, 3.563135e-06, 0.05278178, 0.07485001, 0.0216582, 
    0.02160864, 0.0397453, 0.05898219, 0.01717509, 6.659927e-07, 
    4.158401e-06, 0.119596, 0.08999228, 0.0930577, 0.1081451, 0.05224533, 
    0.07993435, 0.05659706, 0.02426423, 0.03265869, 0.09653558, 0.3216334, 
    0.01529773, 0.05107665, 0.09905766, 0.08110336, 0.0666514, 0.1724028,
  0.4324352, 0.08356422, 0.0008666053, 0.0408709, 0.04261837, 0.06456249, 
    0.0627214, 0.03877186, 0.04781593, 0.1673382, 0.02340631, 0.04065328, 
    0.1198436, 0.07596157, 0.03777084, 0.03854726, 0.03351055, 0.03147386, 
    0.02560381, 0.01704371, 0.07497767, 0.2809402, 0.4766115, 0.03159231, 
    0.001901017, 0.0001472819, 0.06131947, 0.1702331, 0.4891609,
  0.1916912, 0.1517815, 0.01380627, 0.03780842, 0.20868, 0.06253308, 
    0.08665995, 0.05874947, 0.07522856, 0.05502446, 0.02661163, 0.1370975, 
    0.02341736, 0.01450446, 0.01587867, 0.04885165, 0.04054424, 0.02617003, 
    0.02382679, 0.0578797, 0.2228036, 0.3530467, 0.08167151, 0.009046664, 
    0.0007067202, 0.05336004, 0.0361446, 0.09885707, 0.2910571,
  4.502666e-05, 3.182504e-05, 6.648112e-05, 0.01787805, 0.02087585, 
    0.07280958, 0.07488796, 0.03172075, 0.046633, 0.03161348, 0.02330476, 
    0.03037764, 0.04178024, 0.05434901, 0.03704095, 0.04934179, 0.061087, 
    0.07829569, 0.1022222, 0.1228542, 0.1160026, 0.07034612, 0.230157, 
    0.06203469, 0.03159264, 0.03030876, 0.05551388, 0.1130766, -3.640655e-05,
  3.224345e-07, 9.358046e-09, -9.124143e-09, 0.0005801196, 1.061296e-06, 
    0.03092266, 0.01458081, 0.03731893, 0.02994858, 0.04197603, 0.04974676, 
    0.04390139, 0.03225095, 0.04353096, 0.02722992, 0.03152414, 0.02221055, 
    0.04734941, 0.127918, 0.2068977, 0.03682589, 0.1949855, 0.01838249, 
    0.01811753, 0.01581778, 0.03832056, 0.04820181, 0.07228153, 3.162037e-07,
  -5.95708e-06, 0.006253086, 0.0004223113, 5.947359e-05, 0.002336095, 
    6.275662e-08, 0.0006606858, 0.03153214, 0.2632415, 0.009068611, 
    0.1296428, 0.1538363, 0.1291215, 0.09602182, 0.07670337, 0.10759, 
    0.04565534, 0.07656816, 0.1874505, 0.1613873, 0.02126849, 0.03303059, 
    0.03472969, 0.06909891, 0.05262356, 0.03749207, 0.0459822, 0.04529997, 
    0.03321011,
  0.05644422, 0.01934567, 0.06435739, 0.178073, 0.0135901, 0.002220568, 
    0.07317956, 0.00748726, 0.01102622, 0.04414778, 0.1257757, 0.07481763, 
    0.2110886, 0.2437906, 0.2047151, 0.2001905, 0.2315269, 0.3861359, 
    0.2388263, 0.009114778, 0.03067218, 0.05283343, 0.1624718, 0.07597245, 
    0.1682527, 0.1206535, 0.1498324, 0.1140823, 0.07423297,
  0.2183981, 0.2528844, 0.2626098, 0.1662835, 0.1477764, 0.09830964, 
    0.1776295, 0.3174733, 0.1623302, 0.09555257, 0.1205546, 0.3089796, 
    0.2894973, 0.1948872, 0.2412556, 0.3305372, 0.2793694, 0.3228754, 
    0.2539394, 0.1554634, 0.1177894, 0.1774485, 0.3634308, 0.4196057, 
    0.2350368, 0.3184938, 0.3002893, 0.2825084, 0.2414863,
  0.2070254, 0.3337428, 0.3762745, 0.4457955, 0.4467773, 0.3131098, 
    0.4432626, 0.3852917, 0.4587233, 0.4416838, 0.4066511, 0.4910318, 
    0.3174953, 0.2846382, 0.2862666, 0.3808255, 0.5484182, 0.4591794, 
    0.3644729, 0.1637948, 0.2654083, 0.3251871, 0.1913819, 0.4100476, 
    0.385347, 0.2907847, 0.2588117, 0.2868549, 0.2693759,
  0.270853, 0.1737598, 0.2978546, 0.3436362, 0.4042122, 0.3941876, 0.5223766, 
    0.4961926, 0.334288, 0.4249654, 0.3493363, 0.358731, 0.3381287, 
    0.2942737, 0.3558618, 0.5397967, 0.4280435, 0.320076, 0.4320247, 
    0.3673605, 0.4239581, 0.5126194, 0.321766, 0.4622891, 0.2100689, 
    0.4708169, 0.3033182, 0.2433179, 0.3410458,
  0.4241187, 0.378538, 0.4273211, 0.3524684, 0.4441577, 0.4404451, 0.3891426, 
    0.3997532, 0.2549536, 0.4495618, 0.4616265, 0.4611418, 0.4121714, 
    0.3294323, 0.3864809, 0.309162, 0.2776962, 0.2657393, 0.3174525, 
    0.4136677, 0.4475131, 0.3239639, 0.3063167, 0.4267786, 0.2437998, 
    0.1759776, 0.172078, 0.3136386, 0.3360311,
  0.2310605, 0.2238118, 0.216563, 0.2093142, 0.2020655, 0.1948167, 0.1875679, 
    0.1806994, 0.190689, 0.2006785, 0.210668, 0.2206576, 0.2306471, 
    0.2406366, 0.2602654, 0.2613547, 0.2624439, 0.2635331, 0.2646224, 
    0.2657116, 0.2668009, 0.2784723, 0.2746423, 0.2708123, 0.2669823, 
    0.2631522, 0.2593222, 0.2554922, 0.2368596,
  0.3803351, 0.3958192, 0.2437769, 0.1102758, 0.04708398, 0.06026174, 
    0.03500009, 0.00973139, 0.04616051, 0.07752596, 0.1874401, 0.2856665, 
    0.2849966, -0.01380521, 0.04521147, 0.04794109, 0.10548, 0.1259976, 
    0.1155507, 0.1570629, 0.4458366, 0.5118053, 0.4469048, 0.2905331, 
    0.2755714, 0.3308896, 0.1931092, 0.2076293, 0.3657596,
  0.3610727, 0.0695681, 0.08157845, 0.01989396, 0.09074996, 0.1761355, 
    0.02176079, 0.2003063, 0.2071654, 0.1932721, 0.1816157, 0.1462219, 
    0.09783442, 0.1222603, 0.2899882, 0.3364823, 0.3777139, 0.441578, 
    0.4123748, 0.4056663, 0.3923991, 0.3675306, 0.3395383, 0.4781044, 
    0.2320893, 0.4082124, 0.5241556, 0.5260856, 0.5171071,
  0.5597947, 0.533479, 0.5588974, 0.3695709, 0.2791176, 0.3196006, 0.3162708, 
    0.352888, 0.4005498, 0.2897254, 0.22379, 0.2244292, 0.2845149, 0.2707175, 
    0.2167824, 0.2687976, 0.3611018, 0.3942422, 0.3903458, 0.3090373, 
    0.2176204, 0.1743236, 0.2203258, 0.2721776, 0.2746856, 0.3923151, 
    0.4379962, 0.4876584, 0.54108,
  0.4026108, 0.3412088, 0.3430679, 0.2981787, 0.2923093, 0.2890748, 
    0.2670286, 0.2584459, 0.2936658, 0.3010267, 0.2565193, 0.197911, 
    0.1457383, 0.1355316, 0.1389555, 0.2740253, 0.3845075, 0.3681585, 
    0.4039405, 0.3890606, 0.3138701, 0.2639642, 0.207004, 0.1692675, 
    0.0469349, 0.2562914, 0.5324138, 0.3469418, 0.4382662,
  0.2206208, 0.1397049, 0.09539989, 0.1337416, 0.1455474, 0.1584235, 
    0.2158413, 0.264123, 0.2230131, 0.1627489, 0.05753365, 0.03714984, 
    0.0408311, 0.2071976, 0.2489369, 0.2654364, 0.2632126, 0.2286779, 
    0.2203085, 0.1456143, 0.1753089, 0.1810769, 0.150261, 0.245017, 
    0.03666525, 0.1194087, 0.1477247, 0.1129517, 0.2012033,
  0.08690767, 0.08629359, 0.009677663, 0.07554384, 0.116858, 0.1429652, 
    0.08834431, 0.07272176, 0.09719442, 0.006517177, 0.005864269, 
    -4.509593e-05, 0.011415, 0.03270256, 0.1106145, 0.08579957, 0.1061129, 
    0.05943393, 0.1979889, 0.09850532, 0.06991159, 0.03016436, 0.0609746, 
    0.009884887, 0.0318617, 0.1621178, 0.1281306, 0.03045224, 0.1124182,
  0.1695471, 7.36122e-05, -3.811588e-05, 0.02571674, 0.01944635, 0.008346023, 
    0.004721594, 0.01337893, 0.02039605, 0.00587883, 2.996242e-08, 
    -1.05994e-07, 0.04453041, 0.04941241, 0.0335298, 0.07026038, 0.02730367, 
    0.03462704, 0.03380956, 0.0103448, 0.00809125, 0.03373716, 0.1199119, 
    0.02318413, 0.03768375, 0.1016919, 0.03726421, 0.0168407, 0.1206836,
  0.4890782, 0.190849, 0.0003008558, 0.08321707, 0.01839749, 0.02486331, 
    0.03324694, 0.02185496, 0.01204363, 0.03224509, 0.01043566, 0.02170249, 
    0.08710568, 0.02398353, 0.01229116, 0.01650047, 0.005654124, 0.004781575, 
    0.003281303, 0.002394411, 0.01981278, 0.09451485, 0.4401004, 0.02694745, 
    0.0007612836, 5.003715e-05, 0.01257343, 0.05098768, 0.2025438,
  0.1659809, 0.1279447, 0.01281307, 0.03881389, 0.0986384, 0.02203423, 
    0.01678215, 0.02041291, 0.07341768, 0.02549475, 0.004957477, 0.02054021, 
    0.005686906, 0.002402904, 0.003640941, 0.008221706, 0.01102693, 
    0.0138371, 0.007594571, 0.02125591, 0.109708, 0.497777, 0.3734337, 
    0.0051688, 0.0002958559, 0.01435422, 0.006402344, 0.03012902, 0.212348,
  2.43552e-05, 2.700923e-05, 5.621185e-05, 0.01398256, 0.03205284, 
    0.009361638, 0.04728953, 0.01127779, 0.02429774, 0.006285787, 
    0.009928917, 0.01131085, 0.02293274, 0.02856121, 0.02203975, 0.02892125, 
    0.03965618, 0.06415619, 0.06593841, 0.05487514, 0.06685991, 0.03913671, 
    0.2906588, 0.04547868, 0.007951778, 0.01491002, 0.0143977, 0.03812081, 
    -6.436079e-05,
  2.897515e-07, 7.857627e-09, -7.787903e-09, 0.0001141598, 1.817924e-06, 
    0.03397495, 0.01431939, 0.01115122, 0.02233231, 0.01274554, 0.02831288, 
    0.02764878, 0.01064357, 0.0154448, 0.009076747, 0.006592678, 0.004226268, 
    0.02853461, 0.05070076, 0.1185122, 0.04825668, 0.151257, 0.003005421, 
    0.001811703, 0.002722759, 0.00952597, 0.01176374, 0.05433367, 2.830351e-07,
  -6.639639e-06, 0.004657365, 0.0001023451, 0.0003525511, 0.0009645867, 
    4.119391e-08, 0.0004900335, 0.02620674, 0.2367415, 0.008948582, 
    0.0979975, 0.1248916, 0.08769684, 0.06339749, 0.04480304, 0.05959996, 
    0.01442411, 0.03041552, 0.08334754, 0.1603562, 0.01871085, 0.02625787, 
    0.02231076, 0.03411948, 0.02766736, 0.0106085, 0.0171364, 0.01553487, 
    0.03783738,
  0.04316799, 0.01081483, 0.04377692, 0.1734538, 0.003685153, 0.001408508, 
    0.06580482, 0.005541749, 0.008604235, 0.04051725, 0.1254159, 0.05608253, 
    0.1759682, 0.2039471, 0.1693659, 0.1766383, 0.2647589, 0.3853007, 
    0.3471543, 0.008239079, 0.02815577, 0.05006818, 0.1427684, 0.06626269, 
    0.1448451, 0.1023721, 0.1338105, 0.1169967, 0.05334056,
  0.1468977, 0.2590922, 0.2394663, 0.1566105, 0.1197679, 0.08950715, 
    0.1532804, 0.2988761, 0.1439826, 0.09798768, 0.116933, 0.3099183, 
    0.2248392, 0.1532511, 0.1877189, 0.2810943, 0.2360847, 0.3572485, 
    0.299753, 0.178946, 0.1077267, 0.1386081, 0.3199302, 0.4276868, 
    0.2125244, 0.2816591, 0.2497789, 0.2590773, 0.1869276,
  0.1673813, 0.3954862, 0.3790882, 0.4659372, 0.5057385, 0.3250068, 
    0.4185221, 0.3678218, 0.4247935, 0.3835746, 0.3998594, 0.5175208, 
    0.3148512, 0.2206068, 0.1966204, 0.3324983, 0.6108109, 0.4337275, 
    0.4284116, 0.2006099, 0.2937215, 0.2966107, 0.1503872, 0.3683012, 
    0.314012, 0.2552902, 0.2075921, 0.226587, 0.2144469,
  0.2194383, 0.1330295, 0.3053226, 0.2902212, 0.36427, 0.3443404, 0.5965112, 
    0.5447671, 0.3033631, 0.3715716, 0.3734144, 0.3905668, 0.3202656, 
    0.3386223, 0.3492658, 0.4762123, 0.4692856, 0.3406734, 0.4026604, 
    0.2880783, 0.4369906, 0.5747729, 0.4066108, 0.4750756, 0.1532303, 
    0.4469776, 0.3207349, 0.1898454, 0.2833403,
  0.3855137, 0.380996, 0.4571037, 0.3492145, 0.4555629, 0.4263399, 0.3802939, 
    0.4063704, 0.3641038, 0.5178471, 0.5246773, 0.4909732, 0.5019584, 
    0.4334381, 0.4851193, 0.416676, 0.3799258, 0.3781343, 0.4679258, 
    0.5409523, 0.5041812, 0.3023648, 0.2979313, 0.4863889, 0.2150163, 
    0.2012375, 0.1823023, 0.3187691, 0.383112,
  0.1843703, 0.1787973, 0.1732242, 0.1676512, 0.1620781, 0.1565051, 
    0.1509321, 0.1239104, 0.1330797, 0.142249, 0.1514183, 0.1605875, 
    0.1697568, 0.1789261, 0.1949097, 0.1956998, 0.1964899, 0.1972801, 
    0.1980702, 0.1988603, 0.1996505, 0.2186547, 0.2142683, 0.2098819, 
    0.2054955, 0.2011091, 0.1967227, 0.1923364, 0.1888288,
  0.3674456, 0.3804931, 0.2073226, 0.100974, 0.040221, 0.04598275, 0.0159068, 
    0.01315737, 0.03105015, 0.04144007, 0.1080382, 0.2130934, 0.3287604, 
    -0.01132282, 0.06252729, 0.09341342, 0.1951789, 0.164823, 0.1155062, 
    0.1491439, 0.4278047, 0.5110667, 0.3915699, 0.2645764, 0.2428415, 
    0.3683143, 0.1715574, 0.1837407, 0.3480844,
  0.3472968, 0.05959065, 0.07119333, 0.009437041, 0.05043772, 0.141888, 
    0.008407562, 0.1355366, 0.1804211, 0.1555977, 0.1455208, 0.1480114, 
    0.06441573, 0.09909916, 0.3001019, 0.3681021, 0.4213713, 0.4350833, 
    0.3940333, 0.4216258, 0.3716394, 0.3461171, 0.2976855, 0.4554196, 
    0.2293987, 0.4473243, 0.5388594, 0.5050346, 0.4983655,
  0.5201539, 0.4835168, 0.5238839, 0.2943535, 0.2136551, 0.2662957, 
    0.2702444, 0.3023308, 0.3356052, 0.2417916, 0.1885447, 0.1983026, 
    0.2400132, 0.2473758, 0.1775213, 0.2397813, 0.3240568, 0.353164, 
    0.3496068, 0.2755696, 0.1873364, 0.1418523, 0.1875553, 0.2302594, 
    0.2429254, 0.4258634, 0.4390547, 0.4910573, 0.4994695,
  0.3526362, 0.3013011, 0.2677057, 0.2493922, 0.2544954, 0.2309318, 0.220634, 
    0.2105169, 0.2622831, 0.251365, 0.1983642, 0.1644991, 0.1034433, 
    0.09896511, 0.1087583, 0.2550508, 0.3379929, 0.3186949, 0.3444726, 
    0.3383093, 0.259739, 0.1965477, 0.1628107, 0.1301553, 0.03955556, 
    0.2406447, 0.5259184, 0.3145465, 0.4086033,
  0.1763624, 0.1082436, 0.06998944, 0.1193231, 0.1156597, 0.1304398, 
    0.1789312, 0.219084, 0.1875292, 0.116426, 0.03453054, 0.02230081, 
    0.02968293, 0.1444752, 0.2175097, 0.226067, 0.2038602, 0.1849562, 
    0.1934191, 0.1208747, 0.1240897, 0.1366336, 0.1125213, 0.2304128, 
    0.03996313, 0.1030948, 0.1243267, 0.09376052, 0.1721915,
  0.04869201, 0.03747248, 0.005860398, 0.05535527, 0.08437976, 0.09876565, 
    0.04754371, 0.03077762, 0.04337807, 0.003359403, 0.003497594, 
    -0.0001309988, 0.01138634, 0.02463586, 0.07512075, 0.05713753, 
    0.08125684, 0.037462, 0.1573664, 0.07952753, 0.0398223, 0.009264952, 
    0.02649544, 0.006929416, 0.0293077, 0.1142628, 0.1059985, 0.02188911, 
    0.08734886,
  0.07017911, 0.008118604, -2.940913e-05, 0.006350369, 0.005913589, 
    0.004235639, 0.001283863, 0.005140099, 0.009006865, 0.003020234, 
    3.982888e-08, -2.502234e-07, 0.01615676, 0.02092989, 0.01108617, 
    0.04191176, 0.01278012, 0.01402622, 0.01645161, 0.007689633, 0.002876795, 
    0.01327378, 0.05146346, 0.02390958, 0.02341335, 0.08950631, 0.01845926, 
    0.007138616, 0.05807308,
  0.2076699, 0.07599694, 0.0001654736, 0.1246134, 0.004703086, 0.00606602, 
    0.01358597, 0.01084878, 0.002967114, 0.0097594, 0.004394636, 0.003160653, 
    0.04588736, 0.005255544, 0.00333907, 0.005239195, 0.001286942, 
    0.0009972092, 0.001211366, 0.0009405335, 0.007164392, 0.03375256, 
    0.1822033, 0.02441758, 0.0004748927, 2.962171e-05, 0.00326816, 
    0.01813519, 0.07913177,
  0.04499466, 0.1318178, 0.01040391, 0.02788546, 0.01989746, 0.01095339, 
    0.00721772, 0.006492118, 0.06564814, 0.0164575, 0.001512835, 0.00551235, 
    0.001384433, 0.0004615966, 0.001114722, 0.003017348, 0.001477623, 
    0.002404067, 0.0005790727, 0.003538902, 0.03242739, 0.2077613, 0.2433252, 
    0.004198605, 0.0002063266, 0.00419328, 0.001122789, 0.004272378, 
    0.06194205,
  2.074611e-05, 2.355253e-05, 3.635462e-05, 0.008183712, 0.03927974, 
    0.002560124, 0.03289022, 0.004325867, 0.01330209, 0.0007302889, 
    0.004604227, 0.004359439, 0.01078409, 0.0157517, 0.00951029, 0.007182777, 
    0.01751057, 0.03574685, 0.03428929, 0.0153826, 0.03396238, 0.01136175, 
    0.2744969, 0.0298094, 0.003108195, 0.004474614, 0.00381079, 0.006149155, 
    -8.275827e-05,
  2.661796e-07, 6.11496e-09, -5.679788e-09, -9.640782e-06, 8.08998e-07, 
    0.01337258, 0.01471156, 0.0030449, 0.0145702, 0.005006333, 0.01393634, 
    0.008940121, 0.00321128, 0.005088328, 0.002245321, 0.001389688, 
    0.001070645, 0.01034417, 0.0168511, 0.05815528, 0.01239787, 0.1159064, 
    0.001037009, -0.0006076457, 0.0005960524, 0.002802236, 0.004384632, 
    0.0175593, 2.652856e-07,
  -1.040299e-05, 0.002317101, 1.87417e-05, 0.00024262, 0.0002316853, 
    3.659657e-08, 0.000326314, 0.02437291, 0.2107306, 0.009893461, 
    0.07196173, 0.07992462, 0.05054293, 0.02687928, 0.02598886, 0.03222879, 
    0.005778817, 0.01440942, 0.04503158, 0.1154914, 0.01509535, 0.02129225, 
    0.01991332, 0.01230896, 0.0139104, 0.003972383, 0.00657339, 0.006008253, 
    0.03659894,
  0.03595784, 0.004411463, 0.02684577, 0.1701976, 0.000303369, 0.0005913906, 
    0.0534248, 0.003811287, 0.008848034, 0.03534857, 0.1155407, 0.03793374, 
    0.1370728, 0.1707723, 0.1350959, 0.1522944, 0.2576861, 0.3147491, 
    0.2558136, 0.006533776, 0.02563123, 0.04302674, 0.1301015, 0.05917626, 
    0.1104253, 0.08632025, 0.09858607, 0.09145312, 0.03871054,
  0.09227265, 0.2566509, 0.2174132, 0.181699, 0.09653737, 0.08939716, 
    0.1161228, 0.2614377, 0.1139097, 0.08929314, 0.1131321, 0.3034024, 
    0.1811196, 0.1127244, 0.146295, 0.2381112, 0.2040959, 0.3453299, 
    0.3185851, 0.1973673, 0.09764376, 0.1055913, 0.2677889, 0.4203401, 
    0.1840435, 0.2443265, 0.225881, 0.2120584, 0.1373283,
  0.1368573, 0.4035695, 0.3440952, 0.4668694, 0.5227889, 0.3148418, 
    0.3649424, 0.3530752, 0.3772958, 0.3463728, 0.3460941, 0.5078573, 
    0.2971802, 0.1911764, 0.1410553, 0.2865479, 0.6243805, 0.3966365, 
    0.446984, 0.2028955, 0.2807149, 0.2645125, 0.12476, 0.3475529, 0.2559249, 
    0.2159188, 0.1724656, 0.1857956, 0.178352,
  0.1830108, 0.1016776, 0.2994751, 0.2385393, 0.3225996, 0.2932013, 
    0.6317959, 0.553229, 0.2705064, 0.355395, 0.3782237, 0.3693486, 
    0.3283997, 0.2998402, 0.3814027, 0.4107673, 0.5051634, 0.3735882, 
    0.3666481, 0.2271857, 0.4144586, 0.5730149, 0.4513459, 0.5030844, 
    0.1104731, 0.4122053, 0.3433083, 0.1363496, 0.2437192,
  0.3976059, 0.3262284, 0.4631885, 0.3548166, 0.4277827, 0.421524, 0.4320225, 
    0.4407235, 0.4433292, 0.5659149, 0.5563015, 0.5387928, 0.5282356, 
    0.4574879, 0.5177131, 0.5231596, 0.5120499, 0.5678525, 0.6016268, 
    0.6416252, 0.5579097, 0.2790755, 0.3008505, 0.5230861, 0.2041263, 
    0.2164503, 0.1779025, 0.3545901, 0.4409034,
  0.1317762, 0.1260053, 0.1202343, 0.1144634, 0.1086924, 0.1029215, 
    0.09715056, 0.08191349, 0.08672308, 0.09153268, 0.09634227, 0.1011519, 
    0.1059615, 0.110771, 0.1148198, 0.119002, 0.1231843, 0.1273666, 
    0.1315489, 0.1357311, 0.1399134, 0.1624064, 0.1591855, 0.1559646, 
    0.1527437, 0.1495227, 0.1463018, 0.1430809, 0.136393,
  0.3284261, 0.338142, 0.160108, 0.089439, 0.03139071, 0.02992538, 
    0.01089635, 0.01070095, 0.01934653, 0.02251487, 0.0591326, 0.1534093, 
    0.2938079, -0.005874491, 0.09852487, 0.246166, 0.3121945, 0.2324903, 
    0.1180865, 0.1476417, 0.3938483, 0.4974664, 0.3183858, 0.2211862, 
    0.2428679, 0.3884556, 0.1540124, 0.1639387, 0.3215846,
  0.334359, 0.05330861, 0.06295458, 0.007283316, 0.02765848, 0.1103104, 
    0.003974995, 0.09163138, 0.1301154, 0.1177504, 0.1055048, 0.1380834, 
    0.04449311, 0.07958162, 0.2902619, 0.3502942, 0.4081123, 0.4127163, 
    0.3551096, 0.4004053, 0.3108341, 0.3326168, 0.2622356, 0.3983217, 
    0.1976372, 0.4431083, 0.4832699, 0.4547213, 0.4703606,
  0.4500626, 0.3965822, 0.4326918, 0.2192464, 0.1505217, 0.1959615, 
    0.2356386, 0.2453647, 0.2639765, 0.1908628, 0.1528861, 0.151105, 
    0.1994272, 0.2030813, 0.1310562, 0.1918362, 0.257356, 0.306296, 
    0.2959459, 0.2297607, 0.1506011, 0.1190065, 0.1543135, 0.180007, 
    0.2334828, 0.4098641, 0.4135271, 0.4413834, 0.4251314,
  0.313277, 0.2626157, 0.2049747, 0.203299, 0.2091816, 0.1763368, 0.1644337, 
    0.1677815, 0.2102517, 0.1899698, 0.1392154, 0.1145836, 0.05940628, 
    0.06852575, 0.08153842, 0.1976223, 0.2657002, 0.2369453, 0.2621078, 
    0.2568716, 0.1966328, 0.1289346, 0.1089678, 0.09888691, 0.03213805, 
    0.2148406, 0.4558401, 0.2905523, 0.3881733,
  0.1338459, 0.0711989, 0.0506359, 0.1009053, 0.08631094, 0.09222398, 
    0.1223042, 0.158105, 0.1462168, 0.07565964, 0.02324608, 0.01222053, 
    0.02203292, 0.09609912, 0.1789242, 0.1770585, 0.157752, 0.1474494, 
    0.1576957, 0.09669973, 0.08423357, 0.1011226, 0.07903518, 0.2087687, 
    0.03910518, 0.08565578, 0.0961198, 0.07341108, 0.1287077,
  0.02520263, 0.01998213, 0.003853281, 0.03344831, 0.04963613, 0.06421232, 
    0.02454084, 0.01684175, 0.02491746, 0.002122984, 0.001758367, 
    -0.0001708878, 0.00830746, 0.01697376, 0.04691502, 0.03156907, 
    0.05633449, 0.02613626, 0.1238082, 0.05589371, 0.01921193, 0.004088819, 
    0.01336111, 0.004479915, 0.02364826, 0.07276349, 0.07862532, 0.01399568, 
    0.05623953,
  0.03545091, 0.006284441, -1.490964e-05, 0.002562126, 0.0008041187, 
    0.001762357, 0.0006703201, 0.002664239, 0.005250334, 0.001900912, 
    3.734165e-08, -8.387185e-08, 0.006716653, 0.00763438, 0.003657448, 
    0.01510544, 0.005723108, 0.005962552, 0.009452425, 0.003847108, 
    0.001478969, 0.006804011, 0.02794014, 0.0106601, 0.01414648, 0.07746477, 
    0.008006546, 0.003015067, 0.02740223,
  0.102362, 0.02783059, 7.96894e-05, 0.1171264, 0.0008624886, 0.001331649, 
    0.004473642, 0.00383817, 0.001361749, 0.004944838, 0.001614118, 
    0.0008399826, 0.02160618, 0.001919945, 0.001484285, 0.002538208, 
    0.0003342382, 0.0004927638, 0.0007052494, 0.0005189021, 0.003771608, 
    0.01673026, 0.09574892, 0.02247517, 0.0002398507, 1.436758e-05, 
    0.001743266, 0.00913536, 0.0376812,
  0.01874609, 0.1285335, 0.01329319, 0.0177906, 0.008569008, 0.00479023, 
    0.003019282, 0.003389285, 0.05168714, 0.01521254, 0.0008035973, 
    0.00255149, 0.000596556, 0.0002211069, 0.0005216138, 0.001574825, 
    0.0006088225, 0.000408072, 0.0001773291, 0.00118569, 0.01070715, 
    0.09569547, 0.1402947, 0.005655022, 0.0001094171, 0.001963077, 
    0.0002626701, 0.001516658, 0.0265641,
  5.205937e-06, 9.609474e-06, 1.751929e-05, 0.01063258, 0.02862345, 
    0.001324643, 0.01938894, 0.002438826, 0.005629052, 0.0001573419, 
    0.002144854, 0.001798326, 0.004050516, 0.007885753, 0.003582186, 
    0.001824818, 0.006900754, 0.01873297, 0.01935458, 0.005039025, 
    0.01755741, 0.002751053, 0.2184651, 0.02240077, 0.001540552, 0.001360586, 
    0.001602666, 0.002320729, -0.0001732096,
  2.476353e-07, 5.406067e-09, -3.963894e-09, -6.212032e-06, -1.78194e-07, 
    0.005815398, 0.01072631, 0.001404875, 0.01181528, 0.002255111, 
    0.005981207, 0.00279935, 0.001281492, 0.001990365, 0.0005724371, 
    0.0006630686, 0.0004421044, 0.003662545, 0.006564729, 0.03712253, 
    0.005471683, 0.09323296, 0.0005869116, -0.0007551273, 0.0002840651, 
    0.001293169, 0.002318652, 0.009677013, 2.567462e-07,
  -6.664088e-06, 0.002059735, 1.087516e-05, 5.238592e-05, -0.0002041725, 
    3.460148e-08, 0.0001732039, 0.02271132, 0.1866366, 0.005164408, 
    0.04831948, 0.05234104, 0.02821684, 0.01214711, 0.01152964, 0.02212034, 
    0.002197081, 0.007690226, 0.02694866, 0.08314894, 0.01377422, 0.01640621, 
    0.0156104, 0.01318335, 0.004922477, 0.001860272, 0.002757594, 
    0.003026213, 0.03449955,
  0.02647754, 0.001990393, 0.01658354, 0.1634121, -0.0005805494, 
    0.0002992589, 0.03933174, 0.002823959, 0.006190402, 0.03006777, 
    0.1045661, 0.02692069, 0.1052712, 0.1357377, 0.1040547, 0.1224, 
    0.2042726, 0.2257994, 0.1756794, 0.006571854, 0.02215899, 0.03172197, 
    0.106831, 0.04952009, 0.07452352, 0.05180882, 0.06775288, 0.05945178, 
    0.02387006,
  0.05687686, 0.2290998, 0.1822332, 0.1752262, 0.08378954, 0.07335594, 
    0.08657455, 0.2141637, 0.08913453, 0.07505701, 0.1037994, 0.2747622, 
    0.1412649, 0.08081529, 0.1056448, 0.1869399, 0.1740304, 0.3186297, 
    0.2708855, 0.2026128, 0.082629, 0.07753285, 0.2152407, 0.38962, 
    0.1455884, 0.2239735, 0.205284, 0.176686, 0.1023177,
  0.106044, 0.381785, 0.2928179, 0.4302992, 0.4905599, 0.274181, 0.3029695, 
    0.3021569, 0.3158026, 0.2937415, 0.2888223, 0.4662507, 0.2671353, 
    0.1718593, 0.1049206, 0.2376119, 0.6097803, 0.351459, 0.4171115, 
    0.1834332, 0.2541639, 0.2269698, 0.09986743, 0.3086088, 0.21409, 
    0.1752553, 0.146858, 0.1508695, 0.1378374,
  0.1532021, 0.06995106, 0.2885955, 0.1808601, 0.2690092, 0.2340097, 
    0.6074622, 0.4963141, 0.2268698, 0.322467, 0.3706194, 0.366749, 
    0.3436837, 0.2921965, 0.4107405, 0.3515751, 0.4620952, 0.37926, 
    0.3053781, 0.1751672, 0.3755108, 0.5287977, 0.4725415, 0.4740745, 
    0.08807847, 0.3455154, 0.3792543, 0.09961526, 0.2091815,
  0.3763397, 0.2606961, 0.484458, 0.3990683, 0.3846017, 0.4249827, 0.4862723, 
    0.5167097, 0.5516369, 0.5948426, 0.5712769, 0.5726282, 0.5576277, 
    0.4855705, 0.5281685, 0.5790887, 0.5687687, 0.591994, 0.609702, 
    0.6041862, 0.5693883, 0.2779867, 0.3060635, 0.5504619, 0.1826865, 
    0.2121254, 0.1602055, 0.3415973, 0.4367452,
  0.0978635, 0.09329613, 0.08872876, 0.08416137, 0.079594, 0.07502662, 
    0.07045925, 0.05577606, 0.05688602, 0.05799598, 0.05910594, 0.0602159, 
    0.06132586, 0.06243581, 0.06491373, 0.06981672, 0.07471973, 0.07962272, 
    0.08452571, 0.08942872, 0.09433171, 0.1078801, 0.1064346, 0.104989, 
    0.1035434, 0.1020978, 0.1006522, 0.09920666, 0.1015174,
  0.2981948, 0.2801494, 0.1247899, 0.07394078, 0.02773551, 0.01733873, 
    0.004205813, 0.006597324, 0.01510009, 0.01836628, 0.0317625, 0.07218969, 
    0.2025646, -0.00309687, 0.157812, 0.3539811, 0.3801337, 0.2394822, 
    0.1047846, 0.1690127, 0.3463059, 0.5087304, 0.2582676, 0.1695365, 
    0.2353082, 0.4180887, 0.1399607, 0.1397032, 0.2829406,
  0.3061183, 0.04677675, 0.05425525, 0.004588242, 0.01328048, 0.0876986, 
    0.001828512, 0.0675957, 0.07846848, 0.09048283, 0.08308847, 0.1139553, 
    0.03155175, 0.06528261, 0.2665494, 0.3100634, 0.3517935, 0.3508406, 
    0.3146017, 0.34748, 0.2627622, 0.2865821, 0.2148829, 0.3342162, 
    0.1782474, 0.4131449, 0.4016457, 0.3830043, 0.4228344,
  0.3651023, 0.3212055, 0.3421479, 0.1653421, 0.1103316, 0.1426472, 0.189943, 
    0.1889158, 0.206445, 0.1438281, 0.1160079, 0.1115967, 0.15798, 0.1614652, 
    0.09340429, 0.1462697, 0.2016709, 0.2503206, 0.2397658, 0.1763297, 
    0.1140782, 0.09250167, 0.1161149, 0.1308537, 0.1940519, 0.3334509, 
    0.3456255, 0.3653783, 0.3480223,
  0.2688177, 0.211438, 0.164218, 0.1640187, 0.1686747, 0.1307484, 0.1218596, 
    0.1303577, 0.1596379, 0.133945, 0.09431286, 0.07365496, 0.0344093, 
    0.04161798, 0.05413237, 0.1358922, 0.1950647, 0.1534759, 0.1771247, 
    0.1847212, 0.1334197, 0.08276701, 0.068562, 0.07741467, 0.02358185, 
    0.1615305, 0.3765832, 0.2429145, 0.3404449,
  0.09192476, 0.04585771, 0.03593036, 0.06948353, 0.0556216, 0.05912973, 
    0.07763186, 0.1008173, 0.0971604, 0.0471015, 0.01669785, 0.006698298, 
    0.0154023, 0.06293029, 0.1438873, 0.1190429, 0.1071324, 0.1076837, 
    0.116273, 0.07258616, 0.05879556, 0.07259215, 0.04697775, 0.1870093, 
    0.03692335, 0.06270534, 0.0622391, 0.05476601, 0.09112345,
  0.01579104, 0.01201851, 0.002560717, 0.01635391, 0.02396246, 0.03572713, 
    0.01372234, 0.01108772, 0.01703406, 0.001515491, 0.00101729, 
    -0.0001817335, 0.008277256, 0.008828245, 0.03186552, 0.01736013, 
    0.03120599, 0.01614628, 0.07787398, 0.03679192, 0.008024524, 0.002478241, 
    0.008686127, 0.002915242, 0.0176933, 0.04386466, 0.05332222, 0.007615367, 
    0.03177423,
  0.02231628, 0.004130149, -8.719278e-06, 0.001339863, -0.0003873, 
    0.0008041211, 0.0004294013, 0.001680375, 0.003582346, 0.001374412, 
    3.484211e-08, 3.901386e-10, 0.003958547, 0.003017153, 0.002018329, 
    0.005777893, 0.002224955, 0.002687308, 0.005189472, 0.001710319, 
    0.0009338305, 0.004279754, 0.01826392, 0.006747785, 0.007873799, 
    0.06418085, 0.003583132, 0.001709408, 0.01575433,
  0.06194476, 0.01450239, 4.52991e-05, 0.08568439, 0.0002512794, 
    0.0005082314, 0.001410719, 0.001550059, 0.0008568466, 0.003605303, 
    0.0006198414, 0.0004565748, 0.009904698, 0.0008513191, 0.0006832291, 
    0.0009533186, 0.0001819288, 0.0003183514, 0.0004825967, 0.0003399218, 
    0.002427635, 0.01037533, 0.06120391, 0.01912646, 0.0001636613, 
    7.1247e-06, 0.00132957, 0.005712558, 0.02257751,
  0.01029895, 0.109671, 0.01139597, 0.01110671, 0.00520874, 0.002234891, 
    0.001569026, 0.001717714, 0.03542413, 0.01916045, 0.000521863, 
    0.001562341, 0.0003572529, 0.0001302218, 0.0003165179, 0.0009885104, 
    0.000358429, 0.0002139473, 9.375846e-05, 0.0006864617, 0.005574859, 
    0.05532405, 0.09269351, 0.007552759, 5.36505e-05, 0.001176434, 
    0.0001242386, 0.0008313861, 0.01534102,
  -1.982578e-05, 3.304829e-06, 8.952299e-06, 0.01035386, 0.01365192, 
    0.0008518497, 0.01213539, 0.001332714, 0.002485247, 7.997018e-05, 
    0.0008301196, 0.0005403042, 0.001520653, 0.003649571, 0.001202834, 
    0.0005193821, 0.002653282, 0.008676651, 0.00996543, 0.002143854, 
    0.00854174, 0.001087027, 0.1718166, 0.02142044, 0.0008531966, 
    0.0005511045, 0.0007619818, 0.001312077, -0.0001907535,
  2.344654e-07, 5.115377e-09, -2.954218e-09, 4.106879e-06, -1.996068e-08, 
    0.00341884, 0.004752177, 0.0007691525, 0.008669134, 0.001312227, 
    0.002151367, 0.0009677441, 0.0005638561, 0.0008011046, 0.0002349842, 
    0.0004296853, 0.0002890342, 0.001209072, 0.003671726, 0.02603781, 
    0.003255975, 0.0756734, 0.0003896724, -0.000723305, 0.000175896, 
    0.0007989961, 0.001489524, 0.006127322, 2.546411e-07,
  -4.583543e-06, 0.0009304952, -5.830734e-07, -5.355146e-06, -0.0003387972, 
    3.243048e-08, -0.0002159814, 0.02168715, 0.1651162, 0.002488118, 
    0.02545496, 0.03562259, 0.01146127, 0.005288146, 0.005153166, 0.0131534, 
    0.001074769, 0.003918949, 0.01726323, 0.06692601, 0.01148288, 0.01328945, 
    0.01206486, 0.009270994, 0.002178524, 0.001084049, 0.001230091, 
    0.001927979, 0.02756016,
  0.01888506, 0.000955231, 0.01126693, 0.1532099, -0.0006709193, 
    0.0001835362, 0.02784975, 0.002289325, 0.003348467, 0.02337271, 
    0.09133498, 0.01856101, 0.08053114, 0.09960002, 0.07149369, 0.08628626, 
    0.1461625, 0.1470852, 0.1154617, 0.006197933, 0.01634936, 0.02105659, 
    0.07781384, 0.04054002, 0.04666779, 0.02700314, 0.04032043, 0.03544826, 
    0.01283268,
  0.03770996, 0.1902283, 0.1490105, 0.1729531, 0.06476078, 0.05778819, 
    0.06570802, 0.1769171, 0.06950566, 0.06597367, 0.0871615, 0.236819, 
    0.101539, 0.05436192, 0.06967992, 0.128374, 0.1242317, 0.2522314, 
    0.2155662, 0.1934095, 0.06728256, 0.05641314, 0.1684862, 0.3454897, 
    0.1082848, 0.2021562, 0.1687417, 0.138818, 0.0731502,
  0.06732516, 0.3545913, 0.2369485, 0.3821262, 0.4361825, 0.2343039, 
    0.2491593, 0.2453803, 0.2509884, 0.2300998, 0.2302919, 0.4068837, 
    0.2302853, 0.1409511, 0.08014025, 0.185886, 0.5720999, 0.3038399, 
    0.369072, 0.1633393, 0.2229542, 0.1949657, 0.07434878, 0.261106, 
    0.1777393, 0.1416708, 0.1100118, 0.1083638, 0.09243682,
  0.1140269, 0.04424214, 0.2616802, 0.1289168, 0.2183404, 0.1859918, 
    0.5576016, 0.4279901, 0.1956811, 0.2804124, 0.3234188, 0.2947583, 
    0.3345069, 0.262718, 0.3734652, 0.3096317, 0.3796533, 0.3282148, 
    0.2506796, 0.1325192, 0.3229683, 0.4796675, 0.4642808, 0.4440667, 
    0.06815523, 0.2822604, 0.4436505, 0.07426362, 0.1660957,
  0.3671479, 0.2172344, 0.5005611, 0.3876181, 0.3284011, 0.3942732, 
    0.4703867, 0.5023521, 0.5213705, 0.5292102, 0.5329168, 0.5132973, 
    0.5232599, 0.4386528, 0.4400234, 0.5331024, 0.5101004, 0.5486668, 
    0.5447923, 0.5480532, 0.5142328, 0.2572341, 0.3161843, 0.5969811, 
    0.1638901, 0.2076822, 0.1591377, 0.3240464, 0.4070586,
  0.07353182, 0.0707972, 0.06806259, 0.06532797, 0.06259336, 0.05985874, 
    0.05712413, 0.04735678, 0.04762864, 0.0479005, 0.04817236, 0.04844422, 
    0.04871608, 0.04898794, 0.05395816, 0.0567533, 0.05954845, 0.06234359, 
    0.06513873, 0.06793388, 0.07072902, 0.07602466, 0.07569227, 0.07535989, 
    0.0750275, 0.07469511, 0.07436273, 0.07403034, 0.07571951,
  0.2588909, 0.182118, 0.09042493, 0.04775415, 0.01532563, 0.01129966, 
    0.003727751, 0.005896601, 0.01344175, 0.01861492, 0.02188438, 0.03667548, 
    0.1027297, -0.00232925, 0.2324997, 0.336181, 0.3731335, 0.2375143, 
    0.08742282, 0.2016393, 0.3193708, 0.5085735, 0.218387, 0.1368235, 
    0.2193264, 0.4328013, 0.1423308, 0.1193547, 0.2422143,
  0.2687578, 0.03906821, 0.05101308, 0.003231284, 0.01062145, 0.07583566, 
    0.0008814827, 0.05376556, 0.05058232, 0.0760362, 0.07207766, 0.09906364, 
    0.02850992, 0.05215889, 0.2437995, 0.2647872, 0.3005056, 0.3082968, 
    0.2774554, 0.2940773, 0.2079835, 0.2391787, 0.1795987, 0.2899977, 
    0.1652716, 0.3672662, 0.3352773, 0.3223588, 0.3807414,
  0.307341, 0.2615267, 0.2817875, 0.1330974, 0.08617172, 0.1132475, 
    0.1584922, 0.1539057, 0.1711513, 0.1157235, 0.09418043, 0.08897781, 
    0.1282467, 0.1330763, 0.07308196, 0.1185504, 0.1688245, 0.213769, 
    0.2009514, 0.1402287, 0.09169433, 0.07587606, 0.09107599, 0.101108, 
    0.1563541, 0.2643501, 0.2950975, 0.3096748, 0.3040651,
  0.2320249, 0.1746648, 0.1395798, 0.1389416, 0.1430181, 0.1068501, 
    0.1042183, 0.1024005, 0.1231697, 0.1031292, 0.06814917, 0.05148514, 
    0.02289063, 0.02749792, 0.03537395, 0.09291536, 0.1410155, 0.1059815, 
    0.1250027, 0.1354253, 0.09257388, 0.05835935, 0.04777134, 0.06581195, 
    0.01613164, 0.1239068, 0.3062959, 0.203039, 0.2818119,
  0.05939584, 0.02814073, 0.02397615, 0.04748811, 0.03624194, 0.03702, 
    0.05191474, 0.06764505, 0.064622, 0.03242487, 0.01305398, 0.004603665, 
    0.009621531, 0.04286778, 0.1163474, 0.07884233, 0.0723622, 0.07928835, 
    0.07863921, 0.05226068, 0.0394612, 0.05211366, 0.03070951, 0.1675551, 
    0.03633843, 0.04305965, 0.03927423, 0.03792324, 0.0591835,
  0.01150463, 0.008432105, 0.001674996, 0.008742334, 0.01278545, 0.01976439, 
    0.007798833, 0.008244001, 0.01305375, 0.001192552, 0.0007334125, 
    -0.000161299, 0.008008013, 0.005102755, 0.01944092, 0.009662622, 
    0.01628898, 0.01017219, 0.04509715, 0.02299311, 0.004204563, 0.001988904, 
    0.006601001, 0.00229143, 0.01389391, 0.02497243, 0.02787347, 0.004203864, 
    0.01880219,
  0.01628479, 0.002434231, -5.975512e-06, 0.000896481, -0.0004219992, 
    0.0003621278, 0.0003154891, 0.001219003, 0.002730242, 0.001088241, 
    3.377166e-08, 2.405474e-08, 0.002822075, 0.001762686, 0.001421204, 
    0.002889366, 0.001108045, 0.00159543, 0.002663311, 0.0008189504, 
    0.0006780206, 0.003107983, 0.01356484, 0.004906366, 0.005033902, 
    0.05579001, 0.001755412, 0.001208256, 0.01101646,
  0.04433861, 0.009537211, 6.263533e-05, 0.06503224, 0.0001324719, 
    0.0003112252, 0.0005105969, 0.000712816, 0.0006233886, 0.002919202, 
    0.0003992232, 0.000311077, 0.004659931, 0.0005130594, 0.0003896885, 
    0.0004916928, 0.0001640033, 0.0002371764, 0.000368723, 0.0002521529, 
    0.001790091, 0.007460352, 0.04494709, 0.01580288, 0.0005307358, 
    -1.712271e-06, 0.001078866, 0.004120941, 0.01584331,
  0.00690627, 0.08527423, 0.008771955, 0.008132544, 0.003717091, 0.001184871, 
    0.0009919078, 0.0009047341, 0.02547464, 0.02465122, 0.000385993, 
    0.001116985, 0.0002479531, 8.929858e-05, 0.0002208229, 0.0007092379, 
    0.0002506163, 0.0001480197, 6.296132e-05, 0.0004808633, 0.003730776, 
    0.03841103, 0.06899963, 0.003655931, 7.993753e-05, 0.0008269987, 
    0.0001096503, 0.0005601901, 0.0106045,
  -5.938075e-05, 3.089199e-06, 2.504474e-05, 0.009235885, 0.007285913, 
    0.0006230795, 0.009110996, 0.0006481267, 0.001290526, 7.079964e-05, 
    0.0004162277, 0.0002729556, 0.0007300829, 0.001846575, 0.0006018904, 
    0.0002607365, 0.001235009, 0.004010589, 0.00480534, 0.001199836, 
    0.004330689, 0.0005690569, 0.1416133, 0.02358264, 0.0005267687, 
    0.0003255895, 0.0004835487, 0.0008684199, -0.0002036196,
  2.260814e-07, 4.88787e-09, -2.213813e-09, 6.349034e-06, 3.225014e-08, 
    0.002424976, 0.00231338, 0.0004661711, 0.01071807, 0.0009129181, 
    0.0009636256, 0.0005011017, 0.0003503009, 0.0003997482, 0.0001422047, 
    0.0003209359, 0.0002179656, 0.0006712835, 0.00263521, 0.01785916, 
    0.002319103, 0.0639147, 0.000292486, -0.00102652, 0.0001263319, 
    0.0005797701, 0.001091724, 0.004448661, 2.560647e-07,
  -3.243142e-06, 0.0003985599, 4.196362e-05, -1.018345e-05, -0.0003212712, 
    3.050909e-08, -0.000276894, 0.02656086, 0.1526881, 0.001559488, 
    0.01462713, 0.02338882, 0.005887861, 0.002679873, 0.003177298, 
    0.00712962, 0.0007455378, 0.00213713, 0.01134438, 0.05726052, 
    0.009689938, 0.0174653, 0.01145996, 0.002601978, 0.00139646, 0.000792293, 
    0.0007462678, 0.001432364, 0.02198608,
  0.01548786, 0.0004353497, 0.008441875, 0.1459272, -0.0006171078, 
    0.0001338078, 0.02047091, 0.001937984, 0.002167344, 0.018529, 0.08162716, 
    0.01139166, 0.06020585, 0.07337367, 0.05077615, 0.06222657, 0.1008724, 
    0.09421997, 0.0811979, 0.005832065, 0.0129678, 0.01454536, 0.05874323, 
    0.03064784, 0.03079108, 0.01581904, 0.02139275, 0.02344494, 0.008593627,
  0.02697837, 0.1642373, 0.1264756, 0.1566608, 0.05478815, 0.04858059, 
    0.05373282, 0.1522424, 0.06009502, 0.05860719, 0.07814977, 0.2125466, 
    0.07542631, 0.03694956, 0.04981986, 0.08696483, 0.0843339, 0.1887774, 
    0.1680092, 0.1823125, 0.05623182, 0.04563926, 0.1393669, 0.3127192, 
    0.08511309, 0.1720047, 0.1334864, 0.1040279, 0.05319695,
  0.04390235, 0.3322629, 0.2008839, 0.3352933, 0.3967009, 0.2146891, 
    0.2220527, 0.2092093, 0.213477, 0.1952262, 0.1955039, 0.3682514, 
    0.2099121, 0.1229058, 0.06539728, 0.1469469, 0.5322343, 0.2683963, 
    0.33917, 0.1498277, 0.2020357, 0.1736653, 0.0579228, 0.228277, 0.1470261, 
    0.1184271, 0.07900257, 0.07594891, 0.06386989,
  0.07651003, 0.02843624, 0.2465758, 0.09046769, 0.180621, 0.153583, 
    0.5051987, 0.3719451, 0.1859565, 0.2433229, 0.295106, 0.2429571, 
    0.2895272, 0.2139602, 0.3133323, 0.2811646, 0.3352216, 0.2857479, 
    0.205965, 0.1012262, 0.282188, 0.4286365, 0.4168958, 0.4388692, 
    0.05500366, 0.2373458, 0.5367697, 0.06169317, 0.132841,
  0.3532653, 0.1887479, 0.4306717, 0.343051, 0.2824034, 0.3260696, 0.3666997, 
    0.4120115, 0.4219983, 0.3944485, 0.4001576, 0.383187, 0.4092475, 
    0.3123382, 0.3179052, 0.3963382, 0.3718526, 0.3916259, 0.3951079, 
    0.4155212, 0.4274545, 0.2210336, 0.3293791, 0.6268033, 0.1633081, 
    0.1855185, 0.1801411, 0.299632, 0.3431219,
  0.0583335, 0.05671496, 0.05509641, 0.05347787, 0.05185933, 0.05024078, 
    0.04862224, 0.04273539, 0.04302087, 0.04330635, 0.04359183, 0.04387731, 
    0.04416279, 0.04444828, 0.04595651, 0.04805595, 0.05015539, 0.05225483, 
    0.05435426, 0.0564537, 0.05855313, 0.06587194, 0.06510556, 0.06433919, 
    0.06357282, 0.06280645, 0.06204008, 0.0612737, 0.05962834,
  0.2260482, 0.1123141, 0.06302117, 0.03281492, 0.01373502, 0.0153816, 
    0.004152198, 0.006443638, 0.01255577, 0.01834843, 0.01818813, 0.0327837, 
    0.08236566, -0.0009974006, 0.2968249, 0.3119747, 0.3523908, 0.2565878, 
    0.086797, 0.2170917, 0.3090829, 0.4968747, 0.2037497, 0.1261755, 
    0.2280954, 0.4266782, 0.1557137, 0.1086508, 0.2166874,
  0.2570705, 0.04456638, 0.06738605, 0.002867433, 0.009286901, 0.07102343, 
    0.0004939645, 0.05157002, 0.05653138, 0.0735486, 0.07237396, 0.09629852, 
    0.03280165, 0.05180501, 0.2213107, 0.2381861, 0.2805836, 0.285485, 
    0.2534165, 0.2634039, 0.1783519, 0.213673, 0.1654105, 0.2648621, 
    0.1566145, 0.3399073, 0.3001793, 0.2907986, 0.3528565,
  0.2782627, 0.2320283, 0.2536114, 0.1180475, 0.07590669, 0.1003035, 
    0.1460195, 0.1387809, 0.1562532, 0.1012523, 0.08281916, 0.0783516, 
    0.1109741, 0.1173962, 0.06395118, 0.1048218, 0.1467703, 0.1872551, 
    0.1739577, 0.1200978, 0.08065693, 0.06608626, 0.07652603, 0.08525634, 
    0.1301841, 0.2333227, 0.2765751, 0.2783708, 0.2789401,
  0.1893095, 0.1491444, 0.1187609, 0.1179554, 0.1214256, 0.09216114, 
    0.08912623, 0.08535835, 0.1040465, 0.08877119, 0.05510868, 0.04122449, 
    0.01761114, 0.02060851, 0.02717779, 0.07111909, 0.106287, 0.08235857, 
    0.09871565, 0.1043617, 0.0704396, 0.04608795, 0.03730877, 0.07293001, 
    0.01310407, 0.09595509, 0.2508188, 0.1760455, 0.2305393,
  0.04462253, 0.01978422, 0.01829345, 0.03546803, 0.02627538, 0.02729574, 
    0.03697852, 0.04722177, 0.04539493, 0.02541296, 0.00942314, 0.00358147, 
    0.007213186, 0.03191959, 0.1042501, 0.05829611, 0.05301738, 0.05790889, 
    0.05518296, 0.04039302, 0.02890088, 0.03854143, 0.0215814, 0.1627561, 
    0.02923345, 0.02918827, 0.0278219, 0.02638462, 0.04189925,
  0.00913202, 0.006793463, 0.002428833, 0.005654483, 0.007976048, 0.01259238, 
    0.005415424, 0.006850681, 0.0110466, 0.001020073, 0.0005578857, 
    -0.0001326586, 0.01037055, 0.00311858, 0.01091584, 0.006320846, 
    0.009732276, 0.006994917, 0.02914479, 0.01390073, 0.002891954, 
    0.001771451, 0.005570622, 0.001966418, 0.01995195, 0.01592451, 
    0.01537026, 0.002794388, 0.01318033,
  0.01338904, 0.001911813, -2.006173e-05, 0.0007188788, -0.0006621451, 
    0.000217927, 0.0002663566, 0.001012645, 0.002313112, 0.0009335098, 
    3.339507e-08, 4.579431e-08, 0.00230297, 0.001330429, 0.001153668, 
    0.001874505, 0.0007613081, 0.001225964, 0.001544089, 0.0005520291, 
    0.0005567459, 0.0025735, 0.01136286, 0.003967459, 0.01115415, 0.06982367, 
    0.001159578, 0.0009924453, 0.008811688,
  0.03581645, 0.007201626, 0.001134917, 0.06632766, 9.437421e-05, 
    0.0002410527, 0.0003111197, 0.0004589854, 0.0005150983, 0.002233645, 
    0.0003143617, 0.0002495954, 0.002911962, 0.0004005193, 0.0002901848, 
    0.0003479751, 0.0001458427, 0.0001970822, 0.0003124991, 0.0002097791, 
    0.001492782, 0.006117224, 0.03688815, 0.07964802, 0.005144437, 
    0.0002222954, 0.0008766841, 0.003375486, 0.01271703,
  0.005441019, 0.1052245, 0.01103047, 0.007514921, 0.002982606, 0.0008509598, 
    0.0007511057, 0.0006086159, 0.04165777, 0.05087977, 0.000320035, 
    0.0008978654, 0.0001977028, 7.226696e-05, 0.0001794282, 0.0005723594, 
    0.0002006539, 0.0001200571, 5.054344e-05, 0.00038965, 0.002904423, 
    0.03021732, 0.05689847, 0.01014355, 0.002642632, 0.0006740739, 
    0.0001029576, 0.000441451, 0.008384964,
  0.0003446418, 3.586915e-05, 0.0001980299, 0.006981793, 0.004882586, 
    0.0005084914, 0.00532845, 0.0003862486, 0.0002957145, 6.620499e-05, 
    0.0002875785, 0.0001954917, 0.0005024847, 0.001258059, 0.0004203944, 
    0.0001890851, 0.0008240459, 0.002499848, 0.002738979, 0.0009078622, 
    0.002664091, 0.0004141966, 0.2134446, 0.034038, 0.0003983687, 
    0.0002436267, 0.0003758729, 0.0006563382, 0.001942233,
  2.23708e-07, 4.763889e-09, -1.447008e-09, 8.946841e-08, 3.747545e-08, 
    0.001936658, 0.004022856, 0.0003247954, 0.01684215, 0.0004526102, 
    0.0006149578, 0.0003393466, 0.0002678631, 0.0002864295, 0.0001088001, 
    0.000266431, 0.0001758391, 0.0004998129, 0.002154037, 0.01316134, 
    0.001873701, 0.05921913, 0.0002444905, -0.001816886, 0.0001023828, 
    0.0004773688, 0.0008988507, 0.003637352, 2.59726e-07,
  -2.360861e-06, 0.0002676146, 0.000209793, -4.730947e-06, -0.0001701961, 
    2.930715e-08, -2.970029e-05, 0.03946609, 0.1564192, 0.001449793, 
    0.01000279, 0.01426973, 0.003747237, 0.001751554, 0.002442475, 
    0.00479007, 0.0006027939, 0.001542118, 0.008432063, 0.05140975, 
    0.00914278, 0.04837533, 0.01607799, 0.001404072, 0.001109122, 
    0.0006501048, 0.0005753957, 0.001188166, 0.01879296,
  0.01627927, 1.162939e-05, 0.006786316, 0.1467803, -0.0006215295, 
    0.0001107632, 0.01665975, 0.001686955, 0.002194017, 0.01607613, 
    0.09114581, 0.0078495, 0.04526858, 0.05324678, 0.03646534, 0.04244951, 
    0.07235125, 0.05996401, 0.06304246, 0.005466094, 0.0121286, 0.0154953, 
    0.05498049, 0.02345703, 0.02170124, 0.009771402, 0.01323054, 0.01759337, 
    0.006756334,
  0.02070711, 0.1729801, 0.1251534, 0.1529394, 0.04810473, 0.04262268, 
    0.04874251, 0.1504152, 0.06403856, 0.05543299, 0.08691393, 0.218335, 
    0.05992333, 0.02790179, 0.03826609, 0.06173031, 0.06242797, 0.1412251, 
    0.1362336, 0.1885612, 0.05458657, 0.04181542, 0.1468689, 0.3260829, 
    0.07844309, 0.1410263, 0.1028976, 0.07999279, 0.03998089,
  0.03293908, 0.3504344, 0.2091333, 0.3342608, 0.4072826, 0.2203815, 
    0.2256081, 0.2116978, 0.2216749, 0.2080205, 0.1998968, 0.376363, 
    0.213673, 0.1489922, 0.05872401, 0.1257333, 0.5392768, 0.2600694, 
    0.3733394, 0.1489254, 0.2086133, 0.1741424, 0.04914973, 0.2277956, 
    0.1236044, 0.1049041, 0.06157189, 0.05648353, 0.04823103,
  0.06084711, 0.02223907, 0.283794, 0.07155599, 0.1541221, 0.1325914, 
    0.4897065, 0.3554362, 0.205382, 0.2424457, 0.3313121, 0.2314459, 
    0.2619711, 0.1820685, 0.2752486, 0.2673156, 0.3258553, 0.2721536, 
    0.1776364, 0.08334993, 0.2520751, 0.3843696, 0.3908983, 0.4421729, 
    0.04260739, 0.2247707, 0.6008283, 0.06010945, 0.1117945,
  0.3395557, 0.172871, 0.3977808, 0.2976499, 0.2505541, 0.2787052, 0.2930965, 
    0.330079, 0.3396973, 0.3049853, 0.3075298, 0.2919601, 0.314302, 
    0.2261072, 0.2349408, 0.3048034, 0.2902328, 0.3111097, 0.3360042, 
    0.349782, 0.3736839, 0.2087787, 0.343773, 0.6220757, 0.1713524, 
    0.1868394, 0.2054432, 0.3071305, 0.3023108 ;

 average_DT = 730 ;

 average_T1 = 289.5 ;

 average_T2 = 1019.5 ;

 climatology_bounds =
  289.5, 1019.5 ;

 lat = -89.5, -79.5, -69.5, -59.5, -49.5, -39.5, -29.5, -19.5, -9.5, 0.5, 
    10.5, 20.5, 30.5, 40.5, 50.5, 60.5, 70.5, 80.5 ;

 lat_bnds =
  -90, -89,
  -80, -79,
  -70, -69,
  -60, -59,
  -50, -49,
  -40, -39,
  -30, -29,
  -20, -19,
  -10, -9,
  0, 1,
  10, 11,
  20, 21,
  30, 31,
  40, 41,
  50, 51,
  60, 61,
  70, 71,
  80, 81 ;

 lon = 0.625, 13.125, 25.625, 38.125, 50.625, 63.125, 75.625, 88.125, 
    100.625, 113.125, 125.625, 138.125, 150.625, 163.125, 175.625, 188.125, 
    200.625, 213.125, 225.625, 238.125, 250.625, 263.125, 275.625, 288.125, 
    300.625, 313.125, 325.625, 338.125, 350.625 ;

 lon_bnds =
  0, 1.25,
  12.5, 13.75,
  25, 26.25,
  37.5, 38.75,
  50, 51.25,
  62.5, 63.75,
  75, 76.25,
  87.5, 88.75,
  100, 101.25,
  112.5, 113.75,
  125, 126.25,
  137.5, 138.75,
  150, 151.25,
  162.5, 163.75,
  175, 176.25,
  187.5, 188.75,
  200, 201.25,
  212.5, 213.75,
  225, 226.25,
  237.5, 238.75,
  250, 251.25,
  262.5, 263.75,
  275, 276.25,
  287.5, 288.75,
  300, 301.25,
  312.5, 313.75,
  325, 326.25,
  337.5, 338.75,
  350, 351.25 ;

 pfull = 0.0252729048206747, 0.0885404738757409, 0.213072411383256, 
    0.41190537807884, 0.671080828691593, 0.987471468515016, 1.36790961365676, 
    1.82562112064242, 2.38097588033244, 3.06218961364243, 3.90121721567151, 
    4.9296281825995, 6.18008131929323, 7.68875807563375, 9.49537809361575, 
    11.643153995098, 14.1786857151188, 17.1517875598959, 20.6152476986609, 
    24.6245259348741, 29.237386591333, 34.5134757786445, 40.5138467378254, 
    47.3004421634272, 54.9355325495126, 63.4811392623337, 72.9984371159701, 
    83.5471442618119, 95.1849171805989, 107.966767294215, 121.944503506415, 
    137.166169497631, 153.675572970355, 171.511834307961, 190.708985325578, 
    211.295632932361, 233.294677858721, 256.723099608772, 281.591803639405, 
    307.905555737256, 335.66293113824, 364.856338389786, 395.47216160598, 
    427.490864234311, 460.887168786725, 495.630391513078, 531.761718445649, 
    569.289185351388, 607.768705103107, 646.445374671436, 684.792067788697, 
    722.468679913451, 759.124006783627, 794.401045766566, 827.769968639223, 
    858.597822486016, 886.389109609622, 910.841030891388, 931.860653469283, 
    949.549679924174, 964.159924710431, 976.012345333387, 985.470174132691, 
    992.77226220014, 997.948601287575 ;

 time = 0 ;
}
