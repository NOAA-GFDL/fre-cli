netcdf \20030101.grid_spec.tile3 {
dimensions:
	grid_x = 97 ;
	grid_y = 97 ;
	time = UNLIMITED ; // (1 currently)
	grid_xt = 96 ;
	grid_yt = 96 ;
	phalf = 50 ;
variables:
	double grid_x(grid_x) ;
		grid_x:units = "degrees_E" ;
		grid_x:long_name = "cell corner longitude" ;
		grid_x:axis = "X" ;
	double grid_y(grid_y) ;
		grid_y:units = "degrees_N" ;
		grid_y:long_name = "cell corner latitude" ;
		grid_y:axis = "Y" ;
	double time(time) ;
		time:units = "days since 1870-01-01 00:00:00" ;
		time:long_name = "time" ;
		time:axis = "T" ;
		time:calendar_type = "JULIAN" ;
		time:calendar = "julian" ;
	double grid_xt(grid_xt) ;
		grid_xt:units = "degrees_E" ;
		grid_xt:long_name = "T-cell longitude" ;
		grid_xt:axis = "X" ;
	double grid_yt(grid_yt) ;
		grid_yt:units = "degrees_N" ;
		grid_yt:long_name = "T-cell latitude" ;
		grid_yt:axis = "Y" ;
	double phalf(phalf) ;
		phalf:units = "mb" ;
		phalf:long_name = "ref half pressure level" ;
		phalf:axis = "Z" ;
		phalf:positive = "down" ;
	float grid_lon(grid_y, grid_x) ;
		grid_lon:_FillValue = 1.e+20f ;
		grid_lon:missing_value = 1.e+20f ;
		grid_lon:units = "degrees_E" ;
		grid_lon:long_name = "longitude" ;
		grid_lon:cell_methods = "time: point" ;
	float grid_lat(grid_y, grid_x) ;
		grid_lat:_FillValue = 1.e+20f ;
		grid_lat:missing_value = 1.e+20f ;
		grid_lat:units = "degrees_N" ;
		grid_lat:long_name = "latitude" ;
		grid_lat:cell_methods = "time: point" ;
	float grid_lont(grid_yt, grid_xt) ;
		grid_lont:_FillValue = 1.e+20f ;
		grid_lont:missing_value = 1.e+20f ;
		grid_lont:units = "degrees_E" ;
		grid_lont:long_name = "longitude" ;
		grid_lont:cell_methods = "time: point" ;
	float grid_latt(grid_yt, grid_xt) ;
		grid_latt:_FillValue = 1.e+20f ;
		grid_latt:missing_value = 1.e+20f ;
		grid_latt:units = "degrees_N" ;
		grid_latt:long_name = "latitude" ;
		grid_latt:cell_methods = "time: point" ;
	float area(grid_yt, grid_xt) ;
		area:_FillValue = 1.e+20f ;
		area:missing_value = 1.e+20f ;
		area:units = "m**2" ;
		area:long_name = "cell area" ;
		area:cell_methods = "time: point" ;
	float bk(phalf) ;
		bk:_FillValue = 1.e+20f ;
		bk:missing_value = 1.e+20f ;
		bk:long_name = "vertical coordinate sigma value" ;
		bk:cell_methods = "time: point" ;
	float pk(phalf) ;
		pk:_FillValue = 1.e+20f ;
		pk:missing_value = 1.e+20f ;
		pk:units = "pascal" ;
		pk:long_name = "pressure part of the hybrid coordinate" ;
		pk:cell_methods = "time: point" ;
	float sftlf(grid_yt, grid_xt) ;
		sftlf:_FillValue = 1.e+20f ;
		sftlf:missing_value = 1.e+20f ;
		sftlf:units = "1.0" ;
		sftlf:long_name = "Fraction of the Grid Cell Occupied by Land" ;
		sftlf:cell_methods = "time: point" ;
		sftlf:cell_measures = "area: area" ;
		sftlf:standard_name = "land_area_fraction" ;
		sftlf:interp_method = "conserve_order1" ;
	float orog(grid_yt, grid_xt) ;
		orog:_FillValue = 1.e+20f ;
		orog:missing_value = 1.e+20f ;
		orog:units = "m" ;
		orog:long_name = "Surface Altitude" ;
		orog:cell_methods = "time: point" ;
		orog:cell_measures = "area: area" ;
		orog:standard_name = "surface_altitude" ;
		orog:interp_method = "conserve_order1" ;
	float land_mask(grid_yt, grid_xt) ;
		land_mask:_FillValue = 1.e+20f ;
		land_mask:missing_value = 1.e+20f ;
		land_mask:valid_range = -0.01f, 1.01f ;
		land_mask:long_name = "fractional amount of land" ;
		land_mask:cell_methods = "time: point" ;
		land_mask:interp_method = "conserve_order1" ;
	float zsurf(grid_yt, grid_xt) ;
		zsurf:_FillValue = 1.e+20f ;
		zsurf:missing_value = 1.e+20f ;
		zsurf:units = "m" ;
		zsurf:long_name = "surface height" ;
		zsurf:cell_methods = "time: point" ;

// global attributes:
		:title = "ESM4_longamip_D1_am4p2_proto7b_whiteCapsAlbedo_salt_SIS2" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
data:

 grid_x = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19, 
    20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 37, 
    38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 54, 55, 
    56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 72, 73, 
    74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 90, 91, 
    92, 93, 94, 95, 96, 97 ;

 grid_y = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19, 
    20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 37, 
    38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 54, 55, 
    56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 72, 73, 
    74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 90, 91, 
    92, 93, 94, 95, 96, 97 ;

 time = 0 ;

 grid_xt = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19, 
    20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 37, 
    38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 54, 55, 
    56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 72, 73, 
    74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 90, 91, 
    92, 93, 94, 95, 96 ;

 grid_yt = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19, 
    20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 37, 
    38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 54, 55, 
    56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 72, 73, 
    74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 90, 91, 
    92, 93, 94, 95, 96 ;

 phalf = 0.01, 0.0269722, 0.0517136, 0.0889455, 0.142479, 0.2207157, 
    0.3361283, 0.5048096, 0.7479993, 1.0940055, 1.580046, 2.2544108, 
    3.178956, 4.431935, 6.1111558, 8.3374392, 11.2583405, 15.0520759, 
    19.9315829, 26.1486254, 33.997842, 43.820624, 56.0087014, 71.0073115, 
    89.3178242, 111.4997021, 138.1716841, 170.012093, 207.7581856, 
    252.2033875, 304.1464563, 363.9522552, 430.6429622, 501.015122, 
    570.6113482, 635.806353, 694.8286462, 747.1992533, 793.0044191, 
    832.5750255, 866.4443202, 895.1917865, 919.4060705, 939.6860264, 
    956.4664631, 970.1833931, 981.1347983, 989.68, 995.9, 1000 ;

 grid_lon =
  35, 35.78278, 36.57269, 37.36979, 38.17411, 38.98572, 39.80465, 40.63093, 
    41.46459, 42.30565, 43.15412, 44.01001, 44.87331, 45.744, 46.62207, 
    47.50749, 48.40021, 49.30018, 50.20734, 51.12163, 52.04295, 52.97122, 
    53.90633, 54.84815, 55.79657, 56.75144, 57.71262, 58.67992, 59.65319, 
    60.63222, 61.61683, 62.60678, 63.60188, 64.60188, 65.60651, 66.61555, 
    67.62873, 68.64574, 69.66634, 70.69019, 71.71702, 72.7465, 73.77832, 
    74.81216, 75.84769, 76.88457, 77.92248, 78.96107, 80, 81.03893, 82.07752, 
    83.11543, 84.15231, 85.18784, 86.22168, 87.2535, 88.28298, 89.30981, 
    90.33366, 91.35426, 92.37127, 93.38445, 94.39349, 95.39812, 96.39812, 
    97.39321, 98.38318, 99.36778, 100.3468, 101.3201, 102.2874, 103.2486, 
    104.2034, 105.1518, 106.0937, 107.0288, 107.957, 108.8784, 109.7927, 
    110.6998, 111.5998, 112.4925, 113.3779, 114.256, 115.1267, 115.99, 
    116.8459, 117.6944, 118.5354, 119.3691, 120.1954, 121.0143, 121.8259, 
    122.6302, 123.4273, 124.2172, 125,
  34.21722, 35, 35.7905, 36.5888, 37.39495, 38.20903, 39.03109, 39.86116, 
    40.69931, 41.54556, 42.39994, 43.26246, 44.13313, 45.01196, 45.89892, 
    46.794, 47.69717, 48.60838, 49.52757, 50.45469, 51.38964, 52.33234, 
    53.28267, 54.24053, 55.20577, 56.17825, 57.15781, 58.14427, 59.13744, 
    60.13712, 61.14308, 62.15511, 63.17294, 64.19632, 65.22498, 66.25863, 
    67.29697, 68.33968, 69.38647, 70.43697, 71.49085, 72.54777, 73.60736, 
    74.66925, 75.73307, 76.79844, 77.86497, 78.9323, 80, 81.0677, 82.13503, 
    83.20156, 84.26693, 85.33075, 86.39264, 87.45223, 88.50915, 89.56303, 
    90.61353, 91.66032, 92.70303, 93.74137, 94.77502, 95.80368, 96.82706, 
    97.84489, 98.85692, 99.86288, 100.8626, 101.8557, 102.8422, 103.8217, 
    104.7942, 105.7595, 106.7173, 107.6677, 108.6104, 109.5453, 110.4724, 
    111.3916, 112.3028, 113.206, 114.1011, 114.988, 115.8669, 116.7375, 
    117.6001, 118.4544, 119.3007, 120.1388, 120.9689, 121.791, 122.605, 
    123.4112, 124.2095, 125, 125.7828,
  33.42731, 34.2095, 35, 35.79891, 36.6063, 37.42227, 38.24688, 39.0802, 
    39.92228, 40.77319, 41.63295, 42.50162, 43.3792, 44.26571, 45.16115, 
    46.06552, 46.97879, 47.90092, 48.83188, 49.7716, 50.72, 51.677, 52.64248, 
    53.61634, 54.59843, 55.5886, 56.58668, 57.59249, 58.60582, 59.62646, 
    60.65416, 61.68868, 62.72975, 63.77708, 64.83036, 65.88928, 66.95352, 
    68.02271, 69.0965, 70.17452, 71.25639, 72.34169, 73.43002, 74.52098, 
    75.61414, 76.70905, 77.80529, 78.90243, 80, 81.09757, 82.19471, 83.29095, 
    84.38586, 85.47902, 86.56998, 87.65831, 88.74361, 89.82548, 90.9035, 
    91.97729, 93.04648, 94.11072, 95.16964, 96.22292, 97.27025, 98.31132, 
    99.34584, 100.3735, 101.3942, 102.4075, 103.4133, 104.4114, 105.4016, 
    106.3837, 107.3575, 108.323, 109.28, 110.2284, 111.1681, 112.0991, 
    113.0212, 113.9345, 114.8389, 115.7343, 116.6208, 117.4984, 118.367, 
    119.2268, 120.0777, 120.9198, 121.7531, 122.5777, 123.3937, 124.2011, 
    125, 125.7905, 126.5727,
  32.63021, 33.4112, 34.20109, 35, 35.80803, 36.62528, 37.45184, 38.28781, 
    39.13326, 39.98825, 40.85287, 41.72715, 42.61113, 43.50485, 44.40832, 
    45.32156, 46.24454, 47.17727, 48.11968, 49.07174, 50.03338, 51.00451, 
    51.98503, 52.97483, 53.97377, 54.98169, 55.99842, 57.02376, 58.0575, 
    59.09941, 60.14923, 61.20669, 62.2715, 63.34334, 64.42188, 65.50678, 
    66.59766, 67.69415, 68.79581, 69.90228, 71.01307, 72.12776, 73.2459, 
    74.367, 75.49059, 76.61618, 77.74329, 78.87139, 80, 81.12861, 82.25671, 
    83.38382, 84.50941, 85.633, 86.7541, 87.87224, 88.98693, 90.09772, 
    91.20419, 92.30585, 93.40234, 94.49322, 95.57812, 96.65666, 97.72851, 
    98.79331, 99.85078, 100.9006, 101.9425, 102.9762, 104.0016, 105.0183, 
    106.0262, 107.0252, 108.015, 108.9955, 109.9666, 110.9283, 111.8803, 
    112.8227, 113.7555, 114.6784, 115.5917, 116.4951, 117.3889, 118.2729, 
    119.1471, 120.0117, 120.8667, 121.7122, 122.5482, 123.3747, 124.192, 125, 
    125.7989, 126.5888, 127.3698,
  31.82589, 32.60505, 33.3937, 34.19197, 35, 35.8179, 36.6458, 37.4838, 
    38.332, 39.19049, 40.05937, 40.93871, 41.82855, 42.72896, 43.63998, 
    44.56163, 45.49391, 46.43683, 47.39036, 48.35447, 49.32909, 50.31416, 
    51.30958, 52.31524, 53.33099, 54.3567, 55.39217, 56.43721, 57.49159, 
    58.55508, 59.62738, 60.70823, 61.7973, 62.89424, 63.9987, 65.1103, 
    66.22861, 67.35323, 68.4837, 69.61956, 70.76032, 71.90548, 73.05452, 
    74.20692, 75.36213, 76.51961, 77.67879, 78.83911, 80, 81.16089, 82.32121, 
    83.48039, 84.63787, 85.79308, 86.94548, 88.09452, 89.23968, 90.38044, 
    91.5163, 92.64677, 93.77139, 94.8897, 96.0013, 97.10576, 98.20271, 
    99.29177, 100.3726, 101.4449, 102.5084, 103.5628, 104.6078, 105.6433, 
    106.669, 107.6848, 108.6904, 109.6858, 110.6709, 111.6455, 112.6096, 
    113.5632, 114.5061, 115.4384, 116.36, 117.271, 118.1714, 119.0613, 
    119.9406, 120.8095, 121.668, 122.5162, 123.3542, 124.1821, 125, 125.808, 
    126.6063, 127.395, 128.1741,
  31.01428, 31.79097, 32.57773, 33.37472, 34.1821, 35, 35.82858, 36.66796, 
    37.51827, 38.37964, 39.25217, 40.13595, 41.03108, 41.93763, 42.85566, 
    43.78522, 44.72634, 45.67903, 46.64329, 47.6191, 48.60642, 49.60519, 
    50.61533, 51.63671, 52.66924, 53.71273, 54.76702, 55.83191, 56.90716, 
    57.99251, 59.08768, 60.19236, 61.30621, 62.42886, 63.55991, 64.69896, 
    65.84554, 66.99919, 68.15942, 69.3257, 70.4975, 71.67426, 72.85539, 
    74.04031, 75.2284, 76.41905, 77.61163, 78.80549, 80, 81.19451, 82.38837, 
    83.58095, 84.7716, 85.95969, 87.14461, 88.32574, 89.5025, 90.6743, 
    91.84058, 93.00081, 94.15446, 95.30104, 96.44009, 97.57114, 98.69379, 
    99.80763, 100.9123, 102.0075, 103.0928, 104.1681, 105.233, 106.2873, 
    107.3308, 108.3633, 109.3847, 110.3948, 111.3936, 112.3809, 113.3567, 
    114.321, 115.2737, 116.2148, 117.1443, 118.0624, 118.9689, 119.8641, 
    120.7478, 121.6204, 122.4817, 123.332, 124.1714, 125, 125.8179, 126.6253, 
    127.4223, 128.209, 128.9857,
  30.19535, 30.96892, 31.75312, 32.54816, 33.3542, 34.17142, 35, 35.84009, 
    36.69184, 37.55542, 38.43094, 39.31855, 40.21834, 41.13043, 42.0549, 
    42.99183, 43.94127, 44.90327, 45.87783, 46.86496, 47.86464, 48.87683, 
    49.90145, 50.93842, 51.98761, 53.04887, 54.12204, 55.20689, 56.3032, 
    57.41071, 58.52911, 59.65807, 60.79723, 61.94619, 63.10454, 64.27181, 
    65.44752, 66.63114, 67.82214, 69.01993, 70.22392, 71.43348, 72.64796, 
    73.86671, 75.08904, 76.31424, 77.54162, 78.77045, 80, 81.22955, 82.45838, 
    83.68576, 84.91096, 86.13329, 87.35204, 88.56652, 89.77608, 90.98007, 
    92.17786, 93.36886, 94.55248, 95.72819, 96.89545, 98.0538, 99.20277, 
    100.3419, 101.4709, 102.5893, 103.6968, 104.7931, 105.878, 106.9511, 
    108.0124, 109.0616, 110.0985, 111.1232, 112.1354, 113.135, 114.1222, 
    115.0967, 116.0587, 117.0082, 117.9451, 118.8696, 119.7817, 120.6815, 
    121.5691, 122.4446, 123.3082, 124.1599, 125, 125.8286, 126.6458, 
    127.4518, 128.2469, 129.0311, 129.8047,
  29.36907, 30.13884, 30.91981, 31.71219, 32.5162, 33.33204, 34.15991, 35, 
    35.8525, 36.71758, 37.59541, 38.48615, 39.38995, 40.30694, 41.23724, 
    42.18094, 43.13815, 44.10892, 45.0933, 46.09133, 47.10299, 48.12827, 
    49.16711, 50.21945, 51.28517, 52.36414, 53.45618, 54.5611, 55.67866, 
    56.80858, 57.95056, 59.10424, 60.26925, 61.44517, 62.63153, 63.82784, 
    65.03357, 66.24815, 67.47097, 68.70142, 69.93881, 71.18246, 72.43164, 
    73.68562, 74.94361, 76.20486, 77.46854, 78.73386, 80, 81.26614, 82.53146, 
    83.79514, 85.05639, 86.31438, 87.56836, 88.81754, 90.06119, 91.29858, 
    92.52903, 93.75185, 94.96643, 96.17216, 97.36847, 98.55483, 99.73074, 
    100.8958, 102.0494, 103.1914, 104.3213, 105.4389, 106.5438, 107.6359, 
    108.7148, 109.7805, 110.8329, 111.8717, 112.897, 113.9087, 114.9067, 
    115.8911, 116.8618, 117.8191, 118.7628, 119.6931, 120.6101, 121.5138, 
    122.4046, 123.2824, 124.1475, 125, 125.8401, 126.668, 127.4838, 128.2878, 
    129.0802, 129.8612, 130.6309,
  28.53541, 29.30069, 30.07772, 30.86674, 31.668, 32.48173, 33.30816, 
    34.1475, 35, 35.86585, 36.74526, 37.63843, 38.54552, 39.46672, 40.40218, 
    41.35203, 42.31639, 43.29537, 44.28904, 45.29746, 46.32066, 47.35865, 
    48.4114, 49.47886, 50.56093, 51.6575, 52.7684, 53.89345, 55.0324, 
    56.18499, 57.35088, 58.52973, 59.72112, 60.92462, 62.13973, 63.36592, 
    64.6026, 65.84917, 67.10496, 68.36926, 69.64136, 70.92046, 72.20578, 
    73.49648, 74.79169, 76.09055, 77.39217, 78.69563, 80, 81.30437, 82.60783, 
    83.90945, 85.20831, 86.50352, 87.79422, 89.07954, 90.35864, 91.63074, 
    92.89504, 94.15083, 95.3974, 96.63409, 97.86027, 99.07538, 100.2789, 
    101.4703, 102.6491, 103.815, 104.9676, 106.1066, 107.2316, 108.3425, 
    109.4391, 110.5211, 111.5886, 112.6413, 113.6793, 114.7025, 115.711, 
    116.7046, 117.6836, 118.648, 119.5978, 120.5333, 121.4545, 122.3616, 
    123.2547, 124.1341, 125, 125.8525, 126.6918, 127.5183, 128.332, 129.1333, 
    129.9223, 130.6993, 131.4646,
  27.69435, 28.45444, 29.22681, 30.01174, 30.8095, 31.62036, 32.44458, 
    33.28242, 34.13415, 35, 35.88022, 36.77504, 37.68469, 38.60936, 39.54926, 
    40.50455, 41.47541, 42.46196, 43.46433, 44.4826, 45.51685, 46.56712, 
    47.63339, 48.71566, 49.81385, 50.92786, 52.05756, 53.20275, 54.36322, 
    55.53868, 56.72881, 57.93325, 59.15157, 60.3833, 61.62791, 62.88484, 
    64.15346, 65.4331, 66.72302, 68.02248, 69.33064, 70.64666, 71.96964, 
    73.29867, 74.63277, 75.97096, 77.31225, 78.65561, 80, 81.34439, 82.68775, 
    84.02904, 85.36723, 86.70133, 88.03036, 89.35334, 90.66936, 91.97752, 
    93.27698, 94.5669, 95.84654, 97.11516, 98.37209, 99.6167, 100.8484, 
    102.0667, 103.2712, 104.4613, 105.6368, 106.7972, 107.9424, 109.0721, 
    110.1861, 111.2843, 112.3666, 113.4329, 114.4831, 115.5174, 116.5357, 
    117.538, 118.5246, 119.4954, 120.4507, 121.3906, 122.3153, 123.225, 
    124.1198, 125, 125.8659, 126.7176, 127.5554, 128.3796, 129.1905, 
    129.9883, 130.7732, 131.5456, 132.3056,
  26.84588, 27.60006, 28.36704, 29.14713, 29.94063, 30.74784, 31.56906, 
    32.40459, 33.25474, 34.11978, 35, 35.89568, 36.80707, 37.73442, 38.67799, 
    39.63799, 40.61461, 41.60805, 42.61846, 43.64598, 44.69072, 45.75275, 
    46.83212, 47.92883, 49.04284, 50.1741, 51.32246, 52.48778, 53.66984, 
    54.86836, 56.08303, 57.31347, 58.55923, 59.81984, 61.09473, 62.3833, 
    63.68487, 64.9987, 66.32402, 67.65997, 69.00568, 70.36017, 71.72246, 
    73.09153, 74.46629, 75.84566, 77.2285, 78.61367, 80, 81.38633, 82.7715, 
    84.15434, 85.53371, 86.90847, 88.27754, 89.63983, 90.99432, 92.34003, 
    93.67598, 95.0013, 96.31513, 97.6167, 98.90527, 100.1802, 101.4408, 
    102.6865, 103.917, 105.1316, 106.3302, 107.5122, 108.6775, 109.8259, 
    110.9572, 112.0712, 113.1679, 114.2472, 115.3093, 116.354, 117.3815, 
    118.392, 119.3854, 120.362, 121.322, 122.2656, 123.1929, 124.1043, 125, 
    125.8802, 126.7453, 127.5954, 128.4309, 129.2522, 130.0594, 130.8529, 
    131.6329, 132.3999, 133.1541,
  25.98999, 26.73754, 27.49838, 28.27285, 29.0613, 29.86405, 30.68145, 
    31.51385, 32.36157, 33.22496, 34.10432, 35, 35.91229, 36.8415, 37.78791, 
    38.75179, 39.73339, 40.73296, 41.7507, 42.78679, 43.84139, 44.91462, 
    46.00657, 47.11728, 48.24677, 49.39498, 50.56185, 51.74722, 52.95089, 
    54.17262, 55.41209, 56.66891, 57.94265, 59.23279, 60.53875, 61.85987, 
    63.19543, 64.54465, 65.90668, 67.28057, 68.66535, 70.05998, 71.46335, 
    72.87431, 74.29166, 75.71419, 77.14061, 78.56965, 80, 81.43035, 82.85939, 
    84.28581, 85.70834, 87.12569, 88.53665, 89.94002, 91.33465, 92.71943, 
    94.09332, 95.45535, 96.80457, 98.14013, 99.46126, 100.7672, 102.0574, 
    103.3311, 104.5879, 105.8274, 107.0491, 108.2528, 109.4382, 110.605, 
    111.7532, 112.8827, 113.9934, 115.0854, 116.1586, 117.2132, 118.2493, 
    119.267, 120.2666, 121.2482, 122.2121, 123.1585, 124.0877, 125, 125.8957, 
    126.775, 127.6384, 128.4861, 129.3185, 130.136, 130.9387, 131.7271, 
    132.5016, 133.2625, 134.01,
  25.12669, 25.86687, 26.6208, 27.38887, 28.17145, 28.96892, 29.78166, 
    30.61005, 31.45448, 32.31531, 33.19293, 34.08771, 35, 35.93016, 36.87852, 
    37.84542, 38.83117, 39.83604, 40.86031, 41.90422, 42.96797, 44.05175, 
    45.15569, 46.2799, 47.42442, 48.58926, 49.77438, 50.97966, 52.20493, 
    53.44996, 54.71445, 55.99803, 57.30024, 58.62055, 59.95836, 61.31298, 
    62.68364, 64.06949, 65.4696, 66.88296, 68.30848, 69.74501, 71.19135, 
    72.64619, 74.10821, 75.57603, 77.04823, 78.52338, 80, 81.47662, 82.95177, 
    84.42397, 85.89179, 87.35381, 88.80865, 90.25499, 91.69152, 93.11704, 
    94.5304, 95.93051, 97.31636, 98.68702, 100.0416, 101.3794, 102.6998, 
    104.002, 105.2855, 106.55, 107.7951, 109.0203, 110.2256, 111.4107, 
    112.5756, 113.7201, 114.8443, 115.9482, 117.032, 118.0958, 119.1397, 
    120.164, 121.1688, 122.1546, 123.1215, 124.0698, 125, 125.9123, 126.8071, 
    127.6847, 128.5455, 129.39, 130.2183, 131.0311, 131.8286, 132.6111, 
    133.3792, 134.1331, 134.8733,
  24.256, 24.98804, 25.73429, 26.49515, 27.27104, 28.06237, 28.86957, 
    29.69306, 30.53328, 31.39064, 32.26558, 33.1585, 34.06984, 35, 35.94938, 
    36.91836, 37.90731, 38.91659, 39.94653, 40.99742, 42.06955, 43.16315, 
    44.27842, 45.41552, 46.57457, 47.75561, 48.95865, 50.18363, 51.4304, 
    52.69878, 53.98848, 55.29913, 56.63028, 57.9814, 59.35187, 60.74095, 
    62.14783, 63.5716, 65.01125, 66.46568, 67.93371, 69.41405, 70.90537, 
    72.40624, 73.91517, 75.43061, 76.95099, 78.47466, 80, 81.52534, 83.04901, 
    84.56939, 86.08483, 87.59376, 89.09463, 90.58595, 92.06629, 93.53432, 
    94.98875, 96.4284, 97.85217, 99.25905, 100.6481, 102.0186, 103.3697, 
    104.7009, 106.0115, 107.3012, 108.5696, 109.8164, 111.0414, 112.2444, 
    113.4254, 114.5845, 115.7216, 116.8369, 117.9305, 119.0026, 120.0535, 
    121.0834, 122.0927, 123.0816, 124.0506, 125, 125.9302, 126.8415, 
    127.7344, 128.6094, 129.4667, 130.3069, 131.1304, 131.9376, 132.729, 
    133.5049, 134.2657, 135.0119, 135.744,
  23.37793, 24.10108, 24.83885, 25.59168, 26.36002, 27.14434, 27.9451, 
    28.76277, 29.59782, 30.45074, 31.32201, 32.21209, 33.12148, 34.05062, 35, 
    35.97005, 36.96123, 37.97394, 39.00859, 40.06556, 41.14519, 42.24778, 
    43.37363, 44.52294, 45.6959, 46.89263, 48.11319, 49.35756, 50.62568, 
    51.91737, 53.23239, 54.57038, 55.93093, 57.31348, 58.7174, 60.14192, 
    61.58618, 63.04922, 64.52995, 66.02716, 67.53957, 69.06577, 70.60426, 
    72.15347, 73.71172, 75.27731, 76.84843, 78.42329, 80, 81.57671, 83.15157, 
    84.72269, 86.28828, 87.84653, 89.39574, 90.93423, 92.46043, 93.97284, 
    95.47005, 96.95078, 98.41382, 99.85809, 101.2826, 102.6865, 104.0691, 
    105.4296, 106.7676, 108.0826, 109.3743, 110.6424, 111.8868, 113.1074, 
    114.3041, 115.4771, 116.6264, 117.7522, 118.8548, 119.9344, 120.9914, 
    122.0261, 123.0388, 124.0299, 125, 125.9494, 126.8785, 127.7879, 128.678, 
    129.5493, 130.4022, 131.2372, 132.0549, 132.8557, 133.64, 134.4083, 
    135.1611, 135.8989, 136.6221,
  22.49251, 23.206, 23.93448, 24.67844, 25.43838, 26.21478, 27.00817, 
    27.81906, 28.64797, 29.49545, 30.36201, 31.24821, 32.15458, 33.08164, 
    34.02995, 35, 35.99232, 37.00741, 38.04575, 39.10778, 40.19393, 41.30461, 
    42.44015, 43.60088, 44.78704, 45.99885, 47.23642, 48.49981, 49.78901, 
    51.1039, 52.44429, 53.80986, 55.20019, 56.61475, 58.0529, 59.51385, 
    60.9967, 62.50041, 64.02381, 65.56562, 67.12441, 68.69864, 70.28666, 
    71.8867, 73.49693, 75.11539, 76.7401, 78.369, 80, 81.631, 83.2599, 
    84.88461, 86.50307, 88.1133, 89.71334, 91.30136, 92.87559, 94.43438, 
    95.97619, 97.4996, 99.0033, 100.4862, 101.9471, 103.3852, 104.7998, 
    106.1901, 107.5557, 108.8961, 110.211, 111.5002, 112.7636, 114.0012, 
    115.213, 116.3991, 117.5598, 118.6954, 119.8061, 120.8922, 121.9543, 
    122.9926, 124.0077, 125, 125.9701, 126.9184, 127.8454, 128.7518, 129.638, 
    130.5045, 131.352, 132.1809, 132.9918, 133.7852, 134.5616, 135.3216, 
    136.0655, 136.794, 137.5075,
  21.59979, 22.30283, 23.02121, 23.75546, 24.50609, 25.27366, 26.05873, 
    26.86185, 27.68361, 28.52459, 29.38539, 30.2666, 31.16883, 32.09269, 
    33.03877, 34.00768, 35, 36.01632, 37.05721, 38.1232, 39.21481, 40.33253, 
    41.47682, 42.64806, 43.8466, 45.07275, 46.3267, 47.60862, 48.91854, 
    50.25643, 51.62215, 53.01543, 54.43589, 55.88302, 57.35616, 58.85453, 
    60.37718, 61.92302, 63.49079, 65.07911, 66.68642, 68.31102, 69.9511, 
    71.6047, 73.26974, 74.94408, 76.62544, 78.31153, 80, 81.68847, 83.37456, 
    85.05592, 86.73026, 88.3953, 90.0489, 91.68898, 93.31358, 94.92089, 
    96.50921, 98.07699, 99.62282, 101.1455, 102.6438, 104.117, 105.5641, 
    106.9846, 108.3779, 109.7436, 111.0815, 112.3914, 113.6733, 114.9273, 
    116.1534, 117.3519, 118.5232, 119.6675, 120.7852, 121.8768, 122.9428, 
    123.9837, 125, 125.9923, 126.9612, 127.9073, 128.8312, 129.7334, 
    130.6146, 131.4754, 132.3164, 133.1382, 133.9413, 134.7263, 135.4939, 
    136.2445, 136.9788, 137.6972, 138.4002,
  20.69982, 21.39162, 22.09908, 22.82273, 23.56317, 24.32097, 25.09674, 
    25.89108, 26.70463, 27.53804, 28.39195, 29.26704, 30.16396, 31.08341, 
    32.02606, 32.99259, 33.98368, 35, 36.04221, 37.11095, 38.20685, 39.33048, 
    40.4824, 41.66312, 42.8731, 44.11272, 45.38232, 46.68213, 48.0123, 
    49.37288, 50.76379, 52.18483, 53.63569, 55.11587, 56.62475, 58.16152, 
    59.72521, 61.31467, 62.92859, 64.56543, 66.22353, 67.90104, 69.59592, 
    71.30601, 73.02899, 74.76245, 76.50385, 78.25058, 80, 81.74942, 83.49615, 
    85.23755, 86.97101, 88.69399, 90.40408, 92.09896, 93.77647, 95.43457, 
    97.07142, 98.68533, 100.2748, 101.8385, 103.3753, 104.8841, 106.3643, 
    107.8152, 109.2362, 110.6271, 111.9877, 113.3179, 114.6177, 115.8873, 
    117.1269, 118.3369, 119.5176, 120.6695, 121.7932, 122.889, 123.9578, 125, 
    126.0163, 127.0074, 127.9739, 128.9166, 129.836, 130.733, 131.608, 
    132.462, 133.2954, 134.1089, 134.9033, 135.679, 136.4368, 137.1773, 
    137.9009, 138.6084, 139.3002,
  19.79265, 20.47243, 21.16812, 21.88032, 22.60964, 23.35671, 24.12217, 
    24.90669, 25.71096, 26.53567, 27.38154, 28.2493, 29.13969, 30.05347, 
    30.9914, 31.95425, 32.94279, 33.95779, 35, 36.07018, 37.16905, 38.29732, 
    39.45566, 40.6447, 41.86501, 43.11712, 44.40147, 45.71841, 47.06821, 
    48.45102, 49.86686, 51.31562, 52.79705, 54.31071, 55.85601, 57.43214, 
    59.03812, 60.67276, 62.33465, 64.02217, 65.7335, 67.4666, 69.21925, 
    70.98902, 72.77335, 74.5695, 76.37463, 78.18579, 80, 81.81421, 83.62537, 
    85.4305, 87.22665, 89.01098, 90.78075, 92.5334, 94.2665, 95.97783, 
    97.66535, 99.32724, 100.9619, 102.5679, 104.144, 105.6893, 107.2029, 
    108.6844, 110.1331, 111.549, 112.9318, 114.2816, 115.5985, 116.8829, 
    118.135, 119.3553, 120.5443, 121.7027, 122.831, 123.9298, 125, 126.0422, 
    127.0572, 128.0457, 129.0086, 129.9465, 130.8603, 131.7507, 132.6185, 
    133.4643, 134.289, 135.0933, 135.8778, 136.6433, 137.3904, 138.1197, 
    138.8319, 139.5276, 140.2074,
  18.87837, 19.54531, 20.2284, 20.92826, 21.64553, 22.3809, 23.13504, 
    23.90867, 24.70254, 25.5174, 26.35402, 27.21321, 28.09578, 29.00258, 
    29.93444, 30.89222, 31.8768, 32.88905, 33.92982, 35, 36.10043, 37.23193, 
    38.39533, 39.59137, 40.82078, 42.08421, 43.38226, 44.7154, 46.08406, 
    47.48849, 48.92886, 50.40517, 51.91722, 53.4647, 55.04703, 56.66345, 
    58.31297, 59.99436, 61.70615, 63.4466, 65.21374, 67.00535, 68.81896, 
    70.6519, 72.50129, 74.36405, 76.23699, 78.11678, 80, 81.88322, 83.76301, 
    85.63595, 87.49871, 89.3481, 91.18104, 92.99465, 94.78626, 96.55341, 
    98.29385, 100.0056, 101.687, 103.3366, 104.953, 106.5353, 108.0828, 
    109.5948, 111.0711, 112.5115, 113.9159, 115.2846, 116.6177, 117.9158, 
    119.1792, 120.4086, 121.6047, 122.7681, 123.8996, 125, 126.0702, 127.111, 
    128.1232, 129.1078, 130.0656, 130.9974, 131.9042, 132.7868, 133.646, 
    134.4826, 135.2975, 136.0913, 136.865, 137.6191, 138.3545, 139.0717, 
    139.7716, 140.4547, 141.1216,
  17.95705, 18.61036, 19.28, 19.96662, 20.67091, 21.39358, 22.13536, 
    22.89701, 23.67934, 24.48314, 25.30928, 26.15861, 27.03203, 27.93045, 
    28.85481, 29.80607, 30.78519, 31.79315, 32.83095, 33.89957, 35, 36.1332, 
    37.30013, 38.50171, 39.73879, 41.01221, 42.32272, 43.67097, 45.05752, 
    46.48281, 47.94713, 49.45062, 50.99324, 52.57473, 54.19463, 55.8522, 
    57.54649, 59.27624, 61.03991, 62.83566, 64.66137, 66.51461, 68.39268, 
    70.29259, 72.21111, 74.1448, 76.09004, 78.04307, 80, 81.95693, 83.90996, 
    85.8552, 87.78889, 89.70741, 91.60732, 93.48539, 95.33863, 97.16434, 
    98.96009, 100.7238, 102.4535, 104.1478, 105.8054, 107.4253, 109.0068, 
    110.5494, 112.0529, 113.5172, 114.9425, 116.329, 117.6773, 118.9878, 
    120.2612, 121.4983, 122.6999, 123.8668, 125, 126.1004, 127.169, 128.2068, 
    129.2148, 130.1939, 131.1452, 132.0695, 132.968, 133.8414, 134.6907, 
    135.5169, 136.3207, 137.103, 137.8646, 138.6064, 139.3291, 140.0334, 
    140.72, 141.3896, 142.043,
  17.02878, 17.66766, 18.323, 18.99549, 19.68584, 20.39481, 21.12317, 
    21.87173, 22.64135, 23.43288, 24.24725, 25.08538, 25.94825, 26.83685, 
    27.75221, 28.69539, 29.66747, 30.66952, 31.70268, 32.76807, 33.8668, 35, 
    36.16879, 37.37423, 38.6174, 39.89928, 41.22082, 42.58285, 43.98613, 
    45.43129, 46.91879, 48.44895, 50.02188, 51.63745, 53.29532, 54.99484, 
    56.73508, 58.51479, 60.33239, 62.18593, 64.07315, 65.99139, 67.93768, 
    69.9087, 71.90084, 73.91022, 75.93275, 77.96415, 80, 82.03585, 84.06725, 
    86.08978, 88.09916, 90.0913, 92.06232, 94.00861, 95.92685, 97.81406, 
    99.66762, 101.4852, 103.2649, 105.0052, 106.7047, 108.3625, 109.9781, 
    111.551, 113.0812, 114.5687, 116.0139, 117.4172, 118.7792, 120.1007, 
    121.3826, 122.6258, 123.8312, 125, 126.1332, 127.2319, 128.2973, 
    129.3305, 130.3325, 131.3046, 132.2478, 133.1631, 134.0518, 134.9146, 
    135.7527, 136.5671, 137.3587, 138.1283, 138.8768, 139.6052, 140.3142, 
    141.0045, 141.677, 142.3323, 142.9712,
  16.09367, 16.71733, 17.35752, 18.01497, 18.69042, 19.38468, 20.09855, 
    20.83289, 21.5886, 22.36661, 23.16788, 23.99343, 24.84431, 25.72158, 
    26.62638, 27.55985, 28.52318, 29.5176, 30.54434, 31.60467, 32.69987, 
    33.83121, 35, 36.20749, 37.45493, 38.74353, 40.07444, 41.44871, 42.86732, 
    44.33112, 45.8408, 47.39688, 48.99965, 50.64919, 52.34529, 54.08742, 
    55.87473, 57.70599, 59.57961, 61.49355, 63.44538, 65.43224, 67.45084, 
    69.49753, 71.56824, 73.65859, 75.76395, 77.87943, 80, 82.12057, 84.23605, 
    86.34141, 88.43176, 90.50247, 92.54916, 94.56776, 96.55462, 98.50645, 
    100.4204, 102.294, 104.1253, 105.9126, 107.6547, 109.3508, 111.0003, 
    112.6031, 114.1592, 115.6689, 117.1327, 118.5513, 119.9256, 121.2565, 
    122.5451, 123.7925, 125, 126.1688, 127.3001, 128.3953, 129.4557, 
    130.4824, 131.4768, 132.4402, 133.3736, 134.2784, 135.1557, 136.0066, 
    136.8321, 137.6334, 138.4114, 139.1671, 139.9015, 140.6153, 141.3096, 
    141.985, 142.6425, 143.2827, 143.9063,
  15.15185, 15.75947, 16.38366, 17.02517, 17.68477, 18.36328, 19.06158, 
    19.78055, 20.52114, 21.28434, 22.07118, 22.88272, 23.7201, 24.58448, 
    25.47706, 26.39912, 27.35194, 28.33688, 29.3553, 30.40863, 31.49829, 
    32.62577, 33.79251, 35, 36.2497, 37.54304, 38.8814, 40.26611, 41.69838, 
    43.17933, 44.70991, 46.29089, 47.92281, 49.60596, 51.34034, 53.12559, 
    54.96098, 56.84534, 58.77709, 60.75413, 62.77388, 64.83324, 66.92863, 
    69.05596, 71.21069, 73.38788, 75.58224, 77.78819, 80, 82.21181, 84.41776, 
    86.61212, 88.78931, 90.94404, 93.07137, 95.16676, 97.22612, 99.24586, 
    101.2229, 103.1547, 105.039, 106.8744, 108.6597, 110.394, 112.0772, 
    113.7091, 115.2901, 116.8207, 118.3016, 119.7339, 121.1186, 122.457, 
    123.7503, 125, 126.2075, 127.3742, 128.5017, 129.5914, 130.6447, 
    131.6631, 132.6481, 133.6009, 134.5229, 135.4155, 136.2799, 137.1173, 
    137.9288, 138.7157, 139.4789, 140.2195, 140.9384, 141.6367, 142.3152, 
    142.9748, 143.6163, 144.2405, 144.8482,
  14.20343, 14.79423, 15.40157, 16.02623, 16.66901, 17.33076, 18.01239, 
    18.71483, 19.43907, 20.18615, 20.95716, 21.75323, 22.57558, 23.42543, 
    24.3041, 25.21295, 26.1534, 27.1269, 28.13499, 29.17922, 30.26121, 
    31.3826, 32.54507, 33.7503, 35, 36.29585, 37.6395, 39.03254, 40.47651, 
    41.9728, 43.52268, 45.12722, 46.78728, 48.50342, 50.27589, 52.10457, 
    53.98889, 55.92782, 57.91981, 59.96273, 62.05387, 64.18992, 66.36694, 
    68.58039, 70.8252, 73.09575, 75.38602, 77.68964, 80, 82.31036, 84.61398, 
    86.90425, 89.1748, 91.41961, 93.63306, 95.81008, 97.94613, 100.0373, 
    102.0802, 104.0722, 106.0111, 107.8954, 109.7241, 111.4966, 113.2127, 
    114.8728, 116.4773, 118.0272, 119.5235, 120.9675, 122.3605, 123.7042, 
    125, 126.2497, 127.4549, 128.6174, 129.7388, 130.8208, 131.865, 132.8731, 
    133.8466, 134.787, 135.6959, 136.5746, 137.4244, 138.2468, 139.0428, 
    139.8138, 140.5609, 141.2852, 141.9876, 142.6692, 143.331, 143.9738, 
    144.5984, 145.2058, 145.7966,
  13.24856, 13.82175, 14.4114, 15.01831, 15.6433, 16.28727, 16.95113, 
    17.63586, 18.3425, 19.07214, 19.82591, 20.60502, 21.41073, 22.24439, 
    23.10737, 24.00115, 24.92726, 25.88728, 26.88288, 27.91578, 28.98779, 
    30.10072, 31.25647, 32.45696, 33.70415, 35, 36.34645, 37.74542, 39.19877, 
    40.70824, 42.27547, 43.90189, 45.58871, 47.33686, 49.14692, 51.01906, 
    52.95296, 54.94778, 57.00206, 59.11371, 61.2799, 63.4971, 65.76101, 
    68.06663, 70.40823, 72.77946, 75.17344, 77.58282, 80, 82.41718, 84.82656, 
    87.22054, 89.59177, 91.93337, 94.23899, 96.5029, 98.7201, 100.8863, 
    102.9979, 105.0522, 107.047, 108.9809, 110.8531, 112.6631, 114.4113, 
    116.0981, 117.7245, 119.2918, 120.8012, 122.2546, 123.6535, 125, 
    126.2958, 127.543, 128.7435, 129.8993, 131.0122, 132.0842, 133.1171, 
    134.1127, 135.0727, 135.9988, 136.8926, 137.7556, 138.5893, 139.395, 
    140.1741, 140.9279, 141.6575, 142.3641, 143.0489, 143.7127, 144.3567, 
    144.9817, 145.5886, 146.1783, 146.7514,
  12.28739, 12.84219, 13.41332, 14.00158, 14.60783, 15.23297, 15.87796, 
    16.54382, 17.2316, 17.94244, 18.67754, 19.43815, 20.22562, 21.04135, 
    21.88682, 22.76358, 23.6733, 24.61768, 25.59853, 26.61774, 27.67728, 
    28.77918, 29.92556, 31.1186, 32.3605, 33.65355, 35, 36.40213, 37.86216, 
    39.38226, 40.96445, 42.61062, 44.32241, 46.10118, 47.94793, 49.86321, 
    51.84705, 53.89887, 56.01741, 58.20064, 60.44569, 62.74881, 65.10536, 
    67.50979, 69.95567, 72.4358, 74.94226, 77.46661, 80, 82.53339, 85.05774, 
    87.5642, 90.04433, 92.49021, 94.89464, 97.25119, 99.55431, 101.7994, 
    103.9826, 106.1011, 108.153, 110.1368, 112.0521, 113.8988, 115.6776, 
    117.3894, 119.0355, 120.6177, 122.1378, 123.5979, 125, 126.3465, 
    127.6395, 128.8814, 130.0744, 131.2208, 132.3227, 133.3823, 134.4015, 
    135.3823, 136.3267, 137.2364, 138.1132, 138.9586, 139.7744, 140.5618, 
    141.3225, 142.0576, 142.7684, 143.4562, 144.122, 144.767, 145.3922, 
    145.9984, 146.5867, 147.1578, 147.7126,
  11.32008, 11.85573, 12.40751, 12.97624, 13.56279, 14.16809, 14.79311, 
    15.4389, 16.10655, 16.79724, 17.51222, 18.25278, 19.02034, 19.81637, 
    20.64244, 21.50019, 22.39138, 23.31787, 24.28159, 25.28459, 26.32903, 
    27.41715, 28.55129, 29.73389, 30.96746, 32.25458, 33.59787, 35, 36.46361, 
    37.99131, 39.58562, 41.24892, 42.98337, 44.79087, 46.67292, 48.63058, 
    50.66433, 52.77399, 54.95856, 57.21618, 59.54401, 61.93813, 64.39354, 
    66.90412, 69.46265, 72.06094, 74.68987, 77.33966, 80, 82.66034, 85.31013, 
    87.93906, 90.53735, 93.09588, 95.60646, 98.06187, 100.456, 102.7838, 
    105.0414, 107.226, 109.3357, 111.3694, 113.3271, 115.2091, 117.0166, 
    118.7511, 120.4144, 122.0087, 123.5364, 125, 126.4021, 127.7454, 
    129.0325, 130.2661, 131.4487, 132.5829, 133.671, 134.7154, 135.7184, 
    136.6821, 137.6086, 138.4998, 139.3576, 140.1836, 140.9797, 141.7472, 
    142.4878, 143.2028, 143.8934, 144.5611, 145.2069, 145.8319, 146.4372, 
    147.0238, 147.5925, 148.1443, 148.6799,
  10.34682, 10.86256, 11.39418, 11.9425, 12.50841, 13.09284, 13.6968, 
    14.32134, 14.9676, 15.63678, 16.33016, 17.04911, 17.79507, 18.5696, 
    19.37432, 20.21099, 21.08146, 21.9877, 22.93179, 23.91594, 24.94248, 
    26.01387, 27.13268, 28.30161, 29.52349, 30.80123, 32.13784, 33.53639, 35, 
    36.53178, 38.13481, 39.81203, 41.56625, 43.39997, 45.31535, 47.31408, 
    49.39722, 51.56511, 53.8172, 56.15191, 58.5665, 61.05698, 63.618, 
    66.24284, 68.92341, 71.65034, 74.41312, 77.20037, 80, 82.79963, 85.58688, 
    88.34966, 91.07659, 93.75716, 96.382, 98.94302, 101.4335, 103.8481, 
    106.1828, 108.4349, 110.6028, 112.6859, 114.6847, 116.6, 118.4338, 
    120.188, 121.8652, 123.4682, 125, 126.4636, 127.8622, 129.1988, 130.4765, 
    131.6984, 132.8673, 133.9861, 135.0575, 136.0841, 137.0682, 138.0123, 
    138.9185, 139.789, 140.6257, 141.4304, 142.2049, 142.9509, 143.6698, 
    144.3632, 145.0324, 145.6787, 146.3032, 146.9072, 147.4916, 148.0575, 
    148.6058, 149.1374, 149.6532,
  9.367781, 9.862885, 10.37354, 10.90059, 11.44492, 12.00749, 12.58929, 
    13.19142, 13.81502, 14.46132, 15.13164, 15.82738, 16.55004, 17.30122, 
    18.08263, 18.8961, 19.74357, 20.62712, 21.54898, 22.51151, 23.51719, 
    24.56871, 25.66888, 26.82067, 28.0272, 29.29176, 30.61774, 32.00869, 
    33.46822, 35, 36.60772, 38.29502, 40.06539, 41.92211, 43.86813, 45.9059, 
    48.03725, 50.26324, 52.5839, 54.99814, 57.50347, 60.09591, 62.76982, 
    65.51788, 68.33101, 71.19851, 74.10822, 77.04679, 80, 82.95321, 85.89178, 
    88.80149, 91.66899, 94.48212, 97.23017, 99.9041, 102.4965, 105.0019, 
    107.4161, 109.7368, 111.9627, 114.0941, 116.1319, 118.0779, 119.9346, 
    121.705, 123.3923, 125, 126.5318, 127.9913, 129.3823, 130.7083, 131.9728, 
    133.1793, 134.3311, 135.4313, 136.4828, 137.4885, 138.451, 139.3729, 
    140.2564, 141.1039, 141.9174, 142.6988, 143.45, 144.1726, 144.8684, 
    145.5387, 146.185, 146.8086, 147.4107, 147.9925, 148.5551, 149.0994, 
    149.6264, 150.1371, 150.6322,
  8.383177, 8.856917, 9.345838, 9.850773, 10.37261, 10.91231, 11.47089, 
    12.04944, 12.64912, 13.27118, 13.91697, 14.58791, 15.28555, 16.01152, 
    16.76761, 17.55571, 18.37785, 19.23622, 20.13314, 21.07113, 22.05287, 
    23.08121, 24.1592, 25.29009, 26.47732, 27.72453, 29.03555, 30.41438, 
    31.86519, 33.39228, 35, 36.69275, 38.47487, 40.35052, 42.32358, 44.39749, 
    46.57505, 48.85823, 51.24794, 53.74372, 56.34361, 59.04377, 61.83841, 
    64.71956, 67.67712, 70.69882, 73.77054, 76.87655, 80, 83.12345, 86.22946, 
    89.30118, 92.32288, 95.28044, 98.1616, 100.9562, 103.6564, 106.2563, 
    108.7521, 111.1418, 113.4249, 115.6025, 117.6764, 119.6495, 121.5251, 
    123.3072, 125, 126.6077, 128.1348, 129.5856, 130.9644, 132.2755, 
    133.5227, 134.7099, 135.8408, 136.9188, 137.9471, 138.9289, 139.8669, 
    140.7638, 141.6221, 142.4443, 143.2324, 143.9885, 144.7144, 145.4121, 
    146.083, 146.7288, 147.3509, 147.9506, 148.5291, 149.0877, 149.6274, 
    150.1492, 150.6542, 151.1431, 151.6168,
  7.393215, 7.844895, 8.311317, 8.793312, 9.291768, 9.807635, 10.34193, 
    10.89576, 11.47027, 12.06675, 12.68653, 13.33109, 14.00197, 14.70088, 
    15.42961, 16.19014, 16.98457, 17.81517, 18.68438, 19.59484, 20.54938, 
    21.55105, 22.60312, 23.70911, 24.87277, 26.09811, 27.38938, 28.75108, 
    30.18797, 31.70498, 33.30725, 35, 36.78852, 38.67802, 40.67348, 42.77955, 
    45.00024, 47.33874, 49.79707, 52.37581, 55.07372, 57.88741, 60.81107, 
    63.83621, 66.95157, 70.14314, 73.39439, 76.68673, 80, 83.31327, 86.60561, 
    89.85686, 93.04843, 96.16379, 99.18893, 102.1126, 104.9263, 107.6242, 
    110.2029, 112.6613, 114.9998, 117.2204, 119.3265, 121.322, 123.2115, 125, 
    126.6928, 128.295, 129.812, 131.2489, 132.6106, 133.9019, 135.1272, 
    136.2909, 137.3969, 138.449, 139.4506, 140.4052, 141.3156, 142.1848, 
    143.0154, 143.8099, 144.5704, 145.2991, 145.998, 146.6689, 147.3135, 
    147.9333, 148.5297, 149.1042, 149.6581, 150.1924, 150.7082, 151.2067, 
    151.6887, 152.1551, 152.6068,
  6.39812, 6.827063, 7.270251, 7.728505, 8.202703, 8.693789, 9.202773, 
    9.730745, 10.27888, 10.84843, 11.44077, 12.05735, 12.69976, 13.36972, 
    14.06907, 14.79981, 15.56411, 16.36431, 17.20295, 18.08277, 19.00676, 
    19.97812, 21.00035, 22.07719, 23.21272, 24.41129, 25.67759, 27.01663, 
    28.43375, 29.93461, 31.52513, 33.21148, 35, 36.89709, 38.90907, 41.04199, 
    43.30139, 45.69201, 48.2174, 50.87953, 53.67833, 56.6112, 59.6726, 
    62.85364, 66.14191, 69.52138, 72.97269, 76.47366, 80, 83.52634, 87.02731, 
    90.47862, 93.85809, 97.14635, 100.3274, 103.3888, 106.3217, 109.1205, 
    111.7826, 114.308, 116.6986, 118.958, 121.0909, 123.1029, 125, 126.7885, 
    128.4749, 130.0654, 131.5662, 132.9834, 134.3224, 135.5887, 136.7873, 
    137.9228, 138.9996, 140.0219, 140.9932, 141.9172, 142.7971, 143.6357, 
    144.4359, 145.2002, 145.9309, 146.6303, 147.3002, 147.9427, 148.5592, 
    149.1516, 149.7211, 150.2693, 150.7972, 151.3062, 151.7973, 152.2715, 
    152.7298, 153.1729, 153.6019,
  5.398128, 5.80368, 6.222924, 6.656663, 7.105759, 7.57114, 8.053806, 
    8.554832, 9.075379, 9.616703, 10.18016, 10.76721, 11.37945, 12.01859, 
    12.68652, 13.38525, 14.11698, 14.88413, 15.68929, 16.5353, 17.42527, 
    18.36255, 19.35081, 20.39404, 21.49658, 22.66313, 23.89882, 25.20913, 
    26.60003, 28.07789, 29.64948, 31.32199, 33.10291, 35, 37.0211, 39.17396, 
    41.46598, 43.90385, 46.49313, 49.23772, 52.13926, 55.19647, 58.40453, 
    61.75444, 65.23267, 68.82096, 72.49654, 76.23273, 80, 83.76727, 87.50346, 
    91.17904, 94.76733, 98.24556, 101.5955, 104.8035, 107.8607, 110.7623, 
    113.5069, 116.0961, 118.534, 120.826, 122.9789, 125, 126.8971, 128.678, 
    130.3505, 131.9221, 133.4, 134.7909, 136.1012, 137.3369, 138.5034, 
    139.606, 140.6492, 141.6375, 142.5747, 143.4647, 144.3107, 145.1159, 
    145.883, 146.6148, 147.3135, 147.9814, 148.6205, 149.2328, 149.8198, 
    150.3833, 150.9246, 151.4452, 151.9462, 152.4289, 152.8942, 153.3433, 
    153.7771, 154.1963, 154.6019,
  4.393482, 4.775022, 5.16964, 5.578118, 6.001298, 6.440085, 6.895458, 
    7.368472, 7.86027, 8.372087, 8.905264, 9.461254, 10.04164, 10.64813, 
    11.28261, 11.9471, 12.64384, 13.37525, 14.14399, 14.95297, 15.80537, 
    16.70468, 17.65471, 18.65966, 19.7241, 20.85308, 22.05207, 23.32708, 
    24.68465, 26.13187, 27.67642, 29.32652, 31.09093, 32.9789, 35, 37.16397, 
    39.48043, 41.95853, 44.60641, 47.43058, 50.43513, 53.62088, 56.98439, 
    60.51708, 64.2045, 68.02593, 71.95453, 75.958, 80, 84.042, 88.04547, 
    91.97407, 95.7955, 99.48292, 103.0156, 106.3791, 109.5649, 112.5694, 
    115.3936, 118.0415, 120.5196, 122.836, 125, 127.0211, 128.9091, 130.6735, 
    132.3236, 133.8681, 135.3154, 136.6729, 137.9479, 139.1469, 140.2759, 
    141.3403, 142.3453, 143.2953, 144.1946, 145.047, 145.856, 146.6248, 
    147.3562, 148.0529, 148.7174, 149.3519, 149.9584, 150.5387, 151.0947, 
    151.6279, 152.1397, 152.6315, 153.1045, 153.5599, 153.9987, 154.4219, 
    154.8304, 155.225, 155.6065,
  3.384442, 3.741373, 4.110714, 4.49322, 4.889704, 5.301043, 5.728187, 
    6.172163, 6.634083, 7.115158, 7.616698, 8.140132, 8.687016, 9.259048, 
    9.858084, 10.48615, 11.14547, 11.83848, 12.56786, 13.33655, 14.1478, 
    15.00516, 15.91258, 16.87441, 17.89543, 18.98094, 20.13679, 21.36942, 
    22.68592, 24.09411, 25.60251, 27.22045, 28.95801, 30.82604, 32.83603, 35, 
    37.33021, 39.83878, 42.53716, 45.43531, 48.5408, 51.85757, 55.38464, 
    59.11468, 63.03281, 67.11578, 71.33189, 75.64172, 80, 84.35828, 88.66811, 
    92.88422, 96.96719, 100.8853, 104.6154, 108.1424, 111.4592, 114.5647, 
    117.4628, 120.1612, 122.6698, 125, 127.164, 129.174, 131.042, 132.7796, 
    134.3975, 135.9059, 137.3141, 138.6306, 139.8632, 141.0191, 142.1046, 
    143.1256, 144.0874, 144.9948, 145.8522, 146.6635, 147.4321, 148.1615, 
    148.8545, 149.5139, 150.1419, 150.741, 151.313, 151.8599, 152.3833, 
    152.8848, 153.3659, 153.8278, 154.2718, 154.699, 155.1103, 155.5068, 
    155.8893, 156.2586, 156.6156,
  2.371273, 2.703033, 3.046482, 3.402338, 3.771384, 4.154459, 4.55248, 
    4.966434, 5.397398, 5.846539, 6.315132, 6.804565, 7.316357, 7.852167, 
    8.413816, 9.003303, 9.622821, 10.27479, 10.96188, 11.68703, 12.45351, 
    13.26492, 14.12528, 15.03902, 16.01111, 17.04704, 18.15295, 19.33566, 
    20.60278, 21.96275, 23.42495, 24.99976, 26.69861, 28.53402, 30.51957, 
    32.66979, 35, 37.52589, 40.263, 43.22584, 46.42671, 49.8742, 53.5713, 
    57.51336, 61.68604, 66.06376, 70.60912, 75.27358, 80, 84.72642, 89.39088, 
    93.93624, 98.31396, 102.4866, 106.4287, 110.1258, 113.5733, 116.7742, 
    119.737, 122.4741, 125, 127.3302, 129.4804, 131.466, 133.3014, 135.0002, 
    136.5751, 138.0372, 139.3972, 140.6643, 141.847, 142.953, 143.9889, 
    144.961, 145.8747, 146.7351, 147.5465, 148.313, 149.0381, 149.7252, 
    150.3772, 150.9967, 151.5862, 152.1478, 152.6836, 153.1954, 153.6849, 
    154.1535, 154.6026, 155.0336, 155.4475, 155.8455, 156.2286, 156.5977, 
    156.9535, 157.297, 157.6287,
  1.354252, 1.660314, 1.977288, 2.305858, 2.646764, 3.000807, 3.368856, 
    3.751855, 4.150831, 4.566904, 5.001296, 5.455343, 5.930508, 6.428399, 
    6.950779, 7.499593, 8.076985, 8.685326, 9.32724, 10.00564, 10.72376, 
    11.48521, 12.29401, 13.15465, 14.07218, 15.05222, 16.10113, 17.22602, 
    18.43489, 19.73676, 21.14176, 22.66126, 24.30799, 26.09615, 28.04147, 
    30.16122, 32.47411, 35, 37.75941, 40.77262, 44.05833, 47.6318, 51.50228, 
    55.67005, 60.12311, 64.83437, 69.75993, 74.83959, 80, 85.16041, 90.24007, 
    95.16563, 99.87689, 104.33, 108.4977, 112.3682, 115.9417, 119.2274, 
    122.2406, 125, 127.5259, 129.8388, 131.9585, 133.9039, 135.692, 137.3387, 
    138.8582, 140.2632, 141.5651, 142.774, 143.8989, 144.9478, 145.9278, 
    146.8454, 147.706, 148.5148, 149.2762, 149.9944, 150.6728, 151.3147, 
    151.923, 152.5004, 153.0492, 153.5716, 154.0695, 154.5447, 154.9987, 
    155.4331, 155.8492, 156.2481, 156.6311, 156.9992, 157.3532, 157.6941, 
    158.0227, 158.3397, 158.6458,
  0.3336662, 0.6135356, 0.9034941, 1.204182, 1.516293, 1.840581, 2.177862, 
    2.529026, 2.895045, 3.276976, 3.675979, 4.093322, 4.530401, 4.988749, 
    5.470056, 5.976187, 6.50921, 7.071416, 7.665351, 8.293855, 8.960093, 
    9.667614, 10.42039, 11.22291, 12.08019, 12.99794, 13.98259, 15.04144, 
    16.1828, 17.4161, 18.75206, 20.20293, 21.7826, 23.50687, 25.39359, 
    27.46284, 29.73699, 32.24059, 35, 38.04266, 41.39567, 45.08361, 49.1253, 
    53.52949, 58.2898, 63.37957, 68.74813, 74.32022, 80, 85.67978, 91.25187, 
    96.62043, 101.7102, 106.4705, 110.8747, 114.9164, 118.6043, 121.9573, 
    125, 127.7594, 130.263, 132.5372, 134.6064, 136.4931, 138.2174, 139.7971, 
    141.2479, 142.5839, 143.8172, 144.9586, 146.0174, 147.0021, 147.9198, 
    148.7771, 149.5796, 150.3324, 151.0399, 151.7061, 152.3347, 152.9286, 
    153.4908, 154.0238, 154.5299, 155.0112, 155.4696, 155.9067, 156.324, 
    156.723, 157.1049, 157.471, 157.8221, 158.1594, 158.4837, 158.7958, 
    159.0965, 159.3865, 159.6663,
  359.3098, 359.563, 359.8255, 0.09772872, 0.3804374, 0.6742983, 0.9800709, 
    1.298583, 1.630737, 1.977523, 2.340024, 2.719428, 3.117045, 3.534317, 
    3.97284, 4.434379, 4.920894, 5.434566, 5.977829, 6.553403, 7.164339, 
    7.814067, 8.506453, 9.245869, 10.03727, 10.88629, 11.79936, 12.78382, 
    13.84809, 15.00186, 16.25627, 17.62419, 19.12047, 20.76228, 22.56942, 
    24.56469, 26.77416, 29.22738, 31.95734, 35, 38.39312, 42.17395, 46.37541, 
    51.02029, 56.11345, 61.633, 67.52246, 73.68741, 80, 86.31259, 92.47754, 
    98.367, 103.8865, 108.9797, 113.6246, 117.8261, 121.6069, 125, 128.0427, 
    130.7726, 133.2258, 135.4353, 137.4306, 139.2377, 140.8795, 142.3758, 
    143.7437, 144.9981, 146.1519, 147.2162, 148.2006, 149.1137, 149.9627, 
    150.7541, 151.4935, 152.1859, 152.8357, 153.4466, 154.0222, 154.5654, 
    155.0791, 155.5656, 156.0272, 156.4657, 156.8829, 157.2806, 157.66, 
    158.0225, 158.3693, 158.7014, 159.0199, 159.3257, 159.6196, 159.9023, 
    160.1745, 160.437, 160.6902,
  358.283, 358.5092, 358.7436, 358.9869, 359.2397, 359.5025, 359.7761, 
    0.0611895, 0.3586455, 0.6693593, 0.9943273, 1.334645, 1.691522, 2.066292, 
    2.460434, 2.875589, 3.313586, 3.776463, 4.266501, 4.786263, 5.338629, 
    5.926853, 6.554621, 7.226121, 7.946126, 8.720099, 9.554314, 10.45599, 
    11.4335, 12.49653, 13.65639, 14.92628, 16.32167, 17.86074, 19.56487, 
    21.4592, 23.57329, 25.94167, 28.60433, 31.60689, 35, 38.83752, 43.17246, 
    48.04982, 53.49538, 59.50083, 66.00814, 72.89935, 80, 87.10065, 93.99186, 
    100.4992, 106.5046, 111.9502, 116.8275, 121.1625, 125, 128.3931, 
    131.3957, 134.0583, 136.4267, 138.5408, 140.4351, 142.1393, 143.6783, 
    145.0737, 146.3436, 147.5035, 148.5665, 149.544, 150.4457, 151.2799, 
    152.0539, 152.7739, 153.4454, 154.0732, 154.6614, 155.2137, 155.7335, 
    156.2235, 156.6864, 157.1244, 157.5396, 157.9337, 158.3085, 158.6654, 
    159.0057, 159.3306, 159.6414, 159.9388, 160.2239, 160.4975, 160.7603, 
    161.0131, 161.2564, 161.4909, 161.717,
  357.2535, 357.4522, 357.6583, 357.8722, 358.0945, 358.3257, 358.5665, 
    358.8175, 359.0795, 359.3533, 359.6398, 359.94, 0.2549859, 0.5859436, 
    0.9342362, 1.301358, 1.688978, 2.098961, 2.533401, 2.994655, 3.485386, 
    4.008612, 4.567762, 5.166756, 5.810081, 6.502903, 7.25119, 8.061871, 
    8.943019, 9.904095, 10.95623, 12.11259, 13.3888, 14.80353, 16.37912, 
    18.14243, 20.1258, 22.3682, 24.91639, 27.82605, 31.16248, 35, 39.41894, 
    44.49806, 50.29985, 56.84695, 64.09196, 71.89101, 80, 88.10899, 95.90804, 
    103.153, 109.7001, 115.5019, 120.5811, 125, 128.8375, 132.174, 135.0836, 
    137.6318, 139.8742, 141.8576, 143.6209, 145.1965, 146.6112, 147.8874, 
    149.0438, 150.0959, 151.057, 151.9381, 152.7488, 153.4971, 154.1899, 
    154.8332, 155.4322, 155.9914, 156.5146, 157.0053, 157.4666, 157.901, 
    158.311, 158.6986, 159.0658, 159.4141, 159.745, 160.06, 160.3602, 
    160.6467, 160.9205, 161.1825, 161.4335, 161.6743, 161.9055, 162.1278, 
    162.3417, 162.5478, 162.7465,
  356.2217, 356.3926, 356.57, 356.7541, 356.9455, 357.1446, 357.3521, 
    357.5684, 357.7942, 358.0304, 358.2775, 358.5367, 358.8087, 359.0946, 
    359.3958, 359.7133, 0.04889843, 0.4040801, 0.7807565, 1.18104, 1.607323, 
    2.062325, 2.549154, 3.071369, 3.633067, 4.238988, 4.89464, 5.606458, 
    6.381995, 7.230175, 8.161595, 9.188926, 10.3274, 11.59547, 13.01561, 
    14.61536, 16.4287, 18.49772, 20.8747, 23.62459, 26.82754, 30.58106, 35, 
    40.21146, 46.33897, 53.46891, 61.59522, 70.55551, 80, 89.44449, 98.40478, 
    106.5311, 113.661, 119.7885, 125, 129.4189, 133.1725, 136.3754, 139.1253, 
    141.5023, 143.5713, 145.3846, 146.9844, 148.4045, 149.6726, 150.8111, 
    151.8384, 152.7698, 153.618, 154.3935, 155.1054, 155.761, 156.3669, 
    156.9286, 157.4509, 157.9377, 158.3927, 158.819, 159.2192, 159.5959, 
    159.9511, 160.2867, 160.6043, 160.9054, 161.1913, 161.4633, 161.7225, 
    161.9697, 162.2058, 162.4316, 162.648, 162.8554, 163.0545, 163.2459, 
    163.43, 163.6074, 163.7783,
  355.1878, 355.3307, 355.479, 355.633, 355.7931, 355.9597, 356.1333, 
    356.3144, 356.5035, 356.7013, 356.9085, 357.1257, 357.3538, 357.5938, 
    357.8465, 358.1133, 358.3953, 358.694, 359.011, 359.3481, 359.7074, 
    0.09130464, 0.5024734, 0.9440413, 1.419612, 1.933374, 2.490215, 3.09588, 
    3.757156, 4.482118, 5.280438, 6.163786, 7.146357, 8.245557, 9.482918, 
    10.88532, 12.48664, 14.32995, 16.47051, 18.97971, 21.95018, 25.50194, 
    29.78854, 35, 41.354, 49.05843, 58.22134, 68.70457, 80, 91.29543, 
    101.7787, 110.9416, 118.646, 125, 130.2115, 134.4981, 138.0498, 141.0203, 
    143.5295, 145.67, 147.5134, 149.1147, 150.5171, 151.7544, 152.8536, 
    153.8362, 154.7196, 155.5179, 156.2428, 156.9041, 157.5098, 158.0666, 
    158.5804, 159.056, 159.4975, 159.9087, 160.2926, 160.6519, 160.989, 
    161.306, 161.6047, 161.8867, 162.1535, 162.4062, 162.6462, 162.8743, 
    163.0915, 163.2987, 163.4965, 163.6856, 163.8667, 164.0403, 164.2069, 
    164.367, 164.521, 164.6693, 164.8122,
  354.1523, 354.2669, 354.3859, 354.5094, 354.6379, 354.7716, 354.911, 
    355.0564, 355.2083, 355.3672, 355.5337, 355.7083, 355.8918, 356.0848, 
    356.2883, 356.5031, 356.7303, 356.971, 357.2267, 357.4987, 357.7889, 
    358.0992, 358.4318, 358.7893, 359.1748, 359.5918, 0.04433093, 0.5373426, 
    1.076589, 1.668989, 2.322887, 3.048434, 3.858094, 4.767325, 5.795501, 
    6.967195, 8.313965, 9.876889, 11.7102, 13.88655, 16.50462, 19.70015, 
    23.66103, 28.646, 35, 43.14066, 53.45003, 65.97485, 80, 94.02515, 106.55, 
    116.8593, 125, 131.354, 136.339, 140.2999, 143.4954, 146.1134, 148.2898, 
    150.1231, 151.686, 153.0328, 154.2045, 155.2327, 156.1419, 156.9516, 
    157.6771, 158.331, 158.9234, 159.4627, 159.9557, 160.4082, 160.8252, 
    161.2107, 161.5682, 161.9008, 162.2111, 162.5013, 162.7733, 163.029, 
    163.2697, 163.4969, 163.7117, 163.9152, 164.1082, 164.2917, 164.4663, 
    164.6328, 164.7917, 164.9436, 165.089, 165.2284, 165.3621, 165.4906, 
    165.6141, 165.7331, 165.8477,
  353.1154, 353.2016, 353.291, 353.3838, 353.4804, 353.581, 353.6858, 
    353.7951, 353.9095, 354.029, 354.1543, 354.2858, 354.424, 354.5694, 
    354.7227, 354.8846, 355.0559, 355.2375, 355.4305, 355.636, 355.8552, 
    356.0898, 356.3414, 356.6121, 356.9043, 357.2206, 357.5642, 357.9391, 
    358.3497, 358.8015, 359.3012, 359.8569, 0.4786234, 1.179037, 1.974067, 
    2.884218, 3.936238, 5.165633, 6.620432, 8.366995, 10.49917, 13.15305, 
    16.53109, 20.94157, 26.85934, 35, 46.31718, 61.57259, 80, 98.42741, 
    113.6828, 125, 133.1407, 139.0584, 143.4689, 146.847, 149.5008, 151.633, 
    153.3796, 154.8344, 156.0638, 157.1158, 158.0259, 158.821, 159.5214, 
    160.1431, 160.6988, 161.1985, 161.6503, 162.0609, 162.4358, 162.7795, 
    163.0957, 163.3879, 163.6586, 163.9102, 164.1448, 164.3641, 164.5695, 
    164.7625, 164.9441, 165.1154, 165.2773, 165.4306, 165.576, 165.7142, 
    165.8457, 165.971, 166.0906, 166.2048, 166.3142, 166.4191, 166.5196, 
    166.6162, 166.709, 166.7984, 166.8846,
  352.0775, 352.135, 352.1947, 352.2567, 352.3212, 352.3884, 352.4584, 
    352.5315, 352.6078, 352.6877, 352.7715, 352.8594, 352.9518, 353.049, 
    353.1516, 353.2599, 353.3746, 353.4962, 353.6254, 353.763, 353.9099, 
    354.0672, 354.2361, 354.4178, 354.614, 354.8266, 355.0577, 355.3101, 
    355.5869, 355.8918, 356.2295, 356.6056, 357.0273, 357.5034, 358.0455, 
    358.6681, 359.3909, 0.2400689, 1.25187, 2.477536, 3.991861, 5.908033, 
    8.404778, 11.77866, 16.54997, 23.68282, 35, 53.43872, 80, 106.5613, 125, 
    136.3172, 143.45, 148.2213, 151.5952, 154.092, 156.0081, 157.5225, 
    158.7481, 159.7599, 160.6091, 161.3319, 161.9545, 162.4965, 162.9727, 
    163.3944, 163.7705, 164.1082, 164.4131, 164.6899, 164.9423, 165.1734, 
    165.386, 165.5822, 165.7639, 165.9328, 166.09, 166.237, 166.3746, 
    166.5038, 166.6254, 166.7401, 166.8484, 166.951, 167.0482, 167.1406, 
    167.2285, 167.3123, 167.3922, 167.4685, 167.5416, 167.6116, 167.6788, 
    167.7433, 167.8053, 167.865, 167.9225,
  351.0389, 351.0677, 351.0976, 351.1286, 351.1609, 351.1945, 351.2296, 
    351.2661, 351.3044, 351.3444, 351.3863, 351.4304, 351.4766, 351.5253, 
    351.5767, 351.631, 351.6885, 351.7494, 351.8142, 351.8832, 351.9569, 
    352.0359, 352.1206, 352.2118, 352.3104, 352.4172, 352.5334, 352.6603, 
    352.7996, 352.9532, 353.1234, 353.3133, 353.5263, 353.7673, 354.042, 
    354.3583, 354.7264, 355.1604, 355.6798, 356.3126, 357.1006, 358.109, 
    359.4445, 1.295434, 4.025157, 8.427411, 16.56128, 35, 80, 125, 143.4387, 
    151.5726, 155.9748, 158.7046, 160.5555, 161.891, 162.8994, 163.6874, 
    164.3202, 164.8396, 165.2736, 165.6417, 165.958, 166.2327, 166.4737, 
    166.6867, 166.8766, 167.0468, 167.2004, 167.3397, 167.4666, 167.5828, 
    167.6897, 167.7882, 167.8794, 167.9641, 168.0431, 168.1168, 168.1858, 
    168.2506, 168.3115, 168.369, 168.4233, 168.4747, 168.5234, 168.5697, 
    168.6137, 168.6556, 168.6956, 168.7339, 168.7704, 168.8055, 168.8391, 
    168.8714, 168.9024, 168.9323, 168.9611,
  350, 350, 350, 350, 350, 350, 350, 350, 350, 350, 350, 350, 350, 350, 350, 
    350, 350, 350, 350, 350, 350, 350, 350, 350, 350, 350, 350, 350, 350, 
    350, 350, 350, 350, 350, 350, 350, 350, 350, 350, 350, 350, 350, 350, 
    350, 350, 350, 350, 350, 350, 170, 170, 170, 170, 170, 170, 170, 170, 
    170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 
    170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 
    170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170,
  348.9611, 348.9323, 348.9024, 348.8714, 348.8391, 348.8055, 348.7704, 
    348.7339, 348.6956, 348.6556, 348.6137, 348.5696, 348.5234, 348.4747, 
    348.4233, 348.369, 348.3115, 348.2506, 348.1858, 348.1168, 348.0431, 
    347.9641, 347.8794, 347.7882, 347.6896, 347.5828, 347.4666, 347.3397, 
    347.2004, 347.0468, 346.8766, 346.6867, 346.4737, 346.2327, 345.958, 
    345.6417, 345.2736, 344.8396, 344.3202, 343.6874, 342.8994, 341.891, 
    340.5555, 338.7046, 335.9749, 331.5726, 323.4387, 305, 260, 215, 
    196.5613, 188.4274, 184.0252, 181.2954, 179.4445, 178.109, 177.1006, 
    176.3126, 175.6798, 175.1604, 174.7264, 174.3583, 174.042, 173.7673, 
    173.5263, 173.3133, 173.1234, 172.9532, 172.7996, 172.6603, 172.5334, 
    172.4172, 172.3103, 172.2118, 172.1206, 172.0359, 171.9569, 171.8832, 
    171.8142, 171.7494, 171.6885, 171.631, 171.5767, 171.5253, 171.4766, 
    171.4303, 171.3863, 171.3444, 171.3044, 171.2661, 171.2296, 171.1945, 
    171.1609, 171.1286, 171.0976, 171.0677, 171.0389,
  347.9225, 347.865, 347.8053, 347.7433, 347.6788, 347.6116, 347.5416, 
    347.4685, 347.3922, 347.3123, 347.2285, 347.1406, 347.0482, 346.951, 
    346.8484, 346.7401, 346.6254, 346.5038, 346.3746, 346.237, 346.0901, 
    345.9328, 345.7639, 345.5822, 345.386, 345.1734, 344.9423, 344.6899, 
    344.4131, 344.1082, 343.7705, 343.3944, 342.9727, 342.4966, 341.9545, 
    341.3319, 340.6091, 339.7599, 338.7481, 337.5225, 336.0081, 334.092, 
    331.5952, 328.2213, 323.45, 316.3172, 305, 286.5613, 260, 233.4387, 215, 
    203.6828, 196.55, 191.7787, 188.4048, 185.908, 183.9919, 182.4775, 
    181.2519, 180.2401, 179.3909, 178.6681, 178.0455, 177.5035, 177.0273, 
    176.6056, 176.2295, 175.8918, 175.5869, 175.3101, 175.0577, 174.8266, 
    174.614, 174.4178, 174.2361, 174.0672, 173.91, 173.763, 173.6254, 
    173.4962, 173.3746, 173.2599, 173.1516, 173.049, 172.9518, 172.8594, 
    172.7715, 172.6877, 172.6078, 172.5315, 172.4584, 172.3884, 172.3212, 
    172.2567, 172.1947, 172.135, 172.0775,
  346.8846, 346.7984, 346.709, 346.6162, 346.5196, 346.419, 346.3142, 
    346.2049, 346.0905, 345.971, 345.8457, 345.7142, 345.576, 345.4306, 
    345.2773, 345.1154, 344.9441, 344.7625, 344.5695, 344.364, 344.1448, 
    343.9102, 343.6586, 343.3879, 343.0957, 342.7794, 342.4358, 342.0609, 
    341.6503, 341.1985, 340.6988, 340.1431, 339.5214, 338.821, 338.0259, 
    337.1158, 336.0638, 334.8344, 333.3796, 331.633, 329.5008, 326.847, 
    323.4689, 319.0584, 313.1407, 305, 293.6828, 278.4274, 260, 241.5726, 
    226.3172, 215, 206.8593, 200.9416, 196.5311, 193.153, 190.4992, 188.367, 
    186.6204, 185.1656, 183.9362, 182.8842, 181.9741, 181.179, 180.4786, 
    179.8569, 179.3012, 178.8015, 178.3497, 177.9391, 177.5642, 177.2205, 
    176.9043, 176.6121, 176.3414, 176.0898, 175.8552, 175.6359, 175.4305, 
    175.2375, 175.0559, 174.8846, 174.7227, 174.5694, 174.424, 174.2858, 
    174.1543, 174.029, 173.9094, 173.7952, 173.6858, 173.5809, 173.4804, 
    173.3838, 173.291, 173.2016, 173.1154,
  345.8477, 345.7331, 345.6141, 345.4906, 345.3621, 345.2284, 345.089, 
    344.9436, 344.7917, 344.6328, 344.4663, 344.2917, 344.1082, 343.9152, 
    343.7117, 343.4969, 343.2697, 343.029, 342.7733, 342.5013, 342.2111, 
    341.9008, 341.5682, 341.2107, 340.8252, 340.4082, 339.9557, 339.4626, 
    338.9234, 338.331, 337.6771, 336.9516, 336.1419, 335.2327, 334.2045, 
    333.0328, 331.686, 330.1231, 328.2898, 326.1135, 323.4954, 320.2998, 
    316.339, 311.354, 305, 296.8593, 286.55, 274.0251, 260, 245.9748, 233.45, 
    223.1407, 215, 208.646, 203.661, 199.7001, 196.5046, 193.8866, 191.7102, 
    189.8769, 188.314, 186.9672, 185.7955, 184.7673, 183.8581, 183.0484, 
    182.3229, 181.669, 181.0766, 180.5373, 180.0443, 179.5918, 179.1748, 
    178.7893, 178.4318, 178.0992, 177.7889, 177.4987, 177.2267, 176.971, 
    176.7303, 176.5031, 176.2883, 176.0848, 175.8918, 175.7083, 175.5337, 
    175.3672, 175.2083, 175.0564, 174.911, 174.7716, 174.6379, 174.5094, 
    174.3859, 174.2669, 174.1523,
  344.8122, 344.6693, 344.521, 344.367, 344.2069, 344.0403, 343.8667, 
    343.6856, 343.4965, 343.2987, 343.0915, 342.8743, 342.6462, 342.4062, 
    342.1535, 341.8867, 341.6047, 341.306, 340.989, 340.6519, 340.2926, 
    339.9087, 339.4975, 339.056, 338.5804, 338.0666, 337.5098, 336.9041, 
    336.2429, 335.5179, 334.7196, 333.8362, 332.8536, 331.7545, 330.5171, 
    329.1147, 327.5134, 325.67, 323.5295, 321.0203, 318.0498, 314.498, 
    310.2115, 305, 298.646, 290.9416, 281.7787, 271.2954, 260, 248.7046, 
    238.2213, 229.0584, 221.354, 215, 209.7885, 205.5019, 201.9502, 198.9797, 
    196.4705, 194.33, 192.4866, 190.8853, 189.4829, 188.2456, 187.1464, 
    186.1638, 185.2804, 184.4821, 183.7572, 183.0959, 182.4902, 181.9334, 
    181.4196, 180.944, 180.5025, 180.0913, 179.7074, 179.3481, 179.011, 
    178.694, 178.3953, 178.1133, 177.8465, 177.5938, 177.3538, 177.1257, 
    176.9085, 176.7013, 176.5035, 176.3144, 176.1333, 175.9597, 175.7931, 
    175.633, 175.479, 175.3307, 175.1878,
  343.7783, 343.6074, 343.43, 343.2459, 343.0545, 342.8554, 342.6479, 
    342.4316, 342.2058, 341.9696, 341.7225, 341.4633, 341.1913, 340.9054, 
    340.6042, 340.2867, 339.9511, 339.5959, 339.2192, 338.819, 338.3927, 
    337.9377, 337.4508, 336.9286, 336.3669, 335.761, 335.1053, 334.3936, 
    333.618, 332.7698, 331.8384, 330.8111, 329.6726, 328.4045, 326.9844, 
    325.3846, 323.5713, 321.5023, 319.1253, 316.3754, 313.1725, 309.4189, 
    305, 299.7885, 293.661, 286.5311, 278.4048, 269.4445, 260, 250.5555, 
    241.5952, 233.4689, 226.339, 220.2115, 215, 210.5811, 206.8275, 203.6246, 
    200.8747, 198.4977, 196.4287, 194.6154, 193.0156, 191.5955, 190.3274, 
    189.1889, 188.1616, 187.2302, 186.382, 185.6065, 184.8946, 184.239, 
    183.6331, 183.0714, 182.5491, 182.0623, 181.6073, 181.181, 180.7808, 
    180.4041, 180.0489, 179.7133, 179.3957, 179.0946, 178.8087, 178.5367, 
    178.2775, 178.0303, 177.7942, 177.5684, 177.352, 177.1446, 176.9455, 
    176.7541, 176.57, 176.3926, 176.2217,
  342.7465, 342.5478, 342.3417, 342.1278, 341.9055, 341.6743, 341.4335, 
    341.1825, 340.9205, 340.6467, 340.3602, 340.06, 339.745, 339.4141, 
    339.0658, 338.6986, 338.311, 337.901, 337.4666, 337.0053, 336.5146, 
    335.9914, 335.4323, 334.8333, 334.1899, 333.4971, 332.7488, 331.9381, 
    331.057, 330.0959, 329.0438, 327.8874, 326.6112, 325.1965, 323.6209, 
    321.8576, 319.8742, 317.6318, 315.0836, 312.174, 308.8375, 305, 300.5811, 
    295.502, 289.7002, 283.153, 275.908, 268.109, 260, 251.891, 244.092, 
    236.847, 230.2999, 224.4981, 219.4189, 215, 211.1625, 207.826, 204.9164, 
    202.3682, 200.1258, 198.1424, 196.3791, 194.8035, 193.3888, 192.1126, 
    190.9562, 189.9041, 188.943, 188.0619, 187.2512, 186.5029, 185.8101, 
    185.1668, 184.5678, 184.0086, 183.4854, 182.9947, 182.5334, 182.099, 
    181.689, 181.3014, 180.9342, 180.5859, 180.255, 179.94, 179.6398, 
    179.3533, 179.0795, 178.8175, 178.5665, 178.3257, 178.0945, 177.8722, 
    177.6583, 177.4522, 177.2535,
  341.717, 341.4908, 341.2564, 341.0131, 340.7603, 340.4975, 340.2239, 
    339.9388, 339.6414, 339.3306, 339.0057, 338.6653, 338.3085, 337.9337, 
    337.5396, 337.1244, 336.6864, 336.2235, 335.7335, 335.2137, 334.6614, 
    334.0732, 333.4454, 332.7739, 332.0539, 331.2799, 330.4457, 329.544, 
    328.5665, 327.5035, 326.3436, 325.0737, 323.6783, 322.1393, 320.4351, 
    318.5408, 316.4267, 314.0583, 311.3957, 308.3931, 305, 301.1625, 
    296.8275, 291.9502, 286.5046, 280.4992, 273.9919, 267.1006, 260, 
    252.8994, 246.0081, 239.5008, 233.4954, 228.0498, 223.1725, 218.8375, 
    215, 211.6069, 208.6043, 205.9417, 203.5733, 201.4592, 199.5649, 
    197.8607, 196.3217, 194.9263, 193.6564, 192.4965, 191.4335, 190.456, 
    189.5543, 188.7201, 187.9461, 187.2261, 186.5546, 185.9268, 185.3386, 
    184.7863, 184.2665, 183.7765, 183.3136, 182.8756, 182.4604, 182.0663, 
    181.6915, 181.3346, 180.9943, 180.6694, 180.3586, 180.0612, 179.7761, 
    179.5025, 179.2397, 178.9869, 178.7436, 178.5091, 178.283,
  340.6902, 340.437, 340.1745, 339.9023, 339.6196, 339.3257, 339.0199, 
    338.7014, 338.3693, 338.0225, 337.66, 337.2806, 336.883, 336.4657, 
    336.0272, 335.5656, 335.0791, 334.5654, 334.0222, 333.4466, 332.8357, 
    332.1859, 331.4936, 330.7541, 329.9627, 329.1137, 328.2007, 327.2162, 
    326.1519, 324.9981, 323.7437, 322.3758, 320.8795, 319.2377, 317.4306, 
    315.4353, 313.2258, 310.7726, 308.0427, 305, 301.6069, 297.826, 293.6246, 
    288.9797, 283.8865, 278.367, 272.4775, 266.3126, 260, 253.6874, 247.5225, 
    241.633, 236.1134, 231.0203, 226.3754, 222.174, 218.3931, 215, 211.9573, 
    209.2274, 206.7742, 204.5647, 202.5694, 200.7623, 199.1205, 197.6242, 
    196.2563, 195.0019, 193.8481, 192.7838, 191.7994, 190.8863, 190.0373, 
    189.2459, 188.5065, 187.8141, 187.1643, 186.5534, 185.9778, 185.4346, 
    184.9209, 184.4344, 183.9728, 183.5343, 183.1171, 182.7194, 182.34, 
    181.9775, 181.6307, 181.2986, 180.9801, 180.6743, 180.3804, 180.0977, 
    179.8255, 179.563, 179.3098,
  339.6663, 339.3865, 339.0965, 338.7958, 338.4837, 338.1594, 337.8221, 
    337.471, 337.1049, 336.723, 336.324, 335.9067, 335.4696, 335.0113, 
    334.5299, 334.0238, 333.4908, 332.9286, 332.3347, 331.7061, 331.0399, 
    330.3324, 329.5796, 328.7771, 327.9198, 327.0021, 326.0174, 324.9586, 
    323.8172, 322.5839, 321.2479, 319.7971, 318.2174, 316.4931, 314.6064, 
    312.5372, 310.263, 307.7594, 305, 301.9573, 298.6043, 294.9164, 290.8747, 
    286.4705, 281.7102, 276.6204, 271.2519, 265.6798, 260, 254.3202, 
    248.7481, 243.3796, 238.2898, 233.5295, 229.1253, 225.0836, 221.3957, 
    218.0427, 215, 212.2406, 209.737, 207.4628, 205.3936, 203.5069, 201.7826, 
    200.2029, 198.7521, 197.4161, 196.1828, 195.0414, 193.9826, 192.9979, 
    192.0802, 191.2229, 190.4204, 189.6676, 188.9601, 188.2939, 187.6653, 
    187.0714, 186.5092, 185.9762, 185.4701, 184.9888, 184.5304, 184.0933, 
    183.676, 183.277, 182.8951, 182.529, 182.1779, 181.8406, 181.5163, 
    181.2042, 180.9035, 180.6135, 180.3337,
  338.6458, 338.3397, 338.0227, 337.6942, 337.3532, 336.9992, 336.6311, 
    336.2481, 335.8492, 335.4331, 334.9987, 334.5446, 334.0695, 333.5716, 
    333.0492, 332.5004, 331.923, 331.3147, 330.6728, 329.9944, 329.2762, 
    328.5148, 327.706, 326.8453, 325.9278, 324.9478, 323.8989, 322.774, 
    321.5651, 320.2632, 318.8582, 317.3387, 315.692, 313.9038, 311.9585, 
    309.8388, 307.5259, 305, 302.2406, 299.2274, 295.9417, 292.3682, 
    288.4977, 284.33, 279.8769, 275.1656, 270.2401, 265.1604, 260, 254.8396, 
    249.7599, 244.8344, 240.1231, 235.67, 231.5023, 227.6318, 224.0583, 
    220.7726, 217.7594, 215, 212.4741, 210.1612, 208.0415, 206.0961, 204.308, 
    202.6613, 201.1418, 199.7368, 198.4349, 197.226, 196.1011, 195.0522, 
    194.0722, 193.1546, 192.294, 191.4852, 190.7238, 190.0056, 189.3272, 
    188.6853, 188.077, 187.4996, 186.9508, 186.4284, 185.9305, 185.4553, 
    185.0013, 184.5669, 184.1508, 183.7519, 183.3689, 183.0008, 182.6468, 
    182.3059, 181.9773, 181.6603, 181.3542,
  337.6287, 337.297, 336.9535, 336.5977, 336.2286, 335.8456, 335.4475, 
    335.0336, 334.6026, 334.1535, 333.6849, 333.1954, 332.6837, 332.1478, 
    331.5862, 330.9967, 330.3772, 329.7252, 329.0381, 328.313, 327.5465, 
    326.7351, 325.8747, 324.961, 323.9889, 322.953, 321.847, 320.6643, 
    319.3972, 318.0373, 316.575, 315.0002, 313.3014, 311.466, 309.4804, 
    307.3302, 305, 302.4741, 299.737, 296.7742, 293.5733, 290.1258, 286.4287, 
    282.4866, 278.314, 273.9362, 269.3909, 264.7264, 260, 255.2736, 250.6091, 
    246.0638, 241.686, 237.5134, 233.5713, 229.8742, 226.4267, 223.2258, 
    220.263, 217.5259, 215, 212.6698, 210.5196, 208.534, 206.6986, 204.9998, 
    203.4249, 201.9628, 200.6028, 199.3357, 198.153, 197.047, 196.0111, 
    195.039, 194.1253, 193.2649, 192.4535, 191.687, 190.9619, 190.2748, 
    189.6228, 189.0033, 188.4138, 187.8522, 187.3164, 186.8046, 186.3151, 
    185.8465, 185.3974, 184.9664, 184.5525, 184.1545, 183.7714, 183.4023, 
    183.0465, 182.703, 182.3713,
  336.6156, 336.2586, 335.8893, 335.5068, 335.1103, 334.6989, 334.2718, 
    333.8279, 333.3659, 332.8849, 332.3833, 331.8599, 331.313, 330.7409, 
    330.1419, 329.5139, 328.8545, 328.1615, 327.4321, 326.6635, 325.8522, 
    324.9948, 324.0874, 323.1256, 322.1046, 321.019, 319.8632, 318.6306, 
    317.3141, 315.9059, 314.3975, 312.7795, 311.042, 309.174, 307.164, 305, 
    302.6698, 300.1612, 297.4628, 294.5647, 291.4592, 288.1424, 284.6154, 
    280.8853, 276.9672, 272.8842, 268.6681, 264.3583, 260, 255.6417, 
    251.3319, 247.1158, 243.0328, 239.1147, 235.3846, 231.8576, 228.5408, 
    225.4353, 222.5372, 219.8388, 217.3302, 215, 212.836, 210.826, 208.958, 
    207.2204, 205.6025, 204.0941, 202.6859, 201.3694, 200.1368, 198.9809, 
    197.8954, 196.8744, 195.9126, 195.0052, 194.1478, 193.3365, 192.5679, 
    191.8385, 191.1455, 190.4861, 189.8581, 189.259, 188.687, 188.1401, 
    187.6167, 187.1152, 186.6341, 186.1722, 185.7282, 185.301, 184.8897, 
    184.4932, 184.1107, 183.7414, 183.3844,
  335.6065, 335.225, 334.8304, 334.4219, 333.9987, 333.5599, 333.1046, 
    332.6315, 332.1397, 331.6279, 331.0947, 330.5388, 329.9584, 329.3519, 
    328.7174, 328.0529, 327.3562, 326.6248, 325.856, 325.047, 324.1946, 
    323.2953, 322.3453, 321.3403, 320.2759, 319.1469, 317.9479, 316.6729, 
    315.3153, 313.8681, 312.3236, 310.6735, 308.9091, 307.0211, 305, 302.836, 
    300.5196, 298.0415, 295.3936, 292.5694, 289.5649, 286.3791, 283.0156, 
    279.4829, 275.7955, 271.9741, 268.0455, 264.042, 260, 255.958, 251.9545, 
    248.0259, 244.2045, 240.5171, 236.9844, 233.6209, 230.4351, 227.4306, 
    224.6064, 221.9585, 219.4804, 217.164, 215, 212.9789, 211.0909, 209.3265, 
    207.6764, 206.1319, 204.6846, 203.3271, 202.0521, 200.8531, 199.7241, 
    198.6597, 197.6547, 196.7047, 195.8054, 194.953, 194.144, 193.3752, 
    192.6438, 191.9471, 191.2826, 190.6481, 190.0416, 189.4613, 188.9053, 
    188.3721, 187.8603, 187.3685, 186.8955, 186.4401, 186.0013, 185.5781, 
    185.1696, 184.775, 184.3935,
  334.6019, 334.1963, 333.7771, 333.3433, 332.8942, 332.4289, 331.9462, 
    331.4452, 330.9246, 330.3833, 329.8199, 329.2328, 328.6205, 327.9814, 
    327.3135, 326.6147, 325.883, 325.1159, 324.3107, 323.4647, 322.5747, 
    321.6375, 320.6492, 319.606, 318.5034, 317.3369, 316.1012, 314.7909, 
    313.4, 311.9221, 310.3505, 308.678, 306.8971, 305, 302.9789, 300.826, 
    298.534, 296.0962, 293.5069, 290.7623, 287.8607, 284.8035, 281.5955, 
    278.2455, 274.7673, 271.179, 267.5034, 263.7673, 260, 256.2327, 252.4965, 
    248.821, 245.2327, 241.7544, 238.4045, 235.1965, 232.1393, 229.2377, 
    226.4931, 223.9039, 221.466, 219.174, 217.0211, 215, 213.1029, 211.322, 
    209.6495, 208.0779, 206.6, 205.2091, 203.8988, 202.6631, 201.4966, 
    200.394, 199.3508, 198.3625, 197.4253, 196.5353, 195.6893, 194.8841, 
    194.117, 193.3852, 192.6865, 192.0186, 191.3795, 190.7672, 190.1802, 
    189.6167, 189.0754, 188.5548, 188.0538, 187.5711, 187.1058, 186.6567, 
    186.2229, 185.8037, 185.3981,
  333.6019, 333.1729, 332.7297, 332.2715, 331.7973, 331.3062, 330.7972, 
    330.2693, 329.7211, 329.1516, 328.5592, 327.9427, 327.3002, 326.6303, 
    325.9309, 325.2002, 324.4359, 323.6357, 322.7971, 321.9172, 320.9933, 
    320.0219, 318.9997, 317.9228, 316.7873, 315.5887, 314.3224, 312.9834, 
    311.5663, 310.0654, 308.4749, 306.7885, 305, 303.1029, 301.0909, 298.958, 
    296.6986, 294.308, 291.7826, 289.1205, 286.3217, 283.3888, 280.3274, 
    277.1464, 273.8581, 270.4786, 267.0273, 263.5263, 260, 256.4737, 
    252.9727, 249.5214, 246.1419, 242.8536, 239.6726, 236.6112, 233.6783, 
    230.8795, 228.2174, 225.692, 223.3014, 221.042, 218.9091, 216.8971, 215, 
    213.2115, 211.5251, 209.9346, 208.4338, 207.0166, 205.6776, 204.4113, 
    203.2127, 202.0772, 201.0004, 199.9781, 199.0068, 198.0828, 197.2029, 
    196.3643, 195.5641, 194.7998, 194.0691, 193.3697, 192.6998, 192.0573, 
    191.4408, 190.8484, 190.2789, 189.7307, 189.2028, 188.6938, 188.2027, 
    187.7285, 187.2702, 186.8271, 186.3981,
  332.6068, 332.1551, 331.6887, 331.2067, 330.7082, 330.1924, 329.6581, 
    329.1042, 328.5297, 327.9333, 327.3135, 326.6689, 325.998, 325.2991, 
    324.5704, 323.8098, 323.0154, 322.1848, 321.3156, 320.4052, 319.4506, 
    318.4489, 317.3969, 316.2909, 315.1272, 313.9019, 312.6106, 311.2489, 
    309.812, 308.295, 306.6927, 305, 303.2115, 301.322, 299.3265, 297.2205, 
    294.9998, 292.6613, 290.2029, 287.6242, 284.9263, 282.1126, 279.1889, 
    276.1638, 273.0484, 269.8569, 266.6056, 263.3133, 260, 256.6867, 
    253.3944, 250.1431, 246.9516, 243.8362, 240.8111, 237.8874, 235.0737, 
    232.3758, 229.7971, 227.3387, 225.0002, 222.7796, 220.6735, 218.678, 
    216.7885, 215, 213.3073, 211.705, 210.188, 208.7511, 207.3894, 206.0981, 
    204.8728, 203.7091, 202.6031, 201.551, 200.5494, 199.5948, 198.6844, 
    197.8152, 196.9846, 196.1901, 195.4296, 194.7009, 194.002, 193.3311, 
    192.6865, 192.0667, 191.4703, 190.8958, 190.3419, 189.8076, 189.2918, 
    188.7933, 188.3113, 187.8449, 187.3932,
  331.6168, 331.1431, 330.6542, 330.1492, 329.6274, 329.0877, 328.5291, 
    327.9506, 327.3509, 326.7288, 326.083, 325.4121, 324.7144, 323.9885, 
    323.2324, 322.4443, 321.6222, 320.7638, 319.8669, 318.9289, 317.9471, 
    316.9188, 315.8408, 314.7099, 313.5227, 312.2755, 310.9644, 309.5856, 
    308.1348, 306.6077, 305, 303.3073, 301.5251, 299.6495, 297.6764, 
    295.6025, 293.425, 291.1418, 288.7521, 286.2563, 283.6564, 280.9562, 
    278.1616, 275.2804, 272.3229, 269.3012, 266.2295, 263.1234, 260, 
    256.8766, 253.7705, 250.6988, 247.6771, 244.7196, 241.8384, 239.0438, 
    236.3436, 233.7437, 231.2479, 228.8582, 226.5751, 224.3975, 222.3236, 
    220.3505, 218.4749, 216.6927, 215, 213.3923, 211.8652, 210.4144, 
    209.0356, 207.7245, 206.4773, 205.2901, 204.1592, 203.0812, 202.0529, 
    201.0711, 200.1331, 199.2362, 198.3779, 197.5557, 196.7676, 196.0115, 
    195.2856, 194.5879, 193.917, 193.2712, 192.6491, 192.0494, 191.4709, 
    190.9123, 190.3726, 189.8508, 189.3458, 188.8569, 188.3832,
  330.6322, 330.1371, 329.6265, 329.0994, 328.5551, 327.9925, 327.4107, 
    326.8086, 326.185, 325.5387, 324.8683, 324.1726, 323.45, 322.6988, 
    321.9174, 321.1039, 320.2564, 319.3729, 318.451, 317.4885, 316.4828, 
    315.4313, 314.3311, 313.1793, 311.9728, 310.7083, 309.3823, 307.9913, 
    306.5318, 305, 303.3923, 301.705, 299.9346, 298.0779, 296.1319, 294.0941, 
    291.9627, 289.7368, 287.4161, 285.0019, 282.4965, 279.9041, 277.2302, 
    274.4821, 271.669, 268.8015, 265.8918, 262.9532, 260, 257.0468, 254.1082, 
    251.1985, 248.331, 245.5179, 242.7698, 240.0959, 237.5035, 234.9981, 
    232.5839, 230.2632, 228.0372, 225.9059, 223.8681, 221.9221, 220.0654, 
    218.295, 216.6077, 215, 213.4682, 212.0087, 210.6177, 209.2917, 208.0272, 
    206.8207, 205.6689, 204.5687, 203.5172, 202.5115, 201.549, 200.6271, 
    199.7436, 198.8961, 198.0826, 197.3012, 196.55, 195.8274, 195.1316, 
    194.4613, 193.815, 193.1914, 192.5893, 192.0075, 191.4449, 190.9006, 
    190.3736, 189.8629, 189.3678,
  329.6532, 329.1375, 328.6058, 328.0575, 327.4916, 326.9072, 326.3032, 
    325.6786, 325.0324, 324.3632, 323.6698, 322.9509, 322.2049, 321.4304, 
    320.6257, 319.789, 318.9185, 318.0123, 317.0682, 316.084, 315.0575, 
    313.9861, 312.8673, 311.6984, 310.4765, 309.1988, 307.8622, 306.4636, 
    305, 303.4682, 301.8652, 300.188, 298.4337, 296.6, 294.6847, 292.6859, 
    290.6028, 288.4349, 286.1828, 283.8481, 281.4335, 278.943, 276.382, 
    273.7571, 271.0766, 268.3497, 265.5869, 262.7996, 260, 257.2004, 
    254.4131, 251.6503, 248.9234, 246.2428, 243.618, 241.057, 238.5665, 
    236.1519, 233.8172, 231.5651, 229.3972, 227.3141, 225.3154, 223.4, 
    221.5662, 219.812, 218.1348, 216.5318, 215, 213.5364, 212.1378, 210.8012, 
    209.5235, 208.3016, 207.1327, 206.0139, 204.9425, 203.9159, 202.9318, 
    201.9877, 201.0815, 200.211, 199.3743, 198.5696, 197.7951, 197.0491, 
    196.3302, 195.6368, 194.9676, 194.3213, 193.6968, 193.0928, 192.5084, 
    191.9425, 191.3942, 190.8626, 190.3468,
  328.6799, 328.1443, 327.5925, 327.0238, 326.4372, 325.8319, 325.2069, 
    324.5611, 323.8935, 323.2028, 322.4878, 321.7472, 320.9796, 320.1836, 
    319.3576, 318.4998, 317.6086, 316.6821, 315.7184, 314.7154, 313.671, 
    312.5829, 311.4487, 310.2661, 309.0325, 307.7454, 306.4021, 305, 
    303.5364, 302.0087, 300.4144, 298.7511, 297.0166, 295.2091, 293.3271, 
    291.3694, 289.3357, 287.226, 285.0414, 282.7838, 280.456, 278.0619, 
    275.6064, 273.0959, 270.5374, 267.9391, 265.3101, 262.6603, 260, 
    257.3397, 254.6899, 252.0609, 249.4627, 246.9041, 244.3935, 241.9381, 
    239.544, 237.2162, 234.9586, 232.774, 230.6643, 228.6306, 226.6729, 
    224.7909, 222.9834, 221.2489, 219.5856, 217.9913, 216.4636, 215, 
    213.5979, 212.2546, 210.9675, 209.7339, 208.5513, 207.4171, 206.329, 
    205.2846, 204.2816, 203.3179, 202.3914, 201.5002, 200.6424, 199.8164, 
    199.0203, 198.2528, 197.5122, 196.7972, 196.1066, 195.4389, 194.7931, 
    194.1681, 193.5628, 192.9762, 192.4075, 191.8557, 191.3201,
  327.7126, 327.1578, 326.5867, 325.9984, 325.3922, 324.767, 324.122, 
    323.4562, 322.7684, 322.0576, 321.3224, 320.5619, 319.7744, 318.9586, 
    318.1132, 317.2364, 316.3267, 315.3823, 314.4015, 313.3823, 312.3227, 
    311.2208, 310.0744, 308.8814, 307.6395, 306.3465, 305, 303.5979, 
    302.1378, 300.6177, 299.0356, 297.3894, 295.6776, 293.8988, 292.0521, 
    290.1368, 288.153, 286.1011, 283.9826, 281.7993, 279.5543, 277.2512, 
    274.8947, 272.4902, 270.0443, 267.5642, 265.0577, 262.5334, 260, 
    257.4666, 254.9423, 252.4358, 249.9557, 247.5098, 245.1054, 242.7488, 
    240.4457, 238.2006, 236.0174, 233.8989, 231.847, 229.8632, 227.9479, 
    226.1012, 224.3224, 222.6106, 220.9644, 219.3823, 217.8622, 216.4021, 
    215, 213.6535, 212.3605, 211.1186, 209.9256, 208.7792, 207.6773, 
    206.6177, 205.5985, 204.6177, 203.6733, 202.7636, 201.8868, 201.0414, 
    200.2256, 199.4382, 198.6775, 197.9424, 197.2316, 196.5438, 195.878, 
    195.233, 194.6078, 194.0016, 193.4133, 192.8422, 192.2874,
  326.7514, 326.1783, 325.5886, 324.9817, 324.3567, 323.7127, 323.0489, 
    322.3641, 321.6575, 320.9279, 320.1741, 319.395, 318.5893, 317.7556, 
    316.8926, 315.9988, 315.0728, 314.1127, 313.1171, 312.0842, 311.0122, 
    309.8993, 308.7435, 307.543, 306.2958, 305, 303.6535, 302.2546, 300.8012, 
    299.2917, 297.7245, 296.0981, 294.4113, 292.6631, 290.8531, 288.981, 
    287.047, 285.0522, 282.9979, 280.8863, 278.7201, 276.5029, 274.239, 
    271.9334, 269.5918, 267.2206, 264.8266, 262.4172, 260, 257.5828, 
    255.1734, 252.7795, 250.4082, 248.0666, 245.761, 243.4971, 241.2799, 
    239.1137, 237.0021, 234.9478, 232.953, 231.0191, 229.1469, 227.3369, 
    225.5887, 223.9019, 222.2755, 220.7083, 219.1988, 217.7454, 216.3465, 
    215, 213.7041, 212.457, 211.2565, 210.1007, 208.9878, 207.9158, 206.8829, 
    205.8873, 204.9273, 204.0012, 203.1074, 202.2444, 201.4107, 200.605, 
    199.8259, 199.0721, 198.3425, 197.6359, 196.9511, 196.2873, 195.6433, 
    195.0183, 194.4114, 193.8217, 193.2486,
  325.7966, 325.2058, 324.5984, 323.9738, 323.331, 322.6693, 321.9876, 
    321.2852, 320.5609, 319.8138, 319.0428, 318.2468, 317.4244, 316.5746, 
    315.6959, 314.787, 313.8466, 312.8731, 311.865, 310.8208, 309.7388, 
    308.6174, 307.4549, 306.2497, 305, 303.7042, 302.3605, 300.9675, 
    299.5235, 298.0272, 296.4773, 294.8728, 293.2127, 291.4966, 289.7241, 
    287.8954, 286.0111, 284.0722, 282.0802, 280.0373, 277.9461, 275.8101, 
    273.6331, 271.4196, 269.1748, 266.9043, 264.614, 262.3104, 260, 257.6896, 
    255.386, 253.0957, 250.8252, 248.5804, 246.3669, 244.1899, 242.0539, 
    239.9627, 237.9198, 235.9278, 233.9889, 232.1046, 230.2759, 228.5034, 
    226.7873, 225.1272, 223.5227, 221.9728, 220.4765, 219.0325, 217.6395, 
    216.2959, 215, 213.7503, 212.5451, 211.3826, 210.2612, 209.1792, 208.135, 
    207.1269, 206.1534, 205.213, 204.3041, 203.4254, 202.5756, 201.7532, 
    200.9572, 200.1862, 199.4391, 198.7148, 198.0124, 197.3308, 196.669, 
    196.0262, 195.4016, 194.7942, 194.2034,
  324.8481, 324.2405, 323.6163, 322.9748, 322.3152, 321.6367, 320.9384, 
    320.2195, 319.4789, 318.7157, 317.9288, 317.1173, 316.2799, 315.4155, 
    314.5229, 313.6009, 312.648, 311.6631, 310.6447, 309.5914, 308.5017, 
    307.3742, 306.2075, 305, 303.7503, 302.457, 301.1186, 299.7339, 298.3016, 
    296.8207, 295.2901, 293.7091, 292.0772, 290.394, 288.6597, 286.8744, 
    285.039, 283.1547, 281.2229, 279.2459, 277.2261, 275.1667, 273.0714, 
    270.944, 268.7893, 266.6121, 264.4178, 262.2118, 260, 257.7882, 255.5822, 
    253.3879, 251.2107, 249.056, 246.9286, 244.8332, 242.7739, 240.7541, 
    238.7771, 236.8454, 234.961, 233.1256, 231.3403, 229.606, 227.9228, 
    226.2909, 224.7099, 223.1793, 221.6984, 220.2661, 218.8814, 217.543, 
    216.2497, 215, 213.7925, 212.6258, 211.4983, 210.4086, 209.3553, 
    208.3369, 207.3519, 206.3991, 205.4771, 204.5845, 203.7201, 202.8827, 
    202.0712, 201.2843, 200.5211, 199.7805, 199.0616, 198.3633, 197.6848, 
    197.0252, 196.3837, 195.7595, 195.1518,
  323.9063, 323.2827, 322.6425, 321.985, 321.3096, 320.6153, 319.9015, 
    319.1671, 318.4114, 317.6334, 316.8321, 316.0066, 315.1557, 314.2784, 
    313.3736, 312.4402, 311.4768, 310.4824, 309.4557, 308.3953, 307.3001, 
    306.1688, 305, 303.7925, 302.5451, 301.2565, 299.9256, 298.5513, 
    297.1327, 295.6689, 294.1592, 292.6031, 291.0003, 289.3508, 287.6547, 
    285.9126, 284.1253, 282.294, 280.4204, 278.5064, 276.5546, 274.5677, 
    272.5492, 270.5025, 268.4318, 266.3414, 264.2361, 262.1206, 260, 
    257.8794, 255.7639, 253.6586, 251.5682, 249.4975, 247.4509, 245.4322, 
    243.4454, 241.4935, 239.5796, 237.706, 235.8747, 234.0874, 232.3453, 
    230.6492, 228.9996, 227.3969, 225.8408, 224.3311, 222.8673, 221.4487, 
    220.0744, 218.7435, 217.4549, 216.2075, 215, 213.8312, 212.6999, 
    211.6047, 210.5443, 209.5176, 208.5232, 207.5598, 206.6264, 205.7216, 
    204.8443, 203.9934, 203.1679, 202.3666, 201.5886, 200.8329, 200.0985, 
    199.3847, 198.6904, 198.015, 197.3575, 196.7173, 196.0937,
  322.9712, 322.3323, 321.677, 321.0045, 320.3141, 319.6052, 318.8768, 
    318.1283, 317.3586, 316.5671, 315.7527, 314.9146, 314.0518, 313.1631, 
    312.2478, 311.3046, 310.3326, 309.3305, 308.2973, 307.2319, 306.1332, 
    305, 303.8312, 302.6258, 301.3826, 300.1007, 298.7792, 297.4171, 
    296.0139, 294.5687, 293.0812, 291.5511, 289.9781, 288.3625, 286.7047, 
    285.0052, 283.2649, 281.4852, 279.6676, 277.8141, 275.9268, 274.0086, 
    272.0623, 270.0913, 268.0992, 266.0898, 264.0672, 262.0359, 260, 
    257.9641, 255.9328, 253.9102, 251.9008, 249.9087, 247.9377, 245.9914, 
    244.0732, 242.1859, 240.3324, 238.5148, 236.7351, 234.9948, 233.2953, 
    231.6375, 230.0219, 228.449, 226.9188, 225.4313, 223.9861, 222.5829, 
    221.2208, 219.8993, 218.6174, 217.3742, 216.1688, 215, 213.8668, 
    212.7681, 211.7027, 210.6695, 209.6675, 208.6954, 207.7522, 206.8369, 
    205.9482, 205.0854, 204.2473, 203.4329, 202.6413, 201.8717, 201.1232, 
    200.3948, 199.6858, 198.9955, 198.323, 197.6677, 197.0288,
  322.043, 321.3896, 320.72, 320.0334, 319.3291, 318.6064, 317.8647, 317.103, 
    316.3206, 315.5168, 314.6907, 313.8414, 312.968, 312.0695, 311.1452, 
    310.1939, 309.2148, 308.2068, 307.169, 306.1004, 305, 303.8668, 302.6999, 
    301.4983, 300.2612, 298.9878, 297.6773, 296.329, 294.9425, 293.5172, 
    292.0529, 290.5494, 289.0067, 287.4253, 285.8054, 284.1478, 282.4535, 
    280.7238, 278.9601, 277.1643, 275.3386, 273.4854, 271.6073, 269.7074, 
    267.7889, 265.8552, 263.9099, 261.9569, 260, 258.0431, 256.0901, 
    254.1448, 252.2111, 250.2926, 248.3927, 246.5146, 244.6614, 242.8357, 
    241.0399, 239.2762, 237.5465, 235.8522, 234.1946, 232.5747, 230.9932, 
    229.4506, 227.9471, 226.4828, 225.0575, 223.671, 222.3227, 221.0122, 
    219.7388, 218.5017, 217.3001, 216.1332, 215, 213.8996, 212.8309, 
    211.7932, 210.7852, 209.8061, 208.8548, 207.9305, 207.032, 206.1586, 
    205.3093, 204.4831, 203.6793, 202.897, 202.1354, 201.3936, 200.6709, 
    199.9666, 199.28, 198.6104, 197.957,
  321.1216, 320.4547, 319.7716, 319.0717, 318.3545, 317.6191, 316.865, 
    316.0913, 315.2975, 314.4826, 313.646, 312.7868, 311.9042, 310.9974, 
    310.0656, 309.1078, 308.1232, 307.111, 306.0702, 305, 303.8996, 302.7681, 
    301.6047, 300.4086, 299.1792, 297.9158, 296.6177, 295.2846, 293.916, 
    292.5115, 291.0711, 289.5948, 288.0828, 286.5353, 284.953, 283.3365, 
    281.687, 280.0056, 278.2939, 276.5534, 274.7863, 272.9947, 271.181, 
    269.3481, 267.4987, 265.636, 263.763, 261.8832, 260, 258.1168, 256.237, 
    254.3641, 252.5013, 250.6519, 248.819, 247.0053, 245.2137, 243.4466, 
    241.7061, 239.9944, 238.313, 236.6635, 235.047, 233.4647, 231.9172, 
    230.4052, 228.9289, 227.4885, 226.0841, 224.7154, 223.3823, 222.0842, 
    220.8208, 219.5914, 218.3953, 217.2319, 216.1004, 215, 213.9298, 
    212.8891, 211.8768, 210.8922, 209.9344, 209.0026, 208.0958, 207.2132, 
    206.354, 205.5174, 204.7025, 203.9087, 203.135, 202.3809, 201.6455, 
    200.9283, 200.2284, 199.5453, 198.8784,
  320.2073, 319.5276, 318.8319, 318.1197, 317.3904, 316.6433, 315.8778, 
    315.0933, 314.289, 313.4643, 312.6185, 311.7507, 310.8603, 309.9465, 
    309.0086, 308.0457, 307.0572, 306.0422, 305, 303.9298, 302.831, 301.7027, 
    300.5443, 299.3553, 298.135, 296.8829, 295.5985, 294.2816, 292.9318, 
    291.549, 290.1331, 288.6844, 287.2029, 285.6893, 284.144, 282.5679, 
    280.9619, 279.3272, 277.6653, 275.9778, 274.2665, 272.5334, 270.7808, 
    269.011, 267.2267, 265.4305, 263.6254, 261.8142, 260, 258.1858, 256.3746, 
    254.5695, 252.7733, 250.989, 249.2192, 247.4666, 245.7335, 244.0222, 
    242.3347, 240.6728, 239.0381, 237.4321, 235.856, 234.3107, 232.7971, 
    231.3156, 229.8669, 228.451, 227.0682, 225.7184, 224.4015, 223.1171, 
    221.865, 220.6447, 219.4557, 218.2973, 217.1691, 216.0702, 215, 213.9578, 
    212.9428, 211.9543, 210.9914, 210.0535, 209.1397, 208.2493, 207.3815, 
    206.5357, 205.711, 204.9067, 204.1222, 203.3567, 202.6096, 201.8803, 
    201.1681, 200.4724, 199.7926,
  319.3002, 318.6084, 317.9009, 317.1773, 316.4368, 315.679, 314.9033, 
    314.1089, 313.2954, 312.462, 311.6081, 310.733, 309.836, 308.9166, 
    307.9739, 307.0074, 306.0163, 305, 303.9578, 302.889, 301.7932, 300.6695, 
    299.5176, 298.3369, 297.1269, 295.8873, 294.6177, 293.3179, 291.9877, 
    290.6271, 289.2362, 287.8152, 286.3643, 284.8841, 283.3752, 281.8385, 
    280.2748, 278.6853, 277.0714, 275.4346, 273.7765, 272.099, 270.4041, 
    268.694, 266.971, 265.2375, 263.4962, 261.7494, 260, 258.2506, 256.5038, 
    254.7625, 253.029, 251.306, 249.5959, 247.901, 246.2235, 244.5654, 
    242.9286, 241.3147, 239.7252, 238.1615, 236.6248, 235.1159, 233.6357, 
    232.1848, 230.7638, 229.3729, 228.0123, 226.6821, 225.3823, 224.1127, 
    222.8731, 221.6631, 220.4824, 219.3305, 218.2068, 217.1109, 216.0422, 
    215, 213.9837, 212.9926, 212.0261, 211.0834, 210.164, 209.267, 208.392, 
    207.538, 206.7046, 205.8911, 205.0967, 204.321, 203.5632, 202.8227, 
    202.0991, 201.3916, 200.6998,
  318.4002, 317.6972, 316.9788, 316.2445, 315.4939, 314.7263, 313.9413, 
    313.1382, 312.3164, 311.4754, 310.6146, 309.7334, 308.8312, 307.9073, 
    306.9612, 305.9923, 305, 303.9837, 302.9428, 301.8768, 300.7852, 
    299.6674, 298.5232, 297.352, 296.1534, 294.9272, 293.6733, 292.3914, 
    291.0815, 289.7436, 288.3778, 286.9846, 285.5641, 284.117, 282.6438, 
    281.1455, 279.6228, 278.077, 276.5092, 274.9209, 273.3136, 271.689, 
    270.0489, 268.3953, 266.7303, 265.0559, 263.3746, 261.6885, 260, 
    258.3115, 256.6254, 254.9441, 253.2697, 251.6047, 249.9511, 248.311, 
    246.6864, 245.0791, 243.4908, 241.923, 240.3772, 238.8545, 237.3562, 
    235.883, 234.4359, 233.0154, 231.6221, 230.2564, 228.9185, 227.6086, 
    226.3267, 225.0727, 223.8466, 222.6481, 221.4768, 220.3325, 219.2148, 
    218.1232, 217.0572, 216.0163, 215, 214.0077, 213.0388, 212.0927, 
    211.1688, 210.2666, 209.3854, 208.5246, 207.6836, 206.8618, 206.0587, 
    205.2737, 204.5061, 203.7555, 203.0212, 202.3028, 201.5998,
  317.5075, 316.794, 316.0655, 315.3216, 314.5616, 313.7852, 312.9918, 
    312.1809, 311.352, 310.5045, 309.638, 308.7518, 307.8454, 306.9184, 
    305.9701, 305, 304.0077, 302.9926, 301.9543, 300.8922, 299.8061, 
    298.6954, 297.5598, 296.3991, 295.213, 294.0012, 292.7636, 291.5002, 
    290.211, 288.8961, 287.5557, 286.1902, 284.7998, 283.3853, 281.9471, 
    280.4861, 279.0033, 277.4996, 275.9762, 274.4344, 272.8756, 271.3014, 
    269.7133, 268.1133, 266.5031, 264.8846, 263.2599, 261.631, 260, 258.369, 
    256.7401, 255.1154, 253.4969, 251.8867, 250.2867, 248.6986, 247.1244, 
    245.5656, 244.0238, 242.5004, 240.9967, 239.5139, 238.0529, 236.6148, 
    235.2002, 233.8099, 232.4443, 231.1039, 229.789, 228.4998, 227.2364, 
    225.9988, 224.787, 223.6009, 222.4402, 221.3046, 220.1939, 219.1078, 
    218.0457, 217.0074, 215.9923, 215, 214.0299, 213.0816, 212.1546, 
    211.2482, 210.362, 209.4955, 208.648, 207.8191, 207.0082, 206.2148, 
    205.4384, 204.6784, 203.9345, 203.206, 202.4925,
  316.6221, 315.8989, 315.1612, 314.4083, 313.64, 312.8557, 312.0549, 
    311.2372, 310.4022, 309.5493, 308.678, 307.7879, 306.8785, 305.9494, 305, 
    304.0299, 303.0388, 302.0261, 300.9914, 299.9344, 298.8548, 297.7522, 
    296.6264, 295.4771, 294.3041, 293.1074, 291.8868, 290.6424, 289.3743, 
    288.0826, 286.7676, 285.4296, 284.0691, 282.6865, 281.2826, 279.8581, 
    278.4138, 276.9508, 275.4701, 273.9728, 272.4604, 270.9342, 269.3958, 
    267.8465, 266.2883, 264.7227, 263.1516, 261.5767, 260, 258.4233, 
    256.8484, 255.2773, 253.7117, 252.1535, 250.6043, 249.0658, 247.5396, 
    246.0272, 244.5299, 243.0492, 241.5862, 240.1419, 238.7174, 237.3135, 
    235.9309, 234.5704, 233.2324, 231.9174, 230.6257, 229.3576, 228.1132, 
    226.8926, 225.6959, 224.5229, 223.3736, 222.2478, 221.1452, 220.0656, 
    219.0086, 217.9739, 216.9612, 215.9701, 215, 214.0506, 213.1215, 
    212.2121, 211.322, 210.4507, 209.5978, 208.7628, 207.9451, 207.1443, 
    206.36, 205.5917, 204.8389, 204.1011, 203.3779,
  315.744, 315.012, 314.2657, 313.5049, 312.729, 311.9376, 311.1304, 
    310.3069, 309.4667, 308.6094, 307.7344, 306.8415, 305.9301, 305, 
    304.0506, 303.0816, 302.0927, 301.0834, 300.0535, 299.0026, 297.9305, 
    296.8369, 295.7216, 294.5845, 293.4254, 292.2444, 291.0414, 289.8164, 
    288.5696, 287.3012, 286.0115, 284.7009, 283.3697, 282.0186, 280.6481, 
    279.2591, 277.8522, 276.4284, 274.9887, 273.5343, 272.0663, 270.5859, 
    269.0946, 267.5938, 266.0848, 264.5694, 263.049, 261.5253, 260, 258.4747, 
    256.951, 255.4306, 253.9152, 252.4062, 250.9054, 249.4141, 247.9337, 
    246.4657, 245.0112, 243.5716, 242.1478, 240.741, 239.3519, 237.9814, 
    236.6303, 235.2991, 233.9885, 232.6988, 231.4304, 230.1836, 228.9586, 
    227.7556, 226.5746, 225.4155, 224.2784, 223.1631, 222.0695, 220.9974, 
    219.9465, 218.9166, 217.9073, 216.9184, 215.9494, 215, 214.0698, 
    213.1585, 212.2656, 211.3906, 210.5333, 209.6931, 208.8696, 208.0624, 
    207.271, 206.4951, 205.7343, 204.9881, 204.256,
  314.8733, 314.1331, 313.3792, 312.6111, 311.8286, 311.0311, 310.2184, 
    309.39, 308.5455, 307.6847, 306.8071, 305.9123, 305, 304.0699, 303.1215, 
    302.1546, 301.1688, 300.164, 299.1397, 298.0958, 297.032, 295.9482, 
    294.8443, 293.7201, 292.5756, 291.4107, 290.2256, 289.0204, 287.7951, 
    286.55, 285.2856, 284.002, 282.6998, 281.3795, 280.0416, 278.687, 
    277.3163, 275.9305, 274.5304, 273.117, 271.6915, 270.255, 268.8087, 
    267.3538, 265.8918, 264.424, 262.9518, 261.4766, 260, 258.5234, 257.0482, 
    255.576, 254.1082, 252.6462, 251.1913, 249.745, 248.3085, 246.8829, 
    245.4696, 244.0695, 242.6836, 241.313, 239.9584, 238.6205, 237.3002, 
    235.998, 234.7144, 233.45, 232.2049, 230.9797, 229.7744, 228.5893, 
    227.4244, 226.2799, 225.1557, 224.0518, 222.968, 221.9042, 220.8603, 
    219.836, 218.8312, 217.8454, 216.8785, 215.9302, 215, 214.0877, 213.1929, 
    212.3153, 211.4545, 210.61, 209.7817, 208.9689, 208.1714, 207.3889, 
    206.6208, 205.8669, 205.1267,
  314.01, 313.2625, 312.5016, 311.7271, 310.9387, 310.136, 309.3185, 
    308.4861, 307.6384, 306.7751, 305.8957, 305, 304.0877, 303.1585, 
    302.2121, 301.2482, 300.2666, 299.267, 298.2493, 297.2132, 296.1586, 
    295.0854, 293.9934, 292.8827, 291.7532, 290.605, 289.4381, 288.2528, 
    287.0491, 285.8274, 284.5879, 283.3311, 282.0573, 280.7672, 279.4612, 
    278.1401, 276.8046, 275.4554, 274.0933, 272.7194, 271.3347, 269.94, 
    268.5367, 267.1257, 265.7083, 264.2858, 262.8594, 261.4304, 260, 
    258.5696, 257.1406, 255.7142, 254.2917, 252.8743, 251.4633, 250.06, 
    248.6654, 247.2806, 245.9067, 244.5447, 243.1954, 241.8599, 240.5387, 
    239.2328, 237.9427, 236.6689, 235.4121, 234.1726, 232.9509, 231.7472, 
    230.5618, 229.395, 228.2468, 227.1173, 226.0066, 224.9146, 223.8414, 
    222.7868, 221.7507, 220.733, 219.7334, 218.7518, 217.7879, 216.8415, 
    215.9123, 215, 214.1043, 213.225, 212.3616, 211.5139, 210.6815, 209.864, 
    209.0613, 208.2729, 207.4984, 206.7375, 205.99,
  313.1541, 312.3999, 311.633, 310.8529, 310.0594, 309.2522, 308.4309, 
    307.5954, 306.7453, 305.8802, 305, 304.1043, 303.1929, 302.2656, 301.322, 
    300.362, 299.3854, 298.3919, 297.3815, 296.354, 295.3093, 294.2473, 
    293.1679, 292.0712, 290.9572, 289.8259, 288.6776, 287.5122, 286.3302, 
    285.1317, 283.917, 282.6865, 281.4408, 280.1801, 278.9053, 277.6167, 
    276.3151, 275.0013, 273.676, 272.34, 270.9943, 269.6398, 268.2775, 
    266.9085, 265.5337, 264.1543, 262.7715, 261.3863, 260, 258.6137, 
    257.2285, 255.8457, 254.4663, 253.0915, 251.7225, 250.3602, 249.0057, 
    247.66, 246.324, 244.9987, 243.6849, 242.3833, 241.0947, 239.8198, 
    238.5592, 237.3135, 236.083, 234.8684, 233.6698, 232.4878, 231.3225, 
    230.1741, 229.0428, 227.9288, 226.8321, 225.7527, 224.6907, 223.646, 
    222.6185, 221.608, 220.6146, 219.638, 218.678, 217.7344, 216.8071, 
    215.8957, 215, 214.1198, 213.2547, 212.4046, 211.5691, 210.7478, 
    209.9406, 209.1471, 208.3671, 207.6001, 206.8459,
  312.3057, 311.5456, 310.7732, 309.9883, 309.1905, 308.3796, 307.5554, 
    306.7176, 305.8658, 305, 304.1198, 303.2249, 302.3153, 301.3906, 
    300.4507, 299.4955, 298.5246, 297.538, 296.5357, 295.5174, 294.4832, 
    293.4329, 292.3666, 291.2843, 290.1862, 289.0721, 287.9424, 286.7972, 
    285.6368, 284.4613, 283.2712, 282.0667, 280.8484, 279.6167, 278.3721, 
    277.1151, 275.8465, 274.5669, 273.277, 271.9775, 270.6694, 269.3533, 
    268.0304, 266.7013, 265.3672, 264.029, 262.6877, 261.3444, 260, 258.6556, 
    257.3123, 255.971, 254.6328, 253.2987, 251.9697, 250.6467, 249.3306, 
    248.0225, 246.723, 245.4331, 244.1535, 242.8848, 241.6279, 240.3833, 
    239.1516, 237.9333, 236.7288, 235.5387, 234.3632, 233.2028, 232.0576, 
    230.9279, 229.8138, 228.7157, 227.6334, 226.5671, 225.5169, 224.4826, 
    223.4643, 222.462, 221.4754, 220.5045, 219.5493, 218.6094, 217.6847, 
    216.775, 215.8802, 215, 214.1342, 213.2824, 212.4446, 211.6204, 210.8095, 
    210.0117, 209.2268, 208.4544, 207.6944,
  311.4646, 310.6993, 309.9223, 309.1333, 308.332, 307.5183, 306.6918, 
    305.8525, 305, 304.1342, 303.2547, 302.3616, 301.4545, 300.5333, 
    299.5978, 298.648, 297.6836, 296.7046, 295.711, 294.7025, 293.6794, 
    292.6414, 291.5886, 290.5211, 289.4391, 288.3425, 287.2316, 286.1065, 
    284.9676, 283.815, 282.6491, 281.4703, 280.2789, 279.0754, 277.8603, 
    276.6341, 275.3974, 274.1508, 272.8951, 271.6307, 270.3586, 269.0795, 
    267.7942, 266.5035, 265.2083, 263.9095, 262.6078, 261.3044, 260, 
    258.6956, 257.3922, 256.0905, 254.7917, 253.4965, 252.2058, 250.9205, 
    249.6414, 248.3693, 247.1049, 245.8492, 244.6026, 243.3659, 242.1397, 
    240.9246, 239.7211, 238.5297, 237.3509, 236.185, 235.0324, 233.8934, 
    232.7684, 231.6575, 230.5609, 229.4789, 228.4114, 227.3587, 226.3207, 
    225.2975, 224.289, 223.2954, 222.3164, 221.352, 220.4022, 219.4667, 
    218.5455, 217.6384, 216.7453, 215.8658, 215, 214.1475, 213.3082, 
    212.4817, 211.668, 210.8667, 210.0777, 209.3007, 208.5354,
  310.6309, 309.8612, 309.0802, 308.2878, 307.4838, 306.668, 305.8401, 305, 
    304.1475, 303.2824, 302.4046, 301.5139, 300.61, 299.6931, 298.7628, 
    297.8191, 296.8618, 295.8911, 294.9067, 293.9087, 292.897, 291.8717, 
    290.8329, 289.7805, 288.7148, 287.6359, 286.5438, 285.4389, 284.3214, 
    283.1914, 282.0494, 280.8958, 279.7307, 278.5548, 277.3685, 276.1721, 
    274.9664, 273.7519, 272.529, 271.2986, 270.0612, 268.8175, 267.5684, 
    266.3144, 265.0564, 263.7951, 262.5315, 261.2661, 260, 258.7339, 
    257.4685, 256.2049, 254.9436, 253.6856, 252.4316, 251.1825, 249.9388, 
    248.7014, 247.471, 246.2481, 245.0336, 243.8278, 242.6315, 241.4452, 
    240.2693, 239.1042, 237.9506, 236.8086, 235.6787, 234.5611, 233.4562, 
    232.3641, 231.2852, 230.2195, 229.1671, 228.1283, 227.103, 226.0913, 
    225.0933, 224.1089, 223.1382, 222.1809, 221.2372, 220.3069, 219.39, 
    218.4861, 217.5954, 216.7176, 215.8525, 215, 214.1599, 213.332, 212.5162, 
    211.7122, 210.9198, 210.1388, 209.3691,
  309.8047, 309.0311, 308.2469, 307.4518, 306.6458, 305.8286, 305, 304.1599, 
    303.3082, 302.4446, 301.5691, 300.6815, 299.7816, 298.8696, 297.9451, 
    297.0082, 296.0587, 295.0967, 294.1222, 293.135, 292.1353, 291.1232, 
    290.0985, 289.0616, 288.0124, 286.9511, 285.878, 284.7931, 283.6968, 
    282.5893, 281.4709, 280.3419, 279.2028, 278.0538, 276.8954, 275.7282, 
    274.5525, 273.3689, 272.1779, 270.9801, 269.7761, 268.5665, 267.3521, 
    266.1333, 264.911, 263.6858, 262.4584, 261.2296, 260, 258.7704, 257.5416, 
    256.3142, 255.089, 253.8667, 252.648, 251.4335, 250.2239, 249.0199, 
    247.8221, 246.6311, 245.4475, 244.2718, 243.1045, 241.9462, 240.7972, 
    239.6581, 238.5291, 237.4107, 236.3032, 235.2069, 234.122, 233.0489, 
    231.9876, 230.9384, 229.9015, 228.8768, 227.8646, 226.865, 225.8778, 
    224.9033, 223.9413, 222.9918, 222.0549, 221.1304, 220.2183, 219.3185, 
    218.4309, 217.5554, 216.6918, 215.8401, 215, 214.1714, 213.3542, 
    212.5482, 211.7531, 210.9689, 210.1953,
  308.9857, 308.209, 307.4223, 306.6253, 305.8179, 305, 304.1714, 303.332, 
    302.4817, 301.6204, 300.7478, 299.864, 298.9689, 298.0624, 297.1443, 
    296.2148, 295.2737, 294.321, 293.3567, 292.3809, 291.3936, 290.3948, 
    289.3847, 288.3633, 287.3307, 286.2873, 285.233, 284.1681, 283.0928, 
    282.0075, 280.9123, 279.8076, 278.6938, 277.5711, 276.4401, 275.3011, 
    274.1544, 273.0008, 271.8406, 270.6743, 269.5025, 268.3257, 267.1446, 
    265.9597, 264.7716, 263.581, 262.3884, 261.1945, 260, 258.8055, 257.6116, 
    256.419, 255.2284, 254.0403, 252.8554, 251.6743, 250.4975, 249.3257, 
    248.1594, 246.9992, 245.8455, 244.699, 243.5599, 242.4289, 241.3062, 
    240.1924, 239.0877, 237.9925, 236.9072, 235.8319, 234.767, 233.7127, 
    232.6692, 231.6367, 230.6153, 229.6052, 228.6064, 227.6191, 226.6433, 
    225.679, 224.7263, 223.7852, 222.8557, 221.9376, 221.0311, 220.136, 
    219.2522, 218.3796, 217.5183, 216.668, 215.8286, 215, 214.1821, 213.3747, 
    212.5777, 211.791, 211.0143,
  308.1741, 307.395, 306.6063, 305.808, 305, 304.1821, 303.3542, 302.5162, 
    301.668, 300.8095, 299.9406, 299.0613, 298.1714, 297.271, 296.36, 
    295.4384, 294.5061, 293.5632, 292.6096, 291.6455, 290.6709, 289.6859, 
    288.6904, 287.6848, 286.669, 285.6433, 284.6078, 283.5628, 282.5084, 
    281.4449, 280.3726, 279.2918, 278.2027, 277.1058, 276.0013, 274.8897, 
    273.7714, 272.6468, 271.5163, 270.3804, 269.2397, 268.0945, 266.9455, 
    265.7931, 264.6379, 263.4804, 262.3212, 261.1609, 260, 258.8391, 
    257.6788, 256.5196, 255.3621, 254.2069, 253.0545, 251.9055, 250.7603, 
    249.6196, 248.4837, 247.3532, 246.2286, 245.1103, 243.9987, 242.8942, 
    241.7973, 240.7082, 239.6274, 238.5551, 237.4916, 236.4372, 235.3922, 
    234.3567, 233.331, 232.3152, 231.3096, 230.3142, 229.3291, 228.3545, 
    227.3904, 226.4368, 225.4939, 224.5616, 223.64, 222.729, 221.8286, 
    220.9387, 220.0594, 219.1905, 218.332, 217.4838, 216.6458, 215.8179, 215, 
    214.192, 213.3937, 212.605, 211.8259,
  307.3698, 306.5888, 305.7989, 305, 304.192, 303.3747, 302.5482, 301.7122, 
    300.8667, 300.0117, 299.1471, 298.2729, 297.3889, 296.4951, 295.5917, 
    294.6784, 293.7555, 292.8227, 291.8803, 290.9283, 289.9666, 288.9955, 
    288.015, 287.0252, 286.0262, 285.0183, 284.0016, 282.9762, 281.9425, 
    280.9006, 279.8508, 278.7933, 277.7285, 276.6567, 275.5781, 274.4932, 
    273.4023, 272.3058, 271.2042, 270.0977, 268.9869, 267.8722, 266.7541, 
    265.633, 264.5094, 263.3838, 262.2567, 261.1286, 260, 258.8714, 257.7433, 
    256.6162, 255.4906, 254.367, 253.2459, 252.1278, 251.0131, 249.9023, 
    248.7958, 247.6941, 246.5977, 245.5068, 244.4219, 243.3433, 242.2715, 
    241.2067, 240.1492, 239.0994, 238.0575, 237.0238, 235.9984, 234.9817, 
    233.9738, 232.9748, 231.985, 231.0045, 230.0334, 229.0717, 228.1197, 
    227.1773, 226.2445, 225.3216, 224.4083, 223.5049, 222.6111, 221.7271, 
    220.8529, 219.9883, 219.1333, 218.2878, 217.4518, 216.6253, 215.808, 215, 
    214.2011, 213.4112, 212.6302,
  306.5727, 305.7905, 305, 304.2011, 303.3937, 302.5777, 301.7531, 300.9198, 
    300.0777, 299.2268, 298.367, 297.4984, 296.6208, 295.7343, 294.8388, 
    293.9345, 293.0212, 292.0991, 291.1681, 290.2284, 289.28, 288.323, 
    287.3575, 286.3837, 285.4016, 284.4114, 283.4133, 282.4075, 281.3942, 
    280.3735, 279.3458, 278.3113, 277.2703, 276.2229, 275.1696, 274.1107, 
    273.0465, 271.9773, 270.9035, 269.8255, 268.7436, 267.6583, 266.57, 
    265.479, 264.3859, 263.291, 262.1947, 261.0976, 260, 258.9024, 257.8053, 
    256.709, 255.6141, 254.521, 253.43, 252.3417, 251.2564, 250.1745, 
    249.0965, 248.0227, 246.9535, 245.8893, 244.8304, 243.7771, 242.7298, 
    241.6887, 240.6542, 239.6264, 238.6058, 237.5925, 236.5867, 235.5886, 
    234.5984, 233.6163, 232.6425, 231.677, 230.72, 229.7716, 228.8319, 
    227.9009, 226.9788, 226.0655, 225.1611, 224.2657, 223.3792, 222.5016, 
    221.6329, 220.7732, 219.9223, 219.0802, 218.2469, 217.4223, 216.6063, 
    215.7989, 215, 214.2095, 213.4273,
  305.7828, 305, 304.2095, 303.4112, 302.605, 301.791, 300.9689, 300.1388, 
    299.3007, 298.4544, 297.6001, 296.7375, 295.8669, 294.988, 294.1011, 
    293.206, 292.3028, 291.3916, 290.4724, 289.5453, 288.6104, 287.6677, 
    286.7173, 285.7595, 284.7942, 283.8217, 282.8422, 281.8557, 280.8625, 
    279.8629, 278.8569, 277.8449, 276.8271, 275.8037, 274.775, 273.7414, 
    272.703, 271.6603, 270.6135, 269.563, 268.5092, 267.4522, 266.3926, 
    265.3307, 264.2669, 263.2016, 262.135, 261.0677, 260, 258.9323, 257.865, 
    256.7984, 255.7331, 254.6693, 253.6074, 252.5478, 251.4909, 250.437, 
    249.3865, 248.3397, 247.297, 246.2586, 245.225, 244.1963, 243.1729, 
    242.1551, 241.1431, 240.1371, 239.1374, 238.1443, 237.1578, 236.1783, 
    235.2058, 234.2405, 233.2827, 232.3323, 231.3896, 230.4547, 229.5276, 
    228.6084, 227.6972, 226.794, 225.8989, 225.0119, 224.1331, 223.2625, 
    222.3999, 221.5456, 220.6993, 219.8612, 219.0311, 218.209, 217.395, 
    216.5888, 215.7905, 215, 214.2172,
  305, 304.2172, 303.4273, 302.6302, 301.8259, 301.0143, 300.1953, 299.3691, 
    298.5354, 297.6943, 296.8459, 295.99, 295.1267, 294.256, 293.3779, 
    292.4925, 291.5998, 290.6998, 289.7927, 288.8784, 287.957, 287.0288, 
    286.0937, 285.1519, 284.2034, 283.2486, 282.2874, 281.3201, 280.3468, 
    279.3678, 278.3832, 277.3932, 276.3981, 275.3981, 274.3935, 273.3844, 
    272.3713, 271.3542, 270.3337, 269.3098, 268.283, 267.2535, 266.2217, 
    265.1878, 264.1523, 263.1154, 262.0775, 261.0389, 260, 258.9611, 
    257.9225, 256.8846, 255.8477, 254.8122, 253.7783, 252.7465, 251.717, 
    250.6902, 249.6663, 248.6458, 247.6287, 246.6156, 245.6065, 244.6019, 
    243.6019, 242.6068, 241.6168, 240.6322, 239.6532, 238.6799, 237.7126, 
    236.7514, 235.7966, 234.8482, 233.9063, 232.9712, 232.043, 231.1216, 
    230.2074, 229.3002, 228.4002, 227.5075, 226.6221, 225.744, 224.8733, 
    224.01, 223.1541, 222.3056, 221.4646, 220.6309, 219.8047, 218.9857, 
    218.1741, 217.3698, 216.5727, 215.7828, 215 ;

 grid_lat =
  35.26439, 35.62921, 35.98892, 36.34341, 36.69255, 37.03624, 37.37434, 
    37.70675, 38.03334, 38.354, 38.66859, 38.977, 39.27911, 39.57478, 
    39.8639, 40.14635, 40.42199, 40.69072, 40.9524, 41.20691, 41.45414, 
    41.69396, 41.92625, 42.15091, 42.36781, 42.57683, 42.77788, 42.97084, 
    43.1556, 43.33206, 43.50012, 43.65969, 43.81068, 43.95298, 44.08652, 
    44.21122, 44.32701, 44.4338, 44.53154, 44.62016, 44.6996, 44.76982, 
    44.83077, 44.88241, 44.9247, 44.95763, 44.98116, 44.99529, 45, 44.99529, 
    44.98116, 44.95763, 44.9247, 44.88241, 44.83077, 44.76982, 44.6996, 
    44.62016, 44.53154, 44.4338, 44.32701, 44.21122, 44.08652, 43.95298, 
    43.81068, 43.65969, 43.50012, 43.33206, 43.1556, 42.97084, 42.77788, 
    42.57683, 42.36781, 42.15091, 41.92625, 41.69396, 41.45414, 41.20691, 
    40.9524, 40.69072, 40.42199, 40.14635, 39.8639, 39.57478, 39.27911, 
    38.977, 38.66859, 38.354, 38.03334, 37.70675, 37.37434, 37.03624, 
    36.69255, 36.34341, 35.98892, 35.62921, 35.26439,
  35.62921, 36.00579, 36.37735, 36.74377, 37.10492, 37.46067, 37.81089, 
    38.15546, 38.49422, 38.82706, 39.15382, 39.47439, 39.78861, 40.09635, 
    40.39747, 40.69183, 40.97929, 41.25971, 41.53295, 41.79888, 42.05735, 
    42.30823, 42.55138, 42.78666, 43.01395, 43.23311, 43.44402, 43.64655, 
    43.84056, 44.02596, 44.20261, 44.37041, 44.52925, 44.67902, 44.81961, 
    44.95095, 45.07294, 45.18549, 45.28852, 45.38197, 45.46576, 45.53984, 
    45.60415, 45.65865, 45.7033, 45.73805, 45.7629, 45.77781, 45.78278, 
    45.77781, 45.7629, 45.73805, 45.7033, 45.65865, 45.60415, 45.53984, 
    45.46576, 45.38197, 45.28852, 45.18549, 45.07294, 44.95095, 44.81961, 
    44.67902, 44.52925, 44.37041, 44.20261, 44.02596, 43.84056, 43.64655, 
    43.44402, 43.23311, 43.01395, 42.78666, 42.55138, 42.30823, 42.05735, 
    41.79888, 41.53295, 41.25971, 40.97929, 40.69183, 40.39747, 40.09635, 
    39.78861, 39.47439, 39.15382, 38.82706, 38.49422, 38.15546, 37.81089, 
    37.46067, 37.10492, 36.74377, 36.37735, 36.00579, 35.62921,
  35.98892, 36.37735, 36.76087, 37.13935, 37.51265, 37.88063, 38.24314, 
    38.60004, 38.95119, 39.29642, 39.6356, 39.96857, 40.29517, 40.61526, 
    40.92867, 41.23525, 41.53484, 41.82729, 42.11243, 42.39012, 42.66019, 
    42.92249, 43.17686, 43.42315, 43.66121, 43.89089, 44.11203, 44.3245, 
    44.52815, 44.72285, 44.90845, 45.08484, 45.25187, 45.40944, 45.55742, 
    45.6957, 45.82418, 45.94276, 46.05135, 46.14986, 46.23822, 46.31635, 
    46.38419, 46.44169, 46.4888, 46.52548, 46.5517, 46.56744, 46.57269, 
    46.56744, 46.5517, 46.52548, 46.4888, 46.44169, 46.38419, 46.31635, 
    46.23822, 46.14986, 46.05135, 45.94276, 45.82418, 45.6957, 45.55742, 
    45.40944, 45.25187, 45.08484, 44.90845, 44.72285, 44.52815, 44.3245, 
    44.11203, 43.89089, 43.66121, 43.42315, 43.17686, 42.92249, 42.66019, 
    42.39012, 42.11243, 41.82729, 41.53484, 41.23525, 40.92867, 40.61526, 
    40.29517, 39.96857, 39.6356, 39.29642, 38.95119, 38.60004, 38.24314, 
    37.88063, 37.51265, 37.13935, 36.76087, 36.37735, 35.98892,
  36.34341, 36.74377, 37.13935, 37.53001, 37.91559, 38.29594, 38.67091, 
    39.04033, 39.40405, 39.7619, 40.11372, 40.45934, 40.79858, 41.13129, 
    41.45728, 41.77639, 42.08843, 42.39323, 42.69062, 42.98042, 43.26245, 
    43.53653, 43.8025, 44.06018, 44.30939, 44.54997, 44.78174, 45.00454, 
    45.21821, 45.42259, 45.61752, 45.80286, 45.97845, 46.14417, 46.29986, 
    46.4454, 46.58068, 46.70559, 46.82, 46.92382, 47.01697, 47.09935, 
    47.17091, 47.23156, 47.28126, 47.31997, 47.34763, 47.36425, 47.36979, 
    47.36425, 47.34763, 47.31997, 47.28126, 47.23156, 47.17091, 47.09935, 
    47.01697, 46.92382, 46.82, 46.70559, 46.58068, 46.4454, 46.29986, 
    46.14417, 45.97845, 45.80286, 45.61752, 45.42259, 45.21821, 45.00454, 
    44.78174, 44.54997, 44.30939, 44.06018, 43.8025, 43.53653, 43.26245, 
    42.98042, 42.69062, 42.39323, 42.08843, 41.77639, 41.45728, 41.13129, 
    40.79858, 40.45934, 40.11372, 39.7619, 39.40405, 39.04033, 38.67091, 
    38.29594, 37.91559, 37.53001, 37.13935, 36.74377, 36.34341,
  36.69255, 37.10492, 37.51265, 37.91559, 38.31358, 38.70644, 39.09401, 
    39.47613, 39.85261, 40.22328, 40.58796, 40.94647, 41.29861, 41.64421, 
    41.98307, 42.315, 42.6398, 42.95729, 43.26726, 43.56952, 43.86388, 
    44.15013, 44.42807, 44.69753, 44.95829, 45.21016, 45.45296, 45.68649, 
    45.91058, 46.12503, 46.32969, 46.52436, 46.70888, 46.8831, 47.04686, 
    47.20001, 47.34241, 47.47393, 47.59445, 47.70385, 47.80202, 47.88887, 
    47.96432, 48.02829, 48.08072, 48.12155, 48.15074, 48.16827, 48.17411, 
    48.16827, 48.15074, 48.12155, 48.08072, 48.02829, 47.96432, 47.88887, 
    47.80202, 47.70385, 47.59445, 47.47393, 47.34241, 47.20001, 47.04686, 
    46.8831, 46.70888, 46.52436, 46.32969, 46.12503, 45.91058, 45.68649, 
    45.45296, 45.21016, 44.95829, 44.69753, 44.42807, 44.15013, 43.86388, 
    43.56952, 43.26726, 42.95729, 42.6398, 42.315, 41.98307, 41.64421, 
    41.29861, 40.94647, 40.58796, 40.22328, 39.85261, 39.47613, 39.09401, 
    38.70644, 38.31358, 37.91559, 37.51265, 37.10492, 36.69255,
  37.03624, 37.46067, 37.88063, 38.29594, 38.70644, 39.11194, 39.51227, 
    39.90724, 40.29666, 40.68035, 41.0581, 41.42973, 41.79502, 42.15377, 
    42.50578, 42.85083, 43.18871, 43.51921, 43.84211, 44.15719, 44.46423, 
    44.76302, 45.05334, 45.33495, 45.60766, 45.87124, 46.12547, 46.37015, 
    46.60506, 46.83001, 47.04478, 47.24918, 47.44304, 47.62614, 47.79833, 
    47.95944, 48.10929, 48.24775, 48.37467, 48.48992, 48.59336, 48.68491, 
    48.76445, 48.83191, 48.8872, 48.93027, 48.96106, 48.97956, 48.98572, 
    48.97956, 48.96106, 48.93027, 48.8872, 48.83191, 48.76445, 48.68491, 
    48.59336, 48.48992, 48.37467, 48.24775, 48.10929, 47.95944, 47.79833, 
    47.62614, 47.44304, 47.24918, 47.04478, 46.83001, 46.60506, 46.37015, 
    46.12547, 45.87124, 45.60766, 45.33495, 45.05334, 44.76302, 44.46423, 
    44.15719, 43.84211, 43.51921, 43.18871, 42.85083, 42.50578, 42.15377, 
    41.79502, 41.42973, 41.0581, 40.68035, 40.29666, 39.90724, 39.51227, 
    39.11194, 38.70644, 38.29594, 37.88063, 37.46067, 37.03624,
  37.37434, 37.81089, 38.24314, 38.67091, 39.09401, 39.51227, 39.92548, 
    40.33345, 40.73598, 41.13287, 41.52391, 41.90887, 42.28755, 42.65972, 
    43.02515, 43.38362, 43.73489, 44.07872, 44.41489, 44.74314, 45.06325, 
    45.37495, 45.67802, 45.97221, 46.25727, 46.53297, 46.79906, 47.05531, 
    47.30147, 47.53732, 47.76263, 47.97718, 48.18076, 48.37315, 48.55416, 
    48.72359, 48.88126, 49.02699, 49.16062, 49.282, 49.39099, 49.48746, 
    49.57131, 49.64243, 49.70073, 49.74615, 49.77864, 49.79815, 49.80465, 
    49.79815, 49.77864, 49.74615, 49.70073, 49.64243, 49.57131, 49.48746, 
    49.39099, 49.282, 49.16062, 49.02699, 48.88126, 48.72359, 48.55416, 
    48.37315, 48.18076, 47.97718, 47.76263, 47.53732, 47.30147, 47.05531, 
    46.79906, 46.53297, 46.25727, 45.97221, 45.67802, 45.37495, 45.06325, 
    44.74314, 44.41489, 44.07872, 43.73489, 43.38362, 43.02515, 42.65972, 
    42.28755, 41.90887, 41.52391, 41.13287, 40.73598, 40.33345, 39.92548, 
    39.51227, 39.09401, 38.67091, 38.24314, 37.81089, 37.37434,
  37.70675, 38.15546, 38.60004, 39.04033, 39.47613, 39.90724, 40.33345, 
    40.75457, 41.17037, 41.58063, 41.98514, 42.38366, 42.77596, 43.16179, 
    43.54091, 43.91308, 44.27805, 44.63554, 44.98531, 45.3271, 45.66063, 
    45.98564, 46.30186, 46.60902, 46.90686, 47.1951, 47.47348, 47.74172, 
    47.99957, 48.24677, 48.48305, 48.70818, 48.92191, 49.124, 49.31422, 
    49.49236, 49.6582, 49.81155, 49.95222, 50.08005, 50.19486, 50.29652, 
    50.38489, 50.45986, 50.52134, 50.56924, 50.6035, 50.62407, 50.63093, 
    50.62407, 50.6035, 50.56924, 50.52134, 50.45986, 50.38489, 50.29652, 
    50.19486, 50.08005, 49.95222, 49.81155, 49.6582, 49.49236, 49.31422, 
    49.124, 48.92191, 48.70818, 48.48305, 48.24677, 47.99957, 47.74172, 
    47.47348, 47.1951, 46.90686, 46.60902, 46.30186, 45.98564, 45.66063, 
    45.3271, 44.98531, 44.63554, 44.27805, 43.91308, 43.54091, 43.16179, 
    42.77596, 42.38366, 41.98514, 41.58063, 41.17037, 40.75457, 40.33345, 
    39.90724, 39.47613, 39.04033, 38.60004, 38.15546, 37.70675,
  38.03334, 38.49422, 38.95119, 39.40405, 39.85261, 40.29666, 40.73598, 
    41.17037, 41.59958, 42.02338, 42.44154, 42.85382, 43.25996, 43.6597, 
    44.05278, 44.43893, 44.81789, 45.18936, 45.55307, 45.90874, 46.25607, 
    46.59477, 46.92454, 47.24509, 47.55613, 47.85734, 48.14844, 48.42913, 
    48.69912, 48.95811, 49.20582, 49.44197, 49.66629, 49.8785, 50.07836, 
    50.26561, 50.44002, 50.60136, 50.74942, 50.88401, 51.00494, 51.11204, 
    51.20517, 51.2842, 51.34902, 51.39953, 51.43566, 51.45736, 51.46459, 
    51.45736, 51.43566, 51.39953, 51.34902, 51.2842, 51.20517, 51.11204, 
    51.00494, 50.88401, 50.74942, 50.60136, 50.44002, 50.26561, 50.07836, 
    49.8785, 49.66629, 49.44197, 49.20582, 48.95811, 48.69912, 48.42913, 
    48.14844, 47.85734, 47.55613, 47.24509, 46.92454, 46.59477, 46.25607, 
    45.90874, 45.55307, 45.18936, 44.81789, 44.43893, 44.05278, 43.6597, 
    43.25996, 42.85382, 42.44154, 42.02338, 41.59958, 41.17037, 40.73598, 
    40.29666, 39.85261, 39.40405, 38.95119, 38.49422, 38.03334,
  38.354, 38.82706, 39.29642, 39.7619, 40.22328, 40.68035, 41.13287, 
    41.58063, 42.02338, 42.46088, 42.89287, 43.31909, 43.73928, 44.15316, 
    44.56044, 44.96085, 45.35409, 45.73986, 46.11785, 46.48775, 46.84925, 
    47.20202, 47.54575, 47.8801, 48.20476, 48.51939, 48.82367, 49.11726, 
    49.39985, 49.6711, 49.9307, 50.17833, 50.4137, 50.63649, 50.84642, 
    51.04321, 51.22659, 51.39631, 51.55212, 51.69381, 51.82117, 51.934, 
    52.03214, 52.11544, 52.18378, 52.23703, 52.27514, 52.29802, 52.30565, 
    52.29802, 52.27514, 52.23703, 52.18378, 52.11544, 52.03214, 51.934, 
    51.82117, 51.69381, 51.55212, 51.39631, 51.22659, 51.04321, 50.84642, 
    50.63649, 50.4137, 50.17833, 49.9307, 49.6711, 49.39985, 49.11726, 
    48.82367, 48.51939, 48.20476, 47.8801, 47.54575, 47.20202, 46.84925, 
    46.48775, 46.11785, 45.73986, 45.35409, 44.96085, 44.56044, 44.15316, 
    43.73928, 43.31909, 42.89287, 42.46088, 42.02338, 41.58063, 41.13287, 
    40.68035, 40.22328, 39.7619, 39.29642, 38.82706, 38.354,
  38.66859, 39.15382, 39.6356, 40.11372, 40.58796, 41.0581, 41.52391, 
    41.98514, 42.44154, 42.89287, 43.33884, 43.77919, 44.21362, 44.64186, 
    45.0636, 45.47853, 45.88634, 46.28671, 46.67929, 47.06378, 47.43981, 
    47.80704, 48.16513, 48.51371, 48.85243, 49.18093, 49.49884, 49.8058, 
    50.10146, 50.38545, 50.65742, 50.91702, 51.1639, 51.39774, 51.6182, 
    51.82498, 52.01776, 52.19627, 52.36022, 52.50938, 52.64349, 52.76235, 
    52.86576, 52.95356, 53.0256, 53.08176, 53.12194, 53.14607, 53.15412, 
    53.14607, 53.12194, 53.08176, 53.0256, 52.95356, 52.86576, 52.76235, 
    52.64349, 52.50938, 52.36022, 52.19627, 52.01776, 51.82498, 51.6182, 
    51.39774, 51.1639, 50.91702, 50.65742, 50.38545, 50.10146, 49.8058, 
    49.49884, 49.18093, 48.85243, 48.51371, 48.16513, 47.80704, 47.43981, 
    47.06378, 46.67929, 46.28671, 45.88634, 45.47853, 45.0636, 44.64186, 
    44.21362, 43.77919, 43.33884, 42.89287, 42.44154, 41.98514, 41.52391, 
    41.0581, 40.58796, 40.11372, 39.6356, 39.15382, 38.66859,
  38.977, 39.47439, 39.96857, 40.45934, 40.94647, 41.42973, 41.90887, 
    42.38366, 42.85382, 43.31909, 43.77919, 44.23382, 44.68269, 45.1255, 
    45.56192, 45.99162, 46.41428, 46.82954, 47.23705, 47.63646, 48.02739, 
    48.40947, 48.78232, 49.14555, 49.49877, 49.84158, 50.1736, 50.49441, 
    50.80363, 51.10085, 51.38569, 51.65775, 51.91666, 52.16203, 52.39351, 
    52.61073, 52.81337, 53.00109, 53.17359, 53.33059, 53.47181, 53.59702, 
    53.70599, 53.79853, 53.87448, 53.93369, 53.97606, 54.00152, 54.01001, 
    54.00152, 53.97606, 53.93369, 53.87448, 53.79853, 53.70599, 53.59702, 
    53.47181, 53.33059, 53.17359, 53.00109, 52.81337, 52.61073, 52.39351, 
    52.16203, 51.91666, 51.65775, 51.38569, 51.10085, 50.80363, 50.49441, 
    50.1736, 49.84158, 49.49877, 49.14555, 48.78232, 48.40947, 48.02739, 
    47.63646, 47.23705, 46.82954, 46.41428, 45.99162, 45.56192, 45.1255, 
    44.68269, 44.23382, 43.77919, 43.31909, 42.85382, 42.38366, 41.90887, 
    41.42973, 40.94647, 40.45934, 39.96857, 39.47439, 38.977,
  39.27911, 39.78861, 40.29517, 40.79858, 41.29861, 41.79502, 42.28755, 
    42.77596, 43.25996, 43.73928, 44.21362, 44.68269, 45.14617, 45.60374, 
    46.05505, 46.49977, 46.93754, 47.36799, 47.79074, 48.20541, 48.6116, 
    49.00891, 49.39692, 49.77522, 50.14338, 50.50098, 50.84757, 51.18272, 
    51.506, 51.81697, 52.11519, 52.40023, 52.67167, 52.92909, 53.17208, 
    53.40025, 53.61321, 53.81061, 53.99209, 54.15733, 54.30604, 54.43793, 
    54.55275, 54.6503, 54.73037, 54.79281, 54.8375, 54.86435, 54.87331, 
    54.86435, 54.8375, 54.79281, 54.73037, 54.6503, 54.55275, 54.43793, 
    54.30604, 54.15733, 53.99209, 53.81061, 53.61321, 53.40025, 53.17208, 
    52.92909, 52.67167, 52.40023, 52.11519, 51.81697, 51.506, 51.18272, 
    50.84757, 50.50098, 50.14338, 49.77522, 49.39692, 49.00891, 48.6116, 
    48.20541, 47.79074, 47.36799, 46.93754, 46.49977, 46.05505, 45.60374, 
    45.14617, 44.68269, 44.21362, 43.73928, 43.25996, 42.77596, 42.28755, 
    41.79502, 41.29861, 40.79858, 40.29517, 39.78861, 39.27911,
  39.57478, 40.09635, 40.61526, 41.13129, 41.64421, 42.15377, 42.65972, 
    43.16179, 43.6597, 44.15316, 44.64186, 45.1255, 45.60374, 46.07624, 
    46.54266, 47.00262, 47.45575, 47.90166, 48.33995, 48.77021, 49.19202, 
    49.60493, 50.00851, 50.40231, 50.78586, 51.1587, 51.52035, 51.87035, 
    52.2082, 52.53343, 52.84557, 53.14412, 53.42863, 53.69863, 53.95366, 
    54.19329, 54.41708, 54.62463, 54.81555, 54.98947, 55.14605, 55.28499, 
    55.40599, 55.50881, 55.59324, 55.65909, 55.70623, 55.73455, 55.744, 
    55.73455, 55.70623, 55.65909, 55.59324, 55.50881, 55.40599, 55.28499, 
    55.14605, 54.98947, 54.81555, 54.62463, 54.41708, 54.19329, 53.95366, 
    53.69863, 53.42863, 53.14412, 52.84557, 52.53343, 52.2082, 51.87035, 
    51.52035, 51.1587, 50.78586, 50.40231, 50.00851, 49.60493, 49.19202, 
    48.77021, 48.33995, 47.90166, 47.45575, 47.00262, 46.54266, 46.07624, 
    45.60374, 45.1255, 44.64186, 44.15316, 43.6597, 43.16179, 42.65972, 
    42.15377, 41.64421, 41.13129, 40.61526, 40.09635, 39.57478,
  39.8639, 40.39747, 40.92867, 41.45728, 41.98307, 42.50578, 43.02515, 
    43.54091, 44.05278, 44.56044, 45.0636, 45.56192, 46.05505, 46.54266, 
    47.02436, 47.49977, 47.96851, 48.43015, 48.88427, 49.33044, 49.7682, 
    50.19709, 50.61664, 51.02636, 51.42574, 51.8143, 52.1915, 52.55685, 
    52.9098, 53.24984, 53.57643, 53.88906, 54.18719, 54.47033, 54.73795, 
    54.98958, 55.22473, 55.44294, 55.64378, 55.82684, 55.99172, 56.13808, 
    56.26561, 56.374, 56.46303, 56.53249, 56.58222, 56.6121, 56.62207, 
    56.6121, 56.58222, 56.53249, 56.46303, 56.374, 56.26561, 56.13808, 
    55.99172, 55.82684, 55.64378, 55.44294, 55.22473, 54.98958, 54.73795, 
    54.47033, 54.18719, 53.88906, 53.57643, 53.24984, 52.9098, 52.55685, 
    52.1915, 51.8143, 51.42574, 51.02636, 50.61664, 50.19709, 49.7682, 
    49.33044, 48.88427, 48.43015, 47.96851, 47.49977, 47.02436, 46.54266, 
    46.05505, 45.56192, 45.0636, 44.56044, 44.05278, 43.54091, 43.02515, 
    42.50578, 41.98307, 41.45728, 40.92867, 40.39747, 39.8639,
  40.14635, 40.69183, 41.23525, 41.77639, 42.315, 42.85083, 43.38362, 
    43.91308, 44.43893, 44.96085, 45.47853, 45.99162, 46.49977, 47.00262, 
    47.49977, 47.99084, 48.4754, 48.95301, 49.42325, 49.88563, 50.33969, 
    50.78492, 51.22083, 51.64688, 52.06255, 52.46729, 52.86054, 53.24175, 
    53.61034, 53.96573, 54.30735, 54.63462, 54.94697, 55.24382, 55.52462, 
    55.78882, 56.03588, 56.26529, 56.47657, 56.66924, 56.84288, 56.99708, 
    57.13149, 57.24578, 57.33968, 57.41296, 57.46543, 57.49697, 57.50749, 
    57.49697, 57.46543, 57.41296, 57.33968, 57.24578, 57.13149, 56.99708, 
    56.84288, 56.66924, 56.47657, 56.26529, 56.03588, 55.78882, 55.52462, 
    55.24382, 54.94697, 54.63462, 54.30735, 53.96573, 53.61034, 53.24175, 
    52.86054, 52.46729, 52.06255, 51.64688, 51.22083, 50.78492, 50.33969, 
    49.88563, 49.42325, 48.95301, 48.4754, 47.99084, 47.49977, 47.00262, 
    46.49977, 45.99162, 45.47853, 44.96085, 44.43893, 43.91308, 43.38362, 
    42.85083, 42.315, 41.77639, 41.23525, 40.69183, 40.14635,
  40.42199, 40.97929, 41.53484, 42.08843, 42.6398, 43.18871, 43.73489, 
    44.27805, 44.81789, 45.35409, 45.88634, 46.41428, 46.93754, 47.45575, 
    47.96851, 48.4754, 48.97598, 49.46981, 49.95642, 50.43531, 50.90599, 
    51.36792, 51.82056, 52.26337, 52.69576, 53.11716, 53.52696, 53.92455, 
    54.30932, 54.68064, 55.03786, 55.38037, 55.70753, 56.01871, 56.31329, 
    56.59066, 56.85022, 57.09141, 57.31367, 57.51648, 57.69935, 57.86184, 
    58.00352, 58.12405, 58.22311, 58.30043, 58.35581, 58.3891, 58.40021, 
    58.3891, 58.35581, 58.30043, 58.22311, 58.12405, 58.00352, 57.86184, 
    57.69935, 57.51648, 57.31367, 57.09141, 56.85022, 56.59066, 56.31329, 
    56.01871, 55.70753, 55.38037, 55.03786, 54.68064, 54.30932, 53.92455, 
    53.52696, 53.11716, 52.69576, 52.26337, 51.82056, 51.36792, 50.90599, 
    50.43531, 49.95642, 49.46981, 48.97598, 48.4754, 47.96851, 47.45575, 
    46.93754, 46.41428, 45.88634, 45.35409, 44.81789, 44.27805, 43.73489, 
    43.18871, 42.6398, 42.08843, 41.53484, 40.97929, 40.42199,
  40.69072, 41.25971, 41.82729, 42.39323, 42.95729, 43.51921, 44.07872, 
    44.63554, 45.18936, 45.73986, 46.28671, 46.82954, 47.36799, 47.90166, 
    48.43015, 48.95301, 49.46981, 49.98007, 50.48329, 50.97897, 51.46657, 
    51.94554, 52.4153, 52.87527, 53.32483, 53.76335, 54.1902, 54.60471, 
    55.00621, 55.39402, 55.76746, 56.12582, 56.46842, 56.79456, 57.10355, 
    57.39472, 57.66741, 57.92097, 58.1548, 58.36829, 58.56092, 58.73216, 
    58.88156, 59.0087, 59.11322, 59.19484, 59.2533, 59.28845, 59.30018, 
    59.28845, 59.2533, 59.19484, 59.11322, 59.0087, 58.88156, 58.73216, 
    58.56092, 58.36829, 58.1548, 57.92097, 57.66741, 57.39472, 57.10355, 
    56.79456, 56.46842, 56.12582, 55.76746, 55.39402, 55.00621, 54.60471, 
    54.1902, 53.76335, 53.32483, 52.87527, 52.4153, 51.94554, 51.46657, 
    50.97897, 50.48329, 49.98007, 49.46981, 48.95301, 48.43015, 47.90166, 
    47.36799, 46.82954, 46.28671, 45.73986, 45.18936, 44.63554, 44.07872, 
    43.51921, 42.95729, 42.39323, 41.82729, 41.25971, 40.69072,
  40.9524, 41.53295, 42.11243, 42.69062, 43.26726, 43.84211, 44.41489, 
    44.98531, 45.55307, 46.11785, 46.67929, 47.23705, 47.79074, 48.33995, 
    48.88427, 49.42325, 49.95642, 50.48329, 51.00336, 51.51608, 52.0209, 
    52.51723, 53.00447, 53.48199, 53.94915, 54.40527, 54.84966, 55.28162, 
    55.70042, 56.10532, 56.49557, 56.87043, 57.22911, 57.57087, 57.89494, 
    58.20058, 58.48705, 58.75364, 58.99965, 59.22443, 59.42736, 59.60787, 
    59.76543, 59.89958, 60.00991, 60.09608, 60.15783, 60.19496, 60.20734, 
    60.19496, 60.15783, 60.09608, 60.00991, 59.89958, 59.76543, 59.60787, 
    59.42736, 59.22443, 58.99965, 58.75364, 58.48705, 58.20058, 57.89494, 
    57.57087, 57.22911, 56.87043, 56.49557, 56.10532, 55.70042, 55.28162, 
    54.84966, 54.40527, 53.94915, 53.48199, 53.00447, 52.51723, 52.0209, 
    51.51608, 51.00336, 50.48329, 49.95642, 49.42325, 48.88427, 48.33995, 
    47.79074, 47.23705, 46.67929, 46.11785, 45.55307, 44.98531, 44.41489, 
    43.84211, 43.26726, 42.69062, 42.11243, 41.53295, 40.9524,
  41.20691, 41.79888, 42.39012, 42.98042, 43.56952, 44.15719, 44.74314, 
    45.3271, 45.90874, 46.48775, 47.06378, 47.63646, 48.20541, 48.77021, 
    49.33044, 49.88563, 50.43531, 50.97897, 51.51608, 52.04608, 52.56838, 
    53.08239, 53.58745, 54.08292, 54.5681, 55.04227, 55.50471, 55.95465, 
    56.39131, 56.8139, 57.2216, 57.61359, 57.98904, 58.34711, 58.68696, 
    59.00777, 59.30871, 59.589, 59.84786, 60.08456, 60.29839, 60.48872, 
    60.65495, 60.79654, 60.91304, 61.00407, 61.06931, 61.10854, 61.12163, 
    61.10854, 61.06931, 61.00407, 60.91304, 60.79654, 60.65495, 60.48872, 
    60.29839, 60.08456, 59.84786, 59.589, 59.30871, 59.00777, 58.68696, 
    58.34711, 57.98904, 57.61359, 57.2216, 56.8139, 56.39131, 55.95465, 
    55.50471, 55.04227, 54.5681, 54.08292, 53.58745, 53.08239, 52.56838, 
    52.04608, 51.51608, 50.97897, 50.43531, 49.88563, 49.33044, 48.77021, 
    48.20541, 47.63646, 47.06378, 46.48775, 45.90874, 45.3271, 44.74314, 
    44.15719, 43.56952, 42.98042, 42.39012, 41.79888, 41.20691,
  41.45414, 42.05735, 42.66019, 43.26245, 43.86388, 44.46423, 45.06325, 
    45.66063, 46.25607, 46.84925, 47.43981, 48.02739, 48.6116, 49.19202, 
    49.7682, 50.33969, 50.90599, 51.46657, 52.0209, 52.56838, 53.10843, 
    53.64039, 54.16361, 54.67738, 55.18099, 55.67367, 56.15464, 56.62309, 
    57.07819, 57.51908, 57.94487, 58.35467, 58.74758, 59.12267, 59.47903, 
    59.81574, 60.1319, 60.42662, 60.69904, 60.94834, 61.17372, 61.37446, 
    61.54989, 61.6994, 61.82248, 61.91867, 61.98763, 62.02911, 62.04295, 
    62.02911, 61.98763, 61.91867, 61.82248, 61.6994, 61.54989, 61.37446, 
    61.17372, 60.94834, 60.69904, 60.42662, 60.1319, 59.81574, 59.47903, 
    59.12267, 58.74758, 58.35467, 57.94487, 57.51908, 57.07819, 56.62309, 
    56.15464, 55.67367, 55.18099, 54.67738, 54.16361, 53.64039, 53.10843, 
    52.56838, 52.0209, 51.46657, 50.90599, 50.33969, 49.7682, 49.19202, 
    48.6116, 48.02739, 47.43981, 46.84925, 46.25607, 45.66063, 45.06325, 
    44.46423, 43.86388, 43.26245, 42.66019, 42.05735, 41.45414,
  41.69396, 42.30823, 42.92249, 43.53653, 44.15013, 44.76302, 45.37495, 
    45.98564, 46.59477, 47.20202, 47.80704, 48.40947, 49.00891, 49.60493, 
    50.19709, 50.78492, 51.36792, 51.94554, 52.51723, 53.08239, 53.64039, 
    54.19058, 54.73225, 55.26468, 55.78711, 56.29873, 56.79872, 57.28621, 
    57.76032, 58.22011, 58.66464, 59.09295, 59.50403, 59.89689, 60.27053, 
    60.62392, 60.95608, 61.26601, 61.55275, 61.81537, 62.05299, 62.26479, 
    62.45001, 62.60796, 62.73804, 62.83975, 62.91269, 62.95657, 62.97122, 
    62.95657, 62.91269, 62.83975, 62.73804, 62.60796, 62.45001, 62.26479, 
    62.05299, 61.81537, 61.55275, 61.26601, 60.95608, 60.62392, 60.27053, 
    59.89689, 59.50403, 59.09295, 58.66464, 58.22011, 57.76032, 57.28621, 
    56.79872, 56.29873, 55.78711, 55.26468, 54.73225, 54.19058, 53.64039, 
    53.08239, 52.51723, 51.94554, 51.36792, 50.78492, 50.19709, 49.60493, 
    49.00891, 48.40947, 47.80704, 47.20202, 46.59477, 45.98564, 45.37495, 
    44.76302, 44.15013, 43.53653, 42.92249, 42.30823, 41.69396,
  41.92625, 42.55138, 43.17686, 43.8025, 44.42807, 45.05334, 45.67802, 
    46.30186, 46.92454, 47.54575, 48.16513, 48.78232, 49.39692, 50.00851, 
    50.61664, 51.22083, 51.82056, 52.4153, 53.00447, 53.58745, 54.16361, 
    54.73225, 55.29266, 55.84407, 56.38568, 56.91667, 57.43615, 57.9432, 
    58.43688, 58.9162, 59.38013, 59.82764, 60.25764, 60.66905, 61.06076, 
    61.43166, 61.78063, 62.10659, 62.40846, 62.6852, 62.93583, 63.15939, 
    63.35503, 63.52198, 63.65955, 63.76716, 63.84436, 63.89082, 63.90633, 
    63.89082, 63.84436, 63.76716, 63.65955, 63.52198, 63.35503, 63.15939, 
    62.93583, 62.6852, 62.40846, 62.10659, 61.78063, 61.43166, 61.06076, 
    60.66905, 60.25764, 59.82764, 59.38013, 58.9162, 58.43688, 57.9432, 
    57.43615, 56.91667, 56.38568, 55.84407, 55.29266, 54.73225, 54.16361, 
    53.58745, 53.00447, 52.4153, 51.82056, 51.22083, 50.61664, 50.00851, 
    49.39692, 48.78232, 48.16513, 47.54575, 46.92454, 46.30186, 45.67802, 
    45.05334, 44.42807, 43.8025, 43.17686, 42.55138, 41.92625,
  42.15091, 42.78666, 43.42315, 44.06018, 44.69753, 45.33495, 45.97221, 
    46.60902, 47.24509, 47.8801, 48.51371, 49.14555, 49.77522, 50.40231, 
    51.02636, 51.64688, 52.26337, 52.87527, 53.48199, 54.08292, 54.67738, 
    55.26468, 55.84407, 56.41476, 56.97591, 57.52666, 58.06607, 58.59319, 
    59.10701, 59.60646, 60.09047, 60.55789, 61.00757, 61.43833, 61.84895, 
    62.2382, 62.60488, 62.94775, 63.26563, 63.55734, 63.82177, 64.05786, 
    64.26463, 64.4412, 64.58678, 64.70073, 64.7825, 64.83172, 64.84815, 
    64.83172, 64.7825, 64.70073, 64.58678, 64.4412, 64.26463, 64.05786, 
    63.82177, 63.55734, 63.26563, 62.94775, 62.60488, 62.2382, 61.84895, 
    61.43833, 61.00757, 60.55789, 60.09047, 59.60646, 59.10701, 58.59319, 
    58.06607, 57.52666, 56.97591, 56.41476, 55.84407, 55.26468, 54.67738, 
    54.08292, 53.48199, 52.87527, 52.26337, 51.64688, 51.02636, 50.40231, 
    49.77522, 49.14555, 48.51371, 47.8801, 47.24509, 46.60902, 45.97221, 
    45.33495, 44.69753, 44.06018, 43.42315, 42.78666, 42.15091,
  42.36781, 43.01395, 43.66121, 44.30939, 44.95829, 45.60766, 46.25727, 
    46.90686, 47.55613, 48.20476, 48.85243, 49.49877, 50.14338, 50.78586, 
    51.42574, 52.06255, 52.69576, 53.32483, 53.94915, 54.5681, 55.18099, 
    55.78711, 56.38568, 56.97591, 57.55692, 58.1278, 58.68758, 59.23526, 
    59.76975, 60.28995, 60.79469, 61.28276, 61.7529, 62.20383, 62.63423, 
    63.04275, 63.42805, 63.78878, 64.1236, 64.4312, 64.71033, 64.95979, 
    65.17846, 65.36533, 65.51952, 65.64027, 65.72695, 65.77914, 65.79657, 
    65.77914, 65.72695, 65.64027, 65.51952, 65.36533, 65.17846, 64.95979, 
    64.71033, 64.4312, 64.1236, 63.78878, 63.42805, 63.04275, 62.63423, 
    62.20383, 61.7529, 61.28276, 60.79469, 60.28995, 59.76975, 59.23526, 
    58.68758, 58.1278, 57.55692, 56.97591, 56.38568, 55.78711, 55.18099, 
    54.5681, 53.94915, 53.32483, 52.69576, 52.06255, 51.42574, 50.78586, 
    50.14338, 49.49877, 48.85243, 48.20476, 47.55613, 46.90686, 46.25727, 
    45.60766, 44.95829, 44.30939, 43.66121, 43.01395, 42.36781,
  42.57683, 43.23311, 43.89089, 44.54997, 45.21016, 45.87124, 46.53297, 
    47.1951, 47.85734, 48.51939, 49.18093, 49.84158, 50.50098, 51.1587, 
    51.8143, 52.46729, 53.11716, 53.76335, 54.40527, 55.04227, 55.67367, 
    56.29873, 56.91667, 57.52666, 58.1278, 58.71915, 59.2997, 59.86839, 
    60.4241, 60.96564, 61.49178, 62.00122, 62.49262, 62.96457, 63.41565, 
    63.84439, 64.2493, 64.62888, 64.98164, 65.30614, 65.60093, 65.86467, 
    66.09609, 66.29404, 66.45748, 66.58555, 66.67754, 66.73294, 66.75144, 
    66.73294, 66.67754, 66.58555, 66.45748, 66.29404, 66.09609, 65.86467, 
    65.60093, 65.30614, 64.98164, 64.62888, 64.2493, 63.84439, 63.41565, 
    62.96457, 62.49262, 62.00122, 61.49178, 60.96564, 60.4241, 59.86839, 
    59.2997, 58.71915, 58.1278, 57.52666, 56.91667, 56.29873, 55.67367, 
    55.04227, 54.40527, 53.76335, 53.11716, 52.46729, 51.8143, 51.1587, 
    50.50098, 49.84158, 49.18093, 48.51939, 47.85734, 47.1951, 46.53297, 
    45.87124, 45.21016, 44.54997, 43.89089, 43.23311, 42.57683,
  42.77788, 43.44402, 44.11203, 44.78174, 45.45296, 46.12547, 46.79906, 
    47.47348, 48.14844, 48.82367, 49.49884, 50.1736, 50.84757, 51.52035, 
    52.1915, 52.86054, 53.52696, 54.1902, 54.84966, 55.50471, 56.15464, 
    56.79872, 57.43615, 58.06607, 58.68758, 59.2997, 59.90138, 60.49152, 
    61.06895, 61.63241, 62.18061, 62.71215, 63.2256, 63.71946, 64.19215, 
    64.6421, 65.06765, 65.46716, 65.83895, 66.18141, 66.49293, 66.77197, 
    67.01707, 67.22693, 67.40035, 67.53634, 67.63406, 67.69295, 67.71262, 
    67.69295, 67.63406, 67.53634, 67.40035, 67.22693, 67.01707, 66.77197, 
    66.49293, 66.18141, 65.83895, 65.46716, 65.06765, 64.6421, 64.19215, 
    63.71946, 63.2256, 62.71215, 62.18061, 61.63241, 61.06895, 60.49152, 
    59.90138, 59.2997, 58.68758, 58.06607, 57.43615, 56.79872, 56.15464, 
    55.50471, 54.84966, 54.1902, 53.52696, 52.86054, 52.1915, 51.52035, 
    50.84757, 50.1736, 49.49884, 48.82367, 48.14844, 47.47348, 46.79906, 
    46.12547, 45.45296, 44.78174, 44.11203, 43.44402, 42.77788,
  42.97084, 43.64655, 44.3245, 45.00454, 45.68649, 46.37015, 47.05531, 
    47.74172, 48.42913, 49.11726, 49.8058, 50.49441, 51.18272, 51.87035, 
    52.55685, 53.24175, 53.92455, 54.60471, 55.28162, 55.95465, 56.62309, 
    57.28621, 57.9432, 58.59319, 59.23526, 59.86839, 60.49152, 61.1035, 
    61.70312, 62.28906, 62.85994, 63.41431, 63.95062, 64.46726, 64.96255, 
    65.43473, 65.88202, 66.30258, 66.69459, 67.05619, 67.38558, 67.68102, 
    67.94086, 68.16358, 68.3478, 68.49236, 68.59633, 68.65899, 68.67992, 
    68.65899, 68.59633, 68.49236, 68.3478, 68.16358, 67.94086, 67.68102, 
    67.38558, 67.05619, 66.69459, 66.30258, 65.88202, 65.43473, 64.96255, 
    64.46726, 63.95062, 63.41431, 62.85994, 62.28906, 61.70312, 61.1035, 
    60.49152, 59.86839, 59.23526, 58.59319, 57.9432, 57.28621, 56.62309, 
    55.95465, 55.28162, 54.60471, 53.92455, 53.24175, 52.55685, 51.87035, 
    51.18272, 50.49441, 49.8058, 49.11726, 48.42913, 47.74172, 47.05531, 
    46.37015, 45.68649, 45.00454, 44.3245, 43.64655, 42.97084,
  43.1556, 43.84056, 44.52815, 45.21821, 45.91058, 46.60506, 47.30147, 
    47.99957, 48.69912, 49.39985, 50.10146, 50.80363, 51.506, 52.2082, 
    52.9098, 53.61034, 54.30932, 55.00621, 55.70042, 56.39131, 57.07819, 
    57.76032, 58.43688, 59.10701, 59.76975, 60.4241, 61.06895, 61.70312, 
    62.32535, 62.93428, 63.52847, 64.10636, 64.66634, 65.20666, 65.72551, 
    66.22101, 66.69118, 67.13403, 67.54749, 67.9295, 68.27805, 68.59113, 
    68.86686, 69.10349, 69.29943, 69.45333, 69.56409, 69.63087, 69.65318, 
    69.63087, 69.56409, 69.45333, 69.29943, 69.10349, 68.86686, 68.59113, 
    68.27805, 67.9295, 67.54749, 67.13403, 66.69118, 66.22101, 65.72551, 
    65.20666, 64.66634, 64.10636, 63.52847, 62.93428, 62.32535, 61.70312, 
    61.06895, 60.4241, 59.76975, 59.10701, 58.43688, 57.76032, 57.07819, 
    56.39131, 55.70042, 55.00621, 54.30932, 53.61034, 52.9098, 52.2082, 
    51.506, 50.80363, 50.10146, 49.39985, 48.69912, 47.99957, 47.30147, 
    46.60506, 45.91058, 45.21821, 44.52815, 43.84056, 43.1556,
  43.33206, 44.02596, 44.72285, 45.42259, 46.12503, 46.83001, 47.53732, 
    48.24677, 48.95811, 49.6711, 50.38545, 51.10085, 51.81697, 52.53343, 
    53.24984, 53.96573, 54.68064, 55.39402, 56.10532, 56.8139, 57.51908, 
    58.22011, 58.9162, 59.60646, 60.28995, 60.96564, 61.63241, 62.28906, 
    62.93428, 63.56667, 64.18473, 64.78683, 65.37125, 65.93615, 66.47958, 
    66.9995, 67.49377, 67.96017, 68.39644, 68.80025, 69.16933, 69.50142, 
    69.79435, 70.04609, 70.2548, 70.4189, 70.53708, 70.60838, 70.63222, 
    70.60838, 70.53708, 70.4189, 70.2548, 70.04609, 69.79435, 69.50142, 
    69.16933, 68.80025, 68.39644, 67.96017, 67.49377, 66.9995, 66.47958, 
    65.93615, 65.37125, 64.78683, 64.18473, 63.56667, 62.93428, 62.28906, 
    61.63241, 60.96564, 60.28995, 59.60646, 58.9162, 58.22011, 57.51908, 
    56.8139, 56.10532, 55.39402, 54.68064, 53.96573, 53.24984, 52.53343, 
    51.81697, 51.10085, 50.38545, 49.6711, 48.95811, 48.24677, 47.53732, 
    46.83001, 46.12503, 45.42259, 44.72285, 44.02596, 43.33206,
  43.50012, 44.20261, 44.90845, 45.61752, 46.32969, 47.04478, 47.76263, 
    48.48305, 49.20582, 49.9307, 50.65742, 51.38569, 52.11519, 52.84557, 
    53.57643, 54.30735, 55.03786, 55.76746, 56.49557, 57.2216, 57.94487, 
    58.66464, 59.38013, 60.09047, 60.79469, 61.49178, 62.18061, 62.85994, 
    63.52847, 64.18473, 64.82718, 65.45412, 66.06374, 66.65411, 67.22313, 
    67.76861, 68.28822, 68.77954, 69.24005, 69.66718, 70.05833, 70.41093, 
    70.72251, 70.99072, 71.21339, 71.38868, 71.51503, 71.59132, 71.61682, 
    71.59132, 71.51503, 71.38868, 71.21339, 70.99072, 70.72251, 70.41093, 
    70.05833, 69.66718, 69.24005, 68.77954, 68.28822, 67.76861, 67.22313, 
    66.65411, 66.06374, 65.45412, 64.82718, 64.18473, 63.52847, 62.85994, 
    62.18061, 61.49178, 60.79469, 60.09047, 59.38013, 58.66464, 57.94487, 
    57.2216, 56.49557, 55.76746, 55.03786, 54.30735, 53.57643, 52.84557, 
    52.11519, 51.38569, 50.65742, 49.9307, 49.20582, 48.48305, 47.76263, 
    47.04478, 46.32969, 45.61752, 44.90845, 44.20261, 43.50012,
  43.65969, 44.37041, 45.08484, 45.80286, 46.52436, 47.24918, 47.97718, 
    48.70818, 49.44197, 50.17833, 50.91702, 51.65775, 52.40023, 53.14412, 
    53.88906, 54.63462, 55.38037, 56.12582, 56.87043, 57.61359, 58.35467, 
    59.09295, 59.82764, 60.55789, 61.28276, 62.00122, 62.71215, 63.41431, 
    64.10636, 64.78683, 65.45412, 66.10648, 66.74202, 67.3587, 67.95432, 
    68.5265, 69.07276, 69.59042, 70.07672, 70.52879, 70.9437, 71.31852, 
    71.6504, 71.9366, 72.17461, 72.36224, 72.49763, 72.57942, 72.60679, 
    72.57942, 72.49763, 72.36224, 72.17461, 71.9366, 71.6504, 71.31852, 
    70.9437, 70.52879, 70.07672, 69.59042, 69.07276, 68.5265, 67.95432, 
    67.3587, 66.74202, 66.10648, 65.45412, 64.78683, 64.10636, 63.41431, 
    62.71215, 62.00122, 61.28276, 60.55789, 59.82764, 59.09295, 58.35467, 
    57.61359, 56.87043, 56.12582, 55.38037, 54.63462, 53.88906, 53.14412, 
    52.40023, 51.65775, 50.91702, 50.17833, 49.44197, 48.70818, 47.97718, 
    47.24918, 46.52436, 45.80286, 45.08484, 44.37041, 43.65969,
  43.81068, 44.52925, 45.25187, 45.97845, 46.70888, 47.44304, 48.18076, 
    48.92191, 49.66629, 50.4137, 51.1639, 51.91666, 52.67167, 53.42863, 
    54.18719, 54.94697, 55.70753, 56.46842, 57.22911, 57.98904, 58.74758, 
    59.50403, 60.25764, 61.00757, 61.7529, 62.49262, 63.2256, 63.95062, 
    64.66634, 65.37125, 66.06374, 66.74202, 67.40413, 68.04794, 68.67112, 
    69.27117, 69.84539, 70.39089, 70.90462, 71.38338, 71.8239, 72.22283, 
    72.57687, 72.88284, 73.13778, 73.33907, 73.4845, 73.57245, 73.60188, 
    73.57245, 73.4845, 73.33907, 73.13778, 72.88284, 72.57687, 72.22283, 
    71.8239, 71.38338, 70.90462, 70.39089, 69.84539, 69.27117, 68.67112, 
    68.04794, 67.40413, 66.74202, 66.06374, 65.37125, 64.66634, 63.95062, 
    63.2256, 62.49262, 61.7529, 61.00757, 60.25764, 59.50403, 58.74758, 
    57.98904, 57.22911, 56.46842, 55.70753, 54.94697, 54.18719, 53.42863, 
    52.67167, 51.91666, 51.1639, 50.4137, 49.66629, 48.92191, 48.18076, 
    47.44304, 46.70888, 45.97845, 45.25187, 44.52925, 43.81068,
  43.95298, 44.67902, 45.40944, 46.14417, 46.8831, 47.62614, 48.37315, 
    49.124, 49.8785, 50.63649, 51.39774, 52.16203, 52.92909, 53.69863, 
    54.47033, 55.24382, 56.01871, 56.79456, 57.57087, 58.34711, 59.12267, 
    59.89689, 60.66905, 61.43833, 62.20383, 62.96457, 63.71946, 64.46726, 
    65.20666, 65.93615, 66.65411, 67.3587, 68.04794, 68.7196, 69.37128, 
    70.00032, 70.60384, 71.17871, 71.7216, 72.22897, 72.69713, 73.12227, 
    73.50058, 73.82835, 74.10206, 74.31858, 74.47527, 74.57011, 74.60188, 
    74.57011, 74.47527, 74.31858, 74.10206, 73.82835, 73.50058, 73.12227, 
    72.69713, 72.22897, 71.7216, 71.17871, 70.60384, 70.00032, 69.37128, 
    68.7196, 68.04794, 67.3587, 66.65411, 65.93615, 65.20666, 64.46726, 
    63.71946, 62.96457, 62.20383, 61.43833, 60.66905, 59.89689, 59.12267, 
    58.34711, 57.57087, 56.79456, 56.01871, 55.24382, 54.47033, 53.69863, 
    52.92909, 52.16203, 51.39774, 50.63649, 49.8785, 49.124, 48.37315, 
    47.62614, 46.8831, 46.14417, 45.40944, 44.67902, 43.95298,
  44.08652, 44.81961, 45.55742, 46.29986, 47.04686, 47.79833, 48.55416, 
    49.31422, 50.07836, 50.84642, 51.6182, 52.39351, 53.17208, 53.95366, 
    54.73795, 55.52462, 56.31329, 57.10355, 57.89494, 58.68696, 59.47903, 
    60.27053, 61.06076, 61.84895, 62.63423, 63.41565, 64.19215, 64.96255, 
    65.72551, 66.47958, 67.22313, 67.95432, 68.67112, 69.37128, 70.0523, 
    70.7114, 71.34553, 71.95134, 72.5252, 73.06321, 73.56123, 74.01492, 
    74.41991, 74.77181, 75.06647, 75.30009, 75.46947, 75.57212, 75.60651, 
    75.57212, 75.46947, 75.30009, 75.06647, 74.77181, 74.41991, 74.01492, 
    73.56123, 73.06321, 72.5252, 71.95134, 71.34553, 70.7114, 70.0523, 
    69.37128, 68.67112, 67.95432, 67.22313, 66.47958, 65.72551, 64.96255, 
    64.19215, 63.41565, 62.63423, 61.84895, 61.06076, 60.27053, 59.47903, 
    58.68696, 57.89494, 57.10355, 56.31329, 55.52462, 54.73795, 53.95366, 
    53.17208, 52.39351, 51.6182, 50.84642, 50.07836, 49.31422, 48.55416, 
    47.79833, 47.04686, 46.29986, 45.55742, 44.81961, 44.08652,
  44.21122, 44.95095, 45.6957, 46.4454, 47.20001, 47.95944, 48.72359, 
    49.49236, 50.26561, 51.04321, 51.82498, 52.61073, 53.40025, 54.19329, 
    54.98958, 55.78882, 56.59066, 57.39472, 58.20058, 59.00777, 59.81574, 
    60.62392, 61.43166, 62.2382, 63.04275, 63.84439, 64.6421, 65.43473, 
    66.22101, 66.9995, 67.76861, 68.5265, 69.27117, 70.00032, 70.7114, 
    71.40154, 72.06753, 72.70583, 73.31252, 73.88333, 74.41362, 74.8985, 
    75.33289, 75.71165, 76.02982, 76.28278, 76.46657, 76.57815, 76.61555, 
    76.57815, 76.46657, 76.28278, 76.02982, 75.71165, 75.33289, 74.8985, 
    74.41362, 73.88333, 73.31252, 72.70583, 72.06753, 71.40154, 70.7114, 
    70.00032, 69.27117, 68.5265, 67.76861, 66.9995, 66.22101, 65.43473, 
    64.6421, 63.84439, 63.04275, 62.2382, 61.43166, 60.62392, 59.81574, 
    59.00777, 58.20058, 57.39472, 56.59066, 55.78882, 54.98958, 54.19329, 
    53.40025, 52.61073, 51.82498, 51.04321, 50.26561, 49.49236, 48.72359, 
    47.95944, 47.20001, 46.4454, 45.6957, 44.95095, 44.21122,
  44.32701, 45.07294, 45.82418, 46.58068, 47.34241, 48.10929, 48.88126, 
    49.6582, 50.44002, 51.22659, 52.01776, 52.81337, 53.61321, 54.41708, 
    55.22473, 56.03588, 56.85022, 57.66741, 58.48705, 59.30871, 60.1319, 
    60.95608, 61.78063, 62.60488, 63.42805, 64.2493, 65.06765, 65.88202, 
    66.69118, 67.49377, 68.28822, 69.07276, 69.84539, 70.60384, 71.34553, 
    72.06753, 72.76654, 73.43884, 74.08022, 74.68606, 75.25123, 75.77019, 
    76.23708, 76.64588, 76.99059, 77.26559, 77.46595, 77.58782, 77.62873, 
    77.58782, 77.46595, 77.26559, 76.99059, 76.64588, 76.23708, 75.77019, 
    75.25123, 74.68606, 74.08022, 73.43884, 72.76654, 72.06753, 71.34553, 
    70.60384, 69.84539, 69.07276, 68.28822, 67.49377, 66.69118, 65.88202, 
    65.06765, 64.2493, 63.42805, 62.60488, 61.78063, 60.95608, 60.1319, 
    59.30871, 58.48705, 57.66741, 56.85022, 56.03588, 55.22473, 54.41708, 
    53.61321, 52.81337, 52.01776, 51.22659, 50.44002, 49.6582, 48.88126, 
    48.10929, 47.34241, 46.58068, 45.82418, 45.07294, 44.32701,
  44.4338, 45.18549, 45.94276, 46.70559, 47.47393, 48.24775, 49.02699, 
    49.81155, 50.60136, 51.39631, 52.19627, 53.00109, 53.81061, 54.62463, 
    55.44294, 56.26529, 57.09141, 57.92097, 58.75364, 59.589, 60.42662, 
    61.26601, 62.10659, 62.94775, 63.78878, 64.62888, 65.46716, 66.30258, 
    67.13403, 67.96017, 68.77954, 69.59042, 70.39089, 71.17871, 71.95134, 
    72.70583, 73.43884, 74.14648, 74.82438, 75.46753, 76.07032, 76.62655, 
    77.12947, 77.572, 77.94691, 78.24726, 78.46685, 78.60075, 78.64574, 
    78.60075, 78.46685, 78.24726, 77.94691, 77.572, 77.12947, 76.62655, 
    76.07032, 75.46753, 74.82438, 74.14648, 73.43884, 72.70583, 71.95134, 
    71.17871, 70.39089, 69.59042, 68.77954, 67.96017, 67.13403, 66.30258, 
    65.46716, 64.62888, 63.78878, 62.94775, 62.10659, 61.26601, 60.42662, 
    59.589, 58.75364, 57.92097, 57.09141, 56.26529, 55.44294, 54.62463, 
    53.81061, 53.00109, 52.19627, 51.39631, 50.60136, 49.81155, 49.02699, 
    48.24775, 47.47393, 46.70559, 45.94276, 45.18549, 44.4338,
  44.53154, 45.28852, 46.05135, 46.82, 47.59445, 48.37467, 49.16062, 
    49.95222, 50.74942, 51.55212, 52.36022, 53.17359, 53.99209, 54.81555, 
    55.64378, 56.47657, 57.31367, 58.1548, 58.99965, 59.84786, 60.69904, 
    61.55275, 62.40846, 63.26563, 64.1236, 64.98164, 65.83895, 66.69459, 
    67.54749, 68.39644, 69.24005, 70.07672, 70.90462, 71.7216, 72.5252, 
    73.31252, 74.08022, 74.82438, 75.54044, 76.22314, 76.86639, 77.46332, 
    78.00623, 78.4868, 78.89631, 79.22611, 79.46831, 79.61646, 79.66634, 
    79.61646, 79.46831, 79.22611, 78.89631, 78.4868, 78.00623, 77.46332, 
    76.86639, 76.22314, 75.54044, 74.82438, 74.08022, 73.31252, 72.5252, 
    71.7216, 70.90462, 70.07672, 69.24005, 68.39644, 67.54749, 66.69459, 
    65.83895, 64.98164, 64.1236, 63.26563, 62.40846, 61.55275, 60.69904, 
    59.84786, 58.99965, 58.1548, 57.31367, 56.47657, 55.64378, 54.81555, 
    53.99209, 53.17359, 52.36022, 51.55212, 50.74942, 49.95222, 49.16062, 
    48.37467, 47.59445, 46.82, 46.05135, 45.28852, 44.53154,
  44.62016, 45.38197, 46.14986, 46.92382, 47.70385, 48.48992, 49.282, 
    50.08005, 50.88401, 51.69381, 52.50938, 53.33059, 54.15733, 54.98947, 
    55.82684, 56.66924, 57.51648, 58.36829, 59.22443, 60.08456, 60.94834, 
    61.81537, 62.6852, 63.55734, 64.4312, 65.30614, 66.18141, 67.05619, 
    67.9295, 68.80025, 69.66718, 70.52879, 71.38338, 72.22897, 73.06321, 
    73.88333, 74.68606, 75.46753, 76.22314, 76.94742, 77.63395, 78.2752, 
    78.8625, 79.38612, 79.83553, 80.19992, 80.46906, 80.6344, 80.69019, 
    80.6344, 80.46906, 80.19992, 79.83553, 79.38612, 78.8625, 78.2752, 
    77.63395, 76.94742, 76.22314, 75.46753, 74.68606, 73.88333, 73.06321, 
    72.22897, 71.38338, 70.52879, 69.66718, 68.80025, 67.9295, 67.05619, 
    66.18141, 65.30614, 64.4312, 63.55734, 62.6852, 61.81537, 60.94834, 
    60.08456, 59.22443, 58.36829, 57.51648, 56.66924, 55.82684, 54.98947, 
    54.15733, 53.33059, 52.50938, 51.69381, 50.88401, 50.08005, 49.282, 
    48.48992, 47.70385, 46.92382, 46.14986, 45.38197, 44.62016,
  44.6996, 45.46576, 46.23822, 47.01697, 47.80202, 48.59336, 49.39099, 
    50.19486, 51.00494, 51.82117, 52.64349, 53.47181, 54.30604, 55.14605, 
    55.99172, 56.84288, 57.69935, 58.56092, 59.42736, 60.29839, 61.17372, 
    62.05299, 62.93583, 63.82177, 64.71033, 65.60093, 66.49293, 67.38558, 
    68.27805, 69.16933, 70.05833, 70.9437, 71.8239, 72.69713, 73.56123, 
    74.41362, 75.25123, 76.07032, 76.86639, 77.63395, 78.36636, 79.05556, 
    79.69198, 80.2644, 80.76014, 81.16562, 81.46742, 81.65389, 81.71702, 
    81.65389, 81.46742, 81.16562, 80.76014, 80.2644, 79.69198, 79.05556, 
    78.36636, 77.63395, 76.86639, 76.07032, 75.25123, 74.41362, 73.56123, 
    72.69713, 71.8239, 70.9437, 70.05833, 69.16933, 68.27805, 67.38558, 
    66.49293, 65.60093, 64.71033, 63.82177, 62.93583, 62.05299, 61.17372, 
    60.29839, 59.42736, 58.56092, 57.69935, 56.84288, 55.99172, 55.14605, 
    54.30604, 53.47181, 52.64349, 51.82117, 51.00494, 50.19486, 49.39099, 
    48.59336, 47.80202, 47.01697, 46.23822, 45.46576, 44.6996,
  44.76982, 45.53984, 46.31635, 47.09935, 47.88887, 48.68491, 49.48746, 
    50.29652, 51.11204, 51.934, 52.76235, 53.59702, 54.43793, 55.28499, 
    56.13808, 56.99708, 57.86184, 58.73216, 59.60787, 60.48872, 61.37446, 
    62.26479, 63.15939, 64.05786, 64.95979, 65.86467, 66.77197, 67.68102, 
    68.59113, 69.50142, 70.41093, 71.31852, 72.22283, 73.12227, 74.01492, 
    74.8985, 75.77019, 76.62655, 77.46332, 78.2752, 79.05556, 79.7961, 
    80.48651, 81.11414, 81.66392, 82.11877, 82.46091, 82.67403, 82.7465, 
    82.67403, 82.46091, 82.11877, 81.66392, 81.11414, 80.48651, 79.7961, 
    79.05556, 78.2752, 77.46332, 76.62655, 75.77019, 74.8985, 74.01492, 
    73.12227, 72.22283, 71.31852, 70.41093, 69.50142, 68.59113, 67.68102, 
    66.77197, 65.86467, 64.95979, 64.05786, 63.15939, 62.26479, 61.37446, 
    60.48872, 59.60787, 58.73216, 57.86184, 56.99708, 56.13808, 55.28499, 
    54.43793, 53.59702, 52.76235, 51.934, 51.11204, 50.29652, 49.48746, 
    48.68491, 47.88887, 47.09935, 46.31635, 45.53984, 44.76982,
  44.83077, 45.60415, 46.38419, 47.17091, 47.96432, 48.76445, 49.57131, 
    50.38489, 51.20517, 52.03214, 52.86576, 53.70599, 54.55275, 55.40599, 
    56.26561, 57.13149, 58.00352, 58.88156, 59.76543, 60.65495, 61.54989, 
    62.45001, 63.35503, 64.26463, 65.17846, 66.09609, 67.01707, 67.94086, 
    68.86686, 69.79435, 70.72251, 71.6504, 72.57687, 73.50058, 74.41991, 
    75.33289, 76.23708, 77.12947, 78.00623, 78.8625, 79.69198, 80.48651, 
    81.23547, 81.92511, 82.53796, 83.0528, 83.44577, 83.69351, 83.77832, 
    83.69351, 83.44577, 83.0528, 82.53796, 81.92511, 81.23547, 80.48651, 
    79.69198, 78.8625, 78.00623, 77.12947, 76.23708, 75.33289, 74.41991, 
    73.50058, 72.57687, 71.6504, 70.72251, 69.79435, 68.86686, 67.94086, 
    67.01707, 66.09609, 65.17846, 64.26463, 63.35503, 62.45001, 61.54989, 
    60.65495, 59.76543, 58.88156, 58.00352, 57.13149, 56.26561, 55.40599, 
    54.55275, 53.70599, 52.86576, 52.03214, 51.20517, 50.38489, 49.57131, 
    48.76445, 47.96432, 47.17091, 46.38419, 45.60415, 44.83077,
  44.88241, 45.65865, 46.44169, 47.23156, 48.02829, 48.83191, 49.64243, 
    50.45986, 51.2842, 52.11544, 52.95356, 53.79853, 54.6503, 55.50881, 
    56.374, 57.24578, 58.12405, 59.0087, 59.89958, 60.79654, 61.6994, 
    62.60796, 63.52198, 64.4412, 65.36533, 66.29404, 67.22693, 68.16358, 
    69.10349, 70.04609, 70.99072, 71.9366, 72.88284, 73.82835, 74.77181, 
    75.71165, 76.64588, 77.572, 78.4868, 79.38612, 80.2644, 81.11414, 
    81.92511, 82.6832, 83.36916, 83.95731, 84.41584, 84.71027, 84.81216, 
    84.71027, 84.41584, 83.95731, 83.36916, 82.6832, 81.92511, 81.11414, 
    80.2644, 79.38612, 78.4868, 77.572, 76.64588, 75.71165, 74.77181, 
    73.82835, 72.88284, 71.9366, 70.99072, 70.04609, 69.10349, 68.16358, 
    67.22693, 66.29404, 65.36533, 64.4412, 63.52198, 62.60796, 61.6994, 
    60.79654, 59.89958, 59.0087, 58.12405, 57.24578, 56.374, 55.50881, 
    54.6503, 53.79853, 52.95356, 52.11544, 51.2842, 50.45986, 49.64243, 
    48.83191, 48.02829, 47.23156, 46.44169, 45.65865, 44.88241,
  44.9247, 45.7033, 46.4888, 47.28126, 48.08072, 48.8872, 49.70073, 50.52134, 
    51.34902, 52.18378, 53.0256, 53.87448, 54.73037, 55.59324, 56.46303, 
    57.33968, 58.22311, 59.11322, 60.00991, 60.91304, 61.82248, 62.73804, 
    63.65955, 64.58678, 65.51952, 66.45748, 67.40035, 68.3478, 69.29943, 
    70.2548, 71.21339, 72.17461, 73.13778, 74.10206, 75.06647, 76.02982, 
    76.99059, 77.94691, 78.89631, 79.83553, 80.76014, 81.66392, 82.53796, 
    83.36916, 84.13799, 84.81542, 85.36021, 85.72057, 85.84769, 85.72057, 
    85.36021, 84.81542, 84.13799, 83.36916, 82.53796, 81.66392, 80.76014, 
    79.83553, 78.89631, 77.94691, 76.99059, 76.02982, 75.06647, 74.10206, 
    73.13778, 72.17461, 71.21339, 70.2548, 69.29943, 68.3478, 67.40035, 
    66.45748, 65.51952, 64.58678, 63.65955, 62.73804, 61.82248, 60.91304, 
    60.00991, 59.11322, 58.22311, 57.33968, 56.46303, 55.59324, 54.73037, 
    53.87448, 53.0256, 52.18378, 51.34902, 50.52134, 49.70073, 48.8872, 
    48.08072, 47.28126, 46.4888, 45.7033, 44.9247,
  44.95763, 45.73805, 46.52548, 47.31997, 48.12155, 48.93027, 49.74615, 
    50.56924, 51.39953, 52.23703, 53.08176, 53.93369, 54.79281, 55.65909, 
    56.53249, 57.41296, 58.30043, 59.19484, 60.09608, 61.00407, 61.91867, 
    62.83975, 63.76716, 64.70073, 65.64027, 66.58555, 67.53634, 68.49236, 
    69.45333, 70.4189, 71.38868, 72.36224, 73.33907, 74.31858, 75.30009, 
    76.28278, 77.26559, 78.24726, 79.22611, 80.19992, 81.16562, 82.11877, 
    83.0528, 83.95731, 84.81542, 85.59846, 86.25768, 86.71655, 86.88457, 
    86.71655, 86.25768, 85.59846, 84.81542, 83.95731, 83.0528, 82.11877, 
    81.16562, 80.19992, 79.22611, 78.24726, 77.26559, 76.28278, 75.30009, 
    74.31858, 73.33907, 72.36224, 71.38868, 70.4189, 69.45333, 68.49236, 
    67.53634, 66.58555, 65.64027, 64.70073, 63.76716, 62.83975, 61.91867, 
    61.00407, 60.09608, 59.19484, 58.30043, 57.41296, 56.53249, 55.65909, 
    54.79281, 53.93369, 53.08176, 52.23703, 51.39953, 50.56924, 49.74615, 
    48.93027, 48.12155, 47.31997, 46.52548, 45.73805, 44.95763,
  44.98116, 45.7629, 46.5517, 47.34763, 48.15074, 48.96106, 49.77864, 
    50.6035, 51.43566, 52.27514, 53.12194, 53.97606, 54.8375, 55.70623, 
    56.58222, 57.46543, 58.35581, 59.2533, 60.15783, 61.06931, 61.98763, 
    62.91269, 63.84436, 64.7825, 65.72695, 66.67754, 67.63406, 68.59633, 
    69.56409, 70.53708, 71.51503, 72.49763, 73.4845, 74.47527, 75.46947, 
    76.46657, 77.46595, 78.46685, 79.46831, 80.46906, 81.46742, 82.46091, 
    83.44577, 84.41584, 85.36021, 86.25768, 87.06323, 87.6776, 87.92248, 
    87.6776, 87.06323, 86.25768, 85.36021, 84.41584, 83.44577, 82.46091, 
    81.46742, 80.46906, 79.46831, 78.46685, 77.46595, 76.46657, 75.46947, 
    74.47527, 73.4845, 72.49763, 71.51503, 70.53708, 69.56409, 68.59633, 
    67.63406, 66.67754, 65.72695, 64.7825, 63.84436, 62.91269, 61.98763, 
    61.06931, 60.15783, 59.2533, 58.35581, 57.46543, 56.58222, 55.70623, 
    54.8375, 53.97606, 53.12194, 52.27514, 51.43566, 50.6035, 49.77864, 
    48.96106, 48.15074, 47.34763, 46.5517, 45.7629, 44.98116,
  44.99529, 45.77781, 46.56744, 47.36425, 48.16827, 48.97956, 49.79815, 
    50.62407, 51.45736, 52.29802, 53.14607, 54.00152, 54.86435, 55.73455, 
    56.6121, 57.49697, 58.3891, 59.28845, 60.19496, 61.10854, 62.02911, 
    62.95657, 63.89082, 64.83172, 65.77914, 66.73294, 67.69295, 68.65899, 
    69.63087, 70.60838, 71.59132, 72.57942, 73.57245, 74.57011, 75.57212, 
    76.57815, 77.58782, 78.60075, 79.61646, 80.6344, 81.65389, 82.67403, 
    83.69351, 84.71027, 85.72057, 86.71655, 87.6776, 88.53089, 88.96107, 
    88.53089, 87.6776, 86.71655, 85.72057, 84.71027, 83.69351, 82.67403, 
    81.65389, 80.6344, 79.61646, 78.60075, 77.58782, 76.57815, 75.57212, 
    74.57011, 73.57245, 72.57942, 71.59132, 70.60838, 69.63087, 68.65899, 
    67.69295, 66.73294, 65.77914, 64.83172, 63.89082, 62.95657, 62.02911, 
    61.10854, 60.19496, 59.28845, 58.3891, 57.49697, 56.6121, 55.73455, 
    54.86435, 54.00152, 53.14607, 52.29802, 51.45736, 50.62407, 49.79815, 
    48.97956, 48.16827, 47.36425, 46.56744, 45.77781, 44.99529,
  45, 45.78278, 46.57269, 47.36979, 48.17411, 48.98572, 49.80465, 50.63093, 
    51.46459, 52.30565, 53.15412, 54.01001, 54.87331, 55.744, 56.62207, 
    57.50749, 58.40021, 59.30018, 60.20734, 61.12163, 62.04295, 62.97122, 
    63.90633, 64.84815, 65.79657, 66.75144, 67.71262, 68.67992, 69.65318, 
    70.63222, 71.61682, 72.60679, 73.60188, 74.60188, 75.60651, 76.61555, 
    77.62873, 78.64574, 79.66634, 80.69019, 81.71702, 82.7465, 83.77832, 
    84.81216, 85.84769, 86.88457, 87.92248, 88.96107, 90, 88.96107, 87.92248, 
    86.88457, 85.84769, 84.81216, 83.77832, 82.7465, 81.71702, 80.69019, 
    79.66634, 78.64574, 77.62873, 76.61555, 75.60651, 74.60188, 73.60188, 
    72.60679, 71.61682, 70.63222, 69.65318, 68.67992, 67.71262, 66.75144, 
    65.79657, 64.84815, 63.90633, 62.97122, 62.04295, 61.12163, 60.20734, 
    59.30018, 58.40021, 57.50749, 56.62207, 55.744, 54.87331, 54.01001, 
    53.15412, 52.30565, 51.46459, 50.63093, 49.80465, 48.98572, 48.17411, 
    47.36979, 46.57269, 45.78278, 45,
  44.99529, 45.77781, 46.56744, 47.36425, 48.16827, 48.97956, 49.79815, 
    50.62407, 51.45736, 52.29802, 53.14607, 54.00152, 54.86435, 55.73455, 
    56.6121, 57.49697, 58.3891, 59.28845, 60.19496, 61.10854, 62.02911, 
    62.95657, 63.89082, 64.83172, 65.77914, 66.73294, 67.69295, 68.65899, 
    69.63087, 70.60838, 71.59132, 72.57942, 73.57245, 74.57011, 75.57212, 
    76.57815, 77.58782, 78.60075, 79.61646, 80.6344, 81.65389, 82.67403, 
    83.69351, 84.71027, 85.72057, 86.71655, 87.6776, 88.53089, 88.96107, 
    88.53089, 87.6776, 86.71655, 85.72057, 84.71027, 83.69351, 82.67403, 
    81.65389, 80.6344, 79.61646, 78.60075, 77.58782, 76.57815, 75.57212, 
    74.57011, 73.57245, 72.57942, 71.59132, 70.60838, 69.63087, 68.65899, 
    67.69295, 66.73294, 65.77914, 64.83172, 63.89082, 62.95657, 62.02911, 
    61.10854, 60.19496, 59.28845, 58.3891, 57.49697, 56.6121, 55.73455, 
    54.86435, 54.00152, 53.14607, 52.29802, 51.45736, 50.62407, 49.79815, 
    48.97956, 48.16827, 47.36425, 46.56744, 45.77781, 44.99529,
  44.98116, 45.7629, 46.5517, 47.34763, 48.15074, 48.96106, 49.77864, 
    50.6035, 51.43566, 52.27514, 53.12194, 53.97606, 54.8375, 55.70623, 
    56.58222, 57.46543, 58.35581, 59.2533, 60.15783, 61.06931, 61.98763, 
    62.91269, 63.84436, 64.7825, 65.72695, 66.67754, 67.63406, 68.59633, 
    69.56409, 70.53708, 71.51503, 72.49763, 73.4845, 74.47527, 75.46947, 
    76.46657, 77.46595, 78.46685, 79.46831, 80.46906, 81.46742, 82.46091, 
    83.44577, 84.41584, 85.36021, 86.25768, 87.06323, 87.6776, 87.92248, 
    87.6776, 87.06323, 86.25768, 85.36021, 84.41584, 83.44577, 82.46091, 
    81.46742, 80.46906, 79.46831, 78.46685, 77.46595, 76.46657, 75.46947, 
    74.47527, 73.4845, 72.49763, 71.51503, 70.53708, 69.56409, 68.59633, 
    67.63406, 66.67754, 65.72695, 64.7825, 63.84436, 62.91269, 61.98763, 
    61.06931, 60.15783, 59.2533, 58.35581, 57.46543, 56.58222, 55.70623, 
    54.8375, 53.97606, 53.12194, 52.27514, 51.43566, 50.6035, 49.77864, 
    48.96106, 48.15074, 47.34763, 46.5517, 45.7629, 44.98116,
  44.95763, 45.73805, 46.52548, 47.31997, 48.12155, 48.93027, 49.74615, 
    50.56924, 51.39953, 52.23703, 53.08176, 53.93369, 54.79281, 55.65909, 
    56.53249, 57.41296, 58.30043, 59.19484, 60.09608, 61.00407, 61.91867, 
    62.83975, 63.76716, 64.70073, 65.64027, 66.58555, 67.53634, 68.49236, 
    69.45333, 70.4189, 71.38868, 72.36224, 73.33907, 74.31858, 75.30009, 
    76.28278, 77.26559, 78.24726, 79.22611, 80.19992, 81.16562, 82.11877, 
    83.0528, 83.95731, 84.81542, 85.59846, 86.25768, 86.71655, 86.88457, 
    86.71655, 86.25768, 85.59846, 84.81542, 83.95731, 83.0528, 82.11877, 
    81.16562, 80.19992, 79.22611, 78.24726, 77.26559, 76.28278, 75.30009, 
    74.31858, 73.33907, 72.36224, 71.38868, 70.4189, 69.45333, 68.49236, 
    67.53634, 66.58555, 65.64027, 64.70073, 63.76716, 62.83975, 61.91867, 
    61.00407, 60.09608, 59.19484, 58.30043, 57.41296, 56.53249, 55.65909, 
    54.79281, 53.93369, 53.08176, 52.23703, 51.39953, 50.56924, 49.74615, 
    48.93027, 48.12155, 47.31997, 46.52548, 45.73805, 44.95763,
  44.9247, 45.7033, 46.4888, 47.28126, 48.08072, 48.8872, 49.70073, 50.52134, 
    51.34902, 52.18378, 53.0256, 53.87448, 54.73037, 55.59324, 56.46303, 
    57.33968, 58.22311, 59.11322, 60.00991, 60.91304, 61.82248, 62.73804, 
    63.65955, 64.58678, 65.51952, 66.45748, 67.40035, 68.3478, 69.29943, 
    70.2548, 71.21339, 72.17461, 73.13778, 74.10206, 75.06647, 76.02982, 
    76.99059, 77.94691, 78.89631, 79.83553, 80.76014, 81.66392, 82.53796, 
    83.36916, 84.13799, 84.81542, 85.36021, 85.72057, 85.84769, 85.72057, 
    85.36021, 84.81542, 84.13799, 83.36916, 82.53796, 81.66392, 80.76014, 
    79.83553, 78.89631, 77.94691, 76.99059, 76.02982, 75.06647, 74.10206, 
    73.13778, 72.17461, 71.21339, 70.2548, 69.29943, 68.3478, 67.40035, 
    66.45748, 65.51952, 64.58678, 63.65955, 62.73804, 61.82248, 60.91304, 
    60.00991, 59.11322, 58.22311, 57.33968, 56.46303, 55.59324, 54.73037, 
    53.87448, 53.0256, 52.18378, 51.34902, 50.52134, 49.70073, 48.8872, 
    48.08072, 47.28126, 46.4888, 45.7033, 44.9247,
  44.88241, 45.65865, 46.44169, 47.23156, 48.02829, 48.83191, 49.64243, 
    50.45986, 51.2842, 52.11544, 52.95356, 53.79853, 54.6503, 55.50881, 
    56.374, 57.24578, 58.12405, 59.0087, 59.89958, 60.79654, 61.6994, 
    62.60796, 63.52198, 64.4412, 65.36533, 66.29404, 67.22693, 68.16358, 
    69.10349, 70.04609, 70.99072, 71.9366, 72.88284, 73.82835, 74.77181, 
    75.71165, 76.64588, 77.572, 78.4868, 79.38612, 80.2644, 81.11414, 
    81.92511, 82.6832, 83.36916, 83.95731, 84.41584, 84.71027, 84.81216, 
    84.71027, 84.41584, 83.95731, 83.36916, 82.6832, 81.92511, 81.11414, 
    80.2644, 79.38612, 78.4868, 77.572, 76.64588, 75.71165, 74.77181, 
    73.82835, 72.88284, 71.9366, 70.99072, 70.04609, 69.10349, 68.16358, 
    67.22693, 66.29404, 65.36533, 64.4412, 63.52198, 62.60796, 61.6994, 
    60.79654, 59.89958, 59.0087, 58.12405, 57.24578, 56.374, 55.50881, 
    54.6503, 53.79853, 52.95356, 52.11544, 51.2842, 50.45986, 49.64243, 
    48.83191, 48.02829, 47.23156, 46.44169, 45.65865, 44.88241,
  44.83077, 45.60415, 46.38419, 47.17091, 47.96432, 48.76445, 49.57131, 
    50.38489, 51.20517, 52.03214, 52.86576, 53.70599, 54.55275, 55.40599, 
    56.26561, 57.13149, 58.00352, 58.88156, 59.76543, 60.65495, 61.54989, 
    62.45001, 63.35503, 64.26463, 65.17846, 66.09609, 67.01707, 67.94086, 
    68.86686, 69.79435, 70.72251, 71.6504, 72.57687, 73.50058, 74.41991, 
    75.33289, 76.23708, 77.12947, 78.00623, 78.8625, 79.69198, 80.48651, 
    81.23547, 81.92511, 82.53796, 83.0528, 83.44577, 83.69351, 83.77832, 
    83.69351, 83.44577, 83.0528, 82.53796, 81.92511, 81.23547, 80.48651, 
    79.69198, 78.8625, 78.00623, 77.12947, 76.23708, 75.33289, 74.41991, 
    73.50058, 72.57687, 71.6504, 70.72251, 69.79435, 68.86686, 67.94086, 
    67.01707, 66.09609, 65.17846, 64.26463, 63.35503, 62.45001, 61.54989, 
    60.65495, 59.76543, 58.88156, 58.00352, 57.13149, 56.26561, 55.40599, 
    54.55275, 53.70599, 52.86576, 52.03214, 51.20517, 50.38489, 49.57131, 
    48.76445, 47.96432, 47.17091, 46.38419, 45.60415, 44.83077,
  44.76982, 45.53984, 46.31635, 47.09935, 47.88887, 48.68491, 49.48746, 
    50.29652, 51.11204, 51.934, 52.76235, 53.59702, 54.43793, 55.28499, 
    56.13808, 56.99708, 57.86184, 58.73216, 59.60787, 60.48872, 61.37446, 
    62.26479, 63.15939, 64.05786, 64.95979, 65.86467, 66.77197, 67.68102, 
    68.59113, 69.50142, 70.41093, 71.31852, 72.22283, 73.12227, 74.01492, 
    74.8985, 75.77019, 76.62655, 77.46332, 78.2752, 79.05556, 79.7961, 
    80.48651, 81.11414, 81.66392, 82.11877, 82.46091, 82.67403, 82.7465, 
    82.67403, 82.46091, 82.11877, 81.66392, 81.11414, 80.48651, 79.7961, 
    79.05556, 78.2752, 77.46332, 76.62655, 75.77019, 74.8985, 74.01492, 
    73.12227, 72.22283, 71.31852, 70.41093, 69.50142, 68.59113, 67.68102, 
    66.77197, 65.86467, 64.95979, 64.05786, 63.15939, 62.26479, 61.37446, 
    60.48872, 59.60787, 58.73216, 57.86184, 56.99708, 56.13808, 55.28499, 
    54.43793, 53.59702, 52.76235, 51.934, 51.11204, 50.29652, 49.48746, 
    48.68491, 47.88887, 47.09935, 46.31635, 45.53984, 44.76982,
  44.6996, 45.46576, 46.23822, 47.01697, 47.80202, 48.59336, 49.39099, 
    50.19486, 51.00494, 51.82117, 52.64349, 53.47181, 54.30604, 55.14605, 
    55.99172, 56.84288, 57.69935, 58.56092, 59.42736, 60.29839, 61.17372, 
    62.05299, 62.93583, 63.82177, 64.71033, 65.60093, 66.49293, 67.38558, 
    68.27805, 69.16933, 70.05833, 70.9437, 71.8239, 72.69713, 73.56123, 
    74.41362, 75.25123, 76.07032, 76.86639, 77.63395, 78.36636, 79.05556, 
    79.69198, 80.2644, 80.76014, 81.16562, 81.46742, 81.65389, 81.71702, 
    81.65389, 81.46742, 81.16562, 80.76014, 80.2644, 79.69198, 79.05556, 
    78.36636, 77.63395, 76.86639, 76.07032, 75.25123, 74.41362, 73.56123, 
    72.69713, 71.8239, 70.9437, 70.05833, 69.16933, 68.27805, 67.38558, 
    66.49293, 65.60093, 64.71033, 63.82177, 62.93583, 62.05299, 61.17372, 
    60.29839, 59.42736, 58.56092, 57.69935, 56.84288, 55.99172, 55.14605, 
    54.30604, 53.47181, 52.64349, 51.82117, 51.00494, 50.19486, 49.39099, 
    48.59336, 47.80202, 47.01697, 46.23822, 45.46576, 44.6996,
  44.62016, 45.38197, 46.14986, 46.92382, 47.70385, 48.48992, 49.282, 
    50.08005, 50.88401, 51.69381, 52.50938, 53.33059, 54.15733, 54.98947, 
    55.82684, 56.66924, 57.51648, 58.36829, 59.22443, 60.08456, 60.94834, 
    61.81537, 62.6852, 63.55734, 64.4312, 65.30614, 66.18141, 67.05619, 
    67.9295, 68.80025, 69.66718, 70.52879, 71.38338, 72.22897, 73.06321, 
    73.88333, 74.68606, 75.46753, 76.22314, 76.94742, 77.63395, 78.2752, 
    78.8625, 79.38612, 79.83553, 80.19992, 80.46906, 80.6344, 80.69019, 
    80.6344, 80.46906, 80.19992, 79.83553, 79.38612, 78.8625, 78.2752, 
    77.63395, 76.94742, 76.22314, 75.46753, 74.68606, 73.88333, 73.06321, 
    72.22897, 71.38338, 70.52879, 69.66718, 68.80025, 67.9295, 67.05619, 
    66.18141, 65.30614, 64.4312, 63.55734, 62.6852, 61.81537, 60.94834, 
    60.08456, 59.22443, 58.36829, 57.51648, 56.66924, 55.82684, 54.98947, 
    54.15733, 53.33059, 52.50938, 51.69381, 50.88401, 50.08005, 49.282, 
    48.48992, 47.70385, 46.92382, 46.14986, 45.38197, 44.62016,
  44.53154, 45.28852, 46.05135, 46.82, 47.59445, 48.37467, 49.16062, 
    49.95222, 50.74942, 51.55212, 52.36022, 53.17359, 53.99209, 54.81555, 
    55.64378, 56.47657, 57.31367, 58.1548, 58.99965, 59.84786, 60.69904, 
    61.55275, 62.40846, 63.26563, 64.1236, 64.98164, 65.83895, 66.69459, 
    67.54749, 68.39644, 69.24005, 70.07672, 70.90462, 71.7216, 72.5252, 
    73.31252, 74.08022, 74.82438, 75.54044, 76.22314, 76.86639, 77.46332, 
    78.00623, 78.4868, 78.89631, 79.22611, 79.46831, 79.61646, 79.66634, 
    79.61646, 79.46831, 79.22611, 78.89631, 78.4868, 78.00623, 77.46332, 
    76.86639, 76.22314, 75.54044, 74.82438, 74.08022, 73.31252, 72.5252, 
    71.7216, 70.90462, 70.07672, 69.24005, 68.39644, 67.54749, 66.69459, 
    65.83895, 64.98164, 64.1236, 63.26563, 62.40846, 61.55275, 60.69904, 
    59.84786, 58.99965, 58.1548, 57.31367, 56.47657, 55.64378, 54.81555, 
    53.99209, 53.17359, 52.36022, 51.55212, 50.74942, 49.95222, 49.16062, 
    48.37467, 47.59445, 46.82, 46.05135, 45.28852, 44.53154,
  44.4338, 45.18549, 45.94276, 46.70559, 47.47393, 48.24775, 49.02699, 
    49.81155, 50.60136, 51.39631, 52.19627, 53.00109, 53.81061, 54.62463, 
    55.44294, 56.26529, 57.09141, 57.92097, 58.75364, 59.589, 60.42662, 
    61.26601, 62.10659, 62.94775, 63.78878, 64.62888, 65.46716, 66.30258, 
    67.13403, 67.96017, 68.77954, 69.59042, 70.39089, 71.17871, 71.95134, 
    72.70583, 73.43884, 74.14648, 74.82438, 75.46753, 76.07032, 76.62655, 
    77.12947, 77.572, 77.94691, 78.24726, 78.46685, 78.60075, 78.64574, 
    78.60075, 78.46685, 78.24726, 77.94691, 77.572, 77.12947, 76.62655, 
    76.07032, 75.46753, 74.82438, 74.14648, 73.43884, 72.70583, 71.95134, 
    71.17871, 70.39089, 69.59042, 68.77954, 67.96017, 67.13403, 66.30258, 
    65.46716, 64.62888, 63.78878, 62.94775, 62.10659, 61.26601, 60.42662, 
    59.589, 58.75364, 57.92097, 57.09141, 56.26529, 55.44294, 54.62463, 
    53.81061, 53.00109, 52.19627, 51.39631, 50.60136, 49.81155, 49.02699, 
    48.24775, 47.47393, 46.70559, 45.94276, 45.18549, 44.4338,
  44.32701, 45.07294, 45.82418, 46.58068, 47.34241, 48.10929, 48.88126, 
    49.6582, 50.44002, 51.22659, 52.01776, 52.81337, 53.61321, 54.41708, 
    55.22473, 56.03588, 56.85022, 57.66741, 58.48705, 59.30871, 60.1319, 
    60.95608, 61.78063, 62.60488, 63.42805, 64.2493, 65.06765, 65.88202, 
    66.69118, 67.49377, 68.28822, 69.07276, 69.84539, 70.60384, 71.34553, 
    72.06753, 72.76654, 73.43884, 74.08022, 74.68606, 75.25123, 75.77019, 
    76.23708, 76.64588, 76.99059, 77.26559, 77.46595, 77.58782, 77.62873, 
    77.58782, 77.46595, 77.26559, 76.99059, 76.64588, 76.23708, 75.77019, 
    75.25123, 74.68606, 74.08022, 73.43884, 72.76654, 72.06753, 71.34553, 
    70.60384, 69.84539, 69.07276, 68.28822, 67.49377, 66.69118, 65.88202, 
    65.06765, 64.2493, 63.42805, 62.60488, 61.78063, 60.95608, 60.1319, 
    59.30871, 58.48705, 57.66741, 56.85022, 56.03588, 55.22473, 54.41708, 
    53.61321, 52.81337, 52.01776, 51.22659, 50.44002, 49.6582, 48.88126, 
    48.10929, 47.34241, 46.58068, 45.82418, 45.07294, 44.32701,
  44.21122, 44.95095, 45.6957, 46.4454, 47.20001, 47.95944, 48.72359, 
    49.49236, 50.26561, 51.04321, 51.82498, 52.61073, 53.40025, 54.19329, 
    54.98958, 55.78882, 56.59066, 57.39472, 58.20058, 59.00777, 59.81574, 
    60.62392, 61.43166, 62.2382, 63.04275, 63.84439, 64.6421, 65.43473, 
    66.22101, 66.9995, 67.76861, 68.5265, 69.27117, 70.00032, 70.7114, 
    71.40154, 72.06753, 72.70583, 73.31252, 73.88333, 74.41362, 74.8985, 
    75.33289, 75.71165, 76.02982, 76.28278, 76.46657, 76.57815, 76.61555, 
    76.57815, 76.46657, 76.28278, 76.02982, 75.71165, 75.33289, 74.8985, 
    74.41362, 73.88333, 73.31252, 72.70583, 72.06753, 71.40154, 70.7114, 
    70.00032, 69.27117, 68.5265, 67.76861, 66.9995, 66.22101, 65.43473, 
    64.6421, 63.84439, 63.04275, 62.2382, 61.43166, 60.62392, 59.81574, 
    59.00777, 58.20058, 57.39472, 56.59066, 55.78882, 54.98958, 54.19329, 
    53.40025, 52.61073, 51.82498, 51.04321, 50.26561, 49.49236, 48.72359, 
    47.95944, 47.20001, 46.4454, 45.6957, 44.95095, 44.21122,
  44.08652, 44.81961, 45.55742, 46.29986, 47.04686, 47.79833, 48.55416, 
    49.31422, 50.07836, 50.84642, 51.6182, 52.39351, 53.17208, 53.95366, 
    54.73795, 55.52462, 56.31329, 57.10355, 57.89494, 58.68696, 59.47903, 
    60.27053, 61.06076, 61.84895, 62.63423, 63.41565, 64.19215, 64.96255, 
    65.72551, 66.47958, 67.22313, 67.95432, 68.67112, 69.37128, 70.0523, 
    70.7114, 71.34553, 71.95134, 72.5252, 73.06321, 73.56123, 74.01492, 
    74.41991, 74.77181, 75.06647, 75.30009, 75.46947, 75.57212, 75.60651, 
    75.57212, 75.46947, 75.30009, 75.06647, 74.77181, 74.41991, 74.01492, 
    73.56123, 73.06321, 72.5252, 71.95134, 71.34553, 70.7114, 70.0523, 
    69.37128, 68.67112, 67.95432, 67.22313, 66.47958, 65.72551, 64.96255, 
    64.19215, 63.41565, 62.63423, 61.84895, 61.06076, 60.27053, 59.47903, 
    58.68696, 57.89494, 57.10355, 56.31329, 55.52462, 54.73795, 53.95366, 
    53.17208, 52.39351, 51.6182, 50.84642, 50.07836, 49.31422, 48.55416, 
    47.79833, 47.04686, 46.29986, 45.55742, 44.81961, 44.08652,
  43.95298, 44.67902, 45.40944, 46.14417, 46.8831, 47.62614, 48.37315, 
    49.124, 49.8785, 50.63649, 51.39774, 52.16203, 52.92909, 53.69863, 
    54.47033, 55.24382, 56.01871, 56.79456, 57.57087, 58.34711, 59.12267, 
    59.89689, 60.66905, 61.43833, 62.20383, 62.96457, 63.71946, 64.46726, 
    65.20666, 65.93615, 66.65411, 67.3587, 68.04794, 68.7196, 69.37128, 
    70.00032, 70.60384, 71.17871, 71.7216, 72.22897, 72.69713, 73.12227, 
    73.50058, 73.82835, 74.10206, 74.31858, 74.47527, 74.57011, 74.60188, 
    74.57011, 74.47527, 74.31858, 74.10206, 73.82835, 73.50058, 73.12227, 
    72.69713, 72.22897, 71.7216, 71.17871, 70.60384, 70.00032, 69.37128, 
    68.7196, 68.04794, 67.3587, 66.65411, 65.93615, 65.20666, 64.46726, 
    63.71946, 62.96457, 62.20383, 61.43833, 60.66905, 59.89689, 59.12267, 
    58.34711, 57.57087, 56.79456, 56.01871, 55.24382, 54.47033, 53.69863, 
    52.92909, 52.16203, 51.39774, 50.63649, 49.8785, 49.124, 48.37315, 
    47.62614, 46.8831, 46.14417, 45.40944, 44.67902, 43.95298,
  43.81068, 44.52925, 45.25187, 45.97845, 46.70888, 47.44304, 48.18076, 
    48.92191, 49.66629, 50.4137, 51.1639, 51.91666, 52.67167, 53.42863, 
    54.18719, 54.94697, 55.70753, 56.46842, 57.22911, 57.98904, 58.74758, 
    59.50403, 60.25764, 61.00757, 61.7529, 62.49262, 63.2256, 63.95062, 
    64.66634, 65.37125, 66.06374, 66.74202, 67.40413, 68.04794, 68.67112, 
    69.27117, 69.84539, 70.39089, 70.90462, 71.38338, 71.8239, 72.22283, 
    72.57687, 72.88284, 73.13778, 73.33907, 73.4845, 73.57245, 73.60188, 
    73.57245, 73.4845, 73.33907, 73.13778, 72.88284, 72.57687, 72.22283, 
    71.8239, 71.38338, 70.90462, 70.39089, 69.84539, 69.27117, 68.67112, 
    68.04794, 67.40413, 66.74202, 66.06374, 65.37125, 64.66634, 63.95062, 
    63.2256, 62.49262, 61.7529, 61.00757, 60.25764, 59.50403, 58.74758, 
    57.98904, 57.22911, 56.46842, 55.70753, 54.94697, 54.18719, 53.42863, 
    52.67167, 51.91666, 51.1639, 50.4137, 49.66629, 48.92191, 48.18076, 
    47.44304, 46.70888, 45.97845, 45.25187, 44.52925, 43.81068,
  43.65969, 44.37041, 45.08484, 45.80286, 46.52436, 47.24918, 47.97718, 
    48.70818, 49.44197, 50.17833, 50.91702, 51.65775, 52.40023, 53.14412, 
    53.88906, 54.63462, 55.38037, 56.12582, 56.87043, 57.61359, 58.35467, 
    59.09295, 59.82764, 60.55789, 61.28276, 62.00122, 62.71215, 63.41431, 
    64.10636, 64.78683, 65.45412, 66.10648, 66.74202, 67.3587, 67.95432, 
    68.5265, 69.07276, 69.59042, 70.07672, 70.52879, 70.9437, 71.31852, 
    71.6504, 71.9366, 72.17461, 72.36224, 72.49763, 72.57942, 72.60679, 
    72.57942, 72.49763, 72.36224, 72.17461, 71.9366, 71.6504, 71.31852, 
    70.9437, 70.52879, 70.07672, 69.59042, 69.07276, 68.5265, 67.95432, 
    67.3587, 66.74202, 66.10648, 65.45412, 64.78683, 64.10636, 63.41431, 
    62.71215, 62.00122, 61.28276, 60.55789, 59.82764, 59.09295, 58.35467, 
    57.61359, 56.87043, 56.12582, 55.38037, 54.63462, 53.88906, 53.14412, 
    52.40023, 51.65775, 50.91702, 50.17833, 49.44197, 48.70818, 47.97718, 
    47.24918, 46.52436, 45.80286, 45.08484, 44.37041, 43.65969,
  43.50012, 44.20261, 44.90845, 45.61752, 46.32969, 47.04478, 47.76263, 
    48.48305, 49.20582, 49.9307, 50.65742, 51.38569, 52.11519, 52.84557, 
    53.57643, 54.30735, 55.03786, 55.76746, 56.49557, 57.2216, 57.94487, 
    58.66464, 59.38013, 60.09047, 60.79469, 61.49178, 62.18061, 62.85994, 
    63.52847, 64.18473, 64.82718, 65.45412, 66.06374, 66.65411, 67.22313, 
    67.76861, 68.28822, 68.77954, 69.24005, 69.66718, 70.05833, 70.41093, 
    70.72251, 70.99072, 71.21339, 71.38868, 71.51503, 71.59132, 71.61682, 
    71.59132, 71.51503, 71.38868, 71.21339, 70.99072, 70.72251, 70.41093, 
    70.05833, 69.66718, 69.24005, 68.77954, 68.28822, 67.76861, 67.22313, 
    66.65411, 66.06374, 65.45412, 64.82718, 64.18473, 63.52847, 62.85994, 
    62.18061, 61.49178, 60.79469, 60.09047, 59.38013, 58.66464, 57.94487, 
    57.2216, 56.49557, 55.76746, 55.03786, 54.30735, 53.57643, 52.84557, 
    52.11519, 51.38569, 50.65742, 49.9307, 49.20582, 48.48305, 47.76263, 
    47.04478, 46.32969, 45.61752, 44.90845, 44.20261, 43.50012,
  43.33206, 44.02596, 44.72285, 45.42259, 46.12503, 46.83001, 47.53732, 
    48.24677, 48.95811, 49.6711, 50.38545, 51.10085, 51.81697, 52.53343, 
    53.24984, 53.96573, 54.68064, 55.39402, 56.10532, 56.8139, 57.51908, 
    58.22011, 58.9162, 59.60646, 60.28995, 60.96564, 61.63241, 62.28906, 
    62.93428, 63.56667, 64.18473, 64.78683, 65.37125, 65.93615, 66.47958, 
    66.9995, 67.49377, 67.96017, 68.39644, 68.80025, 69.16933, 69.50142, 
    69.79435, 70.04609, 70.2548, 70.4189, 70.53708, 70.60838, 70.63222, 
    70.60838, 70.53708, 70.4189, 70.2548, 70.04609, 69.79435, 69.50142, 
    69.16933, 68.80025, 68.39644, 67.96017, 67.49377, 66.9995, 66.47958, 
    65.93615, 65.37125, 64.78683, 64.18473, 63.56667, 62.93428, 62.28906, 
    61.63241, 60.96564, 60.28995, 59.60646, 58.9162, 58.22011, 57.51908, 
    56.8139, 56.10532, 55.39402, 54.68064, 53.96573, 53.24984, 52.53343, 
    51.81697, 51.10085, 50.38545, 49.6711, 48.95811, 48.24677, 47.53732, 
    46.83001, 46.12503, 45.42259, 44.72285, 44.02596, 43.33206,
  43.1556, 43.84056, 44.52815, 45.21821, 45.91058, 46.60506, 47.30147, 
    47.99957, 48.69912, 49.39985, 50.10146, 50.80363, 51.506, 52.2082, 
    52.9098, 53.61034, 54.30932, 55.00621, 55.70042, 56.39131, 57.07819, 
    57.76032, 58.43688, 59.10701, 59.76975, 60.4241, 61.06895, 61.70312, 
    62.32535, 62.93428, 63.52847, 64.10636, 64.66634, 65.20666, 65.72551, 
    66.22101, 66.69118, 67.13403, 67.54749, 67.9295, 68.27805, 68.59113, 
    68.86686, 69.10349, 69.29943, 69.45333, 69.56409, 69.63087, 69.65318, 
    69.63087, 69.56409, 69.45333, 69.29943, 69.10349, 68.86686, 68.59113, 
    68.27805, 67.9295, 67.54749, 67.13403, 66.69118, 66.22101, 65.72551, 
    65.20666, 64.66634, 64.10636, 63.52847, 62.93428, 62.32535, 61.70312, 
    61.06895, 60.4241, 59.76975, 59.10701, 58.43688, 57.76032, 57.07819, 
    56.39131, 55.70042, 55.00621, 54.30932, 53.61034, 52.9098, 52.2082, 
    51.506, 50.80363, 50.10146, 49.39985, 48.69912, 47.99957, 47.30147, 
    46.60506, 45.91058, 45.21821, 44.52815, 43.84056, 43.1556,
  42.97084, 43.64655, 44.3245, 45.00454, 45.68649, 46.37015, 47.05531, 
    47.74172, 48.42913, 49.11726, 49.8058, 50.49441, 51.18272, 51.87035, 
    52.55685, 53.24175, 53.92455, 54.60471, 55.28162, 55.95465, 56.62309, 
    57.28621, 57.9432, 58.59319, 59.23526, 59.86839, 60.49152, 61.1035, 
    61.70312, 62.28906, 62.85994, 63.41431, 63.95062, 64.46726, 64.96255, 
    65.43473, 65.88202, 66.30258, 66.69459, 67.05619, 67.38558, 67.68102, 
    67.94086, 68.16358, 68.3478, 68.49236, 68.59633, 68.65899, 68.67992, 
    68.65899, 68.59633, 68.49236, 68.3478, 68.16358, 67.94086, 67.68102, 
    67.38558, 67.05619, 66.69459, 66.30258, 65.88202, 65.43473, 64.96255, 
    64.46726, 63.95062, 63.41431, 62.85994, 62.28906, 61.70312, 61.1035, 
    60.49152, 59.86839, 59.23526, 58.59319, 57.9432, 57.28621, 56.62309, 
    55.95465, 55.28162, 54.60471, 53.92455, 53.24175, 52.55685, 51.87035, 
    51.18272, 50.49441, 49.8058, 49.11726, 48.42913, 47.74172, 47.05531, 
    46.37015, 45.68649, 45.00454, 44.3245, 43.64655, 42.97084,
  42.77788, 43.44402, 44.11203, 44.78174, 45.45296, 46.12547, 46.79906, 
    47.47348, 48.14844, 48.82367, 49.49884, 50.1736, 50.84757, 51.52035, 
    52.1915, 52.86054, 53.52696, 54.1902, 54.84966, 55.50471, 56.15464, 
    56.79872, 57.43615, 58.06607, 58.68758, 59.2997, 59.90138, 60.49152, 
    61.06895, 61.63241, 62.18061, 62.71215, 63.2256, 63.71946, 64.19215, 
    64.6421, 65.06765, 65.46716, 65.83895, 66.18141, 66.49293, 66.77197, 
    67.01707, 67.22693, 67.40035, 67.53634, 67.63406, 67.69295, 67.71262, 
    67.69295, 67.63406, 67.53634, 67.40035, 67.22693, 67.01707, 66.77197, 
    66.49293, 66.18141, 65.83895, 65.46716, 65.06765, 64.6421, 64.19215, 
    63.71946, 63.2256, 62.71215, 62.18061, 61.63241, 61.06895, 60.49152, 
    59.90138, 59.2997, 58.68758, 58.06607, 57.43615, 56.79872, 56.15464, 
    55.50471, 54.84966, 54.1902, 53.52696, 52.86054, 52.1915, 51.52035, 
    50.84757, 50.1736, 49.49884, 48.82367, 48.14844, 47.47348, 46.79906, 
    46.12547, 45.45296, 44.78174, 44.11203, 43.44402, 42.77788,
  42.57683, 43.23311, 43.89089, 44.54997, 45.21016, 45.87124, 46.53297, 
    47.1951, 47.85734, 48.51939, 49.18093, 49.84158, 50.50098, 51.1587, 
    51.8143, 52.46729, 53.11716, 53.76335, 54.40527, 55.04227, 55.67367, 
    56.29873, 56.91667, 57.52666, 58.1278, 58.71915, 59.2997, 59.86839, 
    60.4241, 60.96564, 61.49178, 62.00122, 62.49262, 62.96457, 63.41565, 
    63.84439, 64.2493, 64.62888, 64.98164, 65.30614, 65.60093, 65.86467, 
    66.09609, 66.29404, 66.45748, 66.58555, 66.67754, 66.73294, 66.75144, 
    66.73294, 66.67754, 66.58555, 66.45748, 66.29404, 66.09609, 65.86467, 
    65.60093, 65.30614, 64.98164, 64.62888, 64.2493, 63.84439, 63.41565, 
    62.96457, 62.49262, 62.00122, 61.49178, 60.96564, 60.4241, 59.86839, 
    59.2997, 58.71915, 58.1278, 57.52666, 56.91667, 56.29873, 55.67367, 
    55.04227, 54.40527, 53.76335, 53.11716, 52.46729, 51.8143, 51.1587, 
    50.50098, 49.84158, 49.18093, 48.51939, 47.85734, 47.1951, 46.53297, 
    45.87124, 45.21016, 44.54997, 43.89089, 43.23311, 42.57683,
  42.36781, 43.01395, 43.66121, 44.30939, 44.95829, 45.60766, 46.25727, 
    46.90686, 47.55613, 48.20476, 48.85243, 49.49877, 50.14338, 50.78586, 
    51.42574, 52.06255, 52.69576, 53.32483, 53.94915, 54.5681, 55.18099, 
    55.78711, 56.38568, 56.97591, 57.55692, 58.1278, 58.68758, 59.23526, 
    59.76975, 60.28995, 60.79469, 61.28276, 61.7529, 62.20383, 62.63423, 
    63.04275, 63.42805, 63.78878, 64.1236, 64.4312, 64.71033, 64.95979, 
    65.17846, 65.36533, 65.51952, 65.64027, 65.72695, 65.77914, 65.79657, 
    65.77914, 65.72695, 65.64027, 65.51952, 65.36533, 65.17846, 64.95979, 
    64.71033, 64.4312, 64.1236, 63.78878, 63.42805, 63.04275, 62.63423, 
    62.20383, 61.7529, 61.28276, 60.79469, 60.28995, 59.76975, 59.23526, 
    58.68758, 58.1278, 57.55692, 56.97591, 56.38568, 55.78711, 55.18099, 
    54.5681, 53.94915, 53.32483, 52.69576, 52.06255, 51.42574, 50.78586, 
    50.14338, 49.49877, 48.85243, 48.20476, 47.55613, 46.90686, 46.25727, 
    45.60766, 44.95829, 44.30939, 43.66121, 43.01395, 42.36781,
  42.15091, 42.78666, 43.42315, 44.06018, 44.69753, 45.33495, 45.97221, 
    46.60902, 47.24509, 47.8801, 48.51371, 49.14555, 49.77522, 50.40231, 
    51.02636, 51.64688, 52.26337, 52.87527, 53.48199, 54.08292, 54.67738, 
    55.26468, 55.84407, 56.41476, 56.97591, 57.52666, 58.06607, 58.59319, 
    59.10701, 59.60646, 60.09047, 60.55789, 61.00757, 61.43833, 61.84895, 
    62.2382, 62.60488, 62.94775, 63.26563, 63.55734, 63.82177, 64.05786, 
    64.26463, 64.4412, 64.58678, 64.70073, 64.7825, 64.83172, 64.84815, 
    64.83172, 64.7825, 64.70073, 64.58678, 64.4412, 64.26463, 64.05786, 
    63.82177, 63.55734, 63.26563, 62.94775, 62.60488, 62.2382, 61.84895, 
    61.43833, 61.00757, 60.55789, 60.09047, 59.60646, 59.10701, 58.59319, 
    58.06607, 57.52666, 56.97591, 56.41476, 55.84407, 55.26468, 54.67738, 
    54.08292, 53.48199, 52.87527, 52.26337, 51.64688, 51.02636, 50.40231, 
    49.77522, 49.14555, 48.51371, 47.8801, 47.24509, 46.60902, 45.97221, 
    45.33495, 44.69753, 44.06018, 43.42315, 42.78666, 42.15091,
  41.92625, 42.55138, 43.17686, 43.8025, 44.42807, 45.05334, 45.67802, 
    46.30186, 46.92454, 47.54575, 48.16513, 48.78232, 49.39692, 50.00851, 
    50.61664, 51.22083, 51.82056, 52.4153, 53.00447, 53.58745, 54.16361, 
    54.73225, 55.29266, 55.84407, 56.38568, 56.91667, 57.43615, 57.9432, 
    58.43688, 58.9162, 59.38013, 59.82764, 60.25764, 60.66905, 61.06076, 
    61.43166, 61.78063, 62.10659, 62.40846, 62.6852, 62.93583, 63.15939, 
    63.35503, 63.52198, 63.65955, 63.76716, 63.84436, 63.89082, 63.90633, 
    63.89082, 63.84436, 63.76716, 63.65955, 63.52198, 63.35503, 63.15939, 
    62.93583, 62.6852, 62.40846, 62.10659, 61.78063, 61.43166, 61.06076, 
    60.66905, 60.25764, 59.82764, 59.38013, 58.9162, 58.43688, 57.9432, 
    57.43615, 56.91667, 56.38568, 55.84407, 55.29266, 54.73225, 54.16361, 
    53.58745, 53.00447, 52.4153, 51.82056, 51.22083, 50.61664, 50.00851, 
    49.39692, 48.78232, 48.16513, 47.54575, 46.92454, 46.30186, 45.67802, 
    45.05334, 44.42807, 43.8025, 43.17686, 42.55138, 41.92625,
  41.69396, 42.30823, 42.92249, 43.53653, 44.15013, 44.76302, 45.37495, 
    45.98564, 46.59477, 47.20202, 47.80704, 48.40947, 49.00891, 49.60493, 
    50.19709, 50.78492, 51.36792, 51.94554, 52.51723, 53.08239, 53.64039, 
    54.19058, 54.73225, 55.26468, 55.78711, 56.29873, 56.79872, 57.28621, 
    57.76032, 58.22011, 58.66464, 59.09295, 59.50403, 59.89689, 60.27053, 
    60.62392, 60.95608, 61.26601, 61.55275, 61.81537, 62.05299, 62.26479, 
    62.45001, 62.60796, 62.73804, 62.83975, 62.91269, 62.95657, 62.97122, 
    62.95657, 62.91269, 62.83975, 62.73804, 62.60796, 62.45001, 62.26479, 
    62.05299, 61.81537, 61.55275, 61.26601, 60.95608, 60.62392, 60.27053, 
    59.89689, 59.50403, 59.09295, 58.66464, 58.22011, 57.76032, 57.28621, 
    56.79872, 56.29873, 55.78711, 55.26468, 54.73225, 54.19058, 53.64039, 
    53.08239, 52.51723, 51.94554, 51.36792, 50.78492, 50.19709, 49.60493, 
    49.00891, 48.40947, 47.80704, 47.20202, 46.59477, 45.98564, 45.37495, 
    44.76302, 44.15013, 43.53653, 42.92249, 42.30823, 41.69396,
  41.45414, 42.05735, 42.66019, 43.26245, 43.86388, 44.46423, 45.06325, 
    45.66063, 46.25607, 46.84925, 47.43981, 48.02739, 48.6116, 49.19202, 
    49.7682, 50.33969, 50.90599, 51.46657, 52.0209, 52.56838, 53.10843, 
    53.64039, 54.16361, 54.67738, 55.18099, 55.67367, 56.15464, 56.62309, 
    57.07819, 57.51908, 57.94487, 58.35467, 58.74758, 59.12267, 59.47903, 
    59.81574, 60.1319, 60.42662, 60.69904, 60.94834, 61.17372, 61.37446, 
    61.54989, 61.6994, 61.82248, 61.91867, 61.98763, 62.02911, 62.04295, 
    62.02911, 61.98763, 61.91867, 61.82248, 61.6994, 61.54989, 61.37446, 
    61.17372, 60.94834, 60.69904, 60.42662, 60.1319, 59.81574, 59.47903, 
    59.12267, 58.74758, 58.35467, 57.94487, 57.51908, 57.07819, 56.62309, 
    56.15464, 55.67367, 55.18099, 54.67738, 54.16361, 53.64039, 53.10843, 
    52.56838, 52.0209, 51.46657, 50.90599, 50.33969, 49.7682, 49.19202, 
    48.6116, 48.02739, 47.43981, 46.84925, 46.25607, 45.66063, 45.06325, 
    44.46423, 43.86388, 43.26245, 42.66019, 42.05735, 41.45414,
  41.20691, 41.79888, 42.39012, 42.98042, 43.56952, 44.15719, 44.74314, 
    45.3271, 45.90874, 46.48775, 47.06378, 47.63646, 48.20541, 48.77021, 
    49.33044, 49.88563, 50.43531, 50.97897, 51.51608, 52.04608, 52.56838, 
    53.08239, 53.58745, 54.08292, 54.5681, 55.04227, 55.50471, 55.95465, 
    56.39131, 56.8139, 57.2216, 57.61359, 57.98904, 58.34711, 58.68696, 
    59.00777, 59.30871, 59.589, 59.84786, 60.08456, 60.29839, 60.48872, 
    60.65495, 60.79654, 60.91304, 61.00407, 61.06931, 61.10854, 61.12163, 
    61.10854, 61.06931, 61.00407, 60.91304, 60.79654, 60.65495, 60.48872, 
    60.29839, 60.08456, 59.84786, 59.589, 59.30871, 59.00777, 58.68696, 
    58.34711, 57.98904, 57.61359, 57.2216, 56.8139, 56.39131, 55.95465, 
    55.50471, 55.04227, 54.5681, 54.08292, 53.58745, 53.08239, 52.56838, 
    52.04608, 51.51608, 50.97897, 50.43531, 49.88563, 49.33044, 48.77021, 
    48.20541, 47.63646, 47.06378, 46.48775, 45.90874, 45.3271, 44.74314, 
    44.15719, 43.56952, 42.98042, 42.39012, 41.79888, 41.20691,
  40.9524, 41.53295, 42.11243, 42.69062, 43.26726, 43.84211, 44.41489, 
    44.98531, 45.55307, 46.11785, 46.67929, 47.23705, 47.79074, 48.33995, 
    48.88427, 49.42325, 49.95642, 50.48329, 51.00336, 51.51608, 52.0209, 
    52.51723, 53.00447, 53.48199, 53.94915, 54.40527, 54.84966, 55.28162, 
    55.70042, 56.10532, 56.49557, 56.87043, 57.22911, 57.57087, 57.89494, 
    58.20058, 58.48705, 58.75364, 58.99965, 59.22443, 59.42736, 59.60787, 
    59.76543, 59.89958, 60.00991, 60.09608, 60.15783, 60.19496, 60.20734, 
    60.19496, 60.15783, 60.09608, 60.00991, 59.89958, 59.76543, 59.60787, 
    59.42736, 59.22443, 58.99965, 58.75364, 58.48705, 58.20058, 57.89494, 
    57.57087, 57.22911, 56.87043, 56.49557, 56.10532, 55.70042, 55.28162, 
    54.84966, 54.40527, 53.94915, 53.48199, 53.00447, 52.51723, 52.0209, 
    51.51608, 51.00336, 50.48329, 49.95642, 49.42325, 48.88427, 48.33995, 
    47.79074, 47.23705, 46.67929, 46.11785, 45.55307, 44.98531, 44.41489, 
    43.84211, 43.26726, 42.69062, 42.11243, 41.53295, 40.9524,
  40.69072, 41.25971, 41.82729, 42.39323, 42.95729, 43.51921, 44.07872, 
    44.63554, 45.18936, 45.73986, 46.28671, 46.82954, 47.36799, 47.90166, 
    48.43015, 48.95301, 49.46981, 49.98007, 50.48329, 50.97897, 51.46657, 
    51.94554, 52.4153, 52.87527, 53.32483, 53.76335, 54.1902, 54.60471, 
    55.00621, 55.39402, 55.76746, 56.12582, 56.46842, 56.79456, 57.10355, 
    57.39472, 57.66741, 57.92097, 58.1548, 58.36829, 58.56092, 58.73216, 
    58.88156, 59.0087, 59.11322, 59.19484, 59.2533, 59.28845, 59.30018, 
    59.28845, 59.2533, 59.19484, 59.11322, 59.0087, 58.88156, 58.73216, 
    58.56092, 58.36829, 58.1548, 57.92097, 57.66741, 57.39472, 57.10355, 
    56.79456, 56.46842, 56.12582, 55.76746, 55.39402, 55.00621, 54.60471, 
    54.1902, 53.76335, 53.32483, 52.87527, 52.4153, 51.94554, 51.46657, 
    50.97897, 50.48329, 49.98007, 49.46981, 48.95301, 48.43015, 47.90166, 
    47.36799, 46.82954, 46.28671, 45.73986, 45.18936, 44.63554, 44.07872, 
    43.51921, 42.95729, 42.39323, 41.82729, 41.25971, 40.69072,
  40.42199, 40.97929, 41.53484, 42.08843, 42.6398, 43.18871, 43.73489, 
    44.27805, 44.81789, 45.35409, 45.88634, 46.41428, 46.93754, 47.45575, 
    47.96851, 48.4754, 48.97598, 49.46981, 49.95642, 50.43531, 50.90599, 
    51.36792, 51.82056, 52.26337, 52.69576, 53.11716, 53.52696, 53.92455, 
    54.30932, 54.68064, 55.03786, 55.38037, 55.70753, 56.01871, 56.31329, 
    56.59066, 56.85022, 57.09141, 57.31367, 57.51648, 57.69935, 57.86184, 
    58.00352, 58.12405, 58.22311, 58.30043, 58.35581, 58.3891, 58.40021, 
    58.3891, 58.35581, 58.30043, 58.22311, 58.12405, 58.00352, 57.86184, 
    57.69935, 57.51648, 57.31367, 57.09141, 56.85022, 56.59066, 56.31329, 
    56.01871, 55.70753, 55.38037, 55.03786, 54.68064, 54.30932, 53.92455, 
    53.52696, 53.11716, 52.69576, 52.26337, 51.82056, 51.36792, 50.90599, 
    50.43531, 49.95642, 49.46981, 48.97598, 48.4754, 47.96851, 47.45575, 
    46.93754, 46.41428, 45.88634, 45.35409, 44.81789, 44.27805, 43.73489, 
    43.18871, 42.6398, 42.08843, 41.53484, 40.97929, 40.42199,
  40.14635, 40.69183, 41.23525, 41.77639, 42.315, 42.85083, 43.38362, 
    43.91308, 44.43893, 44.96085, 45.47853, 45.99162, 46.49977, 47.00262, 
    47.49977, 47.99084, 48.4754, 48.95301, 49.42325, 49.88563, 50.33969, 
    50.78492, 51.22083, 51.64688, 52.06255, 52.46729, 52.86054, 53.24175, 
    53.61034, 53.96573, 54.30735, 54.63462, 54.94697, 55.24382, 55.52462, 
    55.78882, 56.03588, 56.26529, 56.47657, 56.66924, 56.84288, 56.99708, 
    57.13149, 57.24578, 57.33968, 57.41296, 57.46543, 57.49697, 57.50749, 
    57.49697, 57.46543, 57.41296, 57.33968, 57.24578, 57.13149, 56.99708, 
    56.84288, 56.66924, 56.47657, 56.26529, 56.03588, 55.78882, 55.52462, 
    55.24382, 54.94697, 54.63462, 54.30735, 53.96573, 53.61034, 53.24175, 
    52.86054, 52.46729, 52.06255, 51.64688, 51.22083, 50.78492, 50.33969, 
    49.88563, 49.42325, 48.95301, 48.4754, 47.99084, 47.49977, 47.00262, 
    46.49977, 45.99162, 45.47853, 44.96085, 44.43893, 43.91308, 43.38362, 
    42.85083, 42.315, 41.77639, 41.23525, 40.69183, 40.14635,
  39.8639, 40.39747, 40.92867, 41.45728, 41.98307, 42.50578, 43.02515, 
    43.54091, 44.05278, 44.56044, 45.0636, 45.56192, 46.05505, 46.54266, 
    47.02436, 47.49977, 47.96851, 48.43015, 48.88427, 49.33044, 49.7682, 
    50.19709, 50.61664, 51.02636, 51.42574, 51.8143, 52.1915, 52.55685, 
    52.9098, 53.24984, 53.57643, 53.88906, 54.18719, 54.47033, 54.73795, 
    54.98958, 55.22473, 55.44294, 55.64378, 55.82684, 55.99172, 56.13808, 
    56.26561, 56.374, 56.46303, 56.53249, 56.58222, 56.6121, 56.62207, 
    56.6121, 56.58222, 56.53249, 56.46303, 56.374, 56.26561, 56.13808, 
    55.99172, 55.82684, 55.64378, 55.44294, 55.22473, 54.98958, 54.73795, 
    54.47033, 54.18719, 53.88906, 53.57643, 53.24984, 52.9098, 52.55685, 
    52.1915, 51.8143, 51.42574, 51.02636, 50.61664, 50.19709, 49.7682, 
    49.33044, 48.88427, 48.43015, 47.96851, 47.49977, 47.02436, 46.54266, 
    46.05505, 45.56192, 45.0636, 44.56044, 44.05278, 43.54091, 43.02515, 
    42.50578, 41.98307, 41.45728, 40.92867, 40.39747, 39.8639,
  39.57478, 40.09635, 40.61526, 41.13129, 41.64421, 42.15377, 42.65972, 
    43.16179, 43.6597, 44.15316, 44.64186, 45.1255, 45.60374, 46.07624, 
    46.54266, 47.00262, 47.45575, 47.90166, 48.33995, 48.77021, 49.19202, 
    49.60493, 50.00851, 50.40231, 50.78586, 51.1587, 51.52035, 51.87035, 
    52.2082, 52.53343, 52.84557, 53.14412, 53.42863, 53.69863, 53.95366, 
    54.19329, 54.41708, 54.62463, 54.81555, 54.98947, 55.14605, 55.28499, 
    55.40599, 55.50881, 55.59324, 55.65909, 55.70623, 55.73455, 55.744, 
    55.73455, 55.70623, 55.65909, 55.59324, 55.50881, 55.40599, 55.28499, 
    55.14605, 54.98947, 54.81555, 54.62463, 54.41708, 54.19329, 53.95366, 
    53.69863, 53.42863, 53.14412, 52.84557, 52.53343, 52.2082, 51.87035, 
    51.52035, 51.1587, 50.78586, 50.40231, 50.00851, 49.60493, 49.19202, 
    48.77021, 48.33995, 47.90166, 47.45575, 47.00262, 46.54266, 46.07624, 
    45.60374, 45.1255, 44.64186, 44.15316, 43.6597, 43.16179, 42.65972, 
    42.15377, 41.64421, 41.13129, 40.61526, 40.09635, 39.57478,
  39.27911, 39.78861, 40.29517, 40.79858, 41.29861, 41.79502, 42.28755, 
    42.77596, 43.25996, 43.73928, 44.21362, 44.68269, 45.14617, 45.60374, 
    46.05505, 46.49977, 46.93754, 47.36799, 47.79074, 48.20541, 48.6116, 
    49.00891, 49.39692, 49.77522, 50.14338, 50.50098, 50.84757, 51.18272, 
    51.506, 51.81697, 52.11519, 52.40023, 52.67167, 52.92909, 53.17208, 
    53.40025, 53.61321, 53.81061, 53.99209, 54.15733, 54.30604, 54.43793, 
    54.55275, 54.6503, 54.73037, 54.79281, 54.8375, 54.86435, 54.87331, 
    54.86435, 54.8375, 54.79281, 54.73037, 54.6503, 54.55275, 54.43793, 
    54.30604, 54.15733, 53.99209, 53.81061, 53.61321, 53.40025, 53.17208, 
    52.92909, 52.67167, 52.40023, 52.11519, 51.81697, 51.506, 51.18272, 
    50.84757, 50.50098, 50.14338, 49.77522, 49.39692, 49.00891, 48.6116, 
    48.20541, 47.79074, 47.36799, 46.93754, 46.49977, 46.05505, 45.60374, 
    45.14617, 44.68269, 44.21362, 43.73928, 43.25996, 42.77596, 42.28755, 
    41.79502, 41.29861, 40.79858, 40.29517, 39.78861, 39.27911,
  38.977, 39.47439, 39.96857, 40.45934, 40.94647, 41.42973, 41.90887, 
    42.38366, 42.85382, 43.31909, 43.77919, 44.23382, 44.68269, 45.1255, 
    45.56192, 45.99162, 46.41428, 46.82954, 47.23705, 47.63646, 48.02739, 
    48.40947, 48.78232, 49.14555, 49.49877, 49.84158, 50.1736, 50.49441, 
    50.80363, 51.10085, 51.38569, 51.65775, 51.91666, 52.16203, 52.39351, 
    52.61073, 52.81337, 53.00109, 53.17359, 53.33059, 53.47181, 53.59702, 
    53.70599, 53.79853, 53.87448, 53.93369, 53.97606, 54.00152, 54.01001, 
    54.00152, 53.97606, 53.93369, 53.87448, 53.79853, 53.70599, 53.59702, 
    53.47181, 53.33059, 53.17359, 53.00109, 52.81337, 52.61073, 52.39351, 
    52.16203, 51.91666, 51.65775, 51.38569, 51.10085, 50.80363, 50.49441, 
    50.1736, 49.84158, 49.49877, 49.14555, 48.78232, 48.40947, 48.02739, 
    47.63646, 47.23705, 46.82954, 46.41428, 45.99162, 45.56192, 45.1255, 
    44.68269, 44.23382, 43.77919, 43.31909, 42.85382, 42.38366, 41.90887, 
    41.42973, 40.94647, 40.45934, 39.96857, 39.47439, 38.977,
  38.66859, 39.15382, 39.6356, 40.11372, 40.58796, 41.0581, 41.52391, 
    41.98514, 42.44154, 42.89287, 43.33884, 43.77919, 44.21362, 44.64186, 
    45.0636, 45.47853, 45.88634, 46.28671, 46.67929, 47.06378, 47.43981, 
    47.80704, 48.16513, 48.51371, 48.85243, 49.18093, 49.49884, 49.8058, 
    50.10146, 50.38545, 50.65742, 50.91702, 51.1639, 51.39774, 51.6182, 
    51.82498, 52.01776, 52.19627, 52.36022, 52.50938, 52.64349, 52.76235, 
    52.86576, 52.95356, 53.0256, 53.08176, 53.12194, 53.14607, 53.15412, 
    53.14607, 53.12194, 53.08176, 53.0256, 52.95356, 52.86576, 52.76235, 
    52.64349, 52.50938, 52.36022, 52.19627, 52.01776, 51.82498, 51.6182, 
    51.39774, 51.1639, 50.91702, 50.65742, 50.38545, 50.10146, 49.8058, 
    49.49884, 49.18093, 48.85243, 48.51371, 48.16513, 47.80704, 47.43981, 
    47.06378, 46.67929, 46.28671, 45.88634, 45.47853, 45.0636, 44.64186, 
    44.21362, 43.77919, 43.33884, 42.89287, 42.44154, 41.98514, 41.52391, 
    41.0581, 40.58796, 40.11372, 39.6356, 39.15382, 38.66859,
  38.354, 38.82706, 39.29642, 39.7619, 40.22328, 40.68035, 41.13287, 
    41.58063, 42.02338, 42.46088, 42.89287, 43.31909, 43.73928, 44.15316, 
    44.56044, 44.96085, 45.35409, 45.73986, 46.11785, 46.48775, 46.84925, 
    47.20202, 47.54575, 47.8801, 48.20476, 48.51939, 48.82367, 49.11726, 
    49.39985, 49.6711, 49.9307, 50.17833, 50.4137, 50.63649, 50.84642, 
    51.04321, 51.22659, 51.39631, 51.55212, 51.69381, 51.82117, 51.934, 
    52.03214, 52.11544, 52.18378, 52.23703, 52.27514, 52.29802, 52.30565, 
    52.29802, 52.27514, 52.23703, 52.18378, 52.11544, 52.03214, 51.934, 
    51.82117, 51.69381, 51.55212, 51.39631, 51.22659, 51.04321, 50.84642, 
    50.63649, 50.4137, 50.17833, 49.9307, 49.6711, 49.39985, 49.11726, 
    48.82367, 48.51939, 48.20476, 47.8801, 47.54575, 47.20202, 46.84925, 
    46.48775, 46.11785, 45.73986, 45.35409, 44.96085, 44.56044, 44.15316, 
    43.73928, 43.31909, 42.89287, 42.46088, 42.02338, 41.58063, 41.13287, 
    40.68035, 40.22328, 39.7619, 39.29642, 38.82706, 38.354,
  38.03334, 38.49422, 38.95119, 39.40405, 39.85261, 40.29666, 40.73598, 
    41.17037, 41.59958, 42.02338, 42.44154, 42.85382, 43.25996, 43.6597, 
    44.05278, 44.43893, 44.81789, 45.18936, 45.55307, 45.90874, 46.25607, 
    46.59477, 46.92454, 47.24509, 47.55613, 47.85734, 48.14844, 48.42913, 
    48.69912, 48.95811, 49.20582, 49.44197, 49.66629, 49.8785, 50.07836, 
    50.26561, 50.44002, 50.60136, 50.74942, 50.88401, 51.00494, 51.11204, 
    51.20517, 51.2842, 51.34902, 51.39953, 51.43566, 51.45736, 51.46459, 
    51.45736, 51.43566, 51.39953, 51.34902, 51.2842, 51.20517, 51.11204, 
    51.00494, 50.88401, 50.74942, 50.60136, 50.44002, 50.26561, 50.07836, 
    49.8785, 49.66629, 49.44197, 49.20582, 48.95811, 48.69912, 48.42913, 
    48.14844, 47.85734, 47.55613, 47.24509, 46.92454, 46.59477, 46.25607, 
    45.90874, 45.55307, 45.18936, 44.81789, 44.43893, 44.05278, 43.6597, 
    43.25996, 42.85382, 42.44154, 42.02338, 41.59958, 41.17037, 40.73598, 
    40.29666, 39.85261, 39.40405, 38.95119, 38.49422, 38.03334,
  37.70675, 38.15546, 38.60004, 39.04033, 39.47613, 39.90724, 40.33345, 
    40.75457, 41.17037, 41.58063, 41.98514, 42.38366, 42.77596, 43.16179, 
    43.54091, 43.91308, 44.27805, 44.63554, 44.98531, 45.3271, 45.66063, 
    45.98564, 46.30186, 46.60902, 46.90686, 47.1951, 47.47348, 47.74172, 
    47.99957, 48.24677, 48.48305, 48.70818, 48.92191, 49.124, 49.31422, 
    49.49236, 49.6582, 49.81155, 49.95222, 50.08005, 50.19486, 50.29652, 
    50.38489, 50.45986, 50.52134, 50.56924, 50.6035, 50.62407, 50.63093, 
    50.62407, 50.6035, 50.56924, 50.52134, 50.45986, 50.38489, 50.29652, 
    50.19486, 50.08005, 49.95222, 49.81155, 49.6582, 49.49236, 49.31422, 
    49.124, 48.92191, 48.70818, 48.48305, 48.24677, 47.99957, 47.74172, 
    47.47348, 47.1951, 46.90686, 46.60902, 46.30186, 45.98564, 45.66063, 
    45.3271, 44.98531, 44.63554, 44.27805, 43.91308, 43.54091, 43.16179, 
    42.77596, 42.38366, 41.98514, 41.58063, 41.17037, 40.75457, 40.33345, 
    39.90724, 39.47613, 39.04033, 38.60004, 38.15546, 37.70675,
  37.37434, 37.81089, 38.24314, 38.67091, 39.09401, 39.51227, 39.92548, 
    40.33345, 40.73598, 41.13287, 41.52391, 41.90887, 42.28755, 42.65972, 
    43.02515, 43.38362, 43.73489, 44.07872, 44.41489, 44.74314, 45.06325, 
    45.37495, 45.67802, 45.97221, 46.25727, 46.53297, 46.79906, 47.05531, 
    47.30147, 47.53732, 47.76263, 47.97718, 48.18076, 48.37315, 48.55416, 
    48.72359, 48.88126, 49.02699, 49.16062, 49.282, 49.39099, 49.48746, 
    49.57131, 49.64243, 49.70073, 49.74615, 49.77864, 49.79815, 49.80465, 
    49.79815, 49.77864, 49.74615, 49.70073, 49.64243, 49.57131, 49.48746, 
    49.39099, 49.282, 49.16062, 49.02699, 48.88126, 48.72359, 48.55416, 
    48.37315, 48.18076, 47.97718, 47.76263, 47.53732, 47.30147, 47.05531, 
    46.79906, 46.53297, 46.25727, 45.97221, 45.67802, 45.37495, 45.06325, 
    44.74314, 44.41489, 44.07872, 43.73489, 43.38362, 43.02515, 42.65972, 
    42.28755, 41.90887, 41.52391, 41.13287, 40.73598, 40.33345, 39.92548, 
    39.51227, 39.09401, 38.67091, 38.24314, 37.81089, 37.37434,
  37.03624, 37.46067, 37.88063, 38.29594, 38.70644, 39.11194, 39.51227, 
    39.90724, 40.29666, 40.68035, 41.0581, 41.42973, 41.79502, 42.15377, 
    42.50578, 42.85083, 43.18871, 43.51921, 43.84211, 44.15719, 44.46423, 
    44.76302, 45.05334, 45.33495, 45.60766, 45.87124, 46.12547, 46.37015, 
    46.60506, 46.83001, 47.04478, 47.24918, 47.44304, 47.62614, 47.79833, 
    47.95944, 48.10929, 48.24775, 48.37467, 48.48992, 48.59336, 48.68491, 
    48.76445, 48.83191, 48.8872, 48.93027, 48.96106, 48.97956, 48.98572, 
    48.97956, 48.96106, 48.93027, 48.8872, 48.83191, 48.76445, 48.68491, 
    48.59336, 48.48992, 48.37467, 48.24775, 48.10929, 47.95944, 47.79833, 
    47.62614, 47.44304, 47.24918, 47.04478, 46.83001, 46.60506, 46.37015, 
    46.12547, 45.87124, 45.60766, 45.33495, 45.05334, 44.76302, 44.46423, 
    44.15719, 43.84211, 43.51921, 43.18871, 42.85083, 42.50578, 42.15377, 
    41.79502, 41.42973, 41.0581, 40.68035, 40.29666, 39.90724, 39.51227, 
    39.11194, 38.70644, 38.29594, 37.88063, 37.46067, 37.03624,
  36.69255, 37.10492, 37.51265, 37.91559, 38.31358, 38.70644, 39.09401, 
    39.47613, 39.85261, 40.22328, 40.58796, 40.94647, 41.29861, 41.64421, 
    41.98307, 42.315, 42.6398, 42.95729, 43.26726, 43.56952, 43.86388, 
    44.15013, 44.42807, 44.69753, 44.95829, 45.21016, 45.45296, 45.68649, 
    45.91058, 46.12503, 46.32969, 46.52436, 46.70888, 46.8831, 47.04686, 
    47.20001, 47.34241, 47.47393, 47.59445, 47.70385, 47.80202, 47.88887, 
    47.96432, 48.02829, 48.08072, 48.12155, 48.15074, 48.16827, 48.17411, 
    48.16827, 48.15074, 48.12155, 48.08072, 48.02829, 47.96432, 47.88887, 
    47.80202, 47.70385, 47.59445, 47.47393, 47.34241, 47.20001, 47.04686, 
    46.8831, 46.70888, 46.52436, 46.32969, 46.12503, 45.91058, 45.68649, 
    45.45296, 45.21016, 44.95829, 44.69753, 44.42807, 44.15013, 43.86388, 
    43.56952, 43.26726, 42.95729, 42.6398, 42.315, 41.98307, 41.64421, 
    41.29861, 40.94647, 40.58796, 40.22328, 39.85261, 39.47613, 39.09401, 
    38.70644, 38.31358, 37.91559, 37.51265, 37.10492, 36.69255,
  36.34341, 36.74377, 37.13935, 37.53001, 37.91559, 38.29594, 38.67091, 
    39.04033, 39.40405, 39.7619, 40.11372, 40.45934, 40.79858, 41.13129, 
    41.45728, 41.77639, 42.08843, 42.39323, 42.69062, 42.98042, 43.26245, 
    43.53653, 43.8025, 44.06018, 44.30939, 44.54997, 44.78174, 45.00454, 
    45.21821, 45.42259, 45.61752, 45.80286, 45.97845, 46.14417, 46.29986, 
    46.4454, 46.58068, 46.70559, 46.82, 46.92382, 47.01697, 47.09935, 
    47.17091, 47.23156, 47.28126, 47.31997, 47.34763, 47.36425, 47.36979, 
    47.36425, 47.34763, 47.31997, 47.28126, 47.23156, 47.17091, 47.09935, 
    47.01697, 46.92382, 46.82, 46.70559, 46.58068, 46.4454, 46.29986, 
    46.14417, 45.97845, 45.80286, 45.61752, 45.42259, 45.21821, 45.00454, 
    44.78174, 44.54997, 44.30939, 44.06018, 43.8025, 43.53653, 43.26245, 
    42.98042, 42.69062, 42.39323, 42.08843, 41.77639, 41.45728, 41.13129, 
    40.79858, 40.45934, 40.11372, 39.7619, 39.40405, 39.04033, 38.67091, 
    38.29594, 37.91559, 37.53001, 37.13935, 36.74377, 36.34341,
  35.98892, 36.37735, 36.76087, 37.13935, 37.51265, 37.88063, 38.24314, 
    38.60004, 38.95119, 39.29642, 39.6356, 39.96857, 40.29517, 40.61526, 
    40.92867, 41.23525, 41.53484, 41.82729, 42.11243, 42.39012, 42.66019, 
    42.92249, 43.17686, 43.42315, 43.66121, 43.89089, 44.11203, 44.3245, 
    44.52815, 44.72285, 44.90845, 45.08484, 45.25187, 45.40944, 45.55742, 
    45.6957, 45.82418, 45.94276, 46.05135, 46.14986, 46.23822, 46.31635, 
    46.38419, 46.44169, 46.4888, 46.52548, 46.5517, 46.56744, 46.57269, 
    46.56744, 46.5517, 46.52548, 46.4888, 46.44169, 46.38419, 46.31635, 
    46.23822, 46.14986, 46.05135, 45.94276, 45.82418, 45.6957, 45.55742, 
    45.40944, 45.25187, 45.08484, 44.90845, 44.72285, 44.52815, 44.3245, 
    44.11203, 43.89089, 43.66121, 43.42315, 43.17686, 42.92249, 42.66019, 
    42.39012, 42.11243, 41.82729, 41.53484, 41.23525, 40.92867, 40.61526, 
    40.29517, 39.96857, 39.6356, 39.29642, 38.95119, 38.60004, 38.24314, 
    37.88063, 37.51265, 37.13935, 36.76087, 36.37735, 35.98892,
  35.62921, 36.00579, 36.37735, 36.74377, 37.10492, 37.46067, 37.81089, 
    38.15546, 38.49422, 38.82706, 39.15382, 39.47439, 39.78861, 40.09635, 
    40.39747, 40.69183, 40.97929, 41.25971, 41.53295, 41.79888, 42.05735, 
    42.30823, 42.55138, 42.78666, 43.01395, 43.23311, 43.44402, 43.64655, 
    43.84056, 44.02596, 44.20261, 44.37041, 44.52925, 44.67902, 44.81961, 
    44.95095, 45.07294, 45.18549, 45.28852, 45.38197, 45.46576, 45.53984, 
    45.60415, 45.65865, 45.7033, 45.73805, 45.7629, 45.77781, 45.78278, 
    45.77781, 45.7629, 45.73805, 45.7033, 45.65865, 45.60415, 45.53984, 
    45.46576, 45.38197, 45.28852, 45.18549, 45.07294, 44.95095, 44.81961, 
    44.67902, 44.52925, 44.37041, 44.20261, 44.02596, 43.84056, 43.64655, 
    43.44402, 43.23311, 43.01395, 42.78666, 42.55138, 42.30823, 42.05735, 
    41.79888, 41.53295, 41.25971, 40.97929, 40.69183, 40.39747, 40.09635, 
    39.78861, 39.47439, 39.15382, 38.82706, 38.49422, 38.15546, 37.81089, 
    37.46067, 37.10492, 36.74377, 36.37735, 36.00579, 35.62921,
  35.26439, 35.62921, 35.98892, 36.34341, 36.69255, 37.03624, 37.37434, 
    37.70675, 38.03334, 38.354, 38.66859, 38.977, 39.27911, 39.57478, 
    39.8639, 40.14635, 40.42199, 40.69072, 40.9524, 41.20691, 41.45414, 
    41.69396, 41.92625, 42.15091, 42.36781, 42.57683, 42.77788, 42.97084, 
    43.1556, 43.33206, 43.50012, 43.65969, 43.81068, 43.95298, 44.08652, 
    44.21122, 44.32701, 44.4338, 44.53154, 44.62016, 44.6996, 44.76982, 
    44.83077, 44.88241, 44.9247, 44.95763, 44.98116, 44.99529, 45, 44.99529, 
    44.98116, 44.95763, 44.9247, 44.88241, 44.83077, 44.76982, 44.6996, 
    44.62016, 44.53154, 44.4338, 44.32701, 44.21122, 44.08652, 43.95298, 
    43.81068, 43.65969, 43.50012, 43.33206, 43.1556, 42.97084, 42.77788, 
    42.57683, 42.36781, 42.15091, 41.92625, 41.69396, 41.45414, 41.20691, 
    40.9524, 40.69072, 40.42199, 40.14635, 39.8639, 39.57478, 39.27911, 
    38.977, 38.66859, 38.354, 38.03334, 37.70675, 37.37434, 37.03624, 
    36.69255, 36.34341, 35.98892, 35.62921, 35.26439 ;

 grid_lont =
  35, 35.78653, 36.58051, 37.38202, 38.19109, 39.00779, 39.83216, 40.66424, 
    41.50406, 42.35163, 43.20698, 44.07011, 44.94102, 45.81969, 46.7061, 
    47.60023, 48.50203, 49.41144, 50.32841, 51.25285, 52.18468, 53.1238, 
    54.0701, 55.02345, 55.98371, 56.95073, 57.92436, 58.90441, 59.89069, 
    60.88301, 61.88113, 62.88485, 63.89391, 64.90805, 65.92702, 66.95055, 
    67.97832, 69.01007, 70.04546, 71.08418, 72.12592, 73.17033, 74.21706, 
    75.26579, 76.31613, 77.36775, 78.42029, 79.47337, 80.52663, 81.57971, 
    82.63225, 83.68387, 84.73421, 85.78294, 86.82967, 87.87408, 88.91582, 
    89.95454, 90.98993, 92.02168, 93.04945, 94.07298, 95.09195, 96.10609, 
    97.11515, 98.11887, 99.117, 100.1093, 101.0956, 102.0756, 103.0493, 
    104.0163, 104.9766, 105.9299, 106.8762, 107.8153, 108.7472, 109.6716, 
    110.5886, 111.498, 112.3998, 113.2939, 114.1803, 115.059, 115.9299, 
    116.793, 117.6484, 118.4959, 119.3358, 120.1678, 120.9922, 121.8089, 
    122.618, 123.4195, 124.2135, 125,
  34.21347, 35, 35.79459, 36.59731, 37.40824, 38.22746, 39.05501, 39.89095, 
    40.73534, 41.5882, 42.44957, 43.31946, 44.1979, 45.08487, 45.98036, 
    46.88437, 47.79684, 48.71775, 49.64702, 50.58459, 51.53038, 52.48428, 
    53.44618, 54.41596, 55.39347, 56.37855, 57.37103, 58.37072, 59.37743, 
    60.39091, 61.41096, 62.43731, 63.46969, 64.50784, 65.55144, 66.6002, 
    67.65379, 68.71187, 69.7741, 70.84013, 71.90958, 72.98206, 74.05721, 
    75.13461, 76.21387, 77.29458, 78.37634, 79.45871, 80.54129, 81.62366, 
    82.70542, 83.78613, 84.86539, 85.94279, 87.01794, 88.09042, 89.15987, 
    90.2259, 91.28813, 92.34621, 93.3998, 94.44856, 95.49216, 96.5303, 
    97.56269, 98.58904, 99.60909, 100.6226, 101.6293, 102.629, 103.6215, 
    104.6065, 105.584, 106.5538, 107.5157, 108.4696, 109.4154, 110.353, 
    111.2822, 112.2032, 113.1156, 114.0196, 114.9151, 115.8021, 116.6805, 
    117.5504, 118.4118, 119.2647, 120.109, 120.945, 121.7725, 122.5918, 
    123.4027, 124.2054, 125, 125.7865,
  33.41949, 34.20541, 35, 35.80334, 36.61554, 37.43667, 38.26682, 39.10607, 
    39.95446, 40.81208, 41.67894, 42.55511, 43.44059, 44.33541, 45.23958, 
    46.15308, 47.07589, 48.00798, 48.9493, 49.89978, 50.85935, 51.82791, 
    52.80535, 53.79154, 54.78633, 55.78957, 56.80106, 57.82062, 58.84803, 
    59.88304, 60.92541, 61.97486, 63.03111, 64.09383, 65.16272, 66.23743, 
    67.3176, 68.40284, 69.49279, 70.58703, 71.68514, 72.78671, 73.89129, 
    74.99844, 76.1077, 77.2186, 78.33069, 79.44348, 80.55652, 81.66931, 
    82.7814, 83.8923, 85.00156, 86.10871, 87.21329, 88.31486, 89.41297, 
    90.50721, 91.59716, 92.6824, 93.76257, 94.83728, 95.90617, 96.96889, 
    98.02514, 99.07459, 100.117, 101.152, 102.1794, 103.1989, 104.2104, 
    105.2137, 106.2085, 107.1946, 108.1721, 109.1406, 110.1002, 111.0507, 
    111.992, 112.9241, 113.8469, 114.7604, 115.6646, 116.5594, 117.4449, 
    118.3211, 119.1879, 120.0455, 120.8939, 121.7332, 122.5633, 123.3845, 
    124.1967, 125, 125.7946, 126.5805,
  32.61798, 33.40269, 34.19666, 35, 35.81284, 36.63528, 37.46742, 38.30936, 
    39.16119, 40.02298, 40.89479, 41.77669, 42.66872, 43.57091, 44.4833, 
    45.40587, 46.33863, 47.28156, 48.23462, 49.19776, 50.17091, 51.15397, 
    52.14684, 53.1494, 54.1615, 55.18297, 56.21362, 57.25326, 58.30164, 
    59.35852, 60.42362, 61.49665, 62.5773, 63.66523, 64.76008, 65.86147, 
    66.96902, 68.08229, 69.20087, 70.32429, 71.4521, 72.5838, 73.71891, 
    74.85693, 75.99734, 77.13962, 78.28323, 79.42766, 80.57234, 81.71677, 
    82.86038, 84.00266, 85.14307, 86.28109, 87.4162, 88.5479, 89.67571, 
    90.79913, 91.91771, 93.03098, 94.13853, 95.23992, 96.33477, 97.4227, 
    98.50335, 99.57638, 100.6415, 101.6984, 102.7467, 103.7864, 104.817, 
    105.8385, 106.8506, 107.8532, 108.846, 109.8291, 110.8022, 111.7654, 
    112.7184, 113.6614, 114.5941, 115.5167, 116.4291, 117.3313, 118.2233, 
    119.1052, 119.977, 120.8388, 121.6906, 122.5326, 123.3647, 124.1872, 125, 
    125.8033, 126.5973, 127.382,
  31.80891, 32.59176, 33.38446, 34.18716, 35, 35.8231, 36.65661, 37.50062, 
    38.35526, 39.22061, 40.09678, 40.98385, 41.88187, 42.79092, 43.71102, 
    44.64221, 45.5845, 46.53789, 47.50235, 48.47785, 49.46433, 50.4617, 
    51.46988, 52.48874, 53.51813, 54.55788, 55.60782, 56.66772, 57.73734, 
    58.81642, 59.90467, 61.00177, 62.10738, 63.22114, 64.34265, 65.47151, 
    66.60727, 67.74947, 68.89764, 70.05127, 71.20984, 72.37281, 73.53963, 
    74.70972, 75.88252, 77.05743, 78.23385, 79.41118, 80.58882, 81.76615, 
    82.94257, 84.11748, 85.29028, 86.46037, 87.62719, 88.79016, 89.94873, 
    91.10236, 92.25053, 93.39273, 94.52849, 95.65735, 96.77886, 97.89262, 
    98.99823, 100.0953, 101.1836, 102.2627, 103.3323, 104.3922, 105.4421, 
    106.4819, 107.5113, 108.5301, 109.5383, 110.5357, 111.5221, 112.4977, 
    113.4621, 114.4155, 115.3578, 116.289, 117.2091, 118.1181, 119.0162, 
    119.9032, 120.7794, 121.6447, 122.4994, 123.3434, 124.1769, 125, 
    125.8128, 126.6155, 127.4082, 128.1911,
  30.99221, 31.77254, 32.56333, 33.36472, 34.1769, 35, 35.83419, 36.67962, 
    37.53641, 38.4047, 39.2846, 40.17622, 41.07965, 41.99498, 42.92228, 
    43.86158, 44.81293, 45.77634, 46.75183, 47.73935, 48.73887, 49.75033, 
    50.77364, 51.80869, 52.85532, 53.9134, 54.98272, 56.06305, 57.15416, 
    58.25577, 59.36757, 60.48923, 61.62037, 62.76061, 63.90952, 65.06664, 
    66.2315, 67.40359, 68.58237, 69.76728, 70.95776, 72.15318, 73.35295, 
    74.55641, 75.76292, 76.9718, 78.1824, 79.39402, 80.60598, 81.8176, 
    83.0282, 84.23708, 85.44359, 86.64705, 87.84682, 89.04224, 90.23272, 
    91.41763, 92.59641, 93.7685, 94.93336, 96.09048, 97.2394, 98.37963, 
    99.51077, 100.6324, 101.7442, 102.8458, 103.937, 105.0173, 106.0866, 
    107.1447, 108.1913, 109.2264, 110.2497, 111.2611, 112.2607, 113.2482, 
    114.2237, 115.1871, 116.1384, 117.0777, 118.005, 118.9203, 119.8238, 
    120.7154, 121.5953, 122.4636, 123.3204, 124.1658, 125, 125.8231, 
    126.6353, 127.4367, 128.2274, 129.0078,
  30.16784, 30.94499, 31.73318, 32.53258, 33.34339, 34.16581, 35, 35.84615, 
    36.70441, 37.57496, 38.45793, 39.35345, 40.26167, 41.18267, 42.11657, 
    43.06343, 44.02333, 44.9963, 45.98236, 46.98153, 47.99377, 49.01904, 
    50.05726, 51.10835, 52.17216, 53.24854, 54.33731, 55.43823, 56.55107, 
    57.67552, 58.81128, 59.95797, 61.11523, 62.28261, 63.45966, 64.64589, 
    65.84076, 67.04373, 68.2542, 69.47156, 70.69515, 71.92432, 73.15836, 
    74.39655, 75.63818, 76.88248, 78.12872, 79.37611, 80.62389, 81.87128, 
    83.11752, 84.36182, 85.60345, 86.84164, 88.07568, 89.30485, 90.52844, 
    91.7458, 92.95627, 94.15924, 95.35411, 96.54034, 97.71739, 98.88477, 
    100.042, 101.1887, 102.3245, 103.4489, 104.5618, 105.6627, 106.7515, 
    107.8278, 108.8917, 109.9427, 110.981, 112.0062, 113.0185, 114.0176, 
    115.0037, 115.9767, 116.9366, 117.8834, 118.8173, 119.7383, 120.6465, 
    121.5421, 122.425, 123.2956, 124.1539, 125, 125.8342, 126.6566, 127.4674, 
    128.2668, 129.055, 129.8322,
  29.33576, 30.10905, 30.89393, 31.69064, 32.49938, 33.32038, 34.15385, 35, 
    35.85902, 36.73111, 37.61644, 38.51518, 39.4275, 40.35353, 41.2934, 
    42.24723, 43.2151, 44.1971, 45.19327, 46.20364, 47.22821, 48.26696, 
    49.31985, 50.38678, 51.46764, 52.56229, 53.67054, 54.79218, 55.92694, 
    57.07454, 58.23465, 59.40688, 60.59082, 61.78603, 62.992, 64.20821, 
    65.43406, 66.66897, 67.91226, 69.16328, 70.42128, 71.68554, 72.95527, 
    74.22968, 75.50793, 76.78922, 78.07266, 79.35741, 80.64259, 81.92734, 
    83.21078, 84.49207, 85.77032, 87.04473, 88.31446, 89.57872, 90.83672, 
    92.08774, 93.33103, 94.56594, 95.79179, 97.008, 98.21397, 99.40917, 
    100.5931, 101.7654, 102.9255, 104.0731, 105.2078, 106.3295, 107.4377, 
    108.5324, 109.6132, 110.6802, 111.733, 112.7718, 113.7964, 114.8067, 
    115.8029, 116.7849, 117.7528, 118.7066, 119.6465, 120.5725, 121.4848, 
    122.3836, 123.2689, 124.141, 125, 125.8461, 126.6796, 127.5006, 128.3094, 
    129.1061, 129.8909, 130.6642,
  28.49594, 29.26466, 30.04553, 30.83881, 31.64474, 32.46359, 33.29559, 
    34.14098, 35, 35.87288, 36.75983, 37.66105, 38.57675, 39.5071, 40.45227, 
    41.41241, 42.38765, 43.37809, 44.38382, 45.4049, 46.44137, 47.49323, 
    48.56046, 49.64299, 50.74073, 51.85356, 52.98129, 54.12373, 55.28061, 
    56.45164, 57.63647, 58.83472, 60.04595, 61.26968, 62.50537, 63.75245, 
    65.0103, 66.27824, 67.55556, 68.84151, 70.13531, 71.4361, 72.74305, 
    74.05524, 75.37177, 76.69168, 78.01403, 79.33784, 80.66216, 81.98597, 
    83.30832, 84.62823, 85.94476, 87.25695, 88.5639, 89.86469, 91.15849, 
    92.44444, 93.72176, 94.9897, 96.24755, 97.49463, 98.73032, 99.95405, 
    101.1653, 102.3635, 103.5484, 104.7194, 105.8763, 107.0187, 108.1464, 
    109.2593, 110.357, 111.4395, 112.5068, 113.5586, 114.5951, 115.6162, 
    116.6219, 117.6124, 118.5876, 119.5477, 120.4929, 121.4232, 122.339, 
    123.2402, 124.1271, 125, 125.859, 126.7044, 127.5364, 128.3553, 129.1612, 
    129.9545, 130.7353, 131.5041,
  27.64837, 28.4118, 29.18793, 29.97702, 30.77939, 31.5953, 32.42504, 
    33.26889, 34.12712, 35, 35.88778, 36.79071, 37.70902, 38.64294, 39.59268, 
    40.55842, 41.54034, 42.53858, 43.55327, 44.58451, 45.63238, 46.69691, 
    47.77811, 48.87594, 49.99035, 51.12122, 52.26839, 53.43167, 54.61082, 
    55.80553, 57.01546, 58.2402, 59.4793, 60.73225, 61.99849, 63.27739, 
    64.56827, 65.87041, 67.18303, 68.50529, 69.83633, 71.17522, 72.521, 
    73.87267, 75.2292, 76.58955, 77.95263, 79.31736, 80.68264, 82.04737, 
    83.41045, 84.7708, 86.12733, 87.479, 88.82478, 90.16367, 91.49471, 
    92.81697, 94.12959, 95.43173, 96.72261, 98.00151, 99.26775, 100.5207, 
    101.7598, 102.9845, 104.1945, 105.3892, 106.5683, 107.7316, 108.8788, 
    110.0097, 111.1241, 112.2219, 113.3031, 114.3676, 115.4155, 116.4467, 
    117.4614, 118.4597, 119.4416, 120.4073, 121.3571, 122.291, 123.2093, 
    124.1122, 125, 125.8729, 126.7311, 127.575, 128.4047, 129.2206, 130.023, 
    130.8121, 131.5882, 132.3516,
  26.79302, 27.55043, 28.32106, 29.10521, 29.90322, 30.7154, 31.54207, 
    32.38356, 33.24017, 34.11222, 35, 35.9038, 36.82391, 37.7606, 38.71411, 
    39.68468, 40.67255, 41.67789, 42.70088, 43.74166, 44.80036, 45.87705, 
    46.97178, 48.08456, 49.21534, 50.36406, 51.53057, 52.7147, 53.91622, 
    55.13484, 56.3702, 57.6219, 58.88946, 60.17235, 61.46997, 62.78166, 
    64.10667, 65.44424, 66.7935, 68.15353, 69.52337, 70.902, 72.28835, 
    73.68132, 75.07974, 76.48245, 77.88824, 79.29588, 80.70412, 82.11176, 
    83.51755, 84.92026, 86.31868, 87.71165, 89.098, 90.47663, 91.84647, 
    93.2065, 94.55576, 95.89333, 97.21835, 98.53003, 99.82764, 101.1105, 
    102.3781, 103.6298, 104.8652, 106.0838, 107.2853, 108.4694, 109.6359, 
    110.7847, 111.9154, 113.0282, 114.1229, 115.1996, 116.2583, 117.2991, 
    118.3221, 119.3275, 120.3153, 121.2859, 122.2394, 123.1761, 124.0962, 
    125, 125.8878, 126.7598, 127.6164, 128.4579, 129.2846, 130.0968, 
    130.8948, 131.6789, 132.4496, 133.207,
  25.92989, 26.68054, 27.44489, 28.22331, 29.01615, 29.82378, 30.64655, 
    31.48482, 32.33895, 33.20929, 34.0962, 35, 35.92104, 36.85962, 37.81606, 
    38.79064, 39.78364, 40.79531, 41.82586, 42.8755, 43.94439, 45.03267, 
    46.14042, 47.2677, 48.41451, 49.58081, 50.76651, 51.97144, 53.19539, 
    54.4381, 55.6992, 56.9783, 58.2749, 59.58846, 60.91832, 62.26379, 
    63.62409, 64.99835, 66.38566, 67.785, 69.1953, 70.61546, 72.04426, 
    73.48048, 74.92283, 76.36999, 77.8206, 79.2733, 80.7267, 82.1794, 
    83.63001, 85.07717, 86.51952, 87.95574, 89.38454, 90.8047, 92.215, 
    93.61434, 95.00165, 96.37591, 97.73621, 99.08168, 100.4115, 101.7251, 
    103.0217, 104.3008, 105.5619, 106.8046, 108.0286, 109.2335, 110.4192, 
    111.5855, 112.7323, 113.8596, 114.9673, 116.0556, 117.1245, 118.1741, 
    119.2047, 120.2164, 121.2094, 122.1839, 123.1404, 124.079, 125, 125.9038, 
    126.7907, 127.661, 128.5152, 129.3535, 130.1762, 130.9838, 131.7767, 
    132.5551, 133.3195, 134.0701,
  25.05898, 25.8021, 26.55941, 27.33128, 28.11813, 28.92034, 29.73833, 
    30.5725, 31.42325, 32.29098, 33.17609, 34.07896, 35, 35.93956, 36.89802, 
    37.87572, 38.87298, 39.89013, 40.92743, 41.98516, 43.06353, 44.16273, 
    45.28292, 46.42419, 47.5866, 48.77015, 49.9748, 51.20041, 52.44681, 
    53.71373, 55.00086, 56.30777, 57.63398, 58.9789, 60.34189, 61.72218, 
    63.11895, 64.53126, 65.9581, 67.39838, 68.85094, 70.3145, 71.78777, 
    73.26935, 74.75782, 76.25169, 77.74946, 79.24956, 80.75044, 82.25054, 
    83.74831, 85.24218, 86.73065, 88.21223, 89.6855, 91.14906, 92.60162, 
    94.0419, 95.46874, 96.88105, 98.27782, 99.65811, 101.0211, 102.366, 
    103.6922, 104.9991, 106.2863, 107.5532, 108.7996, 110.0252, 111.2298, 
    112.4134, 113.5758, 114.7171, 115.8373, 116.9365, 118.0148, 119.0726, 
    120.1099, 121.127, 122.1243, 123.102, 124.0604, 125, 125.921, 126.8239, 
    127.709, 128.5768, 129.4275, 130.2617, 131.0797, 131.8819, 132.6687, 
    133.4406, 134.1979, 134.941,
  24.18031, 24.91513, 25.66458, 26.42909, 27.20908, 28.00501, 28.81733, 
    29.64647, 30.4929, 31.35706, 32.2394, 33.14038, 34.06044, 35, 35.9595, 
    36.93934, 37.93993, 38.96163, 40.0048, 41.06976, 42.1568, 43.26619, 
    44.39812, 45.55278, 46.73028, 47.93068, 49.15396, 50.40006, 51.66884, 
    52.96007, 54.27343, 55.60854, 56.96489, 58.34191, 59.7389, 61.15507, 
    62.58954, 64.0413, 65.50926, 66.99223, 68.48891, 69.99794, 71.51784, 
    73.04707, 74.58404, 76.12708, 77.67448, 79.22453, 80.77547, 82.32552, 
    83.87292, 85.41596, 86.95293, 88.48216, 90.00206, 91.51109, 93.00777, 
    94.49074, 95.9587, 97.41046, 98.84492, 100.2611, 101.6581, 103.0351, 
    104.3915, 105.7266, 107.0399, 108.3312, 109.5999, 110.846, 112.0693, 
    113.2697, 114.4472, 115.6019, 116.7338, 117.8432, 118.9302, 119.9952, 
    121.0384, 122.0601, 123.0607, 124.0405, 125, 125.9396, 126.8596, 
    127.7606, 128.6429, 129.5071, 130.3535, 131.1827, 131.995, 132.7909, 
    133.5709, 134.3354, 135.0849, 135.8197,
  23.2939, 24.01964, 24.76042, 25.51671, 26.28898, 27.07773, 27.88343, 
    28.7066, 29.54773, 30.40732, 31.28589, 32.18394, 33.10198, 34.0405, 35, 
    35.98096, 36.98384, 38.00909, 39.05714, 40.1284, 41.22322, 42.34195, 
    43.48486, 44.65221, 45.84418, 47.0609, 48.30243, 49.56874, 50.85976, 
    52.1753, 53.51507, 54.8787, 56.26572, 57.67552, 59.1074, 60.56054, 
    62.03398, 63.52666, 65.03741, 66.56492, 68.10777, 69.66443, 71.23329, 
    72.81264, 74.40068, 75.99556, 77.59536, 79.19812, 80.80188, 82.40464, 
    84.00444, 85.59932, 87.18736, 88.76671, 90.33557, 91.89223, 93.43508, 
    94.96259, 96.47334, 97.96602, 99.43947, 100.8926, 102.3245, 103.7343, 
    105.1213, 106.4849, 107.8247, 109.1402, 110.4313, 111.6976, 112.9391, 
    114.1558, 115.3478, 116.5151, 117.6581, 118.7768, 119.8716, 120.9429, 
    121.9909, 123.0162, 124.019, 125, 125.9595, 126.898, 127.8161, 128.7141, 
    129.5927, 130.4523, 131.2934, 132.1166, 132.9223, 133.711, 134.4833, 
    135.2396, 135.9804, 136.7061,
  22.39977, 23.11563, 23.84692, 24.59413, 25.35779, 26.13842, 26.93657, 
    27.75277, 28.58759, 29.44158, 30.31532, 31.20936, 32.12428, 33.06066, 
    34.01904, 35, 36.00407, 37.03178, 38.08365, 39.16016, 40.26177, 41.38889, 
    42.5419, 43.72113, 44.92685, 46.15928, 47.41854, 48.7047, 50.01773, 
    51.35749, 52.72377, 54.1162, 55.53435, 56.9776, 58.44526, 59.93645, 
    61.4502, 62.98535, 64.54063, 66.11464, 67.70582, 69.31248, 70.93284, 
    72.56498, 74.2069, 75.85651, 77.51168, 79.17019, 80.82981, 82.48832, 
    84.14349, 85.7931, 87.43502, 89.06716, 90.68752, 92.29418, 93.88536, 
    95.45937, 97.01465, 98.5498, 100.0635, 101.5547, 103.0224, 104.4657, 
    105.8838, 107.2762, 108.6425, 109.9823, 111.2953, 112.5815, 113.8407, 
    115.0732, 116.2789, 117.4581, 118.6111, 119.7382, 120.8398, 121.9163, 
    122.9682, 123.9959, 125, 125.981, 126.9393, 127.8757, 128.7906, 129.6847, 
    130.5584, 131.4124, 132.2472, 133.0634, 133.8616, 134.6422, 135.4059, 
    136.1531, 136.8844, 137.6002,
  21.49797, 22.20316, 22.9241, 23.66137, 24.4155, 25.18707, 25.97667, 
    26.7849, 27.61235, 28.45966, 29.32745, 30.21636, 31.12702, 32.06007, 
    33.01616, 33.99593, 35, 36.02899, 37.08351, 38.16413, 39.27141, 40.40586, 
    41.56797, 42.75816, 43.9768, 45.22419, 46.50057, 47.80608, 49.14077, 
    50.50459, 51.89737, 53.31882, 54.76851, 56.24585, 57.75015, 59.28052, 
    60.83591, 62.41513, 64.01681, 65.6394, 67.28123, 68.94042, 70.615, 
    72.30284, 74.00169, 75.70923, 77.42302, 79.14059, 80.85941, 82.57698, 
    84.29077, 85.99831, 87.69716, 89.385, 91.05958, 92.71877, 94.3606, 
    95.98319, 97.58487, 99.16409, 100.7195, 102.2498, 103.7541, 105.2315, 
    106.6812, 108.1026, 109.4954, 110.8592, 112.1939, 113.4994, 114.7758, 
    116.0232, 117.2418, 118.432, 119.5941, 120.7286, 121.8359, 122.9165, 
    123.971, 125, 126.0041, 126.9838, 127.9399, 128.873, 129.7836, 130.6725, 
    131.5403, 132.3876, 133.2151, 134.0233, 134.8129, 135.5845, 136.3386, 
    137.0759, 137.7968, 138.502,
  20.58856, 21.28225, 21.99202, 22.71844, 23.46211, 24.22366, 25.0037, 
    25.8029, 26.62191, 27.46142, 28.32211, 29.20469, 30.10987, 31.03837, 
    31.99091, 32.96822, 33.97101, 35, 36.0559, 37.13938, 38.25111, 39.39172, 
    40.56179, 41.76188, 42.99245, 44.25394, 45.54667, 46.87091, 48.22681, 
    49.6144, 51.03359, 52.48415, 53.96572, 55.47775, 57.01952, 58.59017, 
    60.1886, 61.81356, 63.46357, 65.13697, 66.83192, 68.54638, 70.27814, 
    72.02484, 73.78397, 75.55289, 77.32889, 79.10915, 80.89085, 82.67111, 
    84.44711, 86.21603, 87.97516, 89.72186, 91.45362, 93.16808, 94.86303, 
    96.53644, 98.18644, 99.81139, 101.4098, 102.9805, 104.5223, 106.0343, 
    107.5158, 108.9664, 110.3856, 111.7732, 113.1291, 114.4533, 115.7461, 
    117.0076, 118.2381, 119.4382, 120.6083, 121.7489, 122.8606, 123.9441, 
    125, 126.029, 127.0318, 128.0091, 128.9616, 129.8901, 130.7953, 131.6779, 
    132.5386, 133.3781, 134.1971, 134.9963, 135.7764, 136.5379, 137.2816, 
    138.008, 138.7177, 139.4114,
  19.67159, 20.35298, 21.0507, 21.76538, 22.49765, 23.24817, 24.01764, 
    24.80673, 25.61618, 26.44673, 27.29912, 28.17414, 29.07257, 29.9952, 
    30.94286, 31.91635, 32.91649, 33.9441, 35, 36.08498, 37.19981, 38.34526, 
    39.52203, 40.7308, 41.97219, 43.24675, 44.55494, 45.89714, 47.27363, 
    48.68455, 50.12992, 51.60961, 53.1233, 54.67052, 56.25058, 57.86261, 
    59.50549, 61.17789, 62.87827, 64.60484, 66.35557, 68.12824, 69.9204, 
    71.72941, 73.55246, 75.3866, 77.22873, 79.07571, 80.92429, 82.77127, 
    84.6134, 86.44754, 88.27059, 90.0796, 91.87176, 93.64443, 95.39516, 
    97.12173, 98.82211, 100.4945, 102.1374, 103.7494, 105.3295, 106.8767, 
    108.3904, 109.8701, 111.3155, 112.7264, 114.1029, 115.4451, 116.7533, 
    118.0278, 119.2692, 120.478, 121.6547, 122.8002, 123.915, 125, 126.0559, 
    127.0835, 128.0836, 129.0571, 130.0048, 130.9274, 131.8259, 132.7009, 
    133.5533, 134.3838, 135.1933, 135.9824, 136.7518, 137.5023, 138.2346, 
    138.9493, 139.647, 140.3284,
  18.74715, 19.41541, 20.10022, 20.80224, 21.52215, 22.26065, 23.01847, 
    23.79636, 24.5951, 25.41549, 26.25834, 27.1245, 28.01484, 28.93024, 
    29.8716, 30.83984, 31.83587, 32.86062, 33.91502, 35, 36.11646, 37.26529, 
    38.44734, 39.66344, 40.91436, 42.20078, 43.52334, 44.88256, 46.27887, 
    47.71254, 49.18372, 50.69239, 52.23835, 53.82118, 55.44026, 57.09473, 
    58.78346, 60.5051, 62.25798, 64.04021, 65.84957, 67.68363, 69.53967, 
    71.41476, 73.30575, 75.20929, 77.12191, 79.04002, 80.95998, 82.87809, 
    84.79071, 86.69425, 88.58524, 90.46033, 92.31637, 94.15043, 95.95979, 
    97.74202, 99.4949, 101.2165, 102.9053, 104.5597, 106.1788, 107.7617, 
    109.3076, 110.8163, 112.2875, 113.7211, 115.1174, 116.4767, 117.7992, 
    119.0856, 120.3366, 121.5527, 122.7347, 123.8835, 125, 126.085, 127.1394, 
    128.1641, 129.1602, 130.1284, 131.0698, 131.9852, 132.8755, 133.7417, 
    134.5845, 135.4049, 136.2036, 136.9815, 137.7393, 138.4779, 139.1978, 
    139.8998, 140.5846, 141.2529,
  17.81532, 18.46962, 19.14065, 19.82909, 20.53567, 21.26113, 22.00623, 
    22.77179, 23.55863, 24.36762, 25.19964, 26.05561, 26.93647, 27.8432, 
    28.77678, 29.73823, 30.72859, 31.74889, 32.80019, 33.88354, 35, 36.1506, 
    37.33636, 38.55825, 39.81722, 41.11413, 42.44979, 43.82489, 45.24004, 
    46.69568, 48.19212, 49.72948, 51.30768, 52.92643, 54.58518, 56.28311, 
    58.01911, 59.79178, 61.5994, 63.43991, 65.31096, 67.20985, 69.13358, 
    71.07888, 73.0422, 75.01979, 77.00771, 79.00187, 80.99813, 82.99229, 
    84.98021, 86.9578, 88.92112, 90.86642, 92.79015, 94.68904, 96.56008, 
    98.4006, 100.2082, 101.9809, 103.7169, 105.4148, 107.0736, 108.6923, 
    110.2705, 111.8079, 113.3043, 114.76, 116.1751, 117.5502, 118.8859, 
    120.1828, 121.4417, 122.6636, 123.8494, 125, 126.1165, 127.1998, 
    128.2511, 129.2714, 130.2618, 131.2232, 132.1568, 133.0635, 133.9444, 
    134.8004, 135.6324, 136.4414, 137.2282, 137.9938, 138.7389, 139.4643, 
    140.1709, 140.8594, 141.5304, 142.1847,
  16.8762, 17.51572, 18.17209, 18.84603, 19.53829, 20.24967, 20.98096, 
    21.73304, 22.50677, 23.30309, 24.12295, 24.96733, 25.83727, 26.73381, 
    27.65805, 28.61111, 29.59413, 30.60828, 31.65474, 32.73471, 33.8494, 35, 
    36.1877, 37.41367, 38.67902, 39.98483, 41.3321, 42.72173, 44.15452, 
    45.63113, 47.15206, 48.71761, 50.32788, 51.9827, 53.68164, 55.42397, 
    57.20862, 59.03416, 60.89882, 62.80042, 64.7364, 66.70383, 68.69939, 
    70.71942, 72.75996, 74.81673, 76.88528, 78.96097, 81.03903, 83.11472, 
    85.18327, 87.24004, 89.28058, 91.30061, 93.29617, 95.2636, 97.19958, 
    99.10118, 100.9658, 102.7914, 104.576, 106.3184, 108.0173, 109.6721, 
    111.2824, 112.8479, 114.3689, 115.8455, 117.2783, 118.6679, 120.0152, 
    121.321, 122.5863, 123.8123, 125, 126.1506, 127.2653, 128.3453, 129.3917, 
    130.4059, 131.3889, 132.3419, 133.2662, 134.1627, 135.0327, 135.8771, 
    136.6969, 137.4932, 138.267, 139.019, 139.7503, 140.4617, 141.154, 
    141.8279, 142.4843, 143.1238,
  15.9299, 16.55382, 17.19465, 17.85316, 18.53012, 19.22636, 19.94274, 
    20.68015, 21.43955, 22.22189, 23.02822, 23.85958, 24.71708, 25.60187, 
    26.51514, 27.4581, 28.43203, 29.43821, 30.47797, 31.55266, 32.66364, 
    33.8123, 35, 36.22811, 37.49796, 38.81084, 40.16799, 41.57055, 43.01954, 
    44.51587, 46.06028, 47.65329, 49.29521, 50.98606, 52.72558, 54.51313, 
    56.34774, 58.22799, 60.15207, 62.11768, 64.12208, 66.16206, 68.23397, 
    70.33372, 72.45686, 74.59853, 76.75368, 78.91698, 81.08302, 83.24632, 
    85.40147, 87.54314, 89.66628, 91.76603, 93.83794, 95.87792, 97.88232, 
    99.84793, 101.772, 103.6523, 105.4869, 107.2744, 109.0139, 110.7048, 
    112.3467, 113.9397, 115.4841, 116.9805, 118.4295, 119.832, 121.1892, 
    122.502, 123.7719, 125, 126.1877, 127.3364, 128.4473, 129.522, 130.5618, 
    131.568, 132.5419, 133.4849, 134.3981, 135.2829, 136.1404, 136.9718, 
    137.7781, 138.5605, 139.3198, 140.0573, 140.7736, 141.4699, 142.1469, 
    142.8053, 143.4462, 144.0701,
  14.97656, 15.58404, 16.20846, 16.8506, 17.51126, 18.19131, 18.89165, 
    19.61322, 20.35701, 21.12406, 21.91544, 22.7323, 23.57581, 24.44721, 
    25.34779, 26.27887, 27.24184, 28.23813, 29.2692, 30.33656, 31.44175, 
    32.58633, 33.77189, 35, 36.27223, 37.59011, 38.95514, 40.36873, 41.83219, 
    43.34671, 44.91329, 46.53275, 48.20564, 49.93225, 51.7125, 53.54596, 
    55.43174, 57.36851, 59.35443, 61.38712, 63.46365, 65.58053, 67.73374, 
    69.91871, 72.1304, 74.36336, 76.61176, 78.86954, 81.13046, 83.38824, 
    85.63664, 87.8696, 90.08129, 92.26626, 94.41947, 96.53635, 98.61288, 
    100.6456, 102.6315, 104.5683, 106.454, 108.2875, 110.0677, 111.7944, 
    113.4673, 115.0867, 116.6533, 118.1678, 119.6313, 121.0449, 122.4099, 
    123.7278, 125, 126.2281, 127.4137, 128.5583, 129.6634, 130.7308, 
    131.7619, 132.7582, 133.7211, 134.6522, 135.5528, 136.4242, 137.2677, 
    138.0846, 138.8759, 139.643, 140.3868, 141.1084, 141.8087, 142.4887, 
    143.1494, 143.7915, 144.416, 145.0234,
  14.01629, 14.60653, 15.21367, 15.8385, 16.48187, 17.14467, 17.82784, 
    18.53236, 19.25927, 20.00965, 20.78466, 21.58549, 22.4134, 23.26972, 
    24.15582, 25.07315, 26.0232, 27.00755, 28.02781, 29.08564, 30.18278, 
    31.32098, 32.50204, 33.72777, 35, 36.32053, 37.69115, 39.11358, 40.58944, 
    42.12026, 43.70737, 45.35192, 47.0548, 48.81659, 50.63749, 52.5173, 
    54.45534, 56.45037, 58.50058, 60.60354, 62.75614, 64.95462, 67.19453, 
    69.47079, 71.77771, 74.10908, 76.45824, 78.8182, 81.1818, 83.54176, 
    85.89092, 88.22229, 90.52921, 92.80547, 95.04538, 97.24386, 99.39646, 
    101.4994, 103.5496, 105.5447, 107.4827, 109.3625, 111.1834, 112.9452, 
    114.6481, 116.2926, 117.8797, 119.4106, 120.8864, 122.3088, 123.6795, 
    125, 126.2722, 127.498, 128.679, 129.8172, 130.9144, 131.9722, 132.9924, 
    133.9768, 134.9268, 135.8442, 136.7303, 137.5866, 138.4145, 139.2153, 
    139.9903, 140.7407, 141.4676, 142.1722, 142.8553, 143.5181, 144.1615, 
    144.7863, 145.3935, 145.9837,
  13.04927, 13.62145, 14.21043, 14.81703, 15.44211, 16.0866, 16.75146, 
    17.43771, 18.14644, 18.87879, 19.63594, 20.41919, 21.22985, 22.06932, 
    22.9391, 23.84072, 24.77581, 25.74607, 26.75325, 27.79922, 28.88587, 
    30.01517, 31.18916, 32.40989, 33.67947, 35, 36.37359, 37.80231, 39.28814, 
    40.83299, 42.43859, 44.10649, 45.83797, 47.634, 49.49513, 51.42148, 
    53.41263, 55.46753, 57.58447, 59.76099, 61.99385, 64.27898, 66.61152, 
    68.98579, 71.39537, 73.83317, 76.29155, 78.76245, 81.23755, 83.70845, 
    86.16683, 88.60463, 91.01421, 93.38848, 95.72102, 98.00616, 100.239, 
    102.4155, 104.5325, 106.5874, 108.5785, 110.5049, 112.366, 114.162, 
    115.8935, 117.5614, 119.167, 120.7119, 122.1977, 123.6264, 125, 126.3205, 
    127.5901, 128.8108, 129.9848, 131.1141, 132.2008, 133.2467, 134.2539, 
    135.2242, 136.1593, 137.0609, 137.9307, 138.7702, 139.5808, 140.3641, 
    141.1212, 141.8536, 142.5623, 143.2485, 143.9134, 144.5579, 145.183, 
    145.7896, 146.3785, 146.9507,
  12.07564, 12.62897, 13.19894, 13.78638, 14.39218, 15.01729, 15.66269, 
    16.32946, 17.01871, 17.73161, 18.46943, 19.23349, 20.0252, 20.84604, 
    21.69757, 22.58146, 23.49943, 24.45333, 25.44506, 26.47666, 27.55021, 
    28.66791, 29.83201, 31.04486, 32.30885, 33.62641, 35, 36.43207, 37.92503, 
    39.48121, 41.10281, 42.79184, 44.55008, 46.37894, 48.27946, 50.25218, 
    52.29701, 54.4132, 56.59922, 58.85265, 61.17015, 63.5474, 65.97906, 
    68.4588, 70.97938, 73.53267, 76.10988, 78.70166, 81.29834, 83.89012, 
    86.46733, 89.02062, 91.5412, 94.02094, 96.4526, 98.82985, 101.1473, 
    103.4008, 105.5868, 107.703, 109.7478, 111.7205, 113.6211, 115.4499, 
    117.2082, 118.8972, 120.5188, 122.075, 123.5679, 125, 126.3736, 127.6912, 
    128.9551, 130.168, 131.3321, 132.4498, 133.5233, 134.5549, 135.5467, 
    136.5006, 137.4185, 138.3024, 139.154, 139.9748, 140.7665, 141.5306, 
    142.2684, 142.9813, 143.6705, 144.3373, 144.9827, 145.6078, 146.2136, 
    146.8011, 147.371, 147.9244,
  11.09559, 11.62928, 12.17938, 12.74674, 13.33228, 13.93695, 14.56177, 
    15.20782, 15.87627, 16.56833, 17.2853, 18.02856, 18.79959, 19.59994, 
    20.43126, 21.2953, 22.19392, 23.12908, 24.10286, 25.11744, 26.1751, 
    27.27827, 28.42946, 29.63127, 30.88642, 32.19769, 33.56793, 35, 36.49678, 
    38.06109, 39.69566, 41.40307, 43.18566, 45.04543, 46.98399, 49.0024, 
    51.10109, 53.2797, 55.53698, 57.87068, 60.27742, 62.75264, 65.29052, 
    67.88404, 70.52498, 73.20405, 75.91105, 78.63511, 81.36489, 84.08895, 
    86.79595, 89.47502, 92.11596, 94.70948, 97.24737, 99.72258, 102.1293, 
    104.463, 106.7203, 108.8989, 110.9976, 113.016, 114.9546, 116.8143, 
    118.5969, 120.3043, 121.9389, 123.5032, 125, 126.4321, 127.8023, 
    129.1136, 130.3687, 131.5705, 132.7217, 133.8249, 134.8826, 135.8971, 
    136.8709, 137.8061, 138.7047, 139.5687, 140.4001, 141.2004, 141.9714, 
    142.7147, 143.4317, 144.1237, 144.7922, 145.4382, 146.063, 146.6677, 
    147.2533, 147.8206, 148.3707, 148.9044,
  10.10931, 10.62257, 11.15197, 11.69836, 12.26266, 12.84584, 13.44893, 
    14.07306, 14.71939, 15.38918, 16.08378, 16.80461, 17.55319, 18.33116, 
    19.14024, 19.98227, 20.85923, 21.77319, 22.72637, 23.72113, 24.75996, 
    25.84548, 26.98046, 28.16781, 29.41056, 30.71186, 32.07497, 33.50322, 35, 
    36.56869, 38.21262, 39.93501, 41.73889, 43.62696, 45.60155, 47.66441, 
    49.81659, 52.05832, 54.3888, 56.80604, 59.30675, 61.88618, 64.53806, 
    67.2546, 70.02649, 72.84306, 75.69244, 78.5619, 81.4381, 84.30756, 
    87.15694, 89.97351, 92.7454, 95.46194, 98.11382, 100.6933, 103.194, 
    105.6112, 107.9417, 110.1834, 112.3356, 114.3984, 116.373, 118.2611, 
    120.065, 121.7874, 123.4313, 125, 126.4968, 127.925, 129.2881, 130.5894, 
    131.8322, 133.0195, 134.1545, 135.24, 136.2789, 137.2736, 138.2268, 
    139.1408, 140.0177, 140.8598, 141.6688, 142.4468, 143.1954, 143.9162, 
    144.6108, 145.2806, 145.9269, 146.5511, 147.1542, 147.7373, 148.3016, 
    148.848, 149.3774, 149.8907,
  9.116993, 9.609083, 10.11696, 10.64148, 11.18358, 11.74423, 12.32448, 
    12.92546, 13.54836, 14.19447, 14.86516, 15.5619, 16.28627, 17.03993, 
    17.8247, 18.64251, 19.49541, 20.3856, 21.31545, 22.28746, 23.30432, 
    24.36887, 25.48413, 26.65329, 27.87974, 29.16701, 30.51879, 31.93891, 
    33.43131, 35, 36.64899, 38.38225, 40.20359, 42.11657, 44.12439, 46.22965, 
    48.43428, 50.73925, 53.14442, 55.64827, 58.24773, 60.938, 63.71237, 
    66.56224, 69.47707, 72.44456, 75.45086, 78.48095, 81.51905, 84.54914, 
    87.55544, 90.52293, 93.43776, 96.28763, 99.062, 101.7523, 104.3517, 
    106.8556, 109.2607, 111.5657, 113.7703, 115.8756, 117.8834, 119.7964, 
    121.6178, 123.351, 125, 126.5687, 128.0611, 129.4812, 130.833, 132.1203, 
    133.3467, 134.5159, 135.6311, 136.6957, 137.7125, 138.6846, 139.6144, 
    140.5046, 141.3575, 142.1753, 142.9601, 143.7137, 144.4381, 145.1348, 
    145.8055, 146.4516, 147.0745, 147.6755, 148.2558, 148.8164, 149.3585, 
    149.883, 150.3909, 150.883,
  8.118866, 8.589039, 9.074591, 9.576381, 10.09533, 10.63243, 11.18872, 
    11.76535, 12.36353, 12.98454, 13.6298, 14.3008, 14.99914, 15.72657, 
    16.48493, 17.27624, 18.10262, 18.96641, 19.87008, 20.81628, 21.80788, 
    22.84794, 23.93972, 25.08671, 26.29263, 27.56141, 28.89719, 30.30434, 
    31.78738, 33.35101, 35, 36.73916, 38.57323, 40.50679, 42.54405, 44.68874, 
    46.94384, 49.31137, 51.7921, 54.38524, 57.08818, 59.8962, 62.8023, 
    65.797, 68.8684, 72.00228, 75.1824, 78.39094, 81.60906, 84.8176, 
    87.99772, 91.1316, 94.203, 97.1977, 100.1038, 102.9118, 105.6148, 
    108.2079, 110.6886, 113.0562, 115.3113, 117.4559, 119.4932, 121.4268, 
    123.2608, 125, 126.649, 128.2126, 129.6957, 131.1028, 132.4386, 133.7074, 
    134.9133, 136.0603, 137.1521, 138.1921, 139.1837, 140.1299, 141.0336, 
    141.8974, 142.7238, 143.5151, 144.2734, 145.0009, 145.6992, 146.3702, 
    147.0155, 147.6365, 148.2346, 148.8113, 149.3676, 149.9047, 150.4236, 
    150.9254, 151.411, 151.8811,
  7.115152, 7.562692, 8.025139, 8.503347, 8.998231, 9.510773, 10.04203, 
    10.59312, 11.16528, 11.7598, 12.3781, 13.0217, 13.69223, 14.39146, 
    15.1213, 15.8838, 16.68118, 17.51585, 18.39039, 19.30761, 20.27052, 
    21.28238, 22.3467, 23.46725, 24.64808, 25.89351, 27.20815, 28.59693, 
    30.06499, 31.61775, 33.26084, 35, 36.84104, 38.78968, 40.85144, 43.03135, 
    45.33379, 47.76212, 50.31837, 53.00285, 55.81371, 58.74662, 61.79439, 
    64.94675, 68.19027, 71.50849, 74.88224, 78.29022, 81.70978, 85.11776, 
    88.49151, 91.80973, 95.05325, 98.20561, 101.2534, 104.1863, 106.9972, 
    109.6816, 112.2379, 114.6662, 116.9687, 119.1486, 121.2103, 123.159, 125, 
    126.7392, 128.3822, 129.935, 131.4031, 132.7918, 134.1065, 135.3519, 
    136.5327, 137.6533, 138.7176, 139.7295, 140.6924, 141.6096, 142.4841, 
    143.3188, 144.1162, 144.8787, 145.6085, 146.3078, 146.9783, 147.6219, 
    148.2402, 148.8347, 149.4069, 149.958, 150.4892, 151.0018, 151.4967, 
    151.9749, 152.4373, 152.8848,
  6.106095, 6.530308, 6.968895, 7.422698, 7.892619, 8.379629, 8.884773, 
    9.409175, 9.954047, 10.5207, 11.11054, 11.7251, 12.36602, 13.03511, 
    13.73428, 14.46565, 15.2315, 16.03428, 16.8767, 17.76165, 18.69232, 
    19.67212, 20.70479, 21.79436, 22.9452, 24.16203, 25.44992, 26.81434, 
    28.26111, 29.79641, 31.42676, 33.15896, 35, 36.95695, 39.03682, 41.24627, 
    43.5914, 46.07734, 48.70781, 51.48467, 54.40734, 57.47225, 60.67233, 
    63.99661, 67.43004, 70.95351, 74.5443, 78.17673, 81.82327, 85.4557, 
    89.04649, 92.56996, 96.00339, 99.32767, 102.5277, 105.5927, 108.5153, 
    111.2922, 113.9227, 116.4086, 118.7537, 120.9632, 123.043, 125, 126.841, 
    128.5732, 130.2036, 131.7389, 133.1857, 134.5501, 135.838, 137.0548, 
    138.2056, 139.2952, 140.3279, 141.3077, 142.2383, 143.1233, 143.9657, 
    144.7685, 145.5343, 146.2657, 146.9649, 147.634, 148.2749, 148.8895, 
    149.4793, 150.046, 150.5908, 151.1152, 151.6204, 152.1074, 152.5773, 
    153.0311, 153.4697, 153.8939,
  5.091947, 5.492166, 5.906166, 6.334769, 6.77886, 7.239392, 7.717392, 
    8.213969, 8.730321, 9.267746, 9.827646, 10.41155, 11.0211, 11.65809, 
    12.32448, 13.0224, 13.75415, 14.52226, 15.32948, 16.17882, 17.07357, 
    18.0173, 19.01393, 20.06775, 21.18341, 22.366, 23.62106, 24.95457, 
    26.37304, 27.88343, 29.49321, 31.21031, 33.04305, 35, 37.08991, 39.3214, 
    41.70267, 44.24112, 46.94274, 49.81158, 52.84893, 56.05262, 59.41615, 
    62.92815, 66.57185, 70.32514, 74.16086, 78.04782, 81.95218, 85.83914, 
    89.67486, 93.42815, 97.07185, 100.5838, 103.9474, 107.1511, 110.1884, 
    113.0573, 115.7589, 118.2973, 120.6786, 122.9101, 125, 126.957, 128.7897, 
    130.5068, 132.1166, 133.627, 135.0454, 136.3789, 137.634, 138.8166, 
    139.9323, 140.9861, 141.9827, 142.9264, 143.8212, 144.6705, 145.4777, 
    146.2458, 146.9776, 147.6755, 148.3419, 148.9789, 149.5885, 150.1723, 
    150.7323, 151.2697, 151.786, 152.2826, 152.7606, 153.2211, 153.6652, 
    154.0938, 154.5078, 154.9081,
  4.072974, 4.448562, 4.837277, 5.239919, 5.657345, 6.090485, 6.540341, 
    7.007998, 7.494629, 8.001512, 8.530026, 9.08168, 9.65811, 10.2611, 
    10.8926, 11.55474, 12.24985, 12.98048, 13.74942, 14.55974, 15.41482, 
    16.31836, 17.27442, 18.2875, 19.36251, 20.50487, 21.72053, 23.01601, 
    24.39845, 25.87561, 27.45595, 29.14856, 30.96318, 32.91009, 35, 37.24382, 
    39.65233, 42.23573, 45.00304, 47.96128, 51.11454, 54.46289, 58.00124, 
    61.71825, 65.59562, 69.60771, 73.72196, 77.90008, 82.09992, 86.27804, 
    90.39229, 94.40438, 98.28175, 101.9988, 105.5371, 108.8855, 112.0387, 
    114.997, 117.7643, 120.3477, 122.7562, 125, 127.0899, 129.0368, 130.8514, 
    132.5441, 134.1244, 135.6015, 136.984, 138.2795, 139.4951, 140.6375, 
    141.7125, 142.7256, 143.6816, 144.5852, 145.4403, 146.2506, 147.0195, 
    147.7502, 148.4453, 149.1074, 149.7389, 150.3419, 150.9183, 151.47, 
    151.9985, 152.5054, 152.992, 153.4597, 153.9095, 154.3427, 154.7601, 
    155.1627, 155.5514, 155.927,
  3.049454, 3.399804, 3.762572, 4.138524, 4.528489, 4.933362, 5.354114, 
    5.791796, 6.247549, 6.722614, 7.218343, 7.736207, 8.277816, 8.844927, 
    9.439466, 10.06355, 10.71948, 11.40983, 12.13739, 12.90528, 13.71689, 
    14.57603, 15.48687, 16.45404, 17.48269, 18.57852, 19.74782, 20.9976, 
    22.3356, 23.77035, 25.31126, 26.96865, 28.75373, 30.6786, 32.75618, 35, 
    37.4239, 40.04157, 42.86588, 45.90788, 49.17569, 52.6729, 56.39701, 
    60.33771, 64.47548, 68.78084, 73.21452, 77.72898, 82.27102, 86.78548, 
    91.21916, 95.52452, 99.66229, 103.603, 107.3271, 110.8243, 114.0921, 
    117.1341, 119.9584, 122.5761, 125, 127.2438, 129.3214, 131.2463, 
    133.0314, 134.6887, 136.2296, 137.6644, 139.0024, 140.2522, 141.4215, 
    142.5173, 143.546, 144.5131, 145.424, 146.2831, 147.0947, 147.8626, 
    148.5902, 149.2805, 149.9364, 150.5605, 151.1551, 151.7222, 152.2638, 
    152.7817, 153.2774, 153.7525, 154.2082, 154.6459, 155.0666, 155.4715, 
    155.8615, 156.2374, 156.6002, 156.9505,
  2.021674, 2.346215, 2.682407, 3.030981, 3.392728, 3.768503, 4.159237, 
    4.565938, 4.989704, 5.43173, 5.893324, 6.37591, 6.881052, 7.410462, 
    7.966022, 8.549803, 9.164087, 9.811396, 10.49452, 11.21654, 11.98089, 
    12.79138, 13.65226, 14.56826, 15.54466, 16.58737, 17.70299, 18.89891, 
    20.18341, 21.56572, 23.05616, 24.66621, 26.4086, 28.29732, 30.34767, 
    32.5761, 35, 37.63727, 40.50561, 43.62146, 46.99852, 50.64579, 54.56522, 
    58.74911, 63.17771, 67.8175, 72.62102, 77.52846, 82.47154, 87.37898, 
    92.1825, 96.8223, 101.2509, 105.4348, 109.3542, 113.0015, 116.3785, 
    119.4944, 122.3627, 125, 127.4239, 129.6523, 131.7027, 133.5914, 
    135.3338, 136.9438, 138.4343, 139.8166, 141.1011, 142.297, 143.4126, 
    144.4553, 145.4317, 146.3477, 147.2086, 148.0191, 148.7835, 149.5055, 
    150.1886, 150.8359, 151.4502, 152.034, 152.5895, 153.1189, 153.6241, 
    154.1067, 154.5683, 155.0103, 155.4341, 155.8408, 156.2315, 156.6073, 
    156.969, 157.3176, 157.6538, 157.9783,
  0.989933, 1.28813, 1.597158, 1.917706, 2.250523, 2.596416, 2.956268, 
    3.331035, 3.721762, 4.129589, 4.555761, 5.001646, 5.468743, 5.9587, 
    6.473334, 7.01465, 7.584867, 8.186443, 8.822109, 9.494904, 10.20822, 
    10.96584, 11.77201, 12.63149, 13.54963, 14.53247, 15.5868, 16.7203, 
    17.94168, 19.26074, 20.68863, 22.23788, 23.92266, 25.75888, 27.76427, 
    29.95843, 32.36273, 35, 37.89388, 41.06774, 44.54297, 48.33653, 52.45767, 
    56.90404, 61.65757, 66.6812, 71.91743, 77.29012, 82.70988, 88.08257, 
    93.3188, 98.34243, 103.096, 107.5423, 111.6635, 115.457, 118.9323, 
    122.1061, 125, 127.6373, 130.0416, 132.2357, 134.2411, 136.0773, 
    137.7621, 139.3114, 140.7393, 142.0583, 143.2797, 144.4132, 145.4675, 
    146.4504, 147.3685, 148.228, 149.0342, 149.7918, 150.5051, 151.1779, 
    151.8136, 152.4151, 152.9854, 153.5267, 154.0413, 154.5312, 154.9984, 
    155.4442, 155.8704, 156.2782, 156.669, 157.0437, 157.4036, 157.7495, 
    158.0823, 158.4028, 158.7119, 159.0101,
  359.9545, 0.2258954, 0.5072123, 0.7991334, 1.102355, 1.417635, 1.745796, 
    2.087737, 2.444437, 2.816969, 3.206508, 3.614345, 4.041899, 4.490737, 
    4.962586, 5.459363, 5.983191, 6.536436, 7.121729, 7.742018, 8.4006, 
    9.101182, 9.847935, 10.64557, 11.49942, 12.41553, 13.40078, 14.46302, 
    15.6112, 16.85558, 18.2079, 19.68163, 21.29219, 23.05726, 24.99696, 
    27.13412, 29.49439, 32.10612, 35, 38.20808, 41.76202, 45.6902, 50.01339, 
    54.73909, 59.85475, 65.32144, 71.06998, 77.00205, 82.99795, 88.93002, 
    94.67856, 100.1452, 105.2609, 109.9866, 114.3098, 118.238, 121.7919, 125, 
    127.8939, 130.5056, 132.8659, 135.003, 136.9427, 138.7078, 140.3184, 
    141.7921, 143.1444, 144.3888, 145.537, 146.5992, 147.5845, 148.5006, 
    149.3544, 150.1521, 150.8988, 151.5994, 152.258, 152.8783, 153.4636, 
    154.0168, 154.5406, 155.0374, 155.5093, 155.9581, 156.3857, 156.7935, 
    157.183, 157.5556, 157.9123, 158.2542, 158.5824, 158.8976, 159.2009, 
    159.4928, 159.7741, 160.0455,
  358.9158, 359.1599, 359.413, 359.6757, 359.9487, 0.2327171, 0.5284402, 
    0.8367262, 1.158482, 1.494702, 1.846476, 2.215007, 2.601616, 3.007768, 
    3.435082, 3.885358, 4.360597, 4.863032, 5.395164, 5.959797, 6.560083, 
    7.199584, 7.882326, 8.612883, 9.396461, 10.23901, 11.14735, 12.12932, 
    13.19396, 14.35173, 15.61476, 16.99715, 18.51533, 20.18842, 22.03872, 
    24.09212, 26.37854, 28.93226, 31.79192, 35, 38.60137, 42.64027, 47.1551, 
    52.17041, 57.68631, 63.66663, 70.02966, 76.6468, 83.3532, 89.97034, 
    96.33337, 102.3137, 107.8296, 112.8449, 117.3597, 121.3986, 125, 
    128.2081, 131.0677, 133.6215, 135.9079, 137.9613, 139.8116, 141.4847, 
    143.0029, 144.3852, 145.6483, 146.806, 147.8707, 148.8526, 149.761, 
    150.6035, 151.3871, 152.1177, 152.8004, 153.4399, 154.0402, 154.6048, 
    155.137, 155.6394, 156.1146, 156.5649, 156.9922, 157.3984, 157.785, 
    158.1535, 158.5053, 158.8415, 159.1633, 159.4716, 159.7673, 160.0513, 
    160.3243, 160.587, 160.8401, 161.0842,
  357.8741, 358.0904, 358.3148, 358.5479, 358.7902, 359.0422, 359.3048, 
    359.5787, 359.8647, 0.1636643, 0.4766341, 0.8046976, 1.149067, 1.511083, 
    1.892236, 2.294184, 2.718776, 3.168084, 3.644429, 4.15043, 4.689038, 
    5.263601, 5.877925, 6.536353, 7.243857, 8.006155, 8.829846, 9.722579, 
    10.69325, 11.75227, 12.91182, 14.18629, 15.59266, 17.15107, 18.88546, 
    20.82431, 23.00148, 25.45703, 28.23798, 31.39863, 35, 39.10745, 43.7852, 
    49.08622, 55.03613, 61.6122, 68.72269, 76.1976, 83.8024, 91.27731, 
    98.3878, 104.9639, 110.9138, 116.2148, 120.8926, 125, 128.6014, 131.762, 
    134.543, 136.9985, 139.1757, 141.1145, 142.8489, 144.4073, 145.8137, 
    147.0882, 148.2477, 149.3067, 150.2774, 151.1702, 151.9939, 152.7561, 
    153.4637, 154.1221, 154.7364, 155.311, 155.8496, 156.3556, 156.8319, 
    157.2812, 157.7058, 158.1078, 158.4889, 158.8509, 159.1953, 159.5234, 
    159.8363, 160.1353, 160.4213, 160.6952, 160.9578, 161.2098, 161.4521, 
    161.6852, 161.9096, 162.1259,
  356.8297, 357.0179, 357.2133, 357.4162, 357.6272, 357.8468, 358.0757, 
    358.3145, 358.5639, 358.8248, 359.098, 359.3846, 359.6855, 0.002061171, 
    0.3355702, 0.6875198, 1.05958, 1.453624, 1.87176, 2.31637, 2.790152, 
    3.296174, 3.837941, 4.419468, 5.045379, 5.721019, 6.452599, 7.247366, 
    8.113825, 9.062004, 10.1038, 11.25338, 12.52775, 13.94739, 15.53711, 
    17.3271, 19.35421, 21.66347, 24.3098, 27.35973, 30.89255, 35, 39.78226, 
    45.33723, 51.73862, 59.00039, 67.03291, 75.61138, 84.38862, 92.96709, 
    100.9996, 108.2614, 114.6628, 120.2177, 125, 129.1075, 132.6403, 
    135.6902, 138.3365, 140.6458, 142.6729, 144.4629, 146.0526, 147.4723, 
    148.7466, 149.8962, 150.938, 151.8862, 152.7526, 153.5474, 154.279, 
    154.9546, 155.5805, 156.1621, 156.7038, 157.2099, 157.6836, 158.1282, 
    158.5464, 158.9404, 159.3125, 159.6644, 159.9979, 160.3145, 160.6154, 
    160.902, 161.1752, 161.4361, 161.6855, 161.9243, 162.1532, 162.3728, 
    162.5838, 162.7867, 162.9821, 163.1703,
  355.7829, 355.9428, 356.1087, 356.2811, 356.4604, 356.6471, 356.8416, 
    357.0447, 357.257, 357.479, 357.7116, 357.9557, 358.2122, 358.4822, 
    358.7667, 359.0672, 359.385, 359.7219, 0.07960072, 0.4603243, 0.8664198, 
    1.300613, 1.766029, 2.266261, 2.805467, 3.388479, 4.02094, 4.709482, 
    5.461938, 6.287628, 7.197704, 8.20561, 9.32767, 10.58385, 11.99876, 
    13.60299, 15.43478, 17.54233, 19.9866, 22.8449, 26.2148, 30.21773, 35, 
    40.72601, 47.55444, 55.58445, 64.7672, 74.81406, 85.18594, 95.2328, 
    104.4156, 112.4456, 119.274, 125, 129.7823, 133.7852, 137.1551, 140.0134, 
    142.4577, 144.5652, 146.397, 148.0012, 149.4162, 150.6723, 151.7944, 
    152.8023, 153.7124, 154.5381, 155.2905, 155.9791, 156.6115, 157.1945, 
    157.7337, 158.234, 158.6994, 159.1336, 159.5397, 159.9204, 160.2781, 
    160.615, 160.9328, 161.2333, 161.5178, 161.7878, 162.0443, 162.2883, 
    162.521, 162.743, 162.9553, 163.1584, 163.353, 163.5396, 163.7189, 
    163.8913, 164.0572, 164.2171,
  354.7342, 354.8654, 355.0016, 355.1431, 355.2903, 355.4436, 355.6035, 
    355.7703, 355.9448, 356.1273, 356.3187, 356.5195, 356.7307, 356.9529, 
    357.1873, 357.435, 357.6972, 357.9752, 358.2706, 358.5852, 358.9211, 
    359.2806, 359.6663, 0.08128966, 0.5292088, 1.014209, 1.541195, 2.115962, 
    2.745399, 3.43776, 4.203004, 5.053253, 6.003388, 7.071855, 8.281747, 
    9.662291, 11.25089, 13.09596, 15.26091, 17.82959, 20.91378, 24.66276, 
    29.27399, 35, 42.1372, 50.96407, 61.58201, 73.6667, 86.3333, 98.41799, 
    109.0359, 117.8628, 125, 130.726, 135.3372, 139.0862, 142.1704, 144.7391, 
    146.904, 148.7491, 150.3377, 151.7182, 152.9281, 153.9966, 154.9467, 
    155.797, 156.5622, 157.2546, 157.884, 158.4588, 158.9858, 159.4708, 
    159.9187, 160.3337, 160.7194, 161.0789, 161.4148, 161.7294, 162.0248, 
    162.3028, 162.565, 162.8126, 163.0471, 163.2693, 163.4805, 163.6813, 
    163.8727, 164.0552, 164.2297, 164.3966, 164.5564, 164.7097, 164.8569, 
    164.9984, 165.1346, 165.2658,
  353.6839, 353.7861, 353.8923, 354.0027, 354.1175, 354.2371, 354.3618, 
    354.4921, 354.6282, 354.7708, 354.9203, 355.0772, 355.2422, 355.416, 
    355.5993, 355.7931, 355.9983, 356.216, 356.4475, 356.6942, 356.9578, 
    357.2401, 357.5432, 357.8696, 358.2223, 358.6046, 359.0206, 359.475, 
    359.9735, 0.5229301, 1.131602, 1.809731, 2.569962, 3.428143, 4.404378, 
    5.524519, 6.822294, 8.342426, 10.14525, 12.31369, 14.96387, 18.26138, 
    22.44556, 27.8628, 35, 44.47124, 56.81278, 71.87518, 88.12482, 103.1872, 
    115.5288, 125, 132.1372, 137.5544, 141.7386, 145.0361, 147.6863, 
    149.8548, 151.6576, 153.1777, 154.4755, 155.5956, 156.5719, 157.43, 
    158.1903, 158.8684, 159.4771, 160.0265, 160.525, 160.9794, 161.3954, 
    161.7777, 162.1304, 162.4568, 162.7599, 163.0422, 163.3058, 163.5525, 
    163.784, 164.0017, 164.2069, 164.4007, 164.584, 164.7578, 164.9228, 
    165.0797, 165.2292, 165.3718, 165.5079, 165.6382, 165.7629, 165.8825, 
    165.9973, 166.1077, 166.2139, 166.3161,
  352.6322, 352.7054, 352.7814, 352.8604, 352.9426, 353.0282, 353.1175, 
    353.2108, 353.3083, 353.4105, 353.5175, 353.63, 353.7483, 353.8729, 
    354.0044, 354.1435, 354.2908, 354.4471, 354.6134, 354.7907, 354.9802, 
    355.1833, 355.4015, 355.6366, 355.8909, 356.1668, 356.4673, 356.796, 
    357.157, 357.5555, 357.9977, 358.4915, 359.0465, 359.6749, 0.3922898, 
    1.219163, 2.182494, 3.318798, 4.678558, 6.333375, 8.387803, 10.99961, 
    14.41555, 19.03593, 25.52876, 35, 49.04179, 68.69369, 91.30631, 110.9582, 
    125, 134.4712, 140.9641, 145.5845, 149.0004, 151.6122, 153.6666, 
    155.3214, 156.6812, 157.8175, 158.7808, 159.6077, 160.3251, 160.9535, 
    161.5085, 162.0023, 162.4445, 162.843, 163.204, 163.5327, 163.8332, 
    164.1091, 164.3634, 164.5985, 164.8167, 165.0198, 165.2093, 165.3866, 
    165.5529, 165.7092, 165.8565, 165.9956, 166.1271, 166.2517, 166.37, 
    166.4825, 166.5895, 166.6917, 166.7892, 166.8825, 166.9718, 167.0574, 
    167.1396, 167.2186, 167.2946, 167.3678,
  351.5797, 351.6237, 351.6693, 351.7168, 351.7661, 351.8176, 351.8713, 
    351.9273, 351.986, 352.0474, 352.1118, 352.1794, 352.2505, 352.3255, 
    352.4046, 352.4883, 352.577, 352.6711, 352.7713, 352.8781, 352.9923, 
    353.1147, 353.2463, 353.3882, 353.5418, 353.7085, 353.8901, 354.089, 
    354.3076, 354.5491, 354.8176, 355.1178, 355.4557, 355.8391, 356.278, 
    356.7855, 357.379, 358.0826, 358.93, 359.9703, 1.277307, 2.967087, 
    5.232795, 8.417991, 13.18722, 20.95822, 35, 61.56694, 98.43307, 125, 
    139.0418, 146.8128, 151.582, 154.7672, 157.0329, 158.7227, 160.0297, 
    161.07, 161.9174, 162.621, 163.2145, 163.722, 164.1609, 164.5443, 
    164.8822, 165.1824, 165.4509, 165.6924, 165.9111, 166.1099, 166.2915, 
    166.4582, 166.6118, 166.7537, 166.8853, 167.0077, 167.1219, 167.2287, 
    167.3289, 167.423, 167.5117, 167.5954, 167.6745, 167.7495, 167.8206, 
    167.8882, 167.9526, 168.014, 168.0727, 168.1287, 168.1824, 168.2339, 
    168.2832, 168.3307, 168.3763, 168.4203,
  350.5266, 350.5413, 350.5565, 350.5724, 350.5888, 350.606, 350.6239, 
    350.6426, 350.6621, 350.6826, 350.7041, 350.7267, 350.7505, 350.7755, 
    350.8019, 350.8298, 350.8594, 350.8908, 350.9243, 350.96, 350.9981, 
    351.039, 351.083, 351.1305, 351.1818, 351.2375, 351.2983, 351.3649, 
    351.4381, 351.519, 351.6091, 351.7098, 351.8233, 351.9522, 352.0999, 
    352.271, 352.4716, 352.7099, 352.998, 353.3532, 353.8024, 354.3886, 
    355.1859, 356.3333, 358.1248, 1.30631, 8.433065, 35, 125, 151.5669, 
    158.6937, 161.8752, 163.6667, 164.8141, 165.6114, 166.1976, 166.6468, 
    167.0021, 167.2901, 167.5285, 167.729, 167.9001, 168.0478, 168.1767, 
    168.2902, 168.3909, 168.4809, 168.5619, 168.6351, 168.7017, 168.7625, 
    168.8182, 168.8695, 168.917, 168.961, 169.0019, 169.04, 169.0757, 
    169.1091, 169.1406, 169.1702, 169.1981, 169.2245, 169.2496, 169.2733, 
    169.2959, 169.3174, 169.3378, 169.3574, 169.3761, 169.394, 169.4112, 
    169.4277, 169.4435, 169.4587, 169.4734,
  349.4734, 349.4587, 349.4435, 349.4276, 349.4112, 349.394, 349.3761, 
    349.3574, 349.3379, 349.3174, 349.2959, 349.2733, 349.2495, 349.2245, 
    349.1981, 349.1702, 349.1406, 349.1092, 349.0757, 349.04, 349.0019, 
    348.961, 348.917, 348.8695, 348.8182, 348.7625, 348.7017, 348.6351, 
    348.5619, 348.481, 348.3909, 348.2902, 348.1767, 348.0478, 347.9001, 
    347.729, 347.5284, 347.2901, 347.002, 346.6468, 346.1976, 345.6114, 
    344.8141, 343.6667, 341.8752, 338.6937, 331.5669, 305, 215, 188.4331, 
    181.3063, 178.1248, 176.3333, 175.1859, 174.3886, 173.8024, 173.3532, 
    172.9979, 172.7099, 172.4715, 172.271, 172.0999, 171.9522, 171.8233, 
    171.7098, 171.6091, 171.5191, 171.4381, 171.3649, 171.2983, 171.2375, 
    171.1818, 171.1305, 171.083, 171.039, 170.9981, 170.96, 170.9243, 
    170.8909, 170.8594, 170.8298, 170.8019, 170.7755, 170.7504, 170.7267, 
    170.7041, 170.6826, 170.6622, 170.6426, 170.6239, 170.606, 170.5888, 
    170.5723, 170.5565, 170.5413, 170.5266,
  348.4203, 348.3763, 348.3307, 348.2832, 348.2339, 348.1824, 348.1287, 
    348.0727, 348.014, 347.9526, 347.8882, 347.8206, 347.7495, 347.6745, 
    347.5954, 347.5117, 347.423, 347.3289, 347.2287, 347.1219, 347.0077, 
    346.8853, 346.7537, 346.6118, 346.4582, 346.2915, 346.1099, 345.911, 
    345.6924, 345.4509, 345.1824, 344.8822, 344.5443, 344.1609, 343.722, 
    343.2145, 342.621, 341.9174, 341.07, 340.0297, 338.7227, 337.0329, 
    334.7672, 331.582, 326.8128, 319.0418, 305, 278.4331, 241.5669, 215, 
    200.9582, 193.1872, 188.418, 185.2328, 182.9671, 181.2773, 179.9703, 
    178.93, 178.0826, 177.379, 176.7855, 176.278, 175.8391, 175.4557, 
    175.1178, 174.8176, 174.5491, 174.3076, 174.0889, 173.8901, 173.7085, 
    173.5418, 173.3882, 173.2463, 173.1147, 172.9923, 172.8781, 172.7713, 
    172.6711, 172.577, 172.4883, 172.4046, 172.3255, 172.2505, 172.1794, 
    172.1118, 172.0474, 171.986, 171.9273, 171.8713, 171.8176, 171.7661, 
    171.7168, 171.6693, 171.6237, 171.5797,
  347.3678, 347.2946, 347.2186, 347.1396, 347.0574, 346.9718, 346.8825, 
    346.7892, 346.6917, 346.5895, 346.4825, 346.37, 346.2517, 346.1271, 
    345.9956, 345.8565, 345.7092, 345.5529, 345.3866, 345.2093, 345.0198, 
    344.8167, 344.5985, 344.3634, 344.1091, 343.8332, 343.5327, 343.204, 
    342.843, 342.4445, 342.0023, 341.5085, 340.9535, 340.3251, 339.6077, 
    338.7808, 337.8175, 336.6812, 335.3214, 333.6666, 331.6122, 329.0004, 
    325.5844, 320.9641, 314.4712, 305, 290.9582, 271.3063, 248.6937, 
    229.0418, 215, 205.5288, 199.0359, 194.4155, 190.9996, 188.3878, 
    186.3334, 184.6786, 183.3188, 182.1825, 181.2192, 180.3923, 179.6749, 
    179.0465, 178.4915, 177.9977, 177.5555, 177.157, 176.796, 176.4673, 
    176.1668, 175.8909, 175.6366, 175.4015, 175.1833, 174.9802, 174.7907, 
    174.6134, 174.4471, 174.2908, 174.1435, 174.0044, 173.8729, 173.7483, 
    173.63, 173.5175, 173.4105, 173.3083, 173.2108, 173.1175, 173.0282, 
    172.9426, 172.8604, 172.7814, 172.7054, 172.6322,
  346.3161, 346.2139, 346.1077, 345.9973, 345.8825, 345.7629, 345.6382, 
    345.5079, 345.3718, 345.2292, 345.0797, 344.9228, 344.7578, 344.584, 
    344.4007, 344.2069, 344.0017, 343.784, 343.5525, 343.3058, 343.0422, 
    342.7599, 342.4568, 342.1304, 341.7777, 341.3954, 340.9794, 340.525, 
    340.0265, 339.4771, 338.8684, 338.1903, 337.43, 336.5719, 335.5956, 
    334.4755, 333.1777, 331.6576, 329.8547, 327.6863, 325.0361, 321.7386, 
    317.5544, 312.1372, 305, 295.5288, 283.1872, 268.1248, 251.8752, 
    236.8128, 224.4712, 215, 207.8628, 202.4456, 198.2614, 194.9639, 
    192.3137, 190.1452, 188.3424, 186.8223, 185.5245, 184.4044, 183.4281, 
    182.57, 181.8097, 181.1316, 180.5229, 179.9735, 179.475, 179.0206, 
    178.6046, 178.2223, 177.8696, 177.5432, 177.2401, 176.9578, 176.6942, 
    176.4475, 176.216, 175.9983, 175.7931, 175.5993, 175.416, 175.2422, 
    175.0772, 174.9203, 174.7708, 174.6282, 174.4921, 174.3618, 174.2371, 
    174.1175, 174.0027, 173.8923, 173.7861, 173.6839,
  345.2658, 345.1346, 344.9984, 344.8569, 344.7097, 344.5564, 344.3965, 
    344.2297, 344.0552, 343.8727, 343.6813, 343.4805, 343.2693, 343.0471, 
    342.8127, 342.565, 342.3028, 342.0248, 341.7294, 341.4148, 341.0789, 
    340.7194, 340.3337, 339.9187, 339.4708, 338.9858, 338.4588, 337.884, 
    337.2546, 336.5622, 335.797, 334.9467, 333.9966, 332.9281, 331.7183, 
    330.3377, 328.7491, 326.904, 324.7391, 322.1704, 319.0862, 315.3372, 
    310.726, 305, 297.8628, 289.0359, 278.418, 266.3333, 253.6667, 241.582, 
    230.9641, 222.1372, 215, 209.274, 204.6628, 200.9138, 197.8296, 195.2609, 
    193.096, 191.2509, 189.6623, 188.2818, 187.0719, 186.0034, 185.0533, 
    184.203, 183.4378, 182.7454, 182.116, 181.5412, 181.0142, 180.5292, 
    180.0813, 179.6663, 179.2806, 178.9211, 178.5852, 178.2706, 177.9752, 
    177.6972, 177.435, 177.1874, 176.9529, 176.7307, 176.5195, 176.3187, 
    176.1273, 175.9448, 175.7703, 175.6034, 175.4436, 175.2903, 175.1431, 
    175.0016, 174.8654, 174.7342,
  344.2171, 344.0572, 343.8913, 343.7189, 343.5396, 343.3529, 343.1584, 
    342.9553, 342.743, 342.521, 342.2884, 342.0443, 341.7878, 341.5178, 
    341.2333, 340.9328, 340.615, 340.2781, 339.9204, 339.5397, 339.1336, 
    338.6994, 338.234, 337.7337, 337.1945, 336.6115, 335.9791, 335.2905, 
    334.5381, 333.7124, 332.8023, 331.7944, 330.6723, 329.4161, 328.0012, 
    326.397, 324.5652, 322.4577, 320.0134, 317.1551, 313.7852, 309.7823, 305, 
    299.274, 292.4456, 284.4156, 275.2328, 265.1859, 254.8141, 244.7672, 
    235.5845, 227.5544, 220.726, 215, 210.2177, 206.2148, 202.8449, 199.9866, 
    197.5423, 195.4348, 193.603, 191.9988, 190.5838, 189.3277, 188.2056, 
    187.1977, 186.2876, 185.4619, 184.7095, 184.0209, 183.3885, 182.8055, 
    182.2663, 181.766, 181.3006, 180.8664, 180.4603, 180.0796, 179.7219, 
    179.385, 179.0672, 178.7667, 178.4822, 178.2122, 177.9557, 177.7117, 
    177.479, 177.257, 177.0447, 176.8416, 176.647, 176.4604, 176.2811, 
    176.1087, 175.9428, 175.7829,
  343.1703, 342.9821, 342.7867, 342.5838, 342.3728, 342.1532, 341.9243, 
    341.6855, 341.4361, 341.1752, 340.902, 340.6154, 340.3145, 339.9979, 
    339.6644, 339.3125, 338.9404, 338.5464, 338.1282, 337.6836, 337.2098, 
    336.7038, 336.162, 335.5805, 334.9546, 334.279, 333.5474, 332.7526, 
    331.8862, 330.938, 329.8962, 328.7466, 327.4723, 326.0526, 324.4629, 
    322.6729, 320.6458, 318.3365, 315.6902, 312.6403, 309.1075, 305, 
    300.2177, 294.6628, 288.2614, 280.9996, 272.9671, 264.3886, 255.6114, 
    247.0329, 239.0004, 231.7386, 225.3372, 219.7823, 215, 210.8925, 
    207.3597, 204.3098, 201.6635, 199.3542, 197.3271, 195.5371, 193.9474, 
    192.5277, 191.2534, 190.1038, 189.062, 188.1138, 187.2474, 186.4526, 
    185.721, 185.0454, 184.4195, 183.8379, 183.2962, 182.7901, 182.3164, 
    181.8718, 181.4536, 181.0596, 180.6875, 180.3356, 180.0021, 179.6855, 
    179.3846, 179.098, 178.8248, 178.5639, 178.3145, 178.0757, 177.8468, 
    177.6272, 177.4162, 177.2133, 177.0179, 176.8297,
  342.1259, 341.9096, 341.6852, 341.4521, 341.2098, 340.9578, 340.6952, 
    340.4213, 340.1353, 339.8363, 339.5234, 339.1953, 338.8509, 338.4889, 
    338.1078, 337.7058, 337.2812, 336.8319, 336.3556, 335.8496, 335.311, 
    334.7364, 334.1221, 333.4637, 332.7561, 331.9938, 331.1702, 330.2774, 
    329.3068, 328.2477, 327.0882, 325.8137, 324.4073, 322.8489, 321.1145, 
    319.1757, 316.9985, 314.543, 311.762, 308.6014, 305, 300.8925, 296.2148, 
    290.9138, 284.9639, 278.3878, 271.2773, 263.8024, 256.1976, 248.7227, 
    241.6122, 235.0361, 229.0862, 223.7852, 219.1075, 215, 211.3986, 208.238, 
    205.457, 203.0015, 200.8243, 198.8855, 197.1511, 195.5927, 194.1863, 
    192.9118, 191.7523, 190.6933, 189.7226, 188.8298, 188.0061, 187.2439, 
    186.5363, 185.8779, 185.2636, 184.689, 184.1504, 183.6444, 183.1681, 
    182.7188, 182.2942, 181.8922, 181.5111, 181.1491, 180.8047, 180.4766, 
    180.1637, 179.8647, 179.5787, 179.3048, 179.0422, 178.7902, 178.5479, 
    178.3148, 178.0904, 177.8741,
  341.0842, 340.8401, 340.587, 340.3243, 340.0513, 339.7673, 339.4716, 
    339.1633, 338.8415, 338.5053, 338.1535, 337.785, 337.3984, 336.9922, 
    336.5649, 336.1147, 335.6394, 335.137, 334.6048, 334.0402, 333.4399, 
    332.8004, 332.1177, 331.3871, 330.6035, 329.761, 328.8527, 327.8707, 
    326.806, 325.6483, 324.3853, 323.0028, 321.4847, 319.8116, 317.9613, 
    315.9079, 313.6215, 311.0677, 308.2081, 305, 301.3986, 297.3597, 
    292.8449, 287.8296, 282.3137, 276.3334, 269.9703, 263.3532, 256.6468, 
    250.0297, 243.6666, 237.6863, 232.1704, 227.1551, 222.6403, 218.6014, 
    215, 211.7919, 208.9323, 206.3785, 204.0921, 202.0387, 200.1884, 
    198.5153, 196.9971, 195.6148, 194.3517, 193.194, 192.1293, 191.1474, 
    190.239, 189.3965, 188.6129, 187.8823, 187.1996, 186.5601, 185.9598, 
    185.3952, 184.863, 184.3606, 183.8854, 183.4351, 183.0078, 182.6016, 
    182.215, 181.8465, 181.4947, 181.1585, 180.8367, 180.5284, 180.2327, 
    179.9487, 179.6757, 179.413, 179.1599, 178.9158,
  340.0455, 339.7741, 339.4928, 339.2009, 338.8976, 338.5824, 338.2542, 
    337.9123, 337.5556, 337.183, 336.7935, 336.3857, 335.9581, 335.5093, 
    335.0374, 334.5406, 334.0168, 333.4636, 332.8783, 332.258, 331.5994, 
    330.8988, 330.1521, 329.3544, 328.5006, 327.5845, 326.5992, 325.537, 
    324.3888, 323.1444, 321.7921, 320.3184, 318.7078, 316.9427, 315.0031, 
    312.8659, 310.5056, 307.8939, 305, 301.7919, 298.238, 294.3098, 289.9866, 
    285.2609, 280.1453, 274.6786, 268.93, 262.998, 257.002, 251.07, 245.3214, 
    239.8548, 234.7391, 230.0134, 225.6902, 221.762, 218.2081, 215, 212.1061, 
    209.4944, 207.1341, 204.997, 203.0573, 201.2922, 199.6816, 198.2079, 
    196.8556, 195.6112, 194.463, 193.4008, 192.4155, 191.4994, 190.6456, 
    189.8479, 189.1012, 188.4006, 187.742, 187.1217, 186.5364, 185.9832, 
    185.4594, 184.9626, 184.4907, 184.0419, 183.6143, 183.2065, 182.817, 
    182.4444, 182.0877, 181.7458, 181.4176, 181.1024, 180.7991, 180.5072, 
    180.2259, 179.9545,
  339.0101, 338.7119, 338.4028, 338.0823, 337.7495, 337.4036, 337.0437, 
    336.669, 336.2782, 335.8704, 335.4442, 334.9984, 334.5312, 334.0413, 
    333.5267, 332.9854, 332.4151, 331.8136, 331.1779, 330.5051, 329.7918, 
    329.0341, 328.228, 327.3685, 326.4504, 325.4675, 324.4132, 323.2797, 
    322.0583, 320.7393, 319.3114, 317.7621, 316.0773, 314.2411, 312.2357, 
    310.0416, 307.6373, 305, 302.1061, 298.9323, 295.457, 291.6635, 287.5423, 
    283.096, 278.3424, 273.3188, 268.0826, 262.7099, 257.2901, 251.9174, 
    246.6812, 241.6576, 236.904, 232.4577, 228.3365, 224.543, 221.0677, 
    217.8939, 215, 212.3627, 209.9584, 207.7643, 205.7589, 203.9227, 
    202.2379, 200.6886, 199.2607, 197.9417, 196.7203, 195.5868, 194.5325, 
    193.5496, 192.6315, 191.772, 190.9658, 190.2082, 189.4949, 188.8221, 
    188.1864, 187.5849, 187.0146, 186.4733, 185.9587, 185.4688, 185.0016, 
    184.5558, 184.1296, 183.7218, 183.331, 182.9563, 182.5964, 182.2505, 
    181.9177, 181.5972, 181.2881, 180.9899,
  337.9783, 337.6538, 337.3176, 336.969, 336.6073, 336.2315, 335.8408, 
    335.4341, 335.0103, 334.5683, 334.1067, 333.6241, 333.119, 332.5895, 
    332.034, 331.4502, 330.8359, 330.1886, 329.5055, 328.7834, 328.0191, 
    327.2086, 326.3477, 325.4317, 324.4554, 323.4126, 322.297, 321.1011, 
    319.8166, 318.4343, 316.9438, 315.3338, 313.5914, 311.7027, 309.6523, 
    307.4239, 305, 302.3627, 299.4944, 296.3785, 293.0015, 289.3542, 
    285.4348, 281.2509, 276.8223, 272.1825, 267.379, 262.4716, 257.5284, 
    252.621, 247.8175, 243.1777, 238.7491, 234.5652, 230.6458, 226.9985, 
    223.6215, 220.5056, 217.6373, 215, 212.5761, 210.3477, 208.2973, 
    206.4086, 204.6662, 203.0562, 201.5657, 200.1834, 198.8989, 197.703, 
    196.5874, 195.5447, 194.5683, 193.6523, 192.7914, 191.9809, 191.2165, 
    190.4945, 189.8114, 189.1641, 188.5498, 187.966, 187.4105, 186.8811, 
    186.3759, 185.8933, 185.4317, 184.9897, 184.5659, 184.1592, 183.7685, 
    183.3927, 183.031, 182.6824, 182.3462, 182.0217,
  336.9506, 336.6002, 336.2374, 335.8615, 335.4715, 335.0667, 334.6459, 
    334.2082, 333.7524, 333.2774, 332.7816, 332.2638, 331.7222, 331.1551, 
    330.5605, 329.9365, 329.2805, 328.5902, 327.8626, 327.0947, 326.2831, 
    325.424, 324.5131, 323.546, 322.5173, 321.4215, 320.2522, 319.0024, 
    317.6644, 316.2296, 314.6888, 313.0313, 311.2463, 309.3214, 307.2438, 
    305, 302.5761, 299.9584, 297.1341, 294.0921, 290.8243, 287.3271, 283.603, 
    279.6623, 275.5245, 271.2192, 266.7855, 262.271, 257.729, 253.2145, 
    248.7808, 244.4755, 240.3377, 236.397, 232.6729, 229.1757, 225.9079, 
    222.8659, 220.0416, 217.4239, 215, 212.7562, 210.6786, 208.7537, 
    206.9686, 205.3113, 203.7704, 202.3356, 200.9976, 199.7478, 198.5785, 
    197.4827, 196.454, 195.4869, 194.576, 193.7169, 192.9053, 192.1374, 
    191.4098, 190.7195, 190.0636, 189.4395, 188.8449, 188.2778, 187.7362, 
    187.2183, 186.7226, 186.2475, 185.7918, 185.3541, 184.9334, 184.5285, 
    184.1385, 183.7626, 183.3998, 183.0495,
  335.927, 335.5515, 335.1627, 334.7601, 334.3427, 333.9095, 333.4597, 
    332.992, 332.5054, 331.9985, 331.47, 330.9183, 330.3419, 329.7389, 
    329.1074, 328.4453, 327.7502, 327.0195, 326.2506, 325.4402, 324.5852, 
    323.6816, 322.7256, 321.7125, 320.6375, 319.4951, 318.2795, 316.984, 
    315.6016, 314.1244, 312.544, 310.8514, 309.0368, 307.0899, 305, 302.7562, 
    300.3477, 297.7643, 294.9969, 292.0387, 288.8855, 285.5371, 281.9988, 
    278.2817, 274.4044, 270.3923, 266.278, 262.0999, 257.9001, 253.722, 
    249.6077, 245.5956, 241.7182, 238.0012, 234.4629, 231.1145, 227.9613, 
    225.003, 222.2357, 219.6523, 217.2438, 215, 212.9101, 210.9632, 209.1486, 
    207.4559, 205.8756, 204.3985, 203.016, 201.7205, 200.5049, 199.3625, 
    198.2875, 197.2744, 196.3184, 195.4148, 194.5597, 193.7494, 192.9805, 
    192.2498, 191.5547, 190.8926, 190.2611, 189.6581, 189.0817, 188.53, 
    188.0015, 187.4946, 187.008, 186.5403, 186.0905, 185.6573, 185.2399, 
    184.8373, 184.4486, 184.073,
  334.9081, 334.5078, 334.0938, 333.6652, 333.2211, 332.7606, 332.2826, 
    331.786, 331.2697, 330.7323, 330.1724, 329.5884, 328.9789, 328.3419, 
    327.6755, 326.9776, 326.2458, 325.4778, 324.6705, 323.8212, 322.9264, 
    321.9827, 320.9861, 319.9323, 318.8166, 317.634, 316.3789, 315.0454, 
    313.627, 312.1166, 310.5068, 308.7897, 306.957, 305, 302.9101, 300.6786, 
    298.2973, 295.7589, 293.0573, 290.1884, 287.1511, 283.9474, 280.5839, 
    277.0719, 273.4281, 269.6749, 265.8391, 261.9522, 258.0478, 254.1609, 
    250.3251, 246.5719, 242.9281, 239.4162, 236.0526, 232.8489, 229.8116, 
    226.9427, 224.2411, 221.7027, 219.3214, 217.0899, 215, 213.043, 211.2103, 
    209.4932, 207.8834, 206.373, 204.9546, 203.6211, 202.366, 201.1834, 
    200.0677, 199.0139, 198.0173, 197.0736, 196.1788, 195.3295, 194.5223, 
    193.7542, 193.0224, 192.3245, 191.6581, 191.0211, 190.4115, 189.8277, 
    189.2677, 188.7303, 188.214, 187.7174, 187.2394, 186.7789, 186.3348, 
    185.9062, 185.4922, 185.0919,
  333.8939, 333.4697, 333.0311, 332.5773, 332.1074, 331.6204, 331.1152, 
    330.5908, 330.046, 329.4793, 328.8895, 328.2749, 327.634, 326.9649, 
    326.2657, 325.5343, 324.7685, 323.9657, 323.1233, 322.2383, 321.3077, 
    320.3279, 319.2952, 318.2057, 317.0548, 315.838, 314.5501, 313.1857, 
    311.7389, 310.2036, 308.5732, 306.841, 305, 303.043, 300.9632, 298.7537, 
    296.4086, 293.9227, 291.2922, 288.5153, 285.5927, 282.5277, 279.3277, 
    276.0034, 272.57, 269.0465, 265.4557, 261.8233, 258.1767, 254.5443, 
    250.9535, 247.43, 243.9966, 240.6723, 237.4723, 234.4073, 231.4847, 
    228.7078, 226.0773, 223.5914, 221.2463, 219.0368, 216.957, 215, 213.159, 
    211.4268, 209.7964, 208.2611, 206.8143, 205.4499, 204.162, 202.9452, 
    201.7944, 200.7048, 199.6721, 198.6923, 197.7617, 196.8767, 196.0343, 
    195.2315, 194.4657, 193.7343, 193.0351, 192.366, 191.7251, 191.1105, 
    190.5207, 189.954, 189.4092, 188.8848, 188.3796, 187.8926, 187.4227, 
    186.9689, 186.5303, 186.1061,
  332.8849, 332.4373, 331.9749, 331.4966, 331.0018, 330.4892, 329.958, 
    329.4069, 328.8347, 328.2402, 327.6219, 326.9783, 326.3078, 325.6086, 
    324.8787, 324.1162, 323.3188, 322.4842, 321.6096, 320.6924, 319.7295, 
    318.7176, 317.6533, 316.5327, 315.3519, 314.1065, 312.7918, 311.4031, 
    309.935, 308.3822, 306.7392, 305, 303.159, 301.2103, 299.1486, 296.9687, 
    294.6662, 292.2379, 289.6816, 286.9972, 284.1863, 281.2534, 278.2056, 
    275.0533, 271.8097, 268.4915, 265.1178, 261.7098, 258.2902, 254.8822, 
    251.5085, 248.1903, 244.9467, 241.7944, 238.7466, 235.8137, 233.0029, 
    230.3184, 227.7621, 225.3338, 223.0314, 220.8514, 218.7897, 216.841, 215, 
    213.2608, 211.6178, 210.065, 208.5969, 207.2082, 205.8935, 204.6481, 
    203.4673, 202.3467, 201.2824, 200.2705, 199.3076, 198.3904, 197.5159, 
    196.6812, 195.8838, 195.1213, 194.3915, 193.6922, 193.0217, 192.3781, 
    191.7598, 191.1653, 190.5931, 190.042, 189.5108, 188.9982, 188.5033, 
    188.0251, 187.5627, 187.1152,
  331.8811, 331.4109, 330.9254, 330.4236, 329.9047, 329.3676, 328.8113, 
    328.2346, 327.6365, 327.0155, 326.3702, 325.6992, 325.0009, 324.2734, 
    323.5151, 322.7238, 321.8974, 321.0336, 320.1299, 319.1837, 318.1921, 
    317.1521, 316.0603, 314.9133, 313.7074, 312.4386, 311.1028, 309.6957, 
    308.2126, 306.649, 305, 303.2608, 301.4268, 299.4932, 297.456, 295.3112, 
    293.0562, 290.6886, 288.2079, 285.6147, 282.9118, 280.1038, 277.1977, 
    274.203, 271.1316, 267.9977, 264.8176, 261.6091, 258.3909, 255.1824, 
    252.0023, 248.8684, 245.797, 242.8023, 239.8962, 237.0882, 234.3852, 
    231.7921, 229.3114, 226.9438, 224.6887, 222.5441, 220.5068, 218.5732, 
    216.7392, 215, 213.351, 211.7874, 210.3043, 208.8972, 207.5614, 206.2926, 
    205.0867, 203.9397, 202.8479, 201.8079, 200.8163, 199.8701, 198.9664, 
    198.1026, 197.2762, 196.4849, 195.7266, 194.9991, 194.3008, 193.6298, 
    192.9845, 192.3635, 191.7654, 191.1887, 190.6324, 190.0953, 189.5764, 
    189.0746, 188.589, 188.1189,
  330.883, 330.3909, 329.883, 329.3585, 328.8164, 328.2558, 327.6755, 
    327.0746, 326.4516, 325.8055, 325.1348, 324.4381, 323.7137, 322.9601, 
    322.1753, 321.3575, 320.5046, 319.6144, 318.6845, 317.7125, 316.6957, 
    315.6311, 314.5159, 313.3467, 312.1203, 310.833, 309.4812, 308.0611, 
    306.5687, 305, 303.351, 301.6178, 299.7964, 297.8834, 295.8756, 293.7704, 
    291.5657, 289.2607, 286.8556, 284.3517, 281.7523, 279.062, 276.2876, 
    273.4378, 270.5229, 267.5555, 264.5491, 261.519, 258.481, 255.4509, 
    252.4445, 249.4771, 246.5622, 243.7124, 240.938, 238.2477, 235.6483, 
    233.1444, 230.7393, 228.4343, 226.2296, 224.1244, 222.1166, 220.2036, 
    218.3822, 216.649, 215, 213.4313, 211.9389, 210.5188, 209.167, 207.8797, 
    206.6533, 205.4841, 204.3689, 203.3043, 202.2875, 201.3154, 200.3856, 
    199.4954, 198.6425, 197.8247, 197.0399, 196.2863, 195.5619, 194.8652, 
    194.1945, 193.5484, 192.9255, 192.3245, 191.7442, 191.1836, 190.6415, 
    190.117, 189.6091, 189.117,
  329.8907, 329.3774, 328.848, 328.3016, 327.7373, 327.1542, 326.5511, 
    325.9269, 325.2806, 324.6108, 323.9162, 323.1954, 322.4468, 321.6689, 
    320.8598, 320.0177, 319.1408, 318.2268, 317.2736, 316.2789, 315.2401, 
    314.1545, 313.0195, 311.8322, 310.5894, 309.2881, 307.925, 306.4968, 305, 
    303.4313, 301.7874, 300.065, 298.2611, 296.373, 294.3984, 292.3356, 
    290.1834, 287.9417, 285.6112, 283.194, 280.6932, 278.1138, 275.4619, 
    272.7454, 269.9735, 267.157, 264.3076, 261.4381, 258.5619, 255.6924, 
    252.843, 250.0265, 247.2546, 244.5381, 241.8862, 239.3067, 236.806, 
    234.3888, 232.0583, 229.8166, 227.6644, 225.6015, 223.627, 221.7389, 
    219.935, 218.2126, 216.5687, 215, 213.5032, 212.075, 210.7119, 209.4106, 
    208.1678, 206.9805, 205.8455, 204.76, 203.7211, 202.7264, 201.7732, 
    200.8592, 199.9823, 199.1402, 198.3312, 197.5532, 196.8046, 196.0838, 
    195.3892, 194.7194, 194.0731, 193.4489, 192.8458, 192.2627, 191.6984, 
    191.152, 190.6226, 190.1093,
  328.9044, 328.3707, 327.8206, 327.2533, 326.6677, 326.063, 325.4382, 
    324.7922, 324.1237, 323.4317, 322.7147, 321.9714, 321.2004, 320.4001, 
    319.5688, 318.7047, 317.8061, 316.8709, 315.8971, 314.8826, 313.8249, 
    312.7217, 311.5706, 310.3687, 309.1136, 307.8023, 306.4321, 305, 
    303.5032, 301.9389, 300.3043, 298.5969, 296.8143, 294.9546, 293.016, 
    290.9976, 288.8989, 286.7203, 284.463, 282.1293, 279.7226, 277.2474, 
    274.7095, 272.116, 269.475, 266.796, 264.089, 261.3649, 258.6351, 
    255.9111, 253.204, 250.525, 247.884, 245.2905, 242.7526, 240.2774, 
    237.8707, 235.537, 233.2797, 231.1011, 229.0024, 226.984, 225.0454, 
    223.1857, 221.4031, 219.6957, 218.0611, 216.4968, 215, 213.5679, 
    212.1977, 210.8864, 209.6313, 208.4295, 207.2783, 206.1751, 205.1174, 
    204.1029, 203.1291, 202.1939, 201.2953, 200.4313, 199.5999, 198.7996, 
    198.0286, 197.2853, 196.5683, 195.8763, 195.2078, 194.5618, 193.937, 
    193.3323, 192.7467, 192.1794, 191.6293, 191.0956,
  327.9243, 327.371, 326.8011, 326.2136, 325.6078, 324.9827, 324.3373, 
    323.6705, 322.9813, 322.2684, 321.5306, 320.7665, 319.9748, 319.154, 
    318.3024, 317.4185, 316.5006, 315.5467, 314.5549, 313.5233, 312.4498, 
    311.3321, 310.168, 308.9551, 307.6912, 306.3736, 305, 303.5679, 302.075, 
    300.5188, 298.8972, 297.2082, 295.4499, 293.6211, 291.7205, 289.7478, 
    287.703, 285.5868, 283.4008, 281.1473, 278.8298, 276.4526, 274.0209, 
    271.5412, 269.0206, 266.4673, 263.8901, 261.2983, 258.7017, 256.1099, 
    253.5327, 250.9794, 248.4588, 245.9791, 243.5474, 241.1702, 238.8526, 
    236.5992, 234.4132, 232.297, 230.2522, 228.2795, 226.3789, 224.5501, 
    222.7918, 221.1028, 219.4812, 217.925, 216.4321, 215, 213.6264, 212.3089, 
    211.0449, 209.832, 208.6679, 207.5502, 206.4767, 205.4451, 204.4533, 
    203.4994, 202.5815, 201.6976, 200.846, 200.0252, 199.2335, 198.4694, 
    197.7316, 197.0187, 196.3295, 195.6627, 195.0173, 194.3922, 193.7864, 
    193.1989, 192.629, 192.0756,
  326.9507, 326.3785, 325.7896, 325.183, 324.5579, 323.9134, 323.2485, 
    322.5623, 321.8535, 321.1212, 320.364, 319.5808, 318.7701, 317.9307, 
    317.0609, 316.1593, 315.2242, 314.2539, 313.2467, 312.2008, 311.1141, 
    309.9848, 308.8109, 307.5901, 306.3205, 305, 303.6264, 302.1977, 
    300.7119, 299.167, 297.5614, 295.8935, 294.162, 292.366, 290.5049, 
    288.5785, 286.5874, 284.5325, 282.4155, 280.239, 278.0062, 275.721, 
    273.3885, 271.0142, 268.6046, 266.1668, 263.7085, 261.2375, 258.7625, 
    256.2915, 253.8332, 251.3954, 248.9858, 246.6115, 244.279, 241.9939, 
    239.761, 237.5845, 235.4675, 233.4126, 231.4215, 229.4951, 227.634, 
    225.838, 224.1065, 222.4386, 220.833, 219.2881, 217.8023, 216.3736, 215, 
    213.6795, 212.4099, 211.1892, 210.0152, 208.8859, 207.7992, 206.7533, 
    205.7461, 204.7758, 203.8407, 202.9391, 202.0693, 201.2298, 200.4192, 
    199.6359, 198.8788, 198.1464, 197.4377, 196.7515, 196.0866, 195.4421, 
    194.817, 194.2104, 193.6215, 193.0493,
  325.9837, 325.3935, 324.7863, 324.1615, 323.5181, 322.8553, 322.1721, 
    321.4677, 320.7407, 319.9904, 319.2153, 318.4145, 317.5866, 316.7303, 
    315.8442, 314.9268, 313.9768, 312.9925, 311.9722, 310.9144, 309.8172, 
    308.679, 307.498, 306.2722, 305, 303.6795, 302.3088, 300.8864, 299.4106, 
    297.8797, 296.2926, 294.6481, 292.9452, 291.1834, 289.3625, 287.4827, 
    285.5446, 283.5496, 281.4994, 279.3965, 277.2439, 275.0454, 272.8055, 
    270.5292, 268.2223, 265.8909, 263.5418, 261.1818, 258.8182, 256.4582, 
    254.1091, 251.7777, 249.4708, 247.1945, 244.9546, 242.7561, 240.6035, 
    238.5006, 236.4504, 234.4553, 232.5173, 230.6375, 228.8166, 227.0548, 
    225.3519, 223.7074, 222.1203, 220.5894, 219.1136, 217.6911, 216.3205, 
    215, 213.7278, 212.502, 211.321, 210.1828, 209.0856, 208.0278, 207.0076, 
    206.0232, 205.0732, 204.1558, 203.2697, 202.4134, 201.5855, 200.7847, 
    200.0097, 199.2593, 198.5324, 197.8278, 197.1447, 196.4819, 195.8385, 
    195.2137, 194.6065, 194.0163,
  325.0234, 324.416, 323.7915, 323.1494, 322.4887, 321.8087, 321.1083, 
    320.3868, 319.643, 318.8759, 318.0846, 317.2677, 316.4242, 315.5528, 
    314.6522, 313.7211, 312.7581, 311.7619, 310.7308, 309.6635, 308.5583, 
    307.4137, 306.2281, 305, 303.7278, 302.4099, 301.0449, 299.6313, 
    298.1678, 296.6533, 295.0867, 293.4673, 291.7943, 290.0677, 288.2875, 
    286.454, 284.5683, 282.6315, 280.6456, 278.6129, 276.5363, 274.4195, 
    272.2663, 270.0813, 267.8696, 265.6366, 263.3882, 261.1305, 258.8695, 
    256.6118, 254.3634, 252.1304, 249.9187, 247.7337, 245.5805, 243.4637, 
    241.3871, 239.3544, 237.3685, 235.4317, 233.546, 231.7125, 229.9323, 
    228.2056, 226.5327, 224.9133, 223.3467, 221.8322, 220.3687, 218.9551, 
    217.5901, 216.2722, 215, 213.7719, 212.5863, 211.4417, 210.3366, 
    209.2692, 208.2381, 207.2418, 206.2789, 205.3478, 204.4472, 203.5758, 
    202.7323, 201.9154, 201.1241, 200.357, 199.6132, 198.8916, 198.1913, 
    197.5113, 196.8506, 196.2085, 195.584, 194.9766,
  324.0701, 323.4462, 322.8054, 322.1469, 321.4699, 320.7737, 320.0573, 
    319.3199, 318.5605, 317.7781, 316.9718, 316.1404, 315.2829, 314.3981, 
    313.4849, 312.5419, 311.568, 310.5618, 309.522, 308.4474, 307.3364, 
    306.1877, 305, 303.7719, 302.502, 301.1891, 299.832, 298.4294, 296.9805, 
    295.4841, 293.9397, 292.3467, 290.7048, 289.0139, 287.2744, 285.4869, 
    283.6523, 281.772, 279.8479, 277.8823, 275.8779, 273.838, 271.766, 
    269.6663, 267.5432, 265.4015, 263.2463, 261.083, 258.917, 256.7537, 
    254.5985, 252.4568, 250.3337, 248.234, 246.1621, 244.1221, 242.1177, 
    240.1521, 238.228, 236.3477, 234.5131, 232.7256, 230.9861, 229.2952, 
    227.6533, 226.0603, 224.5159, 223.0195, 221.5705, 220.168, 218.8108, 
    217.498, 216.2281, 215, 213.8123, 212.6637, 211.5527, 210.478, 209.4382, 
    208.432, 207.4581, 206.5151, 205.6019, 204.7171, 203.8596, 203.0282, 
    202.2219, 201.4395, 200.6802, 199.9427, 199.2264, 198.5301, 197.8531, 
    197.1947, 196.5538, 195.9299,
  323.1238, 322.4843, 321.8279, 321.154, 320.4617, 319.7503, 319.019, 
    318.267, 317.4932, 316.6969, 315.877, 315.0327, 314.1627, 313.2662, 
    312.3419, 311.3889, 310.4059, 309.3917, 308.3452, 307.2653, 306.1506, 
    305, 303.8123, 302.5863, 301.321, 300.0152, 298.6679, 297.2783, 295.8455, 
    294.3689, 292.8479, 291.2824, 289.6721, 288.0173, 286.3184, 284.576, 
    282.7914, 280.9659, 279.1012, 277.1996, 275.2636, 273.2962, 271.3006, 
    269.2806, 267.2401, 265.1833, 263.1147, 261.039, 258.961, 256.8853, 
    254.8167, 252.7599, 250.7194, 248.6994, 246.7038, 244.7364, 242.8004, 
    240.8988, 239.0342, 237.2086, 235.424, 233.6816, 231.9827, 230.3279, 
    228.7176, 227.1521, 225.6311, 224.1545, 222.7217, 221.3321, 219.9848, 
    218.679, 217.4137, 216.1877, 215, 213.8494, 212.7347, 211.6547, 210.6083, 
    209.5941, 208.6111, 207.6581, 206.7338, 205.8373, 204.9673, 204.1229, 
    203.3031, 202.5068, 201.733, 200.981, 200.2497, 199.5383, 198.846, 
    198.1721, 197.5157, 196.8762,
  322.1847, 321.5304, 320.8593, 320.1709, 319.4643, 318.7389, 317.9938, 
    317.2282, 316.4414, 315.6324, 314.8004, 313.9444, 313.0635, 312.1568, 
    311.2232, 310.2618, 309.2714, 308.2511, 307.1998, 306.1165, 305, 
    303.8494, 302.6636, 301.4417, 300.1828, 298.8859, 297.5502, 296.1751, 
    294.7599, 293.3043, 291.8079, 290.2705, 288.6923, 287.0736, 285.4148, 
    283.7169, 281.9809, 280.2082, 278.4006, 276.5601, 274.689, 272.7902, 
    270.8664, 268.9211, 266.9578, 264.9802, 262.9923, 260.9981, 259.0019, 
    257.0077, 255.0198, 253.0422, 251.0789, 249.1336, 247.2099, 245.311, 
    243.4399, 241.5994, 239.7918, 238.0191, 236.2831, 234.5852, 232.9264, 
    231.3077, 229.7295, 228.1921, 226.6957, 225.24, 223.8249, 222.4498, 
    221.1141, 219.8172, 218.5583, 217.3363, 216.1506, 215, 213.8835, 
    212.8002, 211.7489, 210.7286, 209.7382, 208.7768, 207.8432, 206.9365, 
    206.0556, 205.1996, 204.3676, 203.5586, 202.7718, 202.0062, 201.2611, 
    200.5357, 199.8291, 199.1406, 198.4696, 197.8153,
  321.2528, 320.5846, 319.8998, 319.1978, 318.4778, 317.7393, 316.9815, 
    316.2036, 315.4049, 314.5845, 313.7417, 312.8755, 311.9852, 311.0698, 
    310.1284, 309.1602, 308.1641, 307.1394, 306.085, 305, 303.8835, 302.7347, 
    301.5526, 300.3365, 299.0856, 297.7992, 296.4767, 295.1174, 293.7211, 
    292.2875, 290.8163, 289.3076, 287.7617, 286.1788, 284.5598, 282.9053, 
    281.2166, 279.4949, 277.742, 275.9598, 274.1504, 272.3164, 270.4603, 
    268.5852, 266.6942, 264.7907, 262.8781, 260.96, 259.04, 257.1219, 
    255.2093, 253.3058, 251.4148, 249.5397, 247.6836, 245.8496, 244.0402, 
    242.258, 240.5051, 238.7835, 237.0947, 235.4403, 233.8212, 232.2383, 
    230.6924, 229.1837, 227.7125, 226.2789, 224.8826, 223.5233, 222.2008, 
    220.9144, 219.6634, 218.4473, 217.2653, 216.1165, 215, 213.915, 212.8606, 
    211.8359, 210.8398, 209.8716, 208.9302, 208.0148, 207.1245, 206.2583, 
    205.4155, 204.5951, 203.7964, 203.0185, 202.2607, 201.5221, 200.8022, 
    200.1002, 199.4154, 198.7471,
  320.3284, 319.647, 318.9493, 318.2346, 317.5023, 316.7518, 315.9824, 
    315.1933, 314.3838, 313.5533, 312.7009, 311.8259, 310.9274, 310.0048, 
    309.0571, 308.0836, 307.0835, 306.0559, 305, 303.915, 302.8002, 301.6548, 
    300.478, 299.2692, 298.0278, 296.7533, 295.4451, 294.1029, 292.7264, 
    291.3155, 289.8701, 288.3904, 286.8767, 285.3295, 283.7494, 282.1374, 
    280.4945, 278.8221, 277.1217, 275.3952, 273.6444, 271.8718, 270.0796, 
    268.2706, 266.4475, 264.6134, 262.7713, 260.9243, 259.0757, 257.2287, 
    255.3866, 253.5525, 251.7294, 249.9204, 248.1282, 246.3556, 244.6048, 
    242.8783, 241.1779, 239.5055, 237.8626, 236.2506, 234.6705, 233.1233, 
    231.6096, 230.1299, 228.6846, 227.2736, 225.8971, 224.5549, 223.2467, 
    221.9722, 220.7308, 219.522, 218.3453, 217.1998, 216.085, 215, 213.9441, 
    212.9165, 211.9164, 210.9429, 209.9952, 209.0726, 208.1741, 207.2991, 
    206.4467, 205.6162, 204.8067, 204.0176, 203.2482, 202.4977, 201.7654, 
    201.0507, 200.353, 199.6716,
  319.4114, 318.7177, 318.008, 317.2816, 316.5379, 315.7763, 314.9963, 
    314.1971, 313.3781, 312.5386, 311.6779, 310.7953, 309.8901, 308.9616, 
    308.0091, 307.0318, 306.029, 305, 303.9441, 302.8606, 301.7489, 300.6083, 
    299.4382, 298.2381, 297.0075, 295.7461, 294.4533, 293.1291, 291.7732, 
    290.3856, 288.9664, 287.5158, 286.0343, 284.5222, 282.9805, 281.4098, 
    279.8114, 278.1864, 276.5364, 274.863, 273.1681, 271.4536, 269.7219, 
    267.9752, 266.216, 264.4471, 262.6711, 260.8908, 259.1092, 257.3289, 
    255.5529, 253.784, 252.0248, 250.2781, 248.5464, 246.8319, 245.137, 
    243.4636, 241.8136, 240.1886, 238.5902, 237.0195, 235.4777, 233.9657, 
    232.4841, 231.0336, 229.6144, 228.2268, 226.8709, 225.5467, 224.2539, 
    222.9924, 221.7619, 220.5618, 219.3917, 218.2511, 217.1394, 216.0559, 
    215, 213.971, 212.9682, 211.9909, 211.0384, 210.1099, 209.2047, 208.3221, 
    207.4614, 206.6219, 205.8029, 205.0037, 204.2236, 203.4621, 202.7184, 
    201.992, 201.2823, 200.5886,
  318.502, 317.7968, 317.0759, 316.3386, 315.5845, 314.8129, 314.0233, 
    313.2151, 312.3876, 311.5403, 310.6725, 309.7836, 308.873, 307.9399, 
    306.9838, 306.0041, 305, 303.971, 302.9165, 301.8359, 300.7286, 299.5941, 
    298.432, 297.2419, 296.0232, 294.7758, 293.4994, 292.1939, 290.8592, 
    289.4954, 288.1026, 286.6812, 285.2315, 283.7542, 282.2498, 280.7195, 
    279.1641, 277.5849, 275.9832, 274.3606, 272.7188, 271.0596, 269.385, 
    267.6972, 265.9983, 264.2908, 262.577, 260.8594, 259.1406, 257.423, 
    255.7092, 254.0017, 252.3028, 250.615, 248.9404, 247.2812, 245.6394, 
    244.0168, 242.4151, 240.8359, 239.2805, 237.7502, 236.2458, 234.7685, 
    233.3188, 231.8974, 230.5046, 229.1408, 227.8061, 226.5006, 225.2242, 
    223.9768, 222.7582, 221.568, 220.4059, 219.2714, 218.1641, 217.0835, 
    216.029, 215, 213.9959, 213.0162, 212.0601, 211.127, 210.2164, 209.3275, 
    208.4597, 207.6124, 206.7849, 205.9767, 205.1871, 204.4155, 203.6614, 
    202.9241, 202.2032, 201.498,
  317.6002, 316.8844, 316.1531, 315.4059, 314.6422, 313.8616, 313.0634, 
    312.2472, 311.4124, 310.5584, 309.6847, 308.7906, 307.8757, 306.9393, 
    305.981, 305, 303.9959, 302.9682, 301.9164, 300.8398, 299.7382, 298.6111, 
    297.4581, 296.2789, 295.0732, 293.8407, 292.5815, 291.2953, 289.9823, 
    288.6425, 287.2762, 285.8838, 284.4657, 283.0224, 281.5547, 280.0635, 
    278.5498, 277.0146, 275.4594, 273.8853, 272.2942, 270.6875, 269.0672, 
    267.435, 265.7931, 264.1435, 262.4883, 260.8298, 259.1702, 257.5117, 
    255.8565, 254.2069, 252.565, 250.9328, 249.3125, 247.7058, 246.1146, 
    244.5406, 242.9854, 241.4502, 239.9364, 238.4453, 236.9776, 235.5343, 
    234.1162, 232.7238, 231.3575, 230.0177, 228.7047, 227.4185, 226.1593, 
    224.9268, 223.7211, 222.5419, 221.3889, 220.2618, 219.1602, 218.0836, 
    217.0318, 216.0041, 215, 214.019, 213.0607, 212.1243, 211.2094, 210.3153, 
    209.4416, 208.5876, 207.7528, 206.9366, 206.1384, 205.3578, 204.5941, 
    203.8469, 203.1156, 202.3998,
  316.7061, 315.9804, 315.2396, 314.4833, 313.711, 312.9223, 312.1166, 
    311.2934, 310.4523, 309.5927, 308.7141, 307.8161, 306.898, 305.9595, 305, 
    304.019, 303.0162, 301.9909, 300.9429, 299.8716, 298.7768, 297.6581, 
    296.5151, 295.3478, 294.1558, 292.9391, 291.6976, 290.4312, 289.1402, 
    287.8247, 286.4849, 285.1213, 283.7343, 282.3245, 280.8926, 279.4395, 
    277.966, 276.4733, 274.9626, 273.4351, 271.8922, 270.3356, 268.7667, 
    267.1873, 265.5993, 264.0044, 262.4046, 260.8019, 259.1981, 257.5954, 
    255.9956, 254.4007, 252.8126, 251.2333, 249.6644, 248.1078, 246.5649, 
    245.0374, 243.5267, 242.034, 240.5605, 239.1074, 237.6755, 236.2657, 
    234.8787, 233.5151, 232.1753, 230.8598, 229.5687, 228.3024, 227.0609, 
    225.8442, 224.6522, 223.4849, 222.3419, 221.2232, 220.1284, 219.0571, 
    218.0091, 216.9838, 215.981, 215, 214.0405, 213.102, 212.1839, 211.2859, 
    210.4073, 209.5477, 208.7066, 207.8834, 207.0777, 206.289, 205.5167, 
    204.7604, 204.0196, 203.2939,
  315.8197, 315.0849, 314.3354, 313.5709, 312.7909, 311.995, 311.1827, 
    310.3535, 309.5071, 308.6429, 307.7606, 306.8596, 305.9396, 305, 
    304.0405, 303.0607, 302.0601, 301.0384, 299.9952, 298.9302, 297.8432, 
    296.7338, 295.6019, 294.4472, 293.2697, 292.0693, 290.846, 289.5999, 
    288.3311, 287.0399, 285.7266, 284.3914, 283.0351, 281.6581, 280.2611, 
    278.8449, 277.4105, 275.9587, 274.4907, 273.0078, 271.5111, 270.0021, 
    268.4822, 266.9529, 265.416, 263.8729, 262.3255, 260.7755, 259.2245, 
    257.6745, 256.1271, 254.584, 253.0471, 251.5178, 249.9979, 248.4889, 
    246.9922, 245.5093, 244.0413, 242.5895, 241.1551, 239.7389, 238.3419, 
    236.9649, 235.6085, 234.2734, 232.9601, 231.6688, 230.4001, 229.154, 
    227.9307, 226.7303, 225.5528, 224.3981, 223.2662, 222.1568, 221.0698, 
    220.0048, 218.9616, 217.9399, 216.9393, 215.9595, 215, 214.0604, 
    213.1404, 212.2394, 211.3571, 210.4929, 209.6465, 208.8173, 208.005, 
    207.2091, 206.4291, 205.6646, 204.9151, 204.1803,
  314.941, 314.1979, 313.4406, 312.6687, 311.8819, 311.0797, 310.2617, 
    309.4275, 308.5768, 307.709, 306.8239, 305.921, 305, 304.0604, 303.102, 
    302.1243, 301.127, 300.1099, 299.0726, 298.0148, 296.9365, 295.8373, 
    294.7171, 293.5758, 292.4134, 291.2299, 290.0252, 288.7996, 287.5532, 
    286.2863, 284.9991, 283.6922, 282.366, 281.0211, 279.6581, 278.2778, 
    276.881, 275.4688, 274.0419, 272.6016, 271.1491, 269.6855, 268.2122, 
    266.7307, 265.2422, 263.7483, 262.2505, 260.7505, 259.2495, 257.7495, 
    256.2517, 254.7578, 253.2693, 251.7878, 250.3145, 248.8509, 247.3984, 
    245.9581, 244.5312, 243.1189, 241.7222, 240.3419, 238.9789, 237.634, 
    236.3078, 235.0009, 233.7137, 232.4468, 231.2004, 229.9748, 228.7702, 
    227.5866, 226.4242, 225.2829, 224.1627, 223.0635, 221.9852, 220.9274, 
    219.8901, 218.873, 217.8757, 216.898, 215.9396, 215, 214.079, 213.1761, 
    212.291, 211.4232, 210.5725, 209.7383, 208.9203, 208.1181, 207.3313, 
    206.5594, 205.8021, 205.059,
  314.0701, 313.3195, 312.5551, 311.7767, 310.9839, 310.1762, 309.3535, 
    308.5152, 307.661, 306.7907, 305.9038, 305, 304.079, 303.1404, 302.1839, 
    301.2094, 300.2164, 299.2047, 298.1741, 297.1245, 296.0556, 294.9673, 
    293.8596, 292.7323, 291.5855, 290.4192, 289.2335, 288.0286, 286.8046, 
    285.5619, 284.3008, 283.0217, 281.7251, 280.4116, 279.0817, 277.7362, 
    276.3759, 275.0016, 273.6143, 272.215, 270.8047, 269.3846, 267.9557, 
    266.5195, 265.0772, 263.63, 262.1794, 260.7267, 259.2733, 257.8206, 
    256.37, 254.9228, 253.4805, 252.0443, 250.6154, 249.1953, 247.785, 
    246.3857, 244.9984, 243.6241, 242.2638, 240.9183, 239.5885, 238.2749, 
    236.9783, 235.6992, 234.4381, 233.1954, 231.9714, 230.7665, 229.5808, 
    228.4145, 227.2677, 226.1404, 225.0327, 223.9444, 222.8755, 221.8259, 
    220.7953, 219.7836, 218.7906, 217.8161, 216.8596, 215.921, 215, 214.0962, 
    213.2093, 212.3389, 211.4848, 210.6465, 209.8238, 209.0162, 208.2233, 
    207.4449, 206.6805, 205.9299,
  313.207, 312.4496, 311.679, 310.8948, 310.0968, 309.2846, 308.4579, 
    307.6164, 306.7598, 305.8878, 305, 304.0962, 303.1761, 302.2394, 
    301.2859, 300.3153, 299.3275, 298.3221, 297.2991, 296.2583, 295.1996, 
    294.123, 293.0282, 291.9154, 290.7847, 289.636, 288.4694, 287.2853, 
    286.0838, 284.8652, 283.6298, 282.3781, 281.1105, 279.8276, 278.53, 
    277.2184, 275.8933, 274.5558, 273.2065, 271.8465, 270.4766, 269.098, 
    267.7116, 266.3187, 264.9203, 263.5175, 262.1118, 260.7041, 259.2959, 
    257.8882, 256.4825, 255.0797, 253.6813, 252.2883, 250.902, 249.5234, 
    248.1535, 246.7935, 245.4442, 244.1067, 242.7817, 241.47, 240.1723, 
    238.8895, 237.6219, 236.3702, 235.1348, 233.9162, 232.7147, 231.5306, 
    230.3641, 229.2153, 228.0846, 226.9718, 225.8771, 224.8004, 223.7417, 
    222.7009, 221.6779, 220.6725, 219.6847, 218.7141, 217.7606, 216.8239, 
    215.9038, 215, 214.1122, 213.2402, 212.3836, 211.5421, 210.7154, 
    209.9032, 209.1052, 208.3211, 207.5504, 206.793,
  312.3516, 311.5882, 310.8121, 310.023, 309.2206, 308.4047, 307.575, 
    306.7311, 305.8729, 305, 304.1122, 303.2093, 302.291, 301.3571, 300.4073, 
    299.4416, 298.4597, 297.4614, 296.4467, 295.4155, 294.3676, 293.3031, 
    292.2219, 291.1241, 290.0096, 288.8788, 287.7316, 286.5683, 285.3892, 
    284.1945, 282.9845, 281.7598, 280.5207, 279.2677, 278.0015, 276.7226, 
    275.4317, 274.1296, 272.817, 271.4947, 270.1637, 268.8248, 267.479, 
    266.1273, 264.7708, 263.4105, 262.0474, 260.6826, 259.3174, 257.9526, 
    256.5895, 255.2292, 253.8727, 252.521, 251.1752, 249.8363, 248.5053, 
    247.183, 245.8704, 244.5683, 243.2774, 241.9985, 240.7323, 239.4793, 
    238.2402, 237.0155, 235.8055, 234.6108, 233.4317, 232.2684, 231.1212, 
    229.9903, 228.8759, 227.7781, 226.6969, 225.6324, 224.5845, 223.5533, 
    222.5386, 221.5403, 220.5584, 219.5927, 218.6429, 217.709, 216.7907, 
    215.8878, 215, 214.1271, 213.2689, 212.425, 211.5953, 210.7794, 209.977, 
    209.1879, 208.4118, 207.6484,
  311.5041, 310.7353, 309.9545, 309.1612, 308.3553, 307.5364, 306.7044, 
    305.859, 305, 304.1271, 303.2402, 302.339, 301.4232, 300.4929, 299.5477, 
    298.5876, 297.6124, 296.6219, 295.6162, 294.5951, 293.5586, 292.5068, 
    291.4395, 290.357, 289.2593, 288.1465, 287.0187, 285.8763, 284.7194, 
    283.5484, 282.3635, 281.1653, 279.954, 278.7303, 277.4946, 276.2476, 
    274.9897, 273.7218, 272.4444, 271.1585, 269.8647, 268.5639, 267.257, 
    265.9448, 264.6282, 263.3083, 261.986, 260.6621, 259.3379, 258.014, 
    256.6917, 255.3718, 254.0552, 252.743, 251.4361, 250.1353, 248.8415, 
    247.5556, 246.2782, 245.0103, 243.7525, 242.5054, 241.2697, 240.046, 
    238.8347, 237.6365, 236.4516, 235.2806, 234.1237, 232.9813, 231.8536, 
    230.7407, 229.643, 228.5605, 227.4932, 226.4414, 225.4049, 224.3838, 
    223.3781, 222.3876, 221.4124, 220.4523, 219.5071, 218.5768, 217.6611, 
    216.7598, 215.8729, 215, 214.141, 213.2956, 212.4636, 211.6447, 210.8388, 
    210.0455, 209.2647, 208.4959,
  310.6642, 309.891, 309.1061, 308.3094, 307.5006, 306.6796, 305.8462, 305, 
    304.141, 303.2689, 302.3836, 301.4848, 300.5725, 299.6465, 298.7066, 
    297.7528, 296.7849, 295.8029, 294.8067, 293.7964, 292.7718, 291.733, 
    290.6801, 289.6132, 288.5323, 287.4377, 286.3295, 285.2078, 284.0731, 
    282.9254, 281.7654, 280.5931, 279.4092, 278.214, 277.008, 275.7918, 
    274.5659, 273.331, 272.0877, 270.8367, 269.5787, 268.3145, 267.0447, 
    265.7703, 264.4921, 263.2108, 261.9273, 260.6426, 259.3574, 258.0727, 
    256.7892, 255.5079, 254.2297, 252.9553, 251.6855, 250.4213, 249.1633, 
    247.9123, 246.669, 245.4341, 244.2082, 242.992, 241.786, 240.5908, 
    239.4069, 238.2346, 237.0745, 235.9269, 234.7922, 233.6705, 232.5623, 
    231.4676, 230.3868, 229.3198, 228.267, 227.2282, 226.2036, 225.1933, 
    224.1971, 223.2151, 222.2472, 221.2934, 220.3535, 219.4275, 218.5152, 
    217.6164, 216.7311, 215.859, 215, 214.1539, 213.3204, 212.4994, 211.6906, 
    210.8939, 210.1091, 209.3358,
  309.8322, 309.055, 308.2668, 307.4674, 306.6566, 305.8342, 305, 304.1538, 
    303.2956, 302.425, 301.5421, 300.6465, 299.7383, 298.8173, 297.8834, 
    296.9366, 295.9767, 295.0037, 294.0176, 293.0185, 292.0062, 290.981, 
    289.9427, 288.8917, 287.8279, 286.7515, 285.6627, 284.5618, 283.4489, 
    282.3245, 281.1887, 280.042, 278.8848, 277.7174, 276.5403, 275.3541, 
    274.1592, 272.9563, 271.7458, 270.5284, 269.3048, 268.0757, 266.8416, 
    265.6035, 264.3618, 263.1175, 261.8713, 260.6239, 259.3761, 258.1287, 
    256.8825, 255.6382, 254.3966, 253.1584, 251.9243, 250.6952, 249.4716, 
    248.2542, 247.0437, 245.8408, 244.6459, 243.4597, 242.2826, 241.1152, 
    239.958, 238.8113, 237.6755, 236.5511, 235.4382, 234.3373, 233.2485, 
    232.1722, 231.1084, 230.0573, 229.019, 227.9938, 226.9815, 225.9824, 
    224.9963, 224.0233, 223.0634, 222.1166, 221.1827, 220.2617, 219.3535, 
    218.4579, 217.575, 216.7044, 215.8461, 215, 214.1658, 213.3434, 212.5326, 
    211.7332, 210.945, 210.1678,
  309.0078, 308.2274, 307.4367, 306.6353, 305.8231, 305, 304.1658, 303.3204, 
    302.4636, 301.5953, 300.7154, 299.8238, 298.9203, 298.005, 297.0777, 
    296.1384, 295.1871, 294.2237, 293.2482, 292.2607, 291.2611, 290.2497, 
    289.2263, 288.1913, 287.1447, 286.0866, 285.0173, 283.937, 282.8458, 
    281.7442, 280.6324, 279.5108, 278.3796, 277.2394, 276.0905, 274.9333, 
    273.7685, 272.5964, 271.4176, 270.2327, 269.0422, 267.8468, 266.6471, 
    265.4436, 264.2371, 263.0282, 261.8176, 260.606, 259.394, 258.1824, 
    256.9718, 255.7629, 254.5564, 253.353, 252.1532, 250.9578, 249.7673, 
    248.5824, 247.4036, 246.2315, 245.0666, 243.9095, 242.7606, 241.6204, 
    240.4892, 239.3676, 238.2558, 237.1542, 236.063, 234.9827, 233.9134, 
    232.8553, 231.8087, 230.7736, 229.7503, 228.7389, 227.7393, 226.7518, 
    225.7764, 224.8129, 223.8616, 222.9223, 221.995, 221.0797, 220.1762, 
    219.2846, 218.4047, 217.5364, 216.6796, 215.8342, 215, 214.1769, 
    213.3647, 212.5633, 211.7726, 210.9922,
  308.1911, 307.4082, 306.6155, 305.8128, 305, 304.1769, 303.3434, 302.4994, 
    301.6447, 300.7794, 299.9032, 299.0161, 298.1181, 297.2091, 296.289, 
    295.3578, 294.4155, 293.4621, 292.4977, 291.5222, 290.5357, 289.5383, 
    288.5301, 287.5113, 286.4819, 285.4421, 284.3922, 283.3323, 282.2627, 
    281.1836, 280.0953, 278.9982, 277.8926, 276.7789, 275.6573, 274.5285, 
    273.3927, 272.2505, 271.1024, 269.9487, 268.7902, 267.6272, 266.4604, 
    265.2903, 264.1175, 262.9426, 261.7661, 260.5888, 259.4112, 258.2339, 
    257.0574, 255.8825, 254.7097, 253.5396, 252.3728, 251.2098, 250.0513, 
    248.8976, 247.7495, 246.6073, 245.4715, 244.3427, 243.2211, 242.1074, 
    241.0018, 239.9047, 238.8164, 237.7373, 236.6677, 235.6078, 234.5579, 
    233.5181, 232.4887, 231.4699, 230.4617, 229.4643, 228.4779, 227.5023, 
    226.5379, 225.5845, 224.6422, 223.711, 222.7909, 221.8819, 220.9838, 
    220.0968, 219.2206, 218.3553, 217.5006, 216.6566, 215.8231, 215, 
    214.1872, 213.3845, 212.5918, 211.8089,
  307.382, 306.5973, 305.8033, 305, 304.1872, 303.3647, 302.5326, 301.6906, 
    300.8388, 299.977, 299.1052, 298.2233, 297.3313, 296.4291, 295.5167, 
    294.5941, 293.6614, 292.7184, 291.7654, 290.8022, 289.8291, 288.846, 
    287.8531, 286.8506, 285.8385, 284.817, 283.7864, 282.7467, 281.6984, 
    280.6415, 279.5764, 278.5034, 277.4227, 276.3348, 275.2399, 274.1385, 
    273.031, 271.9177, 270.7991, 269.6757, 268.5479, 267.4162, 266.2811, 
    265.1431, 264.0027, 262.8604, 261.7168, 260.5724, 259.4276, 258.2832, 
    257.1396, 255.9973, 254.8569, 253.7189, 252.5838, 251.4521, 250.3243, 
    249.2009, 248.0823, 246.969, 245.8615, 244.7601, 243.6652, 242.5773, 
    241.4967, 240.4236, 239.3585, 238.3016, 237.2533, 236.2136, 235.183, 
    234.1615, 233.1494, 232.1469, 231.154, 230.1709, 229.1978, 228.2346, 
    227.2816, 226.3386, 225.4059, 224.4833, 223.5709, 222.6687, 221.7767, 
    220.8948, 220.023, 219.1612, 218.3094, 217.4674, 216.6353, 215.8128, 215, 
    214.1967, 213.4027, 212.618,
  306.5805, 305.7946, 305, 304.1967, 303.3845, 302.5633, 301.7332, 300.8939, 
    300.0455, 299.1879, 298.321, 297.4449, 296.5594, 295.6646, 294.7604, 
    293.8469, 292.9241, 291.992, 291.0507, 290.1002, 289.1407, 288.1721, 
    287.1946, 286.2085, 285.2137, 284.2104, 283.1989, 282.1794, 281.152, 
    280.117, 279.0746, 278.0251, 276.9689, 275.9062, 274.8373, 273.7626, 
    272.6824, 271.5972, 270.5072, 269.413, 268.3148, 267.2133, 266.1087, 
    265.0016, 263.8923, 262.7814, 261.6693, 260.5565, 259.4435, 258.3307, 
    257.2186, 256.1077, 254.9984, 253.8913, 252.7867, 251.6852, 250.587, 
    249.4928, 248.4028, 247.3176, 246.2374, 245.1627, 244.0938, 243.0311, 
    241.9749, 240.9254, 239.883, 238.848, 237.8206, 236.8011, 235.7896, 
    234.7863, 233.7915, 232.8053, 231.8279, 230.8594, 229.8998, 228.9493, 
    228.008, 227.0759, 226.1531, 225.2396, 224.3354, 223.4406, 222.5551, 
    221.6789, 220.8121, 219.9545, 219.1061, 218.2668, 217.4367, 216.6155, 
    215.8033, 215, 214.2054, 213.4195,
  305.7865, 305, 304.2054, 303.4027, 302.5918, 301.7726, 300.945, 300.109, 
    299.2647, 298.4118, 297.5504, 296.6805, 295.8021, 294.9151, 294.0196, 
    293.1156, 292.2032, 291.2823, 290.353, 289.4154, 288.4696, 287.5157, 
    286.5538, 285.584, 284.6065, 283.6215, 282.629, 281.6293, 280.6226, 
    279.6091, 278.5891, 277.5627, 276.5303, 275.4922, 274.4485, 273.3998, 
    272.3462, 271.2881, 270.2259, 269.1599, 268.0904, 267.0179, 265.9428, 
    264.8654, 263.7861, 262.7054, 261.6237, 260.5413, 259.4587, 258.3763, 
    257.2946, 256.2139, 255.1346, 254.0572, 252.9821, 251.9096, 250.8401, 
    249.7741, 248.7119, 247.6538, 246.6002, 245.5514, 244.5078, 243.4697, 
    242.4373, 241.411, 240.3909, 239.3774, 238.3707, 237.371, 236.3785, 
    235.3935, 234.416, 233.4462, 232.4843, 231.5304, 230.5846, 229.647, 
    228.7177, 227.7968, 226.8844, 225.9804, 225.0849, 224.1979, 223.3195, 
    222.4496, 221.5882, 220.7353, 219.8909, 219.055, 218.2274, 217.4082, 
    216.5973, 215.7946, 215, 214.2135,
  305, 304.2135, 303.4195, 302.618, 301.8089, 300.9922, 300.1678, 299.3358, 
    298.4959, 297.6484, 296.793, 295.9299, 295.059, 294.1803, 293.2939, 
    292.3998, 291.498, 290.5886, 289.6716, 288.7472, 287.8153, 286.8762, 
    285.9299, 284.9766, 284.0163, 283.0493, 282.0757, 281.0956, 280.1093, 
    279.117, 278.1189, 277.1151, 276.1061, 275.0919, 274.073, 273.0494, 
    272.0217, 270.9899, 269.9545, 268.9158, 267.8741, 266.8297, 265.7829, 
    264.7342, 263.6839, 262.6322, 261.5797, 260.5266, 259.4734, 258.4203, 
    257.3678, 256.3161, 255.2658, 254.2171, 253.1703, 252.1259, 251.0842, 
    250.0455, 249.0101, 247.9783, 246.9505, 245.927, 244.9081, 243.8939, 
    242.8848, 241.8811, 240.883, 239.8907, 238.9044, 237.9244, 236.9507, 
    235.9837, 235.0234, 234.0701, 233.1238, 232.1847, 231.2529, 230.3284, 
    229.4114, 228.502, 227.6002, 226.7061, 225.8197, 224.941, 224.0701, 
    223.207, 222.3516, 221.5041, 220.6642, 219.8322, 219.0078, 218.1911, 
    217.382, 216.5805, 215.7865, 215 ;

 grid_latt =
  35.63342, 36.0016, 36.36466, 36.72248, 37.07492, 37.42188, 37.76321, 
    38.09881, 38.42853, 38.75225, 39.06984, 39.38117, 39.68611, 39.98453, 
    40.27629, 40.56128, 40.83934, 41.11036, 41.37419, 41.63073, 41.87982, 
    42.12135, 42.35519, 42.58122, 42.7993, 43.00933, 43.21118, 43.40474, 
    43.58989, 43.76653, 43.93454, 44.09382, 44.24429, 44.38583, 44.51836, 
    44.64181, 44.75608, 44.8611, 44.9568, 45.04311, 45.11999, 45.18737, 
    45.24522, 45.29348, 45.33213, 45.36115, 45.3805, 45.39018, 45.39018, 
    45.3805, 45.36115, 45.33213, 45.29348, 45.24522, 45.18737, 45.11999, 
    45.04311, 44.9568, 44.8611, 44.75608, 44.64181, 44.51836, 44.38583, 
    44.24429, 44.09382, 43.93454, 43.76653, 43.58989, 43.40474, 43.21118, 
    43.00933, 42.7993, 42.58122, 42.35519, 42.12135, 41.87982, 41.63073, 
    41.37419, 41.11036, 40.83934, 40.56128, 40.27629, 39.98453, 39.68611, 
    39.38117, 39.06984, 38.75225, 38.42853, 38.09881, 37.76321, 37.42188, 
    37.07492, 36.72248, 36.36466, 36.0016, 35.63342,
  36.0016, 36.38164, 36.75665, 37.12651, 37.49107, 37.8502, 38.20377, 
    38.55162, 38.89363, 39.22964, 39.55952, 39.88312, 40.20029, 40.51088, 
    40.81476, 41.11176, 41.40174, 41.68456, 41.96006, 42.2281, 42.48852, 
    42.74119, 42.98596, 43.22269, 43.45123, 43.67144, 43.8832, 44.08636, 
    44.28079, 44.46637, 44.64297, 44.81047, 44.96877, 45.11773, 45.25727, 
    45.38729, 45.50768, 45.61835, 45.71924, 45.81026, 45.89135, 45.96243, 
    46.02346, 46.07439, 46.11519, 46.14581, 46.16624, 46.17646, 46.17646, 
    46.16624, 46.14581, 46.11519, 46.07439, 46.02346, 45.96243, 45.89135, 
    45.81026, 45.71924, 45.61835, 45.50768, 45.38729, 45.25727, 45.11773, 
    44.96877, 44.81047, 44.64297, 44.46637, 44.28079, 44.08636, 43.8832, 
    43.67144, 43.45123, 43.22269, 42.98596, 42.74119, 42.48852, 42.2281, 
    41.96006, 41.68456, 41.40174, 41.11176, 40.81476, 40.51088, 40.20029, 
    39.88312, 39.55952, 39.22964, 38.89363, 38.55162, 38.20377, 37.8502, 
    37.49107, 37.12651, 36.75665, 36.38164, 36.0016,
  36.36466, 36.75665, 37.14373, 37.52576, 37.90258, 38.27405, 38.64002, 
    39.00033, 39.35483, 39.70337, 40.04577, 40.38189, 40.71156, 41.03462, 
    41.35089, 41.66023, 41.96246, 42.2574, 42.54491, 42.82481, 43.09693, 
    43.36111, 43.61718, 43.86499, 44.10437, 44.33515, 44.55719, 44.77034, 
    44.97443, 45.16932, 45.35488, 45.53096, 45.69742, 45.85415, 46.00101, 
    46.13791, 46.26471, 46.38132, 46.48764, 46.5836, 46.66909, 46.74407, 
    46.80845, 46.86219, 46.90523, 46.93755, 46.95911, 46.96989, 46.96989, 
    46.95911, 46.93755, 46.90523, 46.86219, 46.80845, 46.74407, 46.66909, 
    46.5836, 46.48764, 46.38132, 46.26471, 46.13791, 46.00101, 45.85415, 
    45.69742, 45.53096, 45.35488, 45.16932, 44.97443, 44.77034, 44.55719, 
    44.33515, 44.10437, 43.86499, 43.61718, 43.36111, 43.09693, 42.82481, 
    42.54491, 42.2574, 41.96246, 41.66023, 41.35089, 41.03462, 40.71156, 
    40.38189, 40.04577, 39.70337, 39.35483, 39.00033, 38.64002, 38.27405, 
    37.90258, 37.52576, 37.14373, 36.75665, 36.36466,
  36.72248, 37.12651, 37.52576, 37.92007, 38.30929, 38.69325, 39.07178, 
    39.44474, 39.81194, 40.17321, 40.52837, 40.87727, 41.2197, 41.5555, 
    41.88448, 42.20646, 42.52125, 42.82867, 43.12852, 43.42064, 43.70482, 
    43.98088, 44.24864, 44.50792, 44.75852, 45.00027, 45.23299, 45.45651, 
    45.67065, 45.87524, 46.07014, 46.25516, 46.43016, 46.595, 46.74953, 
    46.89362, 47.02713, 47.14996, 47.26199, 47.36312, 47.45325, 47.53231, 
    47.6002, 47.65689, 47.7023, 47.7364, 47.75915, 47.77053, 47.77053, 
    47.75915, 47.7364, 47.7023, 47.65689, 47.6002, 47.53231, 47.45325, 
    47.36312, 47.26199, 47.14996, 47.02713, 46.89362, 46.74953, 46.595, 
    46.43016, 46.25516, 46.07014, 45.87524, 45.67065, 45.45651, 45.23299, 
    45.00027, 44.75852, 44.50792, 44.24864, 43.98088, 43.70482, 43.42064, 
    43.12852, 42.82867, 42.52125, 42.20646, 41.88448, 41.5555, 41.2197, 
    40.87727, 40.52837, 40.17321, 39.81194, 39.44474, 39.07178, 38.69325, 
    38.30929, 37.92007, 37.52576, 37.12651, 36.72248,
  37.07492, 37.49107, 37.90258, 38.30929, 38.71102, 39.10761, 39.49888, 
    39.88465, 40.26473, 40.63895, 41.00711, 41.36901, 41.72447, 42.07329, 
    42.41526, 42.75019, 43.07787, 43.39809, 43.71065, 44.01534, 44.31195, 
    44.60027, 44.88011, 45.15124, 45.41347, 45.66659, 45.91039, 46.14469, 
    46.36929, 46.58398, 46.7886, 46.98296, 47.16688, 47.34019, 47.50273, 
    47.65435, 47.79491, 47.92425, 48.04226, 48.14882, 48.24382, 48.32716, 
    48.39876, 48.45854, 48.50644, 48.54241, 48.56641, 48.57842, 48.57842, 
    48.56641, 48.54241, 48.50644, 48.45854, 48.39876, 48.32716, 48.24382, 
    48.14882, 48.04226, 47.92425, 47.79491, 47.65435, 47.50273, 47.34019, 
    47.16688, 46.98296, 46.7886, 46.58398, 46.36929, 46.14469, 45.91039, 
    45.66659, 45.41347, 45.15124, 44.88011, 44.60027, 44.31195, 44.01534, 
    43.71065, 43.39809, 43.07787, 42.75019, 42.41526, 42.07329, 41.72447, 
    41.36901, 41.00711, 40.63895, 40.26473, 39.88465, 39.49888, 39.10761, 
    38.71102, 38.30929, 37.90258, 37.49107, 37.07492,
  37.42188, 37.8502, 38.27405, 38.69325, 39.10761, 39.51696, 39.9211, 
    40.31985, 40.71301, 41.10036, 41.48173, 41.85689, 42.22562, 42.58773, 
    42.94299, 43.29116, 43.63205, 43.9654, 44.29101, 44.60864, 44.91806, 
    45.21903, 45.51133, 45.79473, 46.06899, 46.33389, 46.5892, 46.83469, 
    47.07016, 47.29537, 47.51012, 47.71421, 47.90744, 48.08961, 48.26053, 
    48.42004, 48.56796, 48.70414, 48.82842, 48.94068, 49.04079, 49.12864, 
    49.20412, 49.26716, 49.31768, 49.35562, 49.38094, 49.3936, 49.3936, 
    49.38094, 49.35562, 49.31768, 49.26716, 49.20412, 49.12864, 49.04079, 
    48.94068, 48.82842, 48.70414, 48.56796, 48.42004, 48.26053, 48.08961, 
    47.90744, 47.71421, 47.51012, 47.29537, 47.07016, 46.83469, 46.5892, 
    46.33389, 46.06899, 45.79473, 45.51133, 45.21903, 44.91806, 44.60864, 
    44.29101, 43.9654, 43.63205, 43.29116, 42.94299, 42.58773, 42.22562, 
    41.85689, 41.48173, 41.10036, 40.71301, 40.31985, 39.9211, 39.51696, 
    39.10761, 38.69325, 38.27405, 37.8502, 37.42188,
  37.76321, 38.20377, 38.64002, 39.07178, 39.49888, 39.9211, 40.33826, 
    40.75014, 41.15653, 41.55723, 41.95201, 42.34064, 42.7229, 43.09856, 
    43.46738, 43.82911, 44.18351, 44.53034, 44.86935, 45.20028, 45.52287, 
    45.83688, 46.14204, 46.43811, 46.72482, 47.00192, 47.26916, 47.52629, 
    47.77305, 48.0092, 48.23452, 48.44876, 48.6517, 48.84312, 49.02282, 
    49.19058, 49.34622, 49.48956, 49.62043, 49.73867, 49.84415, 49.93674, 
    50.01631, 50.08277, 50.13604, 50.17606, 50.20276, 50.21612, 50.21612, 
    50.20276, 50.17606, 50.13604, 50.08277, 50.01631, 49.93674, 49.84415, 
    49.73867, 49.62043, 49.48956, 49.34622, 49.19058, 49.02282, 48.84312, 
    48.6517, 48.44876, 48.23452, 48.0092, 47.77305, 47.52629, 47.26916, 
    47.00192, 46.72482, 46.43811, 46.14204, 45.83688, 45.52287, 45.20028, 
    44.86935, 44.53034, 44.18351, 43.82911, 43.46738, 43.09856, 42.7229, 
    42.34064, 41.95201, 41.55723, 41.15653, 40.75014, 40.33826, 39.9211, 
    39.49888, 39.07178, 38.64002, 38.20377, 37.76321,
  38.09881, 38.55162, 39.00033, 39.44474, 39.88465, 40.31985, 40.75014, 
    41.17529, 41.59509, 42.0093, 42.41769, 42.82002, 43.21604, 43.60551, 
    43.98816, 44.36374, 44.73198, 45.0926, 45.44535, 45.78994, 46.12609, 
    46.45353, 46.77196, 47.08112, 47.3807, 47.67044, 47.95004, 48.21923, 
    48.47774, 48.72528, 48.9616, 49.18642, 49.39951, 49.6006, 49.78946, 
    49.96586, 50.12959, 50.28045, 50.41822, 50.54276, 50.65387, 50.75143, 
    50.83531, 50.90538, 50.96155, 51.00375, 51.03191, 51.046, 51.046, 
    51.03191, 51.00375, 50.96155, 50.90538, 50.83531, 50.75143, 50.65387, 
    50.54276, 50.41822, 50.28045, 50.12959, 49.96586, 49.78946, 49.6006, 
    49.39951, 49.18642, 48.9616, 48.72528, 48.47774, 48.21923, 47.95004, 
    47.67044, 47.3807, 47.08112, 46.77196, 46.45353, 46.12609, 45.78994, 
    45.44535, 45.0926, 44.73198, 44.36374, 43.98816, 43.60551, 43.21604, 
    42.82002, 42.41769, 42.0093, 41.59509, 41.17529, 40.75014, 40.31985, 
    39.88465, 39.44474, 39.00033, 38.55162, 38.09881,
  38.42853, 38.89363, 39.35483, 39.81194, 40.26473, 40.71301, 41.15653, 
    41.59509, 42.02843, 42.45632, 42.87851, 43.29474, 43.70475, 44.10828, 
    44.50503, 44.89474, 45.27712, 45.65187, 46.0187, 46.37732, 46.72741, 
    47.06866, 47.40077, 47.72343, 48.03632, 48.33913, 48.63155, 48.91327, 
    49.18397, 49.44336, 49.69113, 49.927, 50.15067, 50.36186, 50.56031, 
    50.74577, 50.91797, 51.0767, 51.22174, 51.35287, 51.46992, 51.57272, 
    51.66111, 51.73498, 51.7942, 51.8387, 51.8684, 51.88326, 51.88326, 
    51.8684, 51.8387, 51.7942, 51.73498, 51.66111, 51.57272, 51.46992, 
    51.35287, 51.22174, 51.0767, 50.91797, 50.74577, 50.56031, 50.36186, 
    50.15067, 49.927, 49.69113, 49.44336, 49.18397, 48.91327, 48.63155, 
    48.33913, 48.03632, 47.72343, 47.40077, 47.06866, 46.72741, 46.37732, 
    46.0187, 45.65187, 45.27712, 44.89474, 44.50503, 44.10828, 43.70475, 
    43.29474, 42.87851, 42.45632, 42.02843, 41.59509, 41.15653, 40.71301, 
    40.26473, 39.81194, 39.35483, 38.89363, 38.42853,
  38.75225, 39.22964, 39.70337, 40.17321, 40.63895, 41.10036, 41.55723, 
    42.0093, 42.45632, 42.89805, 43.33421, 43.76454, 44.18875, 44.60656, 
    45.01768, 45.4218, 45.81862, 46.20782, 46.58908, 46.96207, 47.32647, 
    47.68195, 48.02814, 48.36473, 48.69137, 49.00771, 49.3134, 49.6081, 
    49.89148, 50.16318, 50.42288, 50.67025, 50.90497, 51.12672, 51.33521, 
    51.53014, 51.71123, 51.87823, 52.03088, 52.16895, 52.29223, 52.40054, 
    52.4937, 52.57156, 52.63401, 52.68093, 52.71225, 52.72793, 52.72793, 
    52.71225, 52.68093, 52.63401, 52.57156, 52.4937, 52.40054, 52.29223, 
    52.16895, 52.03088, 51.87823, 51.71123, 51.53014, 51.33521, 51.12672, 
    50.90497, 50.67025, 50.42288, 50.16318, 49.89148, 49.6081, 49.3134, 
    49.00771, 48.69137, 48.36473, 48.02814, 47.68195, 47.32647, 46.96207, 
    46.58908, 46.20782, 45.81862, 45.4218, 45.01768, 44.60656, 44.18875, 
    43.76454, 43.33421, 42.89805, 42.45632, 42.0093, 41.55723, 41.10036, 
    40.63895, 40.17321, 39.70337, 39.22964, 38.75225,
  39.06984, 39.55952, 40.04577, 40.52837, 41.00711, 41.48173, 41.95201, 
    42.41769, 42.87851, 43.33421, 43.7845, 44.22911, 44.66773, 45.10006, 
    45.52579, 45.94459, 46.35614, 46.76009, 47.15612, 47.54385, 47.92294, 
    48.29302, 48.65372, 49.00467, 49.3455, 49.67582, 49.99525, 50.30342, 
    50.59995, 50.88446, 51.15658, 51.41594, 51.66219, 51.89498, 52.11396, 
    52.31881, 52.50922, 52.68489, 52.84554, 52.99091, 53.12075, 53.23486, 
    53.33304, 53.41512, 53.48095, 53.53043, 53.56347, 53.58, 53.58, 53.56347, 
    53.53043, 53.48095, 53.41512, 53.33304, 53.23486, 53.12075, 52.99091, 
    52.84554, 52.68489, 52.50922, 52.31881, 52.11396, 51.89498, 51.66219, 
    51.41594, 51.15658, 50.88446, 50.59995, 50.30342, 49.99525, 49.67582, 
    49.3455, 49.00467, 48.65372, 48.29302, 47.92294, 47.54385, 47.15612, 
    46.76009, 46.35614, 45.94459, 45.52579, 45.10006, 44.66773, 44.22911, 
    43.7845, 43.33421, 42.87851, 42.41769, 41.95201, 41.48173, 41.00711, 
    40.52837, 40.04577, 39.55952, 39.06984,
  39.38117, 39.88312, 40.38189, 40.87727, 41.36901, 41.85689, 42.34064, 
    42.82002, 43.29474, 43.76454, 44.22911, 44.68816, 45.14137, 45.58843, 
    46.029, 46.46275, 46.88931, 47.30833, 47.71944, 48.12227, 48.51642, 
    48.9015, 49.27712, 49.64286, 49.99833, 50.34309, 50.67675, 50.99888, 
    51.30906, 51.60688, 51.89192, 52.16379, 52.42207, 52.66639, 52.89635, 
    53.1116, 53.31178, 53.49655, 53.6656, 53.81864, 53.95539, 54.07561, 
    54.17908, 54.26561, 54.33502, 54.3872, 54.42204, 54.43948, 54.43948, 
    54.42204, 54.3872, 54.33502, 54.26561, 54.17908, 54.07561, 53.95539, 
    53.81864, 53.6656, 53.49655, 53.31178, 53.1116, 52.89635, 52.66639, 
    52.42207, 52.16379, 51.89192, 51.60688, 51.30906, 50.99888, 50.67675, 
    50.34309, 49.99833, 49.64286, 49.27712, 48.9015, 48.51642, 48.12227, 
    47.71944, 47.30833, 46.88931, 46.46275, 46.029, 45.58843, 45.14137, 
    44.68816, 44.22911, 43.76454, 43.29474, 42.82002, 42.34064, 41.85689, 
    41.36901, 40.87727, 40.38189, 39.88312, 39.38117,
  39.68611, 40.20029, 40.71156, 41.2197, 41.72447, 42.22562, 42.7229, 
    43.21604, 43.70475, 44.18875, 44.66773, 45.14137, 45.60936, 46.07135, 
    46.52699, 46.97591, 47.41776, 47.85214, 48.27867, 48.69693, 49.10651, 
    49.50698, 49.89793, 50.2789, 50.64946, 51.00915, 51.35751, 51.6941, 
    52.01844, 52.33009, 52.62858, 52.91348, 53.18432, 53.44069, 53.68214, 
    53.90828, 54.1187, 54.31304, 54.49093, 54.65204, 54.79607, 54.92273, 
    55.03177, 55.12299, 55.19618, 55.25121, 55.28796, 55.30635, 55.30635, 
    55.28796, 55.25121, 55.19618, 55.12299, 55.03177, 54.92273, 54.79607, 
    54.65204, 54.49093, 54.31304, 54.1187, 53.90828, 53.68214, 53.44069, 
    53.18432, 52.91348, 52.62858, 52.33009, 52.01844, 51.6941, 51.35751, 
    51.00915, 50.64946, 50.2789, 49.89793, 49.50698, 49.10651, 48.69693, 
    48.27867, 47.85214, 47.41776, 46.97591, 46.52699, 46.07135, 45.60936, 
    45.14137, 44.66773, 44.18875, 43.70475, 43.21604, 42.7229, 42.22562, 
    41.72447, 41.2197, 40.71156, 40.20029, 39.68611,
  39.98453, 40.51088, 41.03462, 41.5555, 42.07329, 42.58773, 43.09856, 
    43.60551, 44.10828, 44.60656, 45.10006, 45.58843, 46.07135, 46.54844, 
    47.01936, 47.4837, 47.94109, 48.39112, 48.83337, 49.2674, 49.69277, 
    50.10903, 50.51572, 50.91235, 51.29846, 51.67355, 52.03711, 52.38867, 
    52.7277, 53.05371, 53.3662, 53.66467, 53.94862, 54.21758, 54.47105, 
    54.70861, 54.92978, 55.13416, 55.32135, 55.49096, 55.64265, 55.7761, 
    55.89104, 55.9872, 56.06439, 56.12244, 56.1612, 56.18061, 56.18061, 
    56.1612, 56.12244, 56.06439, 55.9872, 55.89104, 55.7761, 55.64265, 
    55.49096, 55.32135, 55.13416, 54.92978, 54.70861, 54.47105, 54.21758, 
    53.94862, 53.66467, 53.3662, 53.05371, 52.7277, 52.38867, 52.03711, 
    51.67355, 51.29846, 50.91235, 50.51572, 50.10903, 49.69277, 49.2674, 
    48.83337, 48.39112, 47.94109, 47.4837, 47.01936, 46.54844, 46.07135, 
    45.58843, 45.10006, 44.60656, 44.10828, 43.60551, 43.09856, 42.58773, 
    42.07329, 41.5555, 41.03462, 40.51088, 39.98453,
  40.27629, 40.81476, 41.35089, 41.88448, 42.41526, 42.94299, 43.46738, 
    43.98816, 44.50503, 45.01768, 45.52579, 46.029, 46.52699, 47.01936, 
    47.50573, 47.98571, 48.45889, 48.92484, 49.3831, 49.83323, 50.27475, 
    50.70718, 51.13002, 51.54275, 51.94487, 52.33583, 52.7151, 53.08215, 
    53.43641, 53.77734, 54.10438, 54.41699, 54.71461, 54.99673, 55.2628, 
    55.51231, 55.74477, 55.95971, 56.15667, 56.33524, 56.49501, 56.63563, 
    56.75679, 56.85819, 56.93961, 57.00084, 57.04174, 57.06222, 57.06222, 
    57.04174, 57.00084, 56.93961, 56.85819, 56.75679, 56.63563, 56.49501, 
    56.33524, 56.15667, 55.95971, 55.74477, 55.51231, 55.2628, 54.99673, 
    54.71461, 54.41699, 54.10438, 53.77734, 53.43641, 53.08215, 52.7151, 
    52.33583, 51.94487, 51.54275, 51.13002, 50.70718, 50.27475, 49.83323, 
    49.3831, 48.92484, 48.45889, 47.98571, 47.50573, 47.01936, 46.52699, 
    46.029, 45.52579, 45.01768, 44.50503, 43.98816, 43.46738, 42.94299, 
    42.41526, 41.88448, 41.35089, 40.81476, 40.27629,
  40.56128, 41.11176, 41.66023, 42.20646, 42.75019, 43.29116, 43.82911, 
    44.36374, 44.89474, 45.4218, 45.94459, 46.46275, 46.97591, 47.4837, 
    47.98571, 48.48154, 48.97073, 49.45285, 49.92742, 50.39396, 50.85197, 
    51.30094, 51.74033, 52.16959, 52.58817, 52.9955, 53.39099, 53.77406, 
    54.14409, 54.5005, 54.84268, 55.17002, 55.48191, 55.77778, 56.05703, 
    56.31908, 56.56339, 56.78943, 56.99669, 57.18469, 57.35299, 57.50119, 
    57.62892, 57.73586, 57.82175, 57.88636, 57.92953, 57.95115, 57.95115, 
    57.92953, 57.88636, 57.82175, 57.73586, 57.62892, 57.50119, 57.35299, 
    57.18469, 56.99669, 56.78943, 56.56339, 56.31908, 56.05703, 55.77778, 
    55.48191, 55.17002, 54.84268, 54.5005, 54.14409, 53.77406, 53.39099, 
    52.9955, 52.58817, 52.16959, 51.74033, 51.30094, 50.85197, 50.39396, 
    49.92742, 49.45285, 48.97073, 48.48154, 47.98571, 47.4837, 46.97591, 
    46.46275, 45.94459, 45.4218, 44.89474, 44.36374, 43.82911, 43.29116, 
    42.75019, 42.20646, 41.66023, 41.11176, 40.56128,
  40.83934, 41.40174, 41.96246, 42.52125, 43.07787, 43.63205, 44.18351, 
    44.73198, 45.27712, 45.81862, 46.35614, 46.88931, 47.41776, 47.94109, 
    48.45889, 48.97073, 49.47615, 49.97467, 50.46582, 50.94908, 51.42391, 
    51.88978, 52.34612, 52.79234, 53.22784, 53.65202, 54.06424, 54.46386, 
    54.85024, 55.22271, 55.58062, 55.9233, 56.25008, 56.56032, 56.85336, 
    57.12857, 57.38533, 57.62305, 57.84115, 58.0391, 58.21642, 58.37262, 
    58.50731, 58.62013, 58.71076, 58.77895, 58.82452, 58.84734, 58.84734, 
    58.82452, 58.77895, 58.71076, 58.62013, 58.50731, 58.37262, 58.21642, 
    58.0391, 57.84115, 57.62305, 57.38533, 57.12857, 56.85336, 56.56032, 
    56.25008, 55.9233, 55.58062, 55.22271, 54.85024, 54.46386, 54.06424, 
    53.65202, 53.22784, 52.79234, 52.34612, 51.88978, 51.42391, 50.94908, 
    50.46582, 49.97467, 49.47615, 48.97073, 48.45889, 47.94109, 47.41776, 
    46.88931, 46.35614, 45.81862, 45.27712, 44.73198, 44.18351, 43.63205, 
    43.07787, 42.52125, 41.96246, 41.40174, 40.83934,
  41.11036, 41.68456, 42.2574, 42.82867, 43.39809, 43.9654, 44.53034, 
    45.0926, 45.65187, 46.20782, 46.76009, 47.30833, 47.85214, 48.39112, 
    48.92484, 49.45285, 49.97467, 50.48983, 50.9978, 51.49806, 51.99004, 
    52.47316, 52.94683, 53.41042, 53.8633, 54.30482, 54.73428, 55.15101, 
    55.55429, 55.94343, 56.31768, 56.67633, 57.01865, 57.34391, 57.65139, 
    57.9404, 58.21024, 58.46024, 58.68978, 58.89825, 59.08508, 59.24976, 
    59.39183, 59.51086, 59.60653, 59.67853, 59.72665, 59.75075, 59.75075, 
    59.72665, 59.67853, 59.60653, 59.51086, 59.39183, 59.24976, 59.08508, 
    58.89825, 58.68978, 58.46024, 58.21024, 57.9404, 57.65139, 57.34391, 
    57.01865, 56.67633, 56.31768, 55.94343, 55.55429, 55.15101, 54.73428, 
    54.30482, 53.8633, 53.41042, 52.94683, 52.47316, 51.99004, 51.49806, 
    50.9978, 50.48983, 49.97467, 49.45285, 48.92484, 48.39112, 47.85214, 
    47.30833, 46.76009, 46.20782, 45.65187, 45.0926, 44.53034, 43.9654, 
    43.39809, 42.82867, 42.2574, 41.68456, 41.11036,
  41.37419, 41.96006, 42.54491, 43.12852, 43.71065, 44.29101, 44.86935, 
    45.44535, 46.0187, 46.58908, 47.15612, 47.71944, 48.27867, 48.83337, 
    49.3831, 49.92742, 50.46582, 50.9978, 51.52283, 52.04035, 52.54977, 
    53.05048, 53.54185, 54.02324, 54.49394, 54.95327, 55.40049, 55.83487, 
    56.25565, 56.66205, 57.05328, 57.42855, 57.78707, 58.12803, 58.45065, 
    58.75413, 59.03772, 59.30067, 59.54227, 59.76184, 59.95875, 60.13241, 
    60.2823, 60.40795, 60.50896, 60.58501, 60.63584, 60.6613, 60.6613, 
    60.63584, 60.58501, 60.50896, 60.40795, 60.2823, 60.13241, 59.95875, 
    59.76184, 59.54227, 59.30067, 59.03772, 58.75413, 58.45065, 58.12803, 
    57.78707, 57.42855, 57.05328, 56.66205, 56.25565, 55.83487, 55.40049, 
    54.95327, 54.49394, 54.02324, 53.54185, 53.05048, 52.54977, 52.04035, 
    51.52283, 50.9978, 50.46582, 49.92742, 49.3831, 48.83337, 48.27867, 
    47.71944, 47.15612, 46.58908, 46.0187, 45.44535, 44.86935, 44.29101, 
    43.71065, 43.12852, 42.54491, 41.96006, 41.37419,
  41.63073, 42.2281, 42.82481, 43.42064, 44.01534, 44.60864, 45.20028, 
    45.78994, 46.37732, 46.96207, 47.54385, 48.12227, 48.69693, 49.2674, 
    49.83323, 50.39396, 50.94908, 51.49806, 52.04035, 52.57537, 53.10251, 
    53.62113, 54.13057, 54.63013, 55.11909, 55.59671, 56.06221, 56.51479, 
    56.95364, 57.37793, 57.78679, 58.17936, 58.55478, 58.91215, 59.25061, 
    59.56929, 59.86734, 60.14393, 60.39826, 60.62958, 60.83716, 61.02035, 
    61.17855, 61.31122, 61.41792, 61.49828, 61.55201, 61.57893, 61.57893, 
    61.55201, 61.49828, 61.41792, 61.31122, 61.17855, 61.02035, 60.83716, 
    60.62958, 60.39826, 60.14393, 59.86734, 59.56929, 59.25061, 58.91215, 
    58.55478, 58.17936, 57.78679, 57.37793, 56.95364, 56.51479, 56.06221, 
    55.59671, 55.11909, 54.63013, 54.13057, 53.62113, 53.10251, 52.57537, 
    52.04035, 51.49806, 50.94908, 50.39396, 49.83323, 49.2674, 48.69693, 
    48.12227, 47.54385, 46.96207, 46.37732, 45.78994, 45.20028, 44.60864, 
    44.01534, 43.42064, 42.82481, 42.2281, 41.63073,
  41.87982, 42.48852, 43.09693, 43.70482, 44.31195, 44.91806, 45.52287, 
    46.12609, 46.72741, 47.32647, 47.92294, 48.51642, 49.10651, 49.69277, 
    50.27475, 50.85197, 51.42391, 51.99004, 52.54977, 53.10251, 53.64762, 
    54.18444, 54.71228, 55.2304, 55.73805, 56.23442, 56.7187, 57.19004, 
    57.64757, 58.09037, 58.51752, 58.92809, 59.32111, 59.69563, 60.05069, 
    60.38533, 60.6986, 60.98957, 61.25736, 61.50111, 61.72001, 61.91332, 
    62.08035, 62.22052, 62.33329, 62.41824, 62.47506, 62.50353, 62.50353, 
    62.47506, 62.41824, 62.33329, 62.22052, 62.08035, 61.91332, 61.72001, 
    61.50111, 61.25736, 60.98957, 60.6986, 60.38533, 60.05069, 59.69563, 
    59.32111, 58.92809, 58.51752, 58.09037, 57.64757, 57.19004, 56.7187, 
    56.23442, 55.73805, 55.2304, 54.71228, 54.18444, 53.64762, 53.10251, 
    52.54977, 51.99004, 51.42391, 50.85197, 50.27475, 49.69277, 49.10651, 
    48.51642, 47.92294, 47.32647, 46.72741, 46.12609, 45.52287, 44.91806, 
    44.31195, 43.70482, 43.09693, 42.48852, 41.87982,
  42.12135, 42.74119, 43.36111, 43.98088, 44.60027, 45.21903, 45.83688, 
    46.45353, 47.06866, 47.68195, 48.29302, 48.9015, 49.50698, 50.10903, 
    50.70718, 51.30094, 51.88978, 52.47316, 53.05048, 53.62113, 54.18444, 
    54.73974, 55.28629, 55.82333, 56.35006, 56.86565, 57.36921, 57.85986, 
    58.33664, 58.79859, 59.24471, 59.67398, 60.08537, 60.47782, 60.85027, 
    61.20166, 61.53094, 61.8371, 62.11912, 62.37604, 62.60696, 62.81103, 
    62.98748, 63.13563, 63.25488, 63.34475, 63.40488, 63.43501, 63.43501, 
    63.40488, 63.34475, 63.25488, 63.13563, 62.98748, 62.81103, 62.60696, 
    62.37604, 62.11912, 61.8371, 61.53094, 61.20166, 60.85027, 60.47782, 
    60.08537, 59.67398, 59.24471, 58.79859, 58.33664, 57.85986, 57.36921, 
    56.86565, 56.35006, 55.82333, 55.28629, 54.73974, 54.18444, 53.62113, 
    53.05048, 52.47316, 51.88978, 51.30094, 50.70718, 50.10903, 49.50698, 
    48.9015, 48.29302, 47.68195, 47.06866, 46.45353, 45.83688, 45.21903, 
    44.60027, 43.98088, 43.36111, 42.74119, 42.12135,
  42.35519, 42.98596, 43.61718, 44.24864, 44.88011, 45.51133, 46.14204, 
    46.77196, 47.40077, 48.02814, 48.65372, 49.27712, 49.89793, 50.51572, 
    51.13002, 51.74033, 52.34612, 52.94683, 53.54185, 54.13057, 54.71228, 
    55.28629, 55.85184, 56.40814, 56.95434, 57.48957, 58.01291, 58.52339, 
    59.02002, 59.50176, 59.96754, 60.41625, 60.84677, 61.25794, 61.64861, 
    62.0176, 62.36376, 62.68594, 62.98302, 63.25393, 63.49763, 63.71317, 
    63.89967, 64.05634, 64.18253, 64.27767, 64.34134, 64.37325, 64.37325, 
    64.34134, 64.27767, 64.18253, 64.05634, 63.89967, 63.71317, 63.49763, 
    63.25393, 62.98302, 62.68594, 62.36376, 62.0176, 61.64861, 61.25794, 
    60.84677, 60.41625, 59.96754, 59.50176, 59.02002, 58.52339, 58.01291, 
    57.48957, 56.95434, 56.40814, 55.85184, 55.28629, 54.71228, 54.13057, 
    53.54185, 52.94683, 52.34612, 51.74033, 51.13002, 50.51572, 49.89793, 
    49.27712, 48.65372, 48.02814, 47.40077, 46.77196, 46.14204, 45.51133, 
    44.88011, 44.24864, 43.61718, 42.98596, 42.35519,
  42.58122, 43.22269, 43.86499, 44.50792, 45.15124, 45.79473, 46.43811, 
    47.08112, 47.72343, 48.36473, 49.00467, 49.64286, 50.2789, 50.91235, 
    51.54275, 52.16959, 52.79234, 53.41042, 54.02324, 54.63013, 55.2304, 
    55.82333, 56.40814, 56.98399, 57.55002, 58.1053, 58.64888, 59.17973, 
    59.6968, 60.19897, 60.6851, 61.154, 61.60444, 62.03517, 62.44493, 
    62.83242, 63.19636, 63.53547, 63.84851, 64.13426, 64.39157, 64.61935, 
    64.81659, 64.98241, 65.11604, 65.21684, 65.28431, 65.31813, 65.31813, 
    65.28431, 65.21684, 65.11604, 64.98241, 64.81659, 64.61935, 64.39157, 
    64.13426, 63.84851, 63.53547, 63.19636, 62.83242, 62.44493, 62.03517, 
    61.60444, 61.154, 60.6851, 60.19897, 59.6968, 59.17973, 58.64888, 
    58.1053, 57.55002, 56.98399, 56.40814, 55.82333, 55.2304, 54.63013, 
    54.02324, 53.41042, 52.79234, 52.16959, 51.54275, 50.91235, 50.2789, 
    49.64286, 49.00467, 48.36473, 47.72343, 47.08112, 46.43811, 45.79473, 
    45.15124, 44.50792, 43.86499, 43.22269, 42.58122,
  42.7993, 43.45123, 44.10437, 44.75852, 45.41347, 46.06899, 46.72482, 
    47.3807, 48.03632, 48.69137, 49.3455, 49.99833, 50.64946, 51.29846, 
    51.94487, 52.58817, 53.22784, 53.8633, 54.49394, 55.11909, 55.73805, 
    56.35006, 56.95434, 57.55002, 58.1362, 58.71193, 59.2762, 59.82792, 
    60.36599, 60.88923, 61.39641, 61.88625, 62.35743, 62.80859, 63.23833, 
    63.64526, 64.02795, 64.38497, 64.71494, 65.01648, 65.2883, 65.52915, 
    65.73791, 65.91354, 66.05517, 66.16206, 66.23363, 66.26952, 66.26952, 
    66.23363, 66.16206, 66.05517, 65.91354, 65.73791, 65.52915, 65.2883, 
    65.01648, 64.71494, 64.38497, 64.02795, 63.64526, 63.23833, 62.80859, 
    62.35743, 61.88625, 61.39641, 60.88923, 60.36599, 59.82792, 59.2762, 
    58.71193, 58.1362, 57.55002, 56.95434, 56.35006, 55.73805, 55.11909, 
    54.49394, 53.8633, 53.22784, 52.58817, 51.94487, 51.29846, 50.64946, 
    49.99833, 49.3455, 48.69137, 48.03632, 47.3807, 46.72482, 46.06899, 
    45.41347, 44.75852, 44.10437, 43.45123, 42.7993,
  43.00933, 43.67144, 44.33515, 45.00027, 45.66659, 46.33389, 47.00192, 
    47.67044, 48.33913, 49.00771, 49.67582, 50.34309, 51.00915, 51.67355, 
    52.33583, 52.9955, 53.65202, 54.30482, 54.95327, 55.59671, 56.23442, 
    56.86565, 57.48957, 58.1053, 58.71193, 59.30845, 59.89382, 60.4669, 
    61.02654, 61.57146, 62.10038, 62.61193, 63.10468, 63.57715, 64.02785, 
    64.4552, 64.85765, 65.23363, 65.58157, 65.89993, 66.18724, 66.44211, 
    66.66322, 66.84942, 66.99967, 67.11313, 67.18914, 67.22726, 67.22726, 
    67.18914, 67.11313, 66.99967, 66.84942, 66.66322, 66.44211, 66.18724, 
    65.89993, 65.58157, 65.23363, 64.85765, 64.4552, 64.02785, 63.57715, 
    63.10468, 62.61193, 62.10038, 61.57146, 61.02654, 60.4669, 59.89382, 
    59.30845, 58.71193, 58.1053, 57.48957, 56.86565, 56.23442, 55.59671, 
    54.95327, 54.30482, 53.65202, 52.9955, 52.33583, 51.67355, 51.00915, 
    50.34309, 49.67582, 49.00771, 48.33913, 47.67044, 47.00192, 46.33389, 
    45.66659, 45.00027, 44.33515, 43.67144, 43.00933,
  43.21118, 43.8832, 44.55719, 45.23299, 45.91039, 46.5892, 47.26916, 
    47.95004, 48.63155, 49.3134, 49.99525, 50.67675, 51.35751, 52.03711, 
    52.7151, 53.39099, 54.06424, 54.73428, 55.40049, 56.06221, 56.7187, 
    57.36921, 58.01291, 58.64888, 59.2762, 59.89382, 60.50066, 61.09555, 
    61.67727, 62.2445, 62.79585, 63.32987, 63.84503, 64.33974, 64.81236, 
    65.26118, 65.68449, 66.08053, 66.44756, 66.78387, 67.08776, 67.35767, 
    67.59209, 67.78967, 67.94925, 68.06983, 68.15065, 68.19119, 68.19119, 
    68.15065, 68.06983, 67.94925, 67.78967, 67.59209, 67.35767, 67.08776, 
    66.78387, 66.44756, 66.08053, 65.68449, 65.26118, 64.81236, 64.33974, 
    63.84503, 63.32987, 62.79585, 62.2445, 61.67727, 61.09555, 60.50066, 
    59.89382, 59.2762, 58.64888, 58.01291, 57.36921, 56.7187, 56.06221, 
    55.40049, 54.73428, 54.06424, 53.39099, 52.7151, 52.03711, 51.35751, 
    50.67675, 49.99525, 49.3134, 48.63155, 47.95004, 47.26916, 46.5892, 
    45.91039, 45.23299, 44.55719, 43.8832, 43.21118,
  43.40474, 44.08636, 44.77034, 45.45651, 46.14469, 46.83469, 47.52629, 
    48.21923, 48.91327, 49.6081, 50.30342, 50.99888, 51.6941, 52.38867, 
    53.08215, 53.77406, 54.46386, 55.15101, 55.83487, 56.51479, 57.19004, 
    57.85986, 58.52339, 59.17973, 59.82792, 60.4669, 61.09555, 61.71267, 
    62.31697, 62.90707, 63.48152, 64.03877, 64.57719, 65.09508, 65.59063, 
    66.06201, 66.50732, 66.92463, 67.31198, 67.66744, 67.98912, 68.2752, 
    68.52398, 68.7339, 68.90359, 69.03191, 69.11797, 69.16115, 69.16115, 
    69.11797, 69.03191, 68.90359, 68.7339, 68.52398, 68.2752, 67.98912, 
    67.66744, 67.31198, 66.92463, 66.50732, 66.06201, 65.59063, 65.09508, 
    64.57719, 64.03877, 63.48152, 62.90707, 62.31697, 61.71267, 61.09555, 
    60.4669, 59.82792, 59.17973, 58.52339, 57.85986, 57.19004, 56.51479, 
    55.83487, 55.15101, 54.46386, 53.77406, 53.08215, 52.38867, 51.6941, 
    50.99888, 50.30342, 49.6081, 48.91327, 48.21923, 47.52629, 46.83469, 
    46.14469, 45.45651, 44.77034, 44.08636, 43.40474,
  43.58989, 44.28079, 44.97443, 45.67065, 46.36929, 47.07016, 47.77305, 
    48.47774, 49.18397, 49.89148, 50.59995, 51.30906, 52.01844, 52.7277, 
    53.43641, 54.14409, 54.85024, 55.55429, 56.25565, 56.95364, 57.64757, 
    58.33664, 59.02002, 59.6968, 60.36599, 61.02654, 61.67727, 62.31697, 
    62.94429, 63.55782, 64.15601, 64.73723, 65.29976, 65.84176, 66.36131, 
    66.85638, 67.32491, 67.76476, 68.17374, 68.54969, 68.89046, 69.19399, 
    69.45831, 69.68162, 69.86233, 69.99909, 70.09087, 70.13693, 70.13693, 
    70.09087, 69.99909, 69.86233, 69.68162, 69.45831, 69.19399, 68.89046, 
    68.54969, 68.17374, 67.76476, 67.32491, 66.85638, 66.36131, 65.84176, 
    65.29976, 64.73723, 64.15601, 63.55782, 62.94429, 62.31697, 61.67727, 
    61.02654, 60.36599, 59.6968, 59.02002, 58.33664, 57.64757, 56.95364, 
    56.25565, 55.55429, 54.85024, 54.14409, 53.43641, 52.7277, 52.01844, 
    51.30906, 50.59995, 49.89148, 49.18397, 48.47774, 47.77305, 47.07016, 
    46.36929, 45.67065, 44.97443, 44.28079, 43.58989,
  43.76653, 44.46637, 45.16932, 45.87524, 46.58398, 47.29537, 48.0092, 
    48.72528, 49.44336, 50.16318, 50.88446, 51.60688, 52.33009, 53.05371, 
    53.77734, 54.5005, 55.22271, 55.94343, 56.66205, 57.37793, 58.09037, 
    58.79859, 59.50176, 60.19897, 60.88923, 61.57146, 62.2445, 62.90707, 
    63.55782, 64.19525, 64.81778, 65.42369, 66.01116, 66.57823, 67.12283, 
    67.64278, 68.13581, 68.59956, 69.03159, 69.4295, 69.79082, 70.1132, 
    70.39439, 70.63229, 70.82504, 70.97105, 71.06911, 71.11835, 71.11835, 
    71.06911, 70.97105, 70.82504, 70.63229, 70.39439, 70.1132, 69.79082, 
    69.4295, 69.03159, 68.59956, 68.13581, 67.64278, 67.12283, 66.57823, 
    66.01116, 65.42369, 64.81778, 64.19525, 63.55782, 62.90707, 62.2445, 
    61.57146, 60.88923, 60.19897, 59.50176, 58.79859, 58.09037, 57.37793, 
    56.66205, 55.94343, 55.22271, 54.5005, 53.77734, 53.05371, 52.33009, 
    51.60688, 50.88446, 50.16318, 49.44336, 48.72528, 48.0092, 47.29537, 
    46.58398, 45.87524, 45.16932, 44.46637, 43.76653,
  43.93454, 44.64297, 45.35488, 46.07014, 46.7886, 47.51012, 48.23452, 
    48.9616, 49.69113, 50.42288, 51.15658, 51.89192, 52.62858, 53.3662, 
    54.10438, 54.84268, 55.58062, 56.31768, 57.05328, 57.78679, 58.51752, 
    59.24471, 59.96754, 60.6851, 61.39641, 62.10038, 62.79585, 63.48152, 
    64.15601, 64.81778, 65.46519, 66.09647, 66.70969, 67.30276, 67.8735, 
    68.41954, 68.9384, 69.42749, 69.88412, 70.30556, 70.68905, 71.03188, 
    71.33143, 71.58528, 71.79124, 71.94746, 72.05244, 72.10519, 72.10519, 
    72.05244, 71.94746, 71.79124, 71.58528, 71.33143, 71.03188, 70.68905, 
    70.30556, 69.88412, 69.42749, 68.9384, 68.41954, 67.8735, 67.30276, 
    66.70969, 66.09647, 65.46519, 64.81778, 64.15601, 63.48152, 62.79585, 
    62.10038, 61.39641, 60.6851, 59.96754, 59.24471, 58.51752, 57.78679, 
    57.05328, 56.31768, 55.58062, 54.84268, 54.10438, 53.3662, 52.62858, 
    51.89192, 51.15658, 50.42288, 49.69113, 48.9616, 48.23452, 47.51012, 
    46.7886, 46.07014, 45.35488, 44.64297, 43.93454,
  44.09382, 44.81047, 45.53096, 46.25516, 46.98296, 47.71421, 48.44876, 
    49.18642, 49.927, 50.67025, 51.41594, 52.16379, 52.91348, 53.66467, 
    54.41699, 55.17002, 55.9233, 56.67633, 57.42855, 58.17936, 58.92809, 
    59.67398, 60.41625, 61.154, 61.88625, 62.61193, 63.32987, 64.03877, 
    64.73723, 65.42369, 66.09647, 66.75372, 67.39344, 68.01344, 68.61138, 
    69.18474, 69.73082, 70.24678, 70.72966, 71.17637, 71.5838, 71.94884, 
    72.26848, 72.53986, 72.76041, 72.92789, 73.04058, 73.09724, 73.09724, 
    73.04058, 72.92789, 72.76041, 72.53986, 72.26848, 71.94884, 71.5838, 
    71.17637, 70.72966, 70.24678, 69.73082, 69.18474, 68.61138, 68.01344, 
    67.39344, 66.75372, 66.09647, 65.42369, 64.73723, 64.03877, 63.32987, 
    62.61193, 61.88625, 61.154, 60.41625, 59.67398, 58.92809, 58.17936, 
    57.42855, 56.67633, 55.9233, 55.17002, 54.41699, 53.66467, 52.91348, 
    52.16379, 51.41594, 50.67025, 49.927, 49.18642, 48.44876, 47.71421, 
    46.98296, 46.25516, 45.53096, 44.81047, 44.09382,
  44.24429, 44.96877, 45.69742, 46.43016, 47.16688, 47.90744, 48.6517, 
    49.39951, 50.15067, 50.90497, 51.66219, 52.42207, 53.18432, 53.94862, 
    54.71461, 55.48191, 56.25008, 57.01865, 57.78707, 58.55478, 59.32111, 
    60.08537, 60.84677, 61.60444, 62.35743, 63.10468, 63.84503, 64.57719, 
    65.29976, 66.01116, 66.70969, 67.39344, 68.06035, 68.70814, 69.33433, 
    69.93623, 70.51096, 71.0554, 71.56628, 72.04017, 72.47352, 72.86278, 
    73.20444, 73.49516, 73.73187, 73.91193, 74.03321, 74.09423, 74.09423, 
    74.03321, 73.91193, 73.73187, 73.49516, 73.20444, 72.86278, 72.47352, 
    72.04017, 71.56628, 71.0554, 70.51096, 69.93623, 69.33433, 68.70814, 
    68.06035, 67.39344, 66.70969, 66.01116, 65.29976, 64.57719, 63.84503, 
    63.10468, 62.35743, 61.60444, 60.84677, 60.08537, 59.32111, 58.55478, 
    57.78707, 57.01865, 56.25008, 55.48191, 54.71461, 53.94862, 53.18432, 
    52.42207, 51.66219, 50.90497, 50.15067, 49.39951, 48.6517, 47.90744, 
    47.16688, 46.43016, 45.69742, 44.96877, 44.24429,
  44.38583, 45.11773, 45.85415, 46.595, 47.34019, 48.08961, 48.84312, 
    49.6006, 50.36186, 51.12672, 51.89498, 52.66639, 53.44069, 54.21758, 
    54.99673, 55.77778, 56.56032, 57.34391, 58.12803, 58.91215, 59.69563, 
    60.47782, 61.25794, 62.03517, 62.80859, 63.57715, 64.33974, 65.09508, 
    65.84176, 66.57823, 67.30276, 68.01344, 68.70814, 69.38449, 70.03993, 
    70.67162, 71.27643, 71.85101, 72.39178, 72.89487, 73.35633, 73.77206, 
    74.13797, 74.45013, 74.70488, 74.89902, 75.02998, 75.09593, 75.09593, 
    75.02998, 74.89902, 74.70488, 74.45013, 74.13797, 73.77206, 73.35633, 
    72.89487, 72.39178, 71.85101, 71.27643, 70.67162, 70.03993, 69.38449, 
    68.70814, 68.01344, 67.30276, 66.57823, 65.84176, 65.09508, 64.33974, 
    63.57715, 62.80859, 62.03517, 61.25794, 60.47782, 59.69563, 58.91215, 
    58.12803, 57.34391, 56.56032, 55.77778, 54.99673, 54.21758, 53.44069, 
    52.66639, 51.89498, 51.12672, 50.36186, 49.6006, 48.84312, 48.08961, 
    47.34019, 46.595, 45.85415, 45.11773, 44.38583,
  44.51836, 45.25727, 46.00101, 46.74953, 47.50273, 48.26053, 49.02282, 
    49.78946, 50.56031, 51.33521, 52.11396, 52.89635, 53.68214, 54.47105, 
    55.2628, 56.05703, 56.85336, 57.65139, 58.45065, 59.25061, 60.05069, 
    60.85027, 61.64861, 62.44493, 63.23833, 64.02785, 64.81236, 65.59063, 
    66.36131, 67.12283, 67.8735, 68.61138, 69.33433, 70.03993, 70.72552, 
    71.38813, 72.02446, 72.6309, 73.20351, 73.73804, 74.23001, 74.67474, 
    75.06745, 75.40351, 75.67852, 75.88858, 76.03052, 76.10207, 76.10207, 
    76.03052, 75.88858, 75.67852, 75.40351, 75.06745, 74.67474, 74.23001, 
    73.73804, 73.20351, 72.6309, 72.02446, 71.38813, 70.72552, 70.03993, 
    69.33433, 68.61138, 67.8735, 67.12283, 66.36131, 65.59063, 64.81236, 
    64.02785, 63.23833, 62.44493, 61.64861, 60.85027, 60.05069, 59.25061, 
    58.45065, 57.65139, 56.85336, 56.05703, 55.2628, 54.47105, 53.68214, 
    52.89635, 52.11396, 51.33521, 50.56031, 49.78946, 49.02282, 48.26053, 
    47.50273, 46.74953, 46.00101, 45.25727, 44.51836,
  44.64181, 45.38729, 46.13791, 46.89362, 47.65435, 48.42004, 49.19058, 
    49.96586, 50.74577, 51.53014, 52.31881, 53.1116, 53.90828, 54.70861, 
    55.51231, 56.31908, 57.12857, 57.9404, 58.75413, 59.56929, 60.38533, 
    61.20166, 62.0176, 62.83242, 63.64526, 64.4552, 65.26118, 66.06201, 
    66.85638, 67.64278, 68.41954, 69.18474, 69.93623, 70.67162, 71.38813, 
    72.08273, 72.75193, 73.39191, 73.99841, 74.56674, 75.09187, 75.56844, 
    75.99091, 76.35376, 76.65166, 76.87985, 77.03436, 77.11236, 77.11236, 
    77.03436, 76.87985, 76.65166, 76.35376, 75.99091, 75.56844, 75.09187, 
    74.56674, 73.99841, 73.39191, 72.75193, 72.08273, 71.38813, 70.67162, 
    69.93623, 69.18474, 68.41954, 67.64278, 66.85638, 66.06201, 65.26118, 
    64.4552, 63.64526, 62.83242, 62.0176, 61.20166, 60.38533, 59.56929, 
    58.75413, 57.9404, 57.12857, 56.31908, 55.51231, 54.70861, 53.90828, 
    53.1116, 52.31881, 51.53014, 50.74577, 49.96586, 49.19058, 48.42004, 
    47.65435, 46.89362, 46.13791, 45.38729, 44.64181,
  44.75608, 45.50768, 46.26471, 47.02713, 47.79491, 48.56796, 49.34622, 
    50.12959, 50.91797, 51.71123, 52.50922, 53.31178, 54.1187, 54.92978, 
    55.74477, 56.56339, 57.38533, 58.21024, 59.03772, 59.86734, 60.6986, 
    61.53094, 62.36376, 63.19636, 64.02795, 64.85765, 65.68449, 66.50732, 
    67.32491, 68.13581, 68.9384, 69.73082, 70.51096, 71.27643, 72.02446, 
    72.75193, 73.45528, 74.13045, 74.77289, 75.37749, 75.93864, 76.45026, 
    76.90587, 77.2989, 77.62291, 77.87194, 78.04102, 78.1265, 78.1265, 
    78.04102, 77.87194, 77.62291, 77.2989, 76.90587, 76.45026, 75.93864, 
    75.37749, 74.77289, 74.13045, 73.45528, 72.75193, 72.02446, 71.27643, 
    70.51096, 69.73082, 68.9384, 68.13581, 67.32491, 66.50732, 65.68449, 
    64.85765, 64.02795, 63.19636, 62.36376, 61.53094, 60.6986, 59.86734, 
    59.03772, 58.21024, 57.38533, 56.56339, 55.74477, 54.92978, 54.1187, 
    53.31178, 52.50922, 51.71123, 50.91797, 50.12959, 49.34622, 48.56796, 
    47.79491, 47.02713, 46.26471, 45.50768, 44.75608,
  44.8611, 45.61835, 46.38132, 47.14996, 47.92425, 48.70414, 49.48956, 
    50.28045, 51.0767, 51.87823, 52.68489, 53.49655, 54.31304, 55.13416, 
    55.95971, 56.78943, 57.62305, 58.46024, 59.30067, 60.14393, 60.98957, 
    61.8371, 62.68594, 63.53547, 64.38497, 65.23363, 66.08053, 66.92463, 
    67.76476, 68.59956, 69.42749, 70.24678, 71.0554, 71.85101, 72.6309, 
    73.39191, 74.13045, 74.84232, 75.5227, 76.16611, 76.76637, 77.31655, 
    77.8092, 78.23647, 78.59045, 78.86371, 79.04986, 79.14419, 79.14419, 
    79.04986, 78.86371, 78.59045, 78.23647, 77.8092, 77.31655, 76.76637, 
    76.16611, 75.5227, 74.84232, 74.13045, 73.39191, 72.6309, 71.85101, 
    71.0554, 70.24678, 69.42749, 68.59956, 67.76476, 66.92463, 66.08053, 
    65.23363, 64.38497, 63.53547, 62.68594, 61.8371, 60.98957, 60.14393, 
    59.30067, 58.46024, 57.62305, 56.78943, 55.95971, 55.13416, 54.31304, 
    53.49655, 52.68489, 51.87823, 51.0767, 50.28045, 49.48956, 48.70414, 
    47.92425, 47.14996, 46.38132, 45.61835, 44.8611,
  44.9568, 45.71924, 46.48764, 47.26199, 48.04226, 48.82842, 49.62043, 
    50.41822, 51.22174, 52.03088, 52.84554, 53.6656, 54.49093, 55.32135, 
    56.15667, 56.99669, 57.84115, 58.68978, 59.54227, 60.39826, 61.25736, 
    62.11912, 62.98302, 63.84851, 64.71494, 65.58157, 66.44756, 67.31198, 
    68.17374, 69.03159, 69.88412, 70.72966, 71.56628, 72.39178, 73.20351, 
    73.99841, 74.77289, 75.5227, 76.24287, 76.9276, 77.57013, 78.16277, 
    78.69691, 79.16319, 79.55191, 79.85367, 80.06013, 80.16506, 80.16506, 
    80.06013, 79.85367, 79.55191, 79.16319, 78.69691, 78.16277, 77.57013, 
    76.9276, 76.24287, 75.5227, 74.77289, 73.99841, 73.20351, 72.39178, 
    71.56628, 70.72966, 69.88412, 69.03159, 68.17374, 67.31198, 66.44756, 
    65.58157, 64.71494, 63.84851, 62.98302, 62.11912, 61.25736, 60.39826, 
    59.54227, 58.68978, 57.84115, 56.99669, 56.15667, 55.32135, 54.49093, 
    53.6656, 52.84554, 52.03088, 51.22174, 50.41822, 49.62043, 48.82842, 
    48.04226, 47.26199, 46.48764, 45.71924, 44.9568,
  45.04311, 45.81026, 46.5836, 47.36312, 48.14882, 48.94068, 49.73867, 
    50.54276, 51.35287, 52.16895, 52.99091, 53.81864, 54.65204, 55.49096, 
    56.33524, 57.18469, 58.0391, 58.89825, 59.76184, 60.62958, 61.50111, 
    62.37604, 63.25393, 64.13426, 65.01648, 65.89993, 66.78387, 67.66744, 
    68.54969, 69.4295, 70.30556, 71.17637, 72.04017, 72.89487, 73.73804, 
    74.56674, 75.37749, 76.16611, 76.9276, 77.65593, 78.34393, 78.98316, 
    79.56378, 80.07474, 80.5041, 80.83981, 81.07088, 81.18875, 81.18875, 
    81.07088, 80.83981, 80.5041, 80.07474, 79.56378, 78.98316, 78.34393, 
    77.65593, 76.9276, 76.16611, 75.37749, 74.56674, 73.73804, 72.89487, 
    72.04017, 71.17637, 70.30556, 69.4295, 68.54969, 67.66744, 66.78387, 
    65.89993, 65.01648, 64.13426, 63.25393, 62.37604, 61.50111, 60.62958, 
    59.76184, 58.89825, 58.0391, 57.18469, 56.33524, 55.49096, 54.65204, 
    53.81864, 52.99091, 52.16895, 51.35287, 50.54276, 49.73867, 48.94068, 
    48.14882, 47.36312, 46.5836, 45.81026, 45.04311,
  45.11999, 45.89135, 46.66909, 47.45325, 48.24382, 49.04079, 49.84415, 
    50.65387, 51.46992, 52.29223, 53.12075, 53.95539, 54.79607, 55.64265, 
    56.49501, 57.35299, 58.21642, 59.08508, 59.95875, 60.83716, 61.72001, 
    62.60696, 63.49763, 64.39157, 65.2883, 66.18724, 67.08776, 67.98912, 
    68.89046, 69.79082, 70.68905, 71.5838, 72.47352, 73.35633, 74.23001, 
    75.09187, 75.93864, 76.76637, 77.57013, 78.34393, 79.08037, 79.77036, 
    80.40296, 80.96523, 81.44252, 81.81931, 82.08073, 82.21483, 82.21483, 
    82.08073, 81.81931, 81.44252, 80.96523, 80.40296, 79.77036, 79.08037, 
    78.34393, 77.57013, 76.76637, 75.93864, 75.09187, 74.23001, 73.35633, 
    72.47352, 71.5838, 70.68905, 69.79082, 68.89046, 67.98912, 67.08776, 
    66.18724, 65.2883, 64.39157, 63.49763, 62.60696, 61.72001, 60.83716, 
    59.95875, 59.08508, 58.21642, 57.35299, 56.49501, 55.64265, 54.79607, 
    53.95539, 53.12075, 52.29223, 51.46992, 50.65387, 49.84415, 49.04079, 
    48.24382, 47.45325, 46.66909, 45.89135, 45.11999,
  45.18737, 45.96243, 46.74407, 47.53231, 48.32716, 49.12864, 49.93674, 
    50.75143, 51.57272, 52.40054, 53.23486, 54.07561, 54.92273, 55.7761, 
    56.63563, 57.50119, 58.37262, 59.24976, 60.13241, 61.02035, 61.91332, 
    62.81103, 63.71317, 64.61935, 65.52915, 66.44211, 67.35767, 68.2752, 
    69.19399, 70.1132, 71.03188, 71.94884, 72.86278, 73.77206, 74.67474, 
    75.56844, 76.45026, 77.31655, 78.16277, 78.98316, 79.77036, 80.51504, 
    81.20532, 81.82646, 82.3607, 82.78796, 83.08778, 83.24277, 83.24277, 
    83.08778, 82.78796, 82.3607, 81.82646, 81.20532, 80.51504, 79.77036, 
    78.98316, 78.16277, 77.31655, 76.45026, 75.56844, 74.67474, 73.77206, 
    72.86278, 71.94884, 71.03188, 70.1132, 69.19399, 68.2752, 67.35767, 
    66.44211, 65.52915, 64.61935, 63.71317, 62.81103, 61.91332, 61.02035, 
    60.13241, 59.24976, 58.37262, 57.50119, 56.63563, 55.7761, 54.92273, 
    54.07561, 53.23486, 52.40054, 51.57272, 50.75143, 49.93674, 49.12864, 
    48.32716, 47.53231, 46.74407, 45.96243, 45.18737,
  45.24522, 46.02346, 46.80845, 47.6002, 48.39876, 49.20412, 50.01631, 
    50.83531, 51.66111, 52.4937, 53.33304, 54.17908, 55.03177, 55.89104, 
    56.75679, 57.62892, 58.50731, 59.39183, 60.2823, 61.17855, 62.08035, 
    62.98748, 63.89967, 64.81659, 65.73791, 66.66322, 67.59209, 68.52398, 
    69.45831, 70.39439, 71.33143, 72.26848, 73.20444, 74.13797, 75.06745, 
    75.99091, 76.90587, 77.8092, 78.69691, 79.56378, 80.40296, 81.20532, 
    81.95869, 82.6469, 83.249, 83.73922, 84.08896, 84.27195, 84.27195, 
    84.08896, 83.73922, 83.249, 82.6469, 81.95869, 81.20532, 80.40296, 
    79.56378, 78.69691, 77.8092, 76.90587, 75.99091, 75.06745, 74.13797, 
    73.20444, 72.26848, 71.33143, 70.39439, 69.45831, 68.52398, 67.59209, 
    66.66322, 65.73791, 64.81659, 63.89967, 62.98748, 62.08035, 61.17855, 
    60.2823, 59.39183, 58.50731, 57.62892, 56.75679, 55.89104, 55.03177, 
    54.17908, 53.33304, 52.4937, 51.66111, 50.83531, 50.01631, 49.20412, 
    48.39876, 47.6002, 46.80845, 46.02346, 45.24522,
  45.29348, 46.07439, 46.86219, 47.65689, 48.45854, 49.26716, 50.08277, 
    50.90538, 51.73498, 52.57156, 53.41512, 54.26561, 55.12299, 55.9872, 
    56.85819, 57.73586, 58.62013, 59.51086, 60.40795, 61.31122, 62.22052, 
    63.13563, 64.05634, 64.98241, 65.91354, 66.84942, 67.78967, 68.7339, 
    69.68162, 70.63229, 71.58528, 72.53986, 73.49516, 74.45013, 75.40351, 
    76.35376, 77.2989, 78.23647, 79.16319, 80.07474, 80.96523, 81.82646, 
    82.6469, 83.41006, 84.09252, 84.66222, 85.079, 85.30138, 85.30138, 
    85.079, 84.66222, 84.09252, 83.41006, 82.6469, 81.82646, 80.96523, 
    80.07474, 79.16319, 78.23647, 77.2989, 76.35376, 75.40351, 74.45013, 
    73.49516, 72.53986, 71.58528, 70.63229, 69.68162, 68.7339, 67.78967, 
    66.84942, 65.91354, 64.98241, 64.05634, 63.13563, 62.22052, 61.31122, 
    60.40795, 59.51086, 58.62013, 57.73586, 56.85819, 55.9872, 55.12299, 
    54.26561, 53.41512, 52.57156, 51.73498, 50.90538, 50.08277, 49.26716, 
    48.45854, 47.65689, 46.86219, 46.07439, 45.29348,
  45.33213, 46.11519, 46.90523, 47.7023, 48.50644, 49.31768, 50.13604, 
    50.96155, 51.7942, 52.63401, 53.48095, 54.33502, 55.19618, 56.06439, 
    56.93961, 57.82175, 58.71076, 59.60653, 60.50896, 61.41792, 62.33329, 
    63.25488, 64.18253, 65.11604, 66.05517, 66.99967, 67.94925, 68.90359, 
    69.86233, 70.82504, 71.79124, 72.76041, 73.73187, 74.70488, 75.67852, 
    76.65166, 77.62291, 78.59045, 79.55191, 80.5041, 81.44252, 82.3607, 
    83.249, 84.09252, 84.8678, 85.53786, 86.04778, 86.32938, 86.32938, 
    86.04778, 85.53786, 84.8678, 84.09252, 83.249, 82.3607, 81.44252, 
    80.5041, 79.55191, 78.59045, 77.62291, 76.65166, 75.67852, 74.70488, 
    73.73187, 72.76041, 71.79124, 70.82504, 69.86233, 68.90359, 67.94925, 
    66.99967, 66.05517, 65.11604, 64.18253, 63.25488, 62.33329, 61.41792, 
    60.50896, 59.60653, 58.71076, 57.82175, 56.93961, 56.06439, 55.19618, 
    54.33502, 53.48095, 52.63401, 51.7942, 50.96155, 50.13604, 49.31768, 
    48.50644, 47.7023, 46.90523, 46.11519, 45.33213,
  45.36115, 46.14581, 46.93755, 47.7364, 48.54241, 49.35562, 50.17606, 
    51.00375, 51.8387, 52.68093, 53.53043, 54.3872, 55.25121, 56.12244, 
    57.00084, 57.88636, 58.77895, 59.67853, 60.58501, 61.49828, 62.41824, 
    63.34475, 64.27767, 65.21684, 66.16206, 67.11313, 68.06983, 69.03191, 
    69.99909, 70.97105, 71.94746, 72.92789, 73.91193, 74.89902, 75.88858, 
    76.87985, 77.87194, 78.86371, 79.85367, 80.83981, 81.81931, 82.78796, 
    83.73922, 84.66222, 85.53786, 86.33054, 86.97294, 87.35221, 87.35221, 
    86.97294, 86.33054, 85.53786, 84.66222, 83.73922, 82.78796, 81.81931, 
    80.83981, 79.85367, 78.86371, 77.87194, 76.87985, 75.88858, 74.89902, 
    73.91193, 72.92789, 71.94746, 70.97105, 69.99909, 69.03191, 68.06983, 
    67.11313, 66.16206, 65.21684, 64.27767, 63.34475, 62.41824, 61.49828, 
    60.58501, 59.67853, 58.77895, 57.88636, 57.00084, 56.12244, 55.25121, 
    54.3872, 53.53043, 52.68093, 51.8387, 51.00375, 50.17606, 49.35562, 
    48.54241, 47.7364, 46.93755, 46.14581, 45.36115,
  45.3805, 46.16624, 46.95911, 47.75915, 48.56641, 49.38094, 50.20276, 
    51.03191, 51.8684, 52.71225, 53.56347, 54.42204, 55.28796, 56.1612, 
    57.04174, 57.92953, 58.82452, 59.72665, 60.63584, 61.55201, 62.47506, 
    63.40488, 64.34134, 65.28431, 66.23363, 67.18914, 68.15065, 69.11797, 
    70.09087, 71.06911, 72.05244, 73.04058, 74.03321, 75.02998, 76.03052, 
    77.03436, 78.04102, 79.04986, 80.06013, 81.07088, 82.08073, 83.08778, 
    84.08896, 85.079, 86.04778, 86.97294, 87.79688, 88.35755, 88.35755, 
    87.79688, 86.97294, 86.04778, 85.079, 84.08896, 83.08778, 82.08073, 
    81.07088, 80.06013, 79.04986, 78.04102, 77.03436, 76.03052, 75.02998, 
    74.03321, 73.04058, 72.05244, 71.06911, 70.09087, 69.11797, 68.15065, 
    67.18914, 66.23363, 65.28431, 64.34134, 63.40488, 62.47506, 61.55201, 
    60.63584, 59.72665, 58.82452, 57.92953, 57.04174, 56.1612, 55.28796, 
    54.42204, 53.56347, 52.71225, 51.8684, 51.03191, 50.20276, 49.38094, 
    48.56641, 47.75915, 46.95911, 46.16624, 45.3805,
  45.39018, 46.17646, 46.96989, 47.77053, 48.57842, 49.3936, 50.21612, 
    51.046, 51.88326, 52.72793, 53.58, 54.43948, 55.30635, 56.18061, 
    57.06222, 57.95115, 58.84734, 59.75075, 60.6613, 61.57893, 62.50353, 
    63.43501, 64.37325, 65.31813, 66.26952, 67.22726, 68.19119, 69.16115, 
    70.13693, 71.11835, 72.10519, 73.09724, 74.09423, 75.09593, 76.10207, 
    77.11236, 78.1265, 79.14419, 80.16506, 81.18875, 82.21483, 83.24277, 
    84.27195, 85.30138, 86.32938, 87.35221, 88.35755, 89.26539, 89.26539, 
    88.35755, 87.35221, 86.32938, 85.30138, 84.27195, 83.24277, 82.21483, 
    81.18875, 80.16506, 79.14419, 78.1265, 77.11236, 76.10207, 75.09593, 
    74.09423, 73.09724, 72.10519, 71.11835, 70.13693, 69.16115, 68.19119, 
    67.22726, 66.26952, 65.31813, 64.37325, 63.43501, 62.50353, 61.57893, 
    60.6613, 59.75075, 58.84734, 57.95115, 57.06222, 56.18061, 55.30635, 
    54.43948, 53.58, 52.72793, 51.88326, 51.046, 50.21612, 49.3936, 48.57842, 
    47.77053, 46.96989, 46.17646, 45.39018,
  45.39018, 46.17646, 46.96989, 47.77053, 48.57842, 49.3936, 50.21612, 
    51.046, 51.88326, 52.72793, 53.58, 54.43948, 55.30635, 56.18061, 
    57.06222, 57.95115, 58.84734, 59.75075, 60.6613, 61.57893, 62.50353, 
    63.43501, 64.37325, 65.31813, 66.26952, 67.22726, 68.19119, 69.16115, 
    70.13693, 71.11835, 72.10519, 73.09724, 74.09423, 75.09593, 76.10207, 
    77.11236, 78.1265, 79.14419, 80.16506, 81.18875, 82.21483, 83.24277, 
    84.27195, 85.30138, 86.32938, 87.35221, 88.35755, 89.26539, 89.26539, 
    88.35755, 87.35221, 86.32938, 85.30138, 84.27195, 83.24277, 82.21483, 
    81.18875, 80.16506, 79.14419, 78.1265, 77.11236, 76.10207, 75.09593, 
    74.09423, 73.09724, 72.10519, 71.11835, 70.13693, 69.16115, 68.19119, 
    67.22726, 66.26952, 65.31813, 64.37325, 63.43501, 62.50353, 61.57893, 
    60.6613, 59.75075, 58.84734, 57.95115, 57.06222, 56.18061, 55.30635, 
    54.43948, 53.58, 52.72793, 51.88326, 51.046, 50.21612, 49.3936, 48.57842, 
    47.77053, 46.96989, 46.17646, 45.39018,
  45.3805, 46.16624, 46.95911, 47.75915, 48.56641, 49.38094, 50.20276, 
    51.03191, 51.8684, 52.71225, 53.56347, 54.42204, 55.28796, 56.1612, 
    57.04174, 57.92953, 58.82452, 59.72665, 60.63584, 61.55201, 62.47506, 
    63.40488, 64.34134, 65.28431, 66.23363, 67.18914, 68.15065, 69.11797, 
    70.09087, 71.06911, 72.05244, 73.04058, 74.03321, 75.02998, 76.03052, 
    77.03436, 78.04102, 79.04986, 80.06013, 81.07088, 82.08073, 83.08778, 
    84.08896, 85.079, 86.04778, 86.97294, 87.79688, 88.35755, 88.35755, 
    87.79688, 86.97294, 86.04778, 85.079, 84.08896, 83.08778, 82.08073, 
    81.07088, 80.06013, 79.04986, 78.04102, 77.03436, 76.03052, 75.02998, 
    74.03321, 73.04058, 72.05244, 71.06911, 70.09087, 69.11797, 68.15065, 
    67.18914, 66.23363, 65.28431, 64.34134, 63.40488, 62.47506, 61.55201, 
    60.63584, 59.72665, 58.82452, 57.92953, 57.04174, 56.1612, 55.28796, 
    54.42204, 53.56347, 52.71225, 51.8684, 51.03191, 50.20276, 49.38094, 
    48.56641, 47.75915, 46.95911, 46.16624, 45.3805,
  45.36115, 46.14581, 46.93755, 47.7364, 48.54241, 49.35562, 50.17606, 
    51.00375, 51.8387, 52.68093, 53.53043, 54.3872, 55.25121, 56.12244, 
    57.00084, 57.88636, 58.77895, 59.67853, 60.58501, 61.49828, 62.41824, 
    63.34475, 64.27767, 65.21684, 66.16206, 67.11313, 68.06983, 69.03191, 
    69.99909, 70.97105, 71.94746, 72.92789, 73.91193, 74.89902, 75.88858, 
    76.87985, 77.87194, 78.86371, 79.85367, 80.83981, 81.81931, 82.78796, 
    83.73922, 84.66222, 85.53786, 86.33054, 86.97294, 87.35221, 87.35221, 
    86.97294, 86.33054, 85.53786, 84.66222, 83.73922, 82.78796, 81.81931, 
    80.83981, 79.85367, 78.86371, 77.87194, 76.87985, 75.88858, 74.89902, 
    73.91193, 72.92789, 71.94746, 70.97105, 69.99909, 69.03191, 68.06983, 
    67.11313, 66.16206, 65.21684, 64.27767, 63.34475, 62.41824, 61.49828, 
    60.58501, 59.67853, 58.77895, 57.88636, 57.00084, 56.12244, 55.25121, 
    54.3872, 53.53043, 52.68093, 51.8387, 51.00375, 50.17606, 49.35562, 
    48.54241, 47.7364, 46.93755, 46.14581, 45.36115,
  45.33213, 46.11519, 46.90523, 47.7023, 48.50644, 49.31768, 50.13604, 
    50.96155, 51.7942, 52.63401, 53.48095, 54.33502, 55.19618, 56.06439, 
    56.93961, 57.82175, 58.71076, 59.60653, 60.50896, 61.41792, 62.33329, 
    63.25488, 64.18253, 65.11604, 66.05517, 66.99967, 67.94925, 68.90359, 
    69.86233, 70.82504, 71.79124, 72.76041, 73.73187, 74.70488, 75.67852, 
    76.65166, 77.62291, 78.59045, 79.55191, 80.5041, 81.44252, 82.3607, 
    83.249, 84.09252, 84.8678, 85.53786, 86.04778, 86.32938, 86.32938, 
    86.04778, 85.53786, 84.8678, 84.09252, 83.249, 82.3607, 81.44252, 
    80.5041, 79.55191, 78.59045, 77.62291, 76.65166, 75.67852, 74.70488, 
    73.73187, 72.76041, 71.79124, 70.82504, 69.86233, 68.90359, 67.94925, 
    66.99967, 66.05517, 65.11604, 64.18253, 63.25488, 62.33329, 61.41792, 
    60.50896, 59.60653, 58.71076, 57.82175, 56.93961, 56.06439, 55.19618, 
    54.33502, 53.48095, 52.63401, 51.7942, 50.96155, 50.13604, 49.31768, 
    48.50644, 47.7023, 46.90523, 46.11519, 45.33213,
  45.29348, 46.07439, 46.86219, 47.65689, 48.45854, 49.26716, 50.08277, 
    50.90538, 51.73498, 52.57156, 53.41512, 54.26561, 55.12299, 55.9872, 
    56.85819, 57.73586, 58.62013, 59.51086, 60.40795, 61.31122, 62.22052, 
    63.13563, 64.05634, 64.98241, 65.91354, 66.84942, 67.78967, 68.7339, 
    69.68162, 70.63229, 71.58528, 72.53986, 73.49516, 74.45013, 75.40351, 
    76.35376, 77.2989, 78.23647, 79.16319, 80.07474, 80.96523, 81.82646, 
    82.6469, 83.41006, 84.09252, 84.66222, 85.079, 85.30138, 85.30138, 
    85.079, 84.66222, 84.09252, 83.41006, 82.6469, 81.82646, 80.96523, 
    80.07474, 79.16319, 78.23647, 77.2989, 76.35376, 75.40351, 74.45013, 
    73.49516, 72.53986, 71.58528, 70.63229, 69.68162, 68.7339, 67.78967, 
    66.84942, 65.91354, 64.98241, 64.05634, 63.13563, 62.22052, 61.31122, 
    60.40795, 59.51086, 58.62013, 57.73586, 56.85819, 55.9872, 55.12299, 
    54.26561, 53.41512, 52.57156, 51.73498, 50.90538, 50.08277, 49.26716, 
    48.45854, 47.65689, 46.86219, 46.07439, 45.29348,
  45.24522, 46.02346, 46.80845, 47.6002, 48.39876, 49.20412, 50.01631, 
    50.83531, 51.66111, 52.4937, 53.33304, 54.17908, 55.03177, 55.89104, 
    56.75679, 57.62892, 58.50731, 59.39183, 60.2823, 61.17855, 62.08035, 
    62.98748, 63.89967, 64.81659, 65.73791, 66.66322, 67.59209, 68.52398, 
    69.45831, 70.39439, 71.33143, 72.26848, 73.20444, 74.13797, 75.06745, 
    75.99091, 76.90587, 77.8092, 78.69691, 79.56378, 80.40296, 81.20532, 
    81.95869, 82.6469, 83.249, 83.73922, 84.08896, 84.27195, 84.27195, 
    84.08896, 83.73922, 83.249, 82.6469, 81.95869, 81.20532, 80.40296, 
    79.56378, 78.69691, 77.8092, 76.90587, 75.99091, 75.06745, 74.13797, 
    73.20444, 72.26848, 71.33143, 70.39439, 69.45831, 68.52398, 67.59209, 
    66.66322, 65.73791, 64.81659, 63.89967, 62.98748, 62.08035, 61.17855, 
    60.2823, 59.39183, 58.50731, 57.62892, 56.75679, 55.89104, 55.03177, 
    54.17908, 53.33304, 52.4937, 51.66111, 50.83531, 50.01631, 49.20412, 
    48.39876, 47.6002, 46.80845, 46.02346, 45.24522,
  45.18737, 45.96243, 46.74407, 47.53231, 48.32716, 49.12864, 49.93674, 
    50.75143, 51.57272, 52.40054, 53.23486, 54.07561, 54.92273, 55.7761, 
    56.63563, 57.50119, 58.37262, 59.24976, 60.13241, 61.02035, 61.91332, 
    62.81103, 63.71317, 64.61935, 65.52915, 66.44211, 67.35767, 68.2752, 
    69.19399, 70.1132, 71.03188, 71.94884, 72.86278, 73.77206, 74.67474, 
    75.56844, 76.45026, 77.31655, 78.16277, 78.98316, 79.77036, 80.51504, 
    81.20532, 81.82646, 82.3607, 82.78796, 83.08778, 83.24277, 83.24277, 
    83.08778, 82.78796, 82.3607, 81.82646, 81.20532, 80.51504, 79.77036, 
    78.98316, 78.16277, 77.31655, 76.45026, 75.56844, 74.67474, 73.77206, 
    72.86278, 71.94884, 71.03188, 70.1132, 69.19399, 68.2752, 67.35767, 
    66.44211, 65.52915, 64.61935, 63.71317, 62.81103, 61.91332, 61.02035, 
    60.13241, 59.24976, 58.37262, 57.50119, 56.63563, 55.7761, 54.92273, 
    54.07561, 53.23486, 52.40054, 51.57272, 50.75143, 49.93674, 49.12864, 
    48.32716, 47.53231, 46.74407, 45.96243, 45.18737,
  45.11999, 45.89135, 46.66909, 47.45325, 48.24382, 49.04079, 49.84415, 
    50.65387, 51.46992, 52.29223, 53.12075, 53.95539, 54.79607, 55.64265, 
    56.49501, 57.35299, 58.21642, 59.08508, 59.95875, 60.83716, 61.72001, 
    62.60696, 63.49763, 64.39157, 65.2883, 66.18724, 67.08776, 67.98912, 
    68.89046, 69.79082, 70.68905, 71.5838, 72.47352, 73.35633, 74.23001, 
    75.09187, 75.93864, 76.76637, 77.57013, 78.34393, 79.08037, 79.77036, 
    80.40296, 80.96523, 81.44252, 81.81931, 82.08073, 82.21483, 82.21483, 
    82.08073, 81.81931, 81.44252, 80.96523, 80.40296, 79.77036, 79.08037, 
    78.34393, 77.57013, 76.76637, 75.93864, 75.09187, 74.23001, 73.35633, 
    72.47352, 71.5838, 70.68905, 69.79082, 68.89046, 67.98912, 67.08776, 
    66.18724, 65.2883, 64.39157, 63.49763, 62.60696, 61.72001, 60.83716, 
    59.95875, 59.08508, 58.21642, 57.35299, 56.49501, 55.64265, 54.79607, 
    53.95539, 53.12075, 52.29223, 51.46992, 50.65387, 49.84415, 49.04079, 
    48.24382, 47.45325, 46.66909, 45.89135, 45.11999,
  45.04311, 45.81026, 46.5836, 47.36312, 48.14882, 48.94068, 49.73867, 
    50.54276, 51.35287, 52.16895, 52.99091, 53.81864, 54.65204, 55.49096, 
    56.33524, 57.18469, 58.0391, 58.89825, 59.76184, 60.62958, 61.50111, 
    62.37604, 63.25393, 64.13426, 65.01648, 65.89993, 66.78387, 67.66744, 
    68.54969, 69.4295, 70.30556, 71.17637, 72.04017, 72.89487, 73.73804, 
    74.56674, 75.37749, 76.16611, 76.9276, 77.65593, 78.34393, 78.98316, 
    79.56378, 80.07474, 80.5041, 80.83981, 81.07088, 81.18875, 81.18875, 
    81.07088, 80.83981, 80.5041, 80.07474, 79.56378, 78.98316, 78.34393, 
    77.65593, 76.9276, 76.16611, 75.37749, 74.56674, 73.73804, 72.89487, 
    72.04017, 71.17637, 70.30556, 69.4295, 68.54969, 67.66744, 66.78387, 
    65.89993, 65.01648, 64.13426, 63.25393, 62.37604, 61.50111, 60.62958, 
    59.76184, 58.89825, 58.0391, 57.18469, 56.33524, 55.49096, 54.65204, 
    53.81864, 52.99091, 52.16895, 51.35287, 50.54276, 49.73867, 48.94068, 
    48.14882, 47.36312, 46.5836, 45.81026, 45.04311,
  44.9568, 45.71924, 46.48764, 47.26199, 48.04226, 48.82842, 49.62043, 
    50.41822, 51.22174, 52.03088, 52.84554, 53.6656, 54.49093, 55.32135, 
    56.15667, 56.99669, 57.84115, 58.68978, 59.54227, 60.39826, 61.25736, 
    62.11912, 62.98302, 63.84851, 64.71494, 65.58157, 66.44756, 67.31198, 
    68.17374, 69.03159, 69.88412, 70.72966, 71.56628, 72.39178, 73.20351, 
    73.99841, 74.77289, 75.5227, 76.24287, 76.9276, 77.57013, 78.16277, 
    78.69691, 79.16319, 79.55191, 79.85367, 80.06013, 80.16506, 80.16506, 
    80.06013, 79.85367, 79.55191, 79.16319, 78.69691, 78.16277, 77.57013, 
    76.9276, 76.24287, 75.5227, 74.77289, 73.99841, 73.20351, 72.39178, 
    71.56628, 70.72966, 69.88412, 69.03159, 68.17374, 67.31198, 66.44756, 
    65.58157, 64.71494, 63.84851, 62.98302, 62.11912, 61.25736, 60.39826, 
    59.54227, 58.68978, 57.84115, 56.99669, 56.15667, 55.32135, 54.49093, 
    53.6656, 52.84554, 52.03088, 51.22174, 50.41822, 49.62043, 48.82842, 
    48.04226, 47.26199, 46.48764, 45.71924, 44.9568,
  44.8611, 45.61835, 46.38132, 47.14996, 47.92425, 48.70414, 49.48956, 
    50.28045, 51.0767, 51.87823, 52.68489, 53.49655, 54.31304, 55.13416, 
    55.95971, 56.78943, 57.62305, 58.46024, 59.30067, 60.14393, 60.98957, 
    61.8371, 62.68594, 63.53547, 64.38497, 65.23363, 66.08053, 66.92463, 
    67.76476, 68.59956, 69.42749, 70.24678, 71.0554, 71.85101, 72.6309, 
    73.39191, 74.13045, 74.84232, 75.5227, 76.16611, 76.76637, 77.31655, 
    77.8092, 78.23647, 78.59045, 78.86371, 79.04986, 79.14419, 79.14419, 
    79.04986, 78.86371, 78.59045, 78.23647, 77.8092, 77.31655, 76.76637, 
    76.16611, 75.5227, 74.84232, 74.13045, 73.39191, 72.6309, 71.85101, 
    71.0554, 70.24678, 69.42749, 68.59956, 67.76476, 66.92463, 66.08053, 
    65.23363, 64.38497, 63.53547, 62.68594, 61.8371, 60.98957, 60.14393, 
    59.30067, 58.46024, 57.62305, 56.78943, 55.95971, 55.13416, 54.31304, 
    53.49655, 52.68489, 51.87823, 51.0767, 50.28045, 49.48956, 48.70414, 
    47.92425, 47.14996, 46.38132, 45.61835, 44.8611,
  44.75608, 45.50768, 46.26471, 47.02713, 47.79491, 48.56796, 49.34622, 
    50.12959, 50.91797, 51.71123, 52.50922, 53.31178, 54.1187, 54.92978, 
    55.74477, 56.56339, 57.38533, 58.21024, 59.03772, 59.86734, 60.6986, 
    61.53094, 62.36376, 63.19636, 64.02795, 64.85765, 65.68449, 66.50732, 
    67.32491, 68.13581, 68.9384, 69.73082, 70.51096, 71.27643, 72.02446, 
    72.75193, 73.45528, 74.13045, 74.77289, 75.37749, 75.93864, 76.45026, 
    76.90587, 77.2989, 77.62291, 77.87194, 78.04102, 78.1265, 78.1265, 
    78.04102, 77.87194, 77.62291, 77.2989, 76.90587, 76.45026, 75.93864, 
    75.37749, 74.77289, 74.13045, 73.45528, 72.75193, 72.02446, 71.27643, 
    70.51096, 69.73082, 68.9384, 68.13581, 67.32491, 66.50732, 65.68449, 
    64.85765, 64.02795, 63.19636, 62.36376, 61.53094, 60.6986, 59.86734, 
    59.03772, 58.21024, 57.38533, 56.56339, 55.74477, 54.92978, 54.1187, 
    53.31178, 52.50922, 51.71123, 50.91797, 50.12959, 49.34622, 48.56796, 
    47.79491, 47.02713, 46.26471, 45.50768, 44.75608,
  44.64181, 45.38729, 46.13791, 46.89362, 47.65435, 48.42004, 49.19058, 
    49.96586, 50.74577, 51.53014, 52.31881, 53.1116, 53.90828, 54.70861, 
    55.51231, 56.31908, 57.12857, 57.9404, 58.75413, 59.56929, 60.38533, 
    61.20166, 62.0176, 62.83242, 63.64526, 64.4552, 65.26118, 66.06201, 
    66.85638, 67.64278, 68.41954, 69.18474, 69.93623, 70.67162, 71.38813, 
    72.08273, 72.75193, 73.39191, 73.99841, 74.56674, 75.09187, 75.56844, 
    75.99091, 76.35376, 76.65166, 76.87985, 77.03436, 77.11236, 77.11236, 
    77.03436, 76.87985, 76.65166, 76.35376, 75.99091, 75.56844, 75.09187, 
    74.56674, 73.99841, 73.39191, 72.75193, 72.08273, 71.38813, 70.67162, 
    69.93623, 69.18474, 68.41954, 67.64278, 66.85638, 66.06201, 65.26118, 
    64.4552, 63.64526, 62.83242, 62.0176, 61.20166, 60.38533, 59.56929, 
    58.75413, 57.9404, 57.12857, 56.31908, 55.51231, 54.70861, 53.90828, 
    53.1116, 52.31881, 51.53014, 50.74577, 49.96586, 49.19058, 48.42004, 
    47.65435, 46.89362, 46.13791, 45.38729, 44.64181,
  44.51836, 45.25727, 46.00101, 46.74953, 47.50273, 48.26053, 49.02282, 
    49.78946, 50.56031, 51.33521, 52.11396, 52.89635, 53.68214, 54.47105, 
    55.2628, 56.05703, 56.85336, 57.65139, 58.45065, 59.25061, 60.05069, 
    60.85027, 61.64861, 62.44493, 63.23833, 64.02785, 64.81236, 65.59063, 
    66.36131, 67.12283, 67.8735, 68.61138, 69.33433, 70.03993, 70.72552, 
    71.38813, 72.02446, 72.6309, 73.20351, 73.73804, 74.23001, 74.67474, 
    75.06745, 75.40351, 75.67852, 75.88858, 76.03052, 76.10207, 76.10207, 
    76.03052, 75.88858, 75.67852, 75.40351, 75.06745, 74.67474, 74.23001, 
    73.73804, 73.20351, 72.6309, 72.02446, 71.38813, 70.72552, 70.03993, 
    69.33433, 68.61138, 67.8735, 67.12283, 66.36131, 65.59063, 64.81236, 
    64.02785, 63.23833, 62.44493, 61.64861, 60.85027, 60.05069, 59.25061, 
    58.45065, 57.65139, 56.85336, 56.05703, 55.2628, 54.47105, 53.68214, 
    52.89635, 52.11396, 51.33521, 50.56031, 49.78946, 49.02282, 48.26053, 
    47.50273, 46.74953, 46.00101, 45.25727, 44.51836,
  44.38583, 45.11773, 45.85415, 46.595, 47.34019, 48.08961, 48.84312, 
    49.6006, 50.36186, 51.12672, 51.89498, 52.66639, 53.44069, 54.21758, 
    54.99673, 55.77778, 56.56032, 57.34391, 58.12803, 58.91215, 59.69563, 
    60.47782, 61.25794, 62.03517, 62.80859, 63.57715, 64.33974, 65.09508, 
    65.84176, 66.57823, 67.30276, 68.01344, 68.70814, 69.38449, 70.03993, 
    70.67162, 71.27643, 71.85101, 72.39178, 72.89487, 73.35633, 73.77206, 
    74.13797, 74.45013, 74.70488, 74.89902, 75.02998, 75.09593, 75.09593, 
    75.02998, 74.89902, 74.70488, 74.45013, 74.13797, 73.77206, 73.35633, 
    72.89487, 72.39178, 71.85101, 71.27643, 70.67162, 70.03993, 69.38449, 
    68.70814, 68.01344, 67.30276, 66.57823, 65.84176, 65.09508, 64.33974, 
    63.57715, 62.80859, 62.03517, 61.25794, 60.47782, 59.69563, 58.91215, 
    58.12803, 57.34391, 56.56032, 55.77778, 54.99673, 54.21758, 53.44069, 
    52.66639, 51.89498, 51.12672, 50.36186, 49.6006, 48.84312, 48.08961, 
    47.34019, 46.595, 45.85415, 45.11773, 44.38583,
  44.24429, 44.96877, 45.69742, 46.43016, 47.16688, 47.90744, 48.6517, 
    49.39951, 50.15067, 50.90497, 51.66219, 52.42207, 53.18432, 53.94862, 
    54.71461, 55.48191, 56.25008, 57.01865, 57.78707, 58.55478, 59.32111, 
    60.08537, 60.84677, 61.60444, 62.35743, 63.10468, 63.84503, 64.57719, 
    65.29976, 66.01116, 66.70969, 67.39344, 68.06035, 68.70814, 69.33433, 
    69.93623, 70.51096, 71.0554, 71.56628, 72.04017, 72.47352, 72.86278, 
    73.20444, 73.49516, 73.73187, 73.91193, 74.03321, 74.09423, 74.09423, 
    74.03321, 73.91193, 73.73187, 73.49516, 73.20444, 72.86278, 72.47352, 
    72.04017, 71.56628, 71.0554, 70.51096, 69.93623, 69.33433, 68.70814, 
    68.06035, 67.39344, 66.70969, 66.01116, 65.29976, 64.57719, 63.84503, 
    63.10468, 62.35743, 61.60444, 60.84677, 60.08537, 59.32111, 58.55478, 
    57.78707, 57.01865, 56.25008, 55.48191, 54.71461, 53.94862, 53.18432, 
    52.42207, 51.66219, 50.90497, 50.15067, 49.39951, 48.6517, 47.90744, 
    47.16688, 46.43016, 45.69742, 44.96877, 44.24429,
  44.09382, 44.81047, 45.53096, 46.25516, 46.98296, 47.71421, 48.44876, 
    49.18642, 49.927, 50.67025, 51.41594, 52.16379, 52.91348, 53.66467, 
    54.41699, 55.17002, 55.9233, 56.67633, 57.42855, 58.17936, 58.92809, 
    59.67398, 60.41625, 61.154, 61.88625, 62.61193, 63.32987, 64.03877, 
    64.73723, 65.42369, 66.09647, 66.75372, 67.39344, 68.01344, 68.61138, 
    69.18474, 69.73082, 70.24678, 70.72966, 71.17637, 71.5838, 71.94884, 
    72.26848, 72.53986, 72.76041, 72.92789, 73.04058, 73.09724, 73.09724, 
    73.04058, 72.92789, 72.76041, 72.53986, 72.26848, 71.94884, 71.5838, 
    71.17637, 70.72966, 70.24678, 69.73082, 69.18474, 68.61138, 68.01344, 
    67.39344, 66.75372, 66.09647, 65.42369, 64.73723, 64.03877, 63.32987, 
    62.61193, 61.88625, 61.154, 60.41625, 59.67398, 58.92809, 58.17936, 
    57.42855, 56.67633, 55.9233, 55.17002, 54.41699, 53.66467, 52.91348, 
    52.16379, 51.41594, 50.67025, 49.927, 49.18642, 48.44876, 47.71421, 
    46.98296, 46.25516, 45.53096, 44.81047, 44.09382,
  43.93454, 44.64297, 45.35488, 46.07014, 46.7886, 47.51012, 48.23452, 
    48.9616, 49.69113, 50.42288, 51.15658, 51.89192, 52.62858, 53.3662, 
    54.10438, 54.84268, 55.58062, 56.31768, 57.05328, 57.78679, 58.51752, 
    59.24471, 59.96754, 60.6851, 61.39641, 62.10038, 62.79585, 63.48152, 
    64.15601, 64.81778, 65.46519, 66.09647, 66.70969, 67.30276, 67.8735, 
    68.41954, 68.9384, 69.42749, 69.88412, 70.30556, 70.68905, 71.03188, 
    71.33143, 71.58528, 71.79124, 71.94746, 72.05244, 72.10519, 72.10519, 
    72.05244, 71.94746, 71.79124, 71.58528, 71.33143, 71.03188, 70.68905, 
    70.30556, 69.88412, 69.42749, 68.9384, 68.41954, 67.8735, 67.30276, 
    66.70969, 66.09647, 65.46519, 64.81778, 64.15601, 63.48152, 62.79585, 
    62.10038, 61.39641, 60.6851, 59.96754, 59.24471, 58.51752, 57.78679, 
    57.05328, 56.31768, 55.58062, 54.84268, 54.10438, 53.3662, 52.62858, 
    51.89192, 51.15658, 50.42288, 49.69113, 48.9616, 48.23452, 47.51012, 
    46.7886, 46.07014, 45.35488, 44.64297, 43.93454,
  43.76653, 44.46637, 45.16932, 45.87524, 46.58398, 47.29537, 48.0092, 
    48.72528, 49.44336, 50.16318, 50.88446, 51.60688, 52.33009, 53.05371, 
    53.77734, 54.5005, 55.22271, 55.94343, 56.66205, 57.37793, 58.09037, 
    58.79859, 59.50176, 60.19897, 60.88923, 61.57146, 62.2445, 62.90707, 
    63.55782, 64.19525, 64.81778, 65.42369, 66.01116, 66.57823, 67.12283, 
    67.64278, 68.13581, 68.59956, 69.03159, 69.4295, 69.79082, 70.1132, 
    70.39439, 70.63229, 70.82504, 70.97105, 71.06911, 71.11835, 71.11835, 
    71.06911, 70.97105, 70.82504, 70.63229, 70.39439, 70.1132, 69.79082, 
    69.4295, 69.03159, 68.59956, 68.13581, 67.64278, 67.12283, 66.57823, 
    66.01116, 65.42369, 64.81778, 64.19525, 63.55782, 62.90707, 62.2445, 
    61.57146, 60.88923, 60.19897, 59.50176, 58.79859, 58.09037, 57.37793, 
    56.66205, 55.94343, 55.22271, 54.5005, 53.77734, 53.05371, 52.33009, 
    51.60688, 50.88446, 50.16318, 49.44336, 48.72528, 48.0092, 47.29537, 
    46.58398, 45.87524, 45.16932, 44.46637, 43.76653,
  43.58989, 44.28079, 44.97443, 45.67065, 46.36929, 47.07016, 47.77305, 
    48.47774, 49.18397, 49.89148, 50.59995, 51.30906, 52.01844, 52.7277, 
    53.43641, 54.14409, 54.85024, 55.55429, 56.25565, 56.95364, 57.64757, 
    58.33664, 59.02002, 59.6968, 60.36599, 61.02654, 61.67727, 62.31697, 
    62.94429, 63.55782, 64.15601, 64.73723, 65.29976, 65.84176, 66.36131, 
    66.85638, 67.32491, 67.76476, 68.17374, 68.54969, 68.89046, 69.19399, 
    69.45831, 69.68162, 69.86233, 69.99909, 70.09087, 70.13693, 70.13693, 
    70.09087, 69.99909, 69.86233, 69.68162, 69.45831, 69.19399, 68.89046, 
    68.54969, 68.17374, 67.76476, 67.32491, 66.85638, 66.36131, 65.84176, 
    65.29976, 64.73723, 64.15601, 63.55782, 62.94429, 62.31697, 61.67727, 
    61.02654, 60.36599, 59.6968, 59.02002, 58.33664, 57.64757, 56.95364, 
    56.25565, 55.55429, 54.85024, 54.14409, 53.43641, 52.7277, 52.01844, 
    51.30906, 50.59995, 49.89148, 49.18397, 48.47774, 47.77305, 47.07016, 
    46.36929, 45.67065, 44.97443, 44.28079, 43.58989,
  43.40474, 44.08636, 44.77034, 45.45651, 46.14469, 46.83469, 47.52629, 
    48.21923, 48.91327, 49.6081, 50.30342, 50.99888, 51.6941, 52.38867, 
    53.08215, 53.77406, 54.46386, 55.15101, 55.83487, 56.51479, 57.19004, 
    57.85986, 58.52339, 59.17973, 59.82792, 60.4669, 61.09555, 61.71267, 
    62.31697, 62.90707, 63.48152, 64.03877, 64.57719, 65.09508, 65.59063, 
    66.06201, 66.50732, 66.92463, 67.31198, 67.66744, 67.98912, 68.2752, 
    68.52398, 68.7339, 68.90359, 69.03191, 69.11797, 69.16115, 69.16115, 
    69.11797, 69.03191, 68.90359, 68.7339, 68.52398, 68.2752, 67.98912, 
    67.66744, 67.31198, 66.92463, 66.50732, 66.06201, 65.59063, 65.09508, 
    64.57719, 64.03877, 63.48152, 62.90707, 62.31697, 61.71267, 61.09555, 
    60.4669, 59.82792, 59.17973, 58.52339, 57.85986, 57.19004, 56.51479, 
    55.83487, 55.15101, 54.46386, 53.77406, 53.08215, 52.38867, 51.6941, 
    50.99888, 50.30342, 49.6081, 48.91327, 48.21923, 47.52629, 46.83469, 
    46.14469, 45.45651, 44.77034, 44.08636, 43.40474,
  43.21118, 43.8832, 44.55719, 45.23299, 45.91039, 46.5892, 47.26916, 
    47.95004, 48.63155, 49.3134, 49.99525, 50.67675, 51.35751, 52.03711, 
    52.7151, 53.39099, 54.06424, 54.73428, 55.40049, 56.06221, 56.7187, 
    57.36921, 58.01291, 58.64888, 59.2762, 59.89382, 60.50066, 61.09555, 
    61.67727, 62.2445, 62.79585, 63.32987, 63.84503, 64.33974, 64.81236, 
    65.26118, 65.68449, 66.08053, 66.44756, 66.78387, 67.08776, 67.35767, 
    67.59209, 67.78967, 67.94925, 68.06983, 68.15065, 68.19119, 68.19119, 
    68.15065, 68.06983, 67.94925, 67.78967, 67.59209, 67.35767, 67.08776, 
    66.78387, 66.44756, 66.08053, 65.68449, 65.26118, 64.81236, 64.33974, 
    63.84503, 63.32987, 62.79585, 62.2445, 61.67727, 61.09555, 60.50066, 
    59.89382, 59.2762, 58.64888, 58.01291, 57.36921, 56.7187, 56.06221, 
    55.40049, 54.73428, 54.06424, 53.39099, 52.7151, 52.03711, 51.35751, 
    50.67675, 49.99525, 49.3134, 48.63155, 47.95004, 47.26916, 46.5892, 
    45.91039, 45.23299, 44.55719, 43.8832, 43.21118,
  43.00933, 43.67144, 44.33515, 45.00027, 45.66659, 46.33389, 47.00192, 
    47.67044, 48.33913, 49.00771, 49.67582, 50.34309, 51.00915, 51.67355, 
    52.33583, 52.9955, 53.65202, 54.30482, 54.95327, 55.59671, 56.23442, 
    56.86565, 57.48957, 58.1053, 58.71193, 59.30845, 59.89382, 60.4669, 
    61.02654, 61.57146, 62.10038, 62.61193, 63.10468, 63.57715, 64.02785, 
    64.4552, 64.85765, 65.23363, 65.58157, 65.89993, 66.18724, 66.44211, 
    66.66322, 66.84942, 66.99967, 67.11313, 67.18914, 67.22726, 67.22726, 
    67.18914, 67.11313, 66.99967, 66.84942, 66.66322, 66.44211, 66.18724, 
    65.89993, 65.58157, 65.23363, 64.85765, 64.4552, 64.02785, 63.57715, 
    63.10468, 62.61193, 62.10038, 61.57146, 61.02654, 60.4669, 59.89382, 
    59.30845, 58.71193, 58.1053, 57.48957, 56.86565, 56.23442, 55.59671, 
    54.95327, 54.30482, 53.65202, 52.9955, 52.33583, 51.67355, 51.00915, 
    50.34309, 49.67582, 49.00771, 48.33913, 47.67044, 47.00192, 46.33389, 
    45.66659, 45.00027, 44.33515, 43.67144, 43.00933,
  42.7993, 43.45123, 44.10437, 44.75852, 45.41347, 46.06899, 46.72482, 
    47.3807, 48.03632, 48.69137, 49.3455, 49.99833, 50.64946, 51.29846, 
    51.94487, 52.58817, 53.22784, 53.8633, 54.49394, 55.11909, 55.73805, 
    56.35006, 56.95434, 57.55002, 58.1362, 58.71193, 59.2762, 59.82792, 
    60.36599, 60.88923, 61.39641, 61.88625, 62.35743, 62.80859, 63.23833, 
    63.64526, 64.02795, 64.38497, 64.71494, 65.01648, 65.2883, 65.52915, 
    65.73791, 65.91354, 66.05517, 66.16206, 66.23363, 66.26952, 66.26952, 
    66.23363, 66.16206, 66.05517, 65.91354, 65.73791, 65.52915, 65.2883, 
    65.01648, 64.71494, 64.38497, 64.02795, 63.64526, 63.23833, 62.80859, 
    62.35743, 61.88625, 61.39641, 60.88923, 60.36599, 59.82792, 59.2762, 
    58.71193, 58.1362, 57.55002, 56.95434, 56.35006, 55.73805, 55.11909, 
    54.49394, 53.8633, 53.22784, 52.58817, 51.94487, 51.29846, 50.64946, 
    49.99833, 49.3455, 48.69137, 48.03632, 47.3807, 46.72482, 46.06899, 
    45.41347, 44.75852, 44.10437, 43.45123, 42.7993,
  42.58122, 43.22269, 43.86499, 44.50792, 45.15124, 45.79473, 46.43811, 
    47.08112, 47.72343, 48.36473, 49.00467, 49.64286, 50.2789, 50.91235, 
    51.54275, 52.16959, 52.79234, 53.41042, 54.02324, 54.63013, 55.2304, 
    55.82333, 56.40814, 56.98399, 57.55002, 58.1053, 58.64888, 59.17973, 
    59.6968, 60.19897, 60.6851, 61.154, 61.60444, 62.03517, 62.44493, 
    62.83242, 63.19636, 63.53547, 63.84851, 64.13426, 64.39157, 64.61935, 
    64.81659, 64.98241, 65.11604, 65.21684, 65.28431, 65.31813, 65.31813, 
    65.28431, 65.21684, 65.11604, 64.98241, 64.81659, 64.61935, 64.39157, 
    64.13426, 63.84851, 63.53547, 63.19636, 62.83242, 62.44493, 62.03517, 
    61.60444, 61.154, 60.6851, 60.19897, 59.6968, 59.17973, 58.64888, 
    58.1053, 57.55002, 56.98399, 56.40814, 55.82333, 55.2304, 54.63013, 
    54.02324, 53.41042, 52.79234, 52.16959, 51.54275, 50.91235, 50.2789, 
    49.64286, 49.00467, 48.36473, 47.72343, 47.08112, 46.43811, 45.79473, 
    45.15124, 44.50792, 43.86499, 43.22269, 42.58122,
  42.35519, 42.98596, 43.61718, 44.24864, 44.88011, 45.51133, 46.14204, 
    46.77196, 47.40077, 48.02814, 48.65372, 49.27712, 49.89793, 50.51572, 
    51.13002, 51.74033, 52.34612, 52.94683, 53.54185, 54.13057, 54.71228, 
    55.28629, 55.85184, 56.40814, 56.95434, 57.48957, 58.01291, 58.52339, 
    59.02002, 59.50176, 59.96754, 60.41625, 60.84677, 61.25794, 61.64861, 
    62.0176, 62.36376, 62.68594, 62.98302, 63.25393, 63.49763, 63.71317, 
    63.89967, 64.05634, 64.18253, 64.27767, 64.34134, 64.37325, 64.37325, 
    64.34134, 64.27767, 64.18253, 64.05634, 63.89967, 63.71317, 63.49763, 
    63.25393, 62.98302, 62.68594, 62.36376, 62.0176, 61.64861, 61.25794, 
    60.84677, 60.41625, 59.96754, 59.50176, 59.02002, 58.52339, 58.01291, 
    57.48957, 56.95434, 56.40814, 55.85184, 55.28629, 54.71228, 54.13057, 
    53.54185, 52.94683, 52.34612, 51.74033, 51.13002, 50.51572, 49.89793, 
    49.27712, 48.65372, 48.02814, 47.40077, 46.77196, 46.14204, 45.51133, 
    44.88011, 44.24864, 43.61718, 42.98596, 42.35519,
  42.12135, 42.74119, 43.36111, 43.98088, 44.60027, 45.21903, 45.83688, 
    46.45353, 47.06866, 47.68195, 48.29302, 48.9015, 49.50698, 50.10903, 
    50.70718, 51.30094, 51.88978, 52.47316, 53.05048, 53.62113, 54.18444, 
    54.73974, 55.28629, 55.82333, 56.35006, 56.86565, 57.36921, 57.85986, 
    58.33664, 58.79859, 59.24471, 59.67398, 60.08537, 60.47782, 60.85027, 
    61.20166, 61.53094, 61.8371, 62.11912, 62.37604, 62.60696, 62.81103, 
    62.98748, 63.13563, 63.25488, 63.34475, 63.40488, 63.43501, 63.43501, 
    63.40488, 63.34475, 63.25488, 63.13563, 62.98748, 62.81103, 62.60696, 
    62.37604, 62.11912, 61.8371, 61.53094, 61.20166, 60.85027, 60.47782, 
    60.08537, 59.67398, 59.24471, 58.79859, 58.33664, 57.85986, 57.36921, 
    56.86565, 56.35006, 55.82333, 55.28629, 54.73974, 54.18444, 53.62113, 
    53.05048, 52.47316, 51.88978, 51.30094, 50.70718, 50.10903, 49.50698, 
    48.9015, 48.29302, 47.68195, 47.06866, 46.45353, 45.83688, 45.21903, 
    44.60027, 43.98088, 43.36111, 42.74119, 42.12135,
  41.87982, 42.48852, 43.09693, 43.70482, 44.31195, 44.91806, 45.52287, 
    46.12609, 46.72741, 47.32647, 47.92294, 48.51642, 49.10651, 49.69277, 
    50.27475, 50.85197, 51.42391, 51.99004, 52.54977, 53.10251, 53.64762, 
    54.18444, 54.71228, 55.2304, 55.73805, 56.23442, 56.7187, 57.19004, 
    57.64757, 58.09037, 58.51752, 58.92809, 59.32111, 59.69563, 60.05069, 
    60.38533, 60.6986, 60.98957, 61.25736, 61.50111, 61.72001, 61.91332, 
    62.08035, 62.22052, 62.33329, 62.41824, 62.47506, 62.50353, 62.50353, 
    62.47506, 62.41824, 62.33329, 62.22052, 62.08035, 61.91332, 61.72001, 
    61.50111, 61.25736, 60.98957, 60.6986, 60.38533, 60.05069, 59.69563, 
    59.32111, 58.92809, 58.51752, 58.09037, 57.64757, 57.19004, 56.7187, 
    56.23442, 55.73805, 55.2304, 54.71228, 54.18444, 53.64762, 53.10251, 
    52.54977, 51.99004, 51.42391, 50.85197, 50.27475, 49.69277, 49.10651, 
    48.51642, 47.92294, 47.32647, 46.72741, 46.12609, 45.52287, 44.91806, 
    44.31195, 43.70482, 43.09693, 42.48852, 41.87982,
  41.63073, 42.2281, 42.82481, 43.42064, 44.01534, 44.60864, 45.20028, 
    45.78994, 46.37732, 46.96207, 47.54385, 48.12227, 48.69693, 49.2674, 
    49.83323, 50.39396, 50.94908, 51.49806, 52.04035, 52.57537, 53.10251, 
    53.62113, 54.13057, 54.63013, 55.11909, 55.59671, 56.06221, 56.51479, 
    56.95364, 57.37793, 57.78679, 58.17936, 58.55478, 58.91215, 59.25061, 
    59.56929, 59.86734, 60.14393, 60.39826, 60.62958, 60.83716, 61.02035, 
    61.17855, 61.31122, 61.41792, 61.49828, 61.55201, 61.57893, 61.57893, 
    61.55201, 61.49828, 61.41792, 61.31122, 61.17855, 61.02035, 60.83716, 
    60.62958, 60.39826, 60.14393, 59.86734, 59.56929, 59.25061, 58.91215, 
    58.55478, 58.17936, 57.78679, 57.37793, 56.95364, 56.51479, 56.06221, 
    55.59671, 55.11909, 54.63013, 54.13057, 53.62113, 53.10251, 52.57537, 
    52.04035, 51.49806, 50.94908, 50.39396, 49.83323, 49.2674, 48.69693, 
    48.12227, 47.54385, 46.96207, 46.37732, 45.78994, 45.20028, 44.60864, 
    44.01534, 43.42064, 42.82481, 42.2281, 41.63073,
  41.37419, 41.96006, 42.54491, 43.12852, 43.71065, 44.29101, 44.86935, 
    45.44535, 46.0187, 46.58908, 47.15612, 47.71944, 48.27867, 48.83337, 
    49.3831, 49.92742, 50.46582, 50.9978, 51.52283, 52.04035, 52.54977, 
    53.05048, 53.54185, 54.02324, 54.49394, 54.95327, 55.40049, 55.83487, 
    56.25565, 56.66205, 57.05328, 57.42855, 57.78707, 58.12803, 58.45065, 
    58.75413, 59.03772, 59.30067, 59.54227, 59.76184, 59.95875, 60.13241, 
    60.2823, 60.40795, 60.50896, 60.58501, 60.63584, 60.6613, 60.6613, 
    60.63584, 60.58501, 60.50896, 60.40795, 60.2823, 60.13241, 59.95875, 
    59.76184, 59.54227, 59.30067, 59.03772, 58.75413, 58.45065, 58.12803, 
    57.78707, 57.42855, 57.05328, 56.66205, 56.25565, 55.83487, 55.40049, 
    54.95327, 54.49394, 54.02324, 53.54185, 53.05048, 52.54977, 52.04035, 
    51.52283, 50.9978, 50.46582, 49.92742, 49.3831, 48.83337, 48.27867, 
    47.71944, 47.15612, 46.58908, 46.0187, 45.44535, 44.86935, 44.29101, 
    43.71065, 43.12852, 42.54491, 41.96006, 41.37419,
  41.11036, 41.68456, 42.2574, 42.82867, 43.39809, 43.9654, 44.53034, 
    45.0926, 45.65187, 46.20782, 46.76009, 47.30833, 47.85214, 48.39112, 
    48.92484, 49.45285, 49.97467, 50.48983, 50.9978, 51.49806, 51.99004, 
    52.47316, 52.94683, 53.41042, 53.8633, 54.30482, 54.73428, 55.15101, 
    55.55429, 55.94343, 56.31768, 56.67633, 57.01865, 57.34391, 57.65139, 
    57.9404, 58.21024, 58.46024, 58.68978, 58.89825, 59.08508, 59.24976, 
    59.39183, 59.51086, 59.60653, 59.67853, 59.72665, 59.75075, 59.75075, 
    59.72665, 59.67853, 59.60653, 59.51086, 59.39183, 59.24976, 59.08508, 
    58.89825, 58.68978, 58.46024, 58.21024, 57.9404, 57.65139, 57.34391, 
    57.01865, 56.67633, 56.31768, 55.94343, 55.55429, 55.15101, 54.73428, 
    54.30482, 53.8633, 53.41042, 52.94683, 52.47316, 51.99004, 51.49806, 
    50.9978, 50.48983, 49.97467, 49.45285, 48.92484, 48.39112, 47.85214, 
    47.30833, 46.76009, 46.20782, 45.65187, 45.0926, 44.53034, 43.9654, 
    43.39809, 42.82867, 42.2574, 41.68456, 41.11036,
  40.83934, 41.40174, 41.96246, 42.52125, 43.07787, 43.63205, 44.18351, 
    44.73198, 45.27712, 45.81862, 46.35614, 46.88931, 47.41776, 47.94109, 
    48.45889, 48.97073, 49.47615, 49.97467, 50.46582, 50.94908, 51.42391, 
    51.88978, 52.34612, 52.79234, 53.22784, 53.65202, 54.06424, 54.46386, 
    54.85024, 55.22271, 55.58062, 55.9233, 56.25008, 56.56032, 56.85336, 
    57.12857, 57.38533, 57.62305, 57.84115, 58.0391, 58.21642, 58.37262, 
    58.50731, 58.62013, 58.71076, 58.77895, 58.82452, 58.84734, 58.84734, 
    58.82452, 58.77895, 58.71076, 58.62013, 58.50731, 58.37262, 58.21642, 
    58.0391, 57.84115, 57.62305, 57.38533, 57.12857, 56.85336, 56.56032, 
    56.25008, 55.9233, 55.58062, 55.22271, 54.85024, 54.46386, 54.06424, 
    53.65202, 53.22784, 52.79234, 52.34612, 51.88978, 51.42391, 50.94908, 
    50.46582, 49.97467, 49.47615, 48.97073, 48.45889, 47.94109, 47.41776, 
    46.88931, 46.35614, 45.81862, 45.27712, 44.73198, 44.18351, 43.63205, 
    43.07787, 42.52125, 41.96246, 41.40174, 40.83934,
  40.56128, 41.11176, 41.66023, 42.20646, 42.75019, 43.29116, 43.82911, 
    44.36374, 44.89474, 45.4218, 45.94459, 46.46275, 46.97591, 47.4837, 
    47.98571, 48.48154, 48.97073, 49.45285, 49.92742, 50.39396, 50.85197, 
    51.30094, 51.74033, 52.16959, 52.58817, 52.9955, 53.39099, 53.77406, 
    54.14409, 54.5005, 54.84268, 55.17002, 55.48191, 55.77778, 56.05703, 
    56.31908, 56.56339, 56.78943, 56.99669, 57.18469, 57.35299, 57.50119, 
    57.62892, 57.73586, 57.82175, 57.88636, 57.92953, 57.95115, 57.95115, 
    57.92953, 57.88636, 57.82175, 57.73586, 57.62892, 57.50119, 57.35299, 
    57.18469, 56.99669, 56.78943, 56.56339, 56.31908, 56.05703, 55.77778, 
    55.48191, 55.17002, 54.84268, 54.5005, 54.14409, 53.77406, 53.39099, 
    52.9955, 52.58817, 52.16959, 51.74033, 51.30094, 50.85197, 50.39396, 
    49.92742, 49.45285, 48.97073, 48.48154, 47.98571, 47.4837, 46.97591, 
    46.46275, 45.94459, 45.4218, 44.89474, 44.36374, 43.82911, 43.29116, 
    42.75019, 42.20646, 41.66023, 41.11176, 40.56128,
  40.27629, 40.81476, 41.35089, 41.88448, 42.41526, 42.94299, 43.46738, 
    43.98816, 44.50503, 45.01768, 45.52579, 46.029, 46.52699, 47.01936, 
    47.50573, 47.98571, 48.45889, 48.92484, 49.3831, 49.83323, 50.27475, 
    50.70718, 51.13002, 51.54275, 51.94487, 52.33583, 52.7151, 53.08215, 
    53.43641, 53.77734, 54.10438, 54.41699, 54.71461, 54.99673, 55.2628, 
    55.51231, 55.74477, 55.95971, 56.15667, 56.33524, 56.49501, 56.63563, 
    56.75679, 56.85819, 56.93961, 57.00084, 57.04174, 57.06222, 57.06222, 
    57.04174, 57.00084, 56.93961, 56.85819, 56.75679, 56.63563, 56.49501, 
    56.33524, 56.15667, 55.95971, 55.74477, 55.51231, 55.2628, 54.99673, 
    54.71461, 54.41699, 54.10438, 53.77734, 53.43641, 53.08215, 52.7151, 
    52.33583, 51.94487, 51.54275, 51.13002, 50.70718, 50.27475, 49.83323, 
    49.3831, 48.92484, 48.45889, 47.98571, 47.50573, 47.01936, 46.52699, 
    46.029, 45.52579, 45.01768, 44.50503, 43.98816, 43.46738, 42.94299, 
    42.41526, 41.88448, 41.35089, 40.81476, 40.27629,
  39.98453, 40.51088, 41.03462, 41.5555, 42.07329, 42.58773, 43.09856, 
    43.60551, 44.10828, 44.60656, 45.10006, 45.58843, 46.07135, 46.54844, 
    47.01936, 47.4837, 47.94109, 48.39112, 48.83337, 49.2674, 49.69277, 
    50.10903, 50.51572, 50.91235, 51.29846, 51.67355, 52.03711, 52.38867, 
    52.7277, 53.05371, 53.3662, 53.66467, 53.94862, 54.21758, 54.47105, 
    54.70861, 54.92978, 55.13416, 55.32135, 55.49096, 55.64265, 55.7761, 
    55.89104, 55.9872, 56.06439, 56.12244, 56.1612, 56.18061, 56.18061, 
    56.1612, 56.12244, 56.06439, 55.9872, 55.89104, 55.7761, 55.64265, 
    55.49096, 55.32135, 55.13416, 54.92978, 54.70861, 54.47105, 54.21758, 
    53.94862, 53.66467, 53.3662, 53.05371, 52.7277, 52.38867, 52.03711, 
    51.67355, 51.29846, 50.91235, 50.51572, 50.10903, 49.69277, 49.2674, 
    48.83337, 48.39112, 47.94109, 47.4837, 47.01936, 46.54844, 46.07135, 
    45.58843, 45.10006, 44.60656, 44.10828, 43.60551, 43.09856, 42.58773, 
    42.07329, 41.5555, 41.03462, 40.51088, 39.98453,
  39.68611, 40.20029, 40.71156, 41.2197, 41.72447, 42.22562, 42.7229, 
    43.21604, 43.70475, 44.18875, 44.66773, 45.14137, 45.60936, 46.07135, 
    46.52699, 46.97591, 47.41776, 47.85214, 48.27867, 48.69693, 49.10651, 
    49.50698, 49.89793, 50.2789, 50.64946, 51.00915, 51.35751, 51.6941, 
    52.01844, 52.33009, 52.62858, 52.91348, 53.18432, 53.44069, 53.68214, 
    53.90828, 54.1187, 54.31304, 54.49093, 54.65204, 54.79607, 54.92273, 
    55.03177, 55.12299, 55.19618, 55.25121, 55.28796, 55.30635, 55.30635, 
    55.28796, 55.25121, 55.19618, 55.12299, 55.03177, 54.92273, 54.79607, 
    54.65204, 54.49093, 54.31304, 54.1187, 53.90828, 53.68214, 53.44069, 
    53.18432, 52.91348, 52.62858, 52.33009, 52.01844, 51.6941, 51.35751, 
    51.00915, 50.64946, 50.2789, 49.89793, 49.50698, 49.10651, 48.69693, 
    48.27867, 47.85214, 47.41776, 46.97591, 46.52699, 46.07135, 45.60936, 
    45.14137, 44.66773, 44.18875, 43.70475, 43.21604, 42.7229, 42.22562, 
    41.72447, 41.2197, 40.71156, 40.20029, 39.68611,
  39.38117, 39.88312, 40.38189, 40.87727, 41.36901, 41.85689, 42.34064, 
    42.82002, 43.29474, 43.76454, 44.22911, 44.68816, 45.14137, 45.58843, 
    46.029, 46.46275, 46.88931, 47.30833, 47.71944, 48.12227, 48.51642, 
    48.9015, 49.27712, 49.64286, 49.99833, 50.34309, 50.67675, 50.99888, 
    51.30906, 51.60688, 51.89192, 52.16379, 52.42207, 52.66639, 52.89635, 
    53.1116, 53.31178, 53.49655, 53.6656, 53.81864, 53.95539, 54.07561, 
    54.17908, 54.26561, 54.33502, 54.3872, 54.42204, 54.43948, 54.43948, 
    54.42204, 54.3872, 54.33502, 54.26561, 54.17908, 54.07561, 53.95539, 
    53.81864, 53.6656, 53.49655, 53.31178, 53.1116, 52.89635, 52.66639, 
    52.42207, 52.16379, 51.89192, 51.60688, 51.30906, 50.99888, 50.67675, 
    50.34309, 49.99833, 49.64286, 49.27712, 48.9015, 48.51642, 48.12227, 
    47.71944, 47.30833, 46.88931, 46.46275, 46.029, 45.58843, 45.14137, 
    44.68816, 44.22911, 43.76454, 43.29474, 42.82002, 42.34064, 41.85689, 
    41.36901, 40.87727, 40.38189, 39.88312, 39.38117,
  39.06984, 39.55952, 40.04577, 40.52837, 41.00711, 41.48173, 41.95201, 
    42.41769, 42.87851, 43.33421, 43.7845, 44.22911, 44.66773, 45.10006, 
    45.52579, 45.94459, 46.35614, 46.76009, 47.15612, 47.54385, 47.92294, 
    48.29302, 48.65372, 49.00467, 49.3455, 49.67582, 49.99525, 50.30342, 
    50.59995, 50.88446, 51.15658, 51.41594, 51.66219, 51.89498, 52.11396, 
    52.31881, 52.50922, 52.68489, 52.84554, 52.99091, 53.12075, 53.23486, 
    53.33304, 53.41512, 53.48095, 53.53043, 53.56347, 53.58, 53.58, 53.56347, 
    53.53043, 53.48095, 53.41512, 53.33304, 53.23486, 53.12075, 52.99091, 
    52.84554, 52.68489, 52.50922, 52.31881, 52.11396, 51.89498, 51.66219, 
    51.41594, 51.15658, 50.88446, 50.59995, 50.30342, 49.99525, 49.67582, 
    49.3455, 49.00467, 48.65372, 48.29302, 47.92294, 47.54385, 47.15612, 
    46.76009, 46.35614, 45.94459, 45.52579, 45.10006, 44.66773, 44.22911, 
    43.7845, 43.33421, 42.87851, 42.41769, 41.95201, 41.48173, 41.00711, 
    40.52837, 40.04577, 39.55952, 39.06984,
  38.75225, 39.22964, 39.70337, 40.17321, 40.63895, 41.10036, 41.55723, 
    42.0093, 42.45632, 42.89805, 43.33421, 43.76454, 44.18875, 44.60656, 
    45.01768, 45.4218, 45.81862, 46.20782, 46.58908, 46.96207, 47.32647, 
    47.68195, 48.02814, 48.36473, 48.69137, 49.00771, 49.3134, 49.6081, 
    49.89148, 50.16318, 50.42288, 50.67025, 50.90497, 51.12672, 51.33521, 
    51.53014, 51.71123, 51.87823, 52.03088, 52.16895, 52.29223, 52.40054, 
    52.4937, 52.57156, 52.63401, 52.68093, 52.71225, 52.72793, 52.72793, 
    52.71225, 52.68093, 52.63401, 52.57156, 52.4937, 52.40054, 52.29223, 
    52.16895, 52.03088, 51.87823, 51.71123, 51.53014, 51.33521, 51.12672, 
    50.90497, 50.67025, 50.42288, 50.16318, 49.89148, 49.6081, 49.3134, 
    49.00771, 48.69137, 48.36473, 48.02814, 47.68195, 47.32647, 46.96207, 
    46.58908, 46.20782, 45.81862, 45.4218, 45.01768, 44.60656, 44.18875, 
    43.76454, 43.33421, 42.89805, 42.45632, 42.0093, 41.55723, 41.10036, 
    40.63895, 40.17321, 39.70337, 39.22964, 38.75225,
  38.42853, 38.89363, 39.35483, 39.81194, 40.26473, 40.71301, 41.15653, 
    41.59509, 42.02843, 42.45632, 42.87851, 43.29474, 43.70475, 44.10828, 
    44.50503, 44.89474, 45.27712, 45.65187, 46.0187, 46.37732, 46.72741, 
    47.06866, 47.40077, 47.72343, 48.03632, 48.33913, 48.63155, 48.91327, 
    49.18397, 49.44336, 49.69113, 49.927, 50.15067, 50.36186, 50.56031, 
    50.74577, 50.91797, 51.0767, 51.22174, 51.35287, 51.46992, 51.57272, 
    51.66111, 51.73498, 51.7942, 51.8387, 51.8684, 51.88326, 51.88326, 
    51.8684, 51.8387, 51.7942, 51.73498, 51.66111, 51.57272, 51.46992, 
    51.35287, 51.22174, 51.0767, 50.91797, 50.74577, 50.56031, 50.36186, 
    50.15067, 49.927, 49.69113, 49.44336, 49.18397, 48.91327, 48.63155, 
    48.33913, 48.03632, 47.72343, 47.40077, 47.06866, 46.72741, 46.37732, 
    46.0187, 45.65187, 45.27712, 44.89474, 44.50503, 44.10828, 43.70475, 
    43.29474, 42.87851, 42.45632, 42.02843, 41.59509, 41.15653, 40.71301, 
    40.26473, 39.81194, 39.35483, 38.89363, 38.42853,
  38.09881, 38.55162, 39.00033, 39.44474, 39.88465, 40.31985, 40.75014, 
    41.17529, 41.59509, 42.0093, 42.41769, 42.82002, 43.21604, 43.60551, 
    43.98816, 44.36374, 44.73198, 45.0926, 45.44535, 45.78994, 46.12609, 
    46.45353, 46.77196, 47.08112, 47.3807, 47.67044, 47.95004, 48.21923, 
    48.47774, 48.72528, 48.9616, 49.18642, 49.39951, 49.6006, 49.78946, 
    49.96586, 50.12959, 50.28045, 50.41822, 50.54276, 50.65387, 50.75143, 
    50.83531, 50.90538, 50.96155, 51.00375, 51.03191, 51.046, 51.046, 
    51.03191, 51.00375, 50.96155, 50.90538, 50.83531, 50.75143, 50.65387, 
    50.54276, 50.41822, 50.28045, 50.12959, 49.96586, 49.78946, 49.6006, 
    49.39951, 49.18642, 48.9616, 48.72528, 48.47774, 48.21923, 47.95004, 
    47.67044, 47.3807, 47.08112, 46.77196, 46.45353, 46.12609, 45.78994, 
    45.44535, 45.0926, 44.73198, 44.36374, 43.98816, 43.60551, 43.21604, 
    42.82002, 42.41769, 42.0093, 41.59509, 41.17529, 40.75014, 40.31985, 
    39.88465, 39.44474, 39.00033, 38.55162, 38.09881,
  37.76321, 38.20377, 38.64002, 39.07178, 39.49888, 39.9211, 40.33826, 
    40.75014, 41.15653, 41.55723, 41.95201, 42.34064, 42.7229, 43.09856, 
    43.46738, 43.82911, 44.18351, 44.53034, 44.86935, 45.20028, 45.52287, 
    45.83688, 46.14204, 46.43811, 46.72482, 47.00192, 47.26916, 47.52629, 
    47.77305, 48.0092, 48.23452, 48.44876, 48.6517, 48.84312, 49.02282, 
    49.19058, 49.34622, 49.48956, 49.62043, 49.73867, 49.84415, 49.93674, 
    50.01631, 50.08277, 50.13604, 50.17606, 50.20276, 50.21612, 50.21612, 
    50.20276, 50.17606, 50.13604, 50.08277, 50.01631, 49.93674, 49.84415, 
    49.73867, 49.62043, 49.48956, 49.34622, 49.19058, 49.02282, 48.84312, 
    48.6517, 48.44876, 48.23452, 48.0092, 47.77305, 47.52629, 47.26916, 
    47.00192, 46.72482, 46.43811, 46.14204, 45.83688, 45.52287, 45.20028, 
    44.86935, 44.53034, 44.18351, 43.82911, 43.46738, 43.09856, 42.7229, 
    42.34064, 41.95201, 41.55723, 41.15653, 40.75014, 40.33826, 39.9211, 
    39.49888, 39.07178, 38.64002, 38.20377, 37.76321,
  37.42188, 37.8502, 38.27405, 38.69325, 39.10761, 39.51696, 39.9211, 
    40.31985, 40.71301, 41.10036, 41.48173, 41.85689, 42.22562, 42.58773, 
    42.94299, 43.29116, 43.63205, 43.9654, 44.29101, 44.60864, 44.91806, 
    45.21903, 45.51133, 45.79473, 46.06899, 46.33389, 46.5892, 46.83469, 
    47.07016, 47.29537, 47.51012, 47.71421, 47.90744, 48.08961, 48.26053, 
    48.42004, 48.56796, 48.70414, 48.82842, 48.94068, 49.04079, 49.12864, 
    49.20412, 49.26716, 49.31768, 49.35562, 49.38094, 49.3936, 49.3936, 
    49.38094, 49.35562, 49.31768, 49.26716, 49.20412, 49.12864, 49.04079, 
    48.94068, 48.82842, 48.70414, 48.56796, 48.42004, 48.26053, 48.08961, 
    47.90744, 47.71421, 47.51012, 47.29537, 47.07016, 46.83469, 46.5892, 
    46.33389, 46.06899, 45.79473, 45.51133, 45.21903, 44.91806, 44.60864, 
    44.29101, 43.9654, 43.63205, 43.29116, 42.94299, 42.58773, 42.22562, 
    41.85689, 41.48173, 41.10036, 40.71301, 40.31985, 39.9211, 39.51696, 
    39.10761, 38.69325, 38.27405, 37.8502, 37.42188,
  37.07492, 37.49107, 37.90258, 38.30929, 38.71102, 39.10761, 39.49888, 
    39.88465, 40.26473, 40.63895, 41.00711, 41.36901, 41.72447, 42.07329, 
    42.41526, 42.75019, 43.07787, 43.39809, 43.71065, 44.01534, 44.31195, 
    44.60027, 44.88011, 45.15124, 45.41347, 45.66659, 45.91039, 46.14469, 
    46.36929, 46.58398, 46.7886, 46.98296, 47.16688, 47.34019, 47.50273, 
    47.65435, 47.79491, 47.92425, 48.04226, 48.14882, 48.24382, 48.32716, 
    48.39876, 48.45854, 48.50644, 48.54241, 48.56641, 48.57842, 48.57842, 
    48.56641, 48.54241, 48.50644, 48.45854, 48.39876, 48.32716, 48.24382, 
    48.14882, 48.04226, 47.92425, 47.79491, 47.65435, 47.50273, 47.34019, 
    47.16688, 46.98296, 46.7886, 46.58398, 46.36929, 46.14469, 45.91039, 
    45.66659, 45.41347, 45.15124, 44.88011, 44.60027, 44.31195, 44.01534, 
    43.71065, 43.39809, 43.07787, 42.75019, 42.41526, 42.07329, 41.72447, 
    41.36901, 41.00711, 40.63895, 40.26473, 39.88465, 39.49888, 39.10761, 
    38.71102, 38.30929, 37.90258, 37.49107, 37.07492,
  36.72248, 37.12651, 37.52576, 37.92007, 38.30929, 38.69325, 39.07178, 
    39.44474, 39.81194, 40.17321, 40.52837, 40.87727, 41.2197, 41.5555, 
    41.88448, 42.20646, 42.52125, 42.82867, 43.12852, 43.42064, 43.70482, 
    43.98088, 44.24864, 44.50792, 44.75852, 45.00027, 45.23299, 45.45651, 
    45.67065, 45.87524, 46.07014, 46.25516, 46.43016, 46.595, 46.74953, 
    46.89362, 47.02713, 47.14996, 47.26199, 47.36312, 47.45325, 47.53231, 
    47.6002, 47.65689, 47.7023, 47.7364, 47.75915, 47.77053, 47.77053, 
    47.75915, 47.7364, 47.7023, 47.65689, 47.6002, 47.53231, 47.45325, 
    47.36312, 47.26199, 47.14996, 47.02713, 46.89362, 46.74953, 46.595, 
    46.43016, 46.25516, 46.07014, 45.87524, 45.67065, 45.45651, 45.23299, 
    45.00027, 44.75852, 44.50792, 44.24864, 43.98088, 43.70482, 43.42064, 
    43.12852, 42.82867, 42.52125, 42.20646, 41.88448, 41.5555, 41.2197, 
    40.87727, 40.52837, 40.17321, 39.81194, 39.44474, 39.07178, 38.69325, 
    38.30929, 37.92007, 37.52576, 37.12651, 36.72248,
  36.36466, 36.75665, 37.14373, 37.52576, 37.90258, 38.27405, 38.64002, 
    39.00033, 39.35483, 39.70337, 40.04577, 40.38189, 40.71156, 41.03462, 
    41.35089, 41.66023, 41.96246, 42.2574, 42.54491, 42.82481, 43.09693, 
    43.36111, 43.61718, 43.86499, 44.10437, 44.33515, 44.55719, 44.77034, 
    44.97443, 45.16932, 45.35488, 45.53096, 45.69742, 45.85415, 46.00101, 
    46.13791, 46.26471, 46.38132, 46.48764, 46.5836, 46.66909, 46.74407, 
    46.80845, 46.86219, 46.90523, 46.93755, 46.95911, 46.96989, 46.96989, 
    46.95911, 46.93755, 46.90523, 46.86219, 46.80845, 46.74407, 46.66909, 
    46.5836, 46.48764, 46.38132, 46.26471, 46.13791, 46.00101, 45.85415, 
    45.69742, 45.53096, 45.35488, 45.16932, 44.97443, 44.77034, 44.55719, 
    44.33515, 44.10437, 43.86499, 43.61718, 43.36111, 43.09693, 42.82481, 
    42.54491, 42.2574, 41.96246, 41.66023, 41.35089, 41.03462, 40.71156, 
    40.38189, 40.04577, 39.70337, 39.35483, 39.00033, 38.64002, 38.27405, 
    37.90258, 37.52576, 37.14373, 36.75665, 36.36466,
  36.0016, 36.38164, 36.75665, 37.12651, 37.49107, 37.8502, 38.20377, 
    38.55162, 38.89363, 39.22964, 39.55952, 39.88312, 40.20029, 40.51088, 
    40.81476, 41.11176, 41.40174, 41.68456, 41.96006, 42.2281, 42.48852, 
    42.74119, 42.98596, 43.22269, 43.45123, 43.67144, 43.8832, 44.08636, 
    44.28079, 44.46637, 44.64297, 44.81047, 44.96877, 45.11773, 45.25727, 
    45.38729, 45.50768, 45.61835, 45.71924, 45.81026, 45.89135, 45.96243, 
    46.02346, 46.07439, 46.11519, 46.14581, 46.16624, 46.17646, 46.17646, 
    46.16624, 46.14581, 46.11519, 46.07439, 46.02346, 45.96243, 45.89135, 
    45.81026, 45.71924, 45.61835, 45.50768, 45.38729, 45.25727, 45.11773, 
    44.96877, 44.81047, 44.64297, 44.46637, 44.28079, 44.08636, 43.8832, 
    43.67144, 43.45123, 43.22269, 42.98596, 42.74119, 42.48852, 42.2281, 
    41.96006, 41.68456, 41.40174, 41.11176, 40.81476, 40.51088, 40.20029, 
    39.88312, 39.55952, 39.22964, 38.89363, 38.55162, 38.20377, 37.8502, 
    37.49107, 37.12651, 36.75665, 36.38164, 36.0016,
  35.63342, 36.0016, 36.36466, 36.72248, 37.07492, 37.42188, 37.76321, 
    38.09881, 38.42853, 38.75225, 39.06984, 39.38117, 39.68611, 39.98453, 
    40.27629, 40.56128, 40.83934, 41.11036, 41.37419, 41.63073, 41.87982, 
    42.12135, 42.35519, 42.58122, 42.7993, 43.00933, 43.21118, 43.40474, 
    43.58989, 43.76653, 43.93454, 44.09382, 44.24429, 44.38583, 44.51836, 
    44.64181, 44.75608, 44.8611, 44.9568, 45.04311, 45.11999, 45.18737, 
    45.24522, 45.29348, 45.33213, 45.36115, 45.3805, 45.39018, 45.39018, 
    45.3805, 45.36115, 45.33213, 45.29348, 45.24522, 45.18737, 45.11999, 
    45.04311, 44.9568, 44.8611, 44.75608, 44.64181, 44.51836, 44.38583, 
    44.24429, 44.09382, 43.93454, 43.76653, 43.58989, 43.40474, 43.21118, 
    43.00933, 42.7993, 42.58122, 42.35519, 42.12135, 41.87982, 41.63073, 
    41.37419, 41.11036, 40.83934, 40.56128, 40.27629, 39.98453, 39.68611, 
    39.38117, 39.06984, 38.75225, 38.42853, 38.09881, 37.76321, 37.42188, 
    37.07492, 36.72248, 36.36466, 36.0016, 35.63342 ;

 area =
  5.832426e+09, 5.885548e+09, 5.937712e+09, 5.988909e+09, 6.039129e+09, 
    6.088361e+09, 6.136596e+09, 6.183825e+09, 6.230037e+09, 6.275223e+09, 
    6.319373e+09, 6.362479e+09, 6.404531e+09, 6.445522e+09, 6.485442e+09, 
    6.524282e+09, 6.562035e+09, 6.598693e+09, 6.634248e+09, 6.668692e+09, 
    6.702019e+09, 6.734221e+09, 6.76529e+09, 6.795221e+09, 6.824007e+09, 
    6.851641e+09, 6.878117e+09, 6.903431e+09, 6.927576e+09, 6.950547e+09, 
    6.972339e+09, 6.992947e+09, 7.012366e+09, 7.030593e+09, 7.047623e+09, 
    7.063453e+09, 7.078078e+09, 7.091497e+09, 7.103705e+09, 7.1147e+09, 
    7.124479e+09, 7.133041e+09, 7.140384e+09, 7.146505e+09, 7.151404e+09, 
    7.155078e+09, 7.157529e+09, 7.158754e+09, 7.158754e+09, 7.157529e+09, 
    7.155078e+09, 7.151404e+09, 7.146505e+09, 7.140384e+09, 7.133041e+09, 
    7.124479e+09, 7.1147e+09, 7.103705e+09, 7.091497e+09, 7.078078e+09, 
    7.063453e+09, 7.047623e+09, 7.030593e+09, 7.012366e+09, 6.992947e+09, 
    6.972339e+09, 6.950547e+09, 6.927576e+09, 6.903431e+09, 6.878117e+09, 
    6.851641e+09, 6.824007e+09, 6.795221e+09, 6.76529e+09, 6.734221e+09, 
    6.702019e+09, 6.668692e+09, 6.634248e+09, 6.598693e+09, 6.562035e+09, 
    6.524282e+09, 6.485442e+09, 6.445522e+09, 6.404531e+09, 6.362479e+09, 
    6.319373e+09, 6.275223e+09, 6.230037e+09, 6.183825e+09, 6.136596e+09, 
    6.088361e+09, 6.039129e+09, 5.988909e+09, 5.937712e+09, 5.885548e+09, 
    5.832426e+09,
  5.885548e+09, 5.942029e+09, 5.99757e+09, 6.052155e+09, 6.105772e+09, 
    6.158404e+09, 6.210038e+09, 6.260659e+09, 6.310255e+09, 6.35881e+09, 
    6.406312e+09, 6.452746e+09, 6.4981e+09, 6.54236e+09, 6.585513e+09, 
    6.627547e+09, 6.668449e+09, 6.708208e+09, 6.74681e+09, 6.784244e+09, 
    6.8205e+09, 6.855565e+09, 6.889429e+09, 6.922081e+09, 6.953512e+09, 
    6.98371e+09, 7.012667e+09, 7.040374e+09, 7.066821e+09, 7.092e+09, 
    7.115902e+09, 7.138521e+09, 7.159848e+09, 7.179877e+09, 7.198601e+09, 
    7.216014e+09, 7.23211e+09, 7.246883e+09, 7.260329e+09, 7.272444e+09, 
    7.283223e+09, 7.292662e+09, 7.30076e+09, 7.307511e+09, 7.312915e+09, 
    7.316969e+09, 7.319673e+09, 7.321026e+09, 7.321026e+09, 7.319673e+09, 
    7.316969e+09, 7.312915e+09, 7.307511e+09, 7.30076e+09, 7.292662e+09, 
    7.283223e+09, 7.272444e+09, 7.260329e+09, 7.246883e+09, 7.23211e+09, 
    7.216014e+09, 7.198601e+09, 7.179877e+09, 7.159848e+09, 7.138521e+09, 
    7.115902e+09, 7.092e+09, 7.066821e+09, 7.040374e+09, 7.012667e+09, 
    6.98371e+09, 6.953512e+09, 6.922081e+09, 6.889429e+09, 6.855565e+09, 
    6.8205e+09, 6.784244e+09, 6.74681e+09, 6.708208e+09, 6.668449e+09, 
    6.627547e+09, 6.585513e+09, 6.54236e+09, 6.4981e+09, 6.452746e+09, 
    6.406312e+09, 6.35881e+09, 6.310255e+09, 6.260659e+09, 6.210038e+09, 
    6.158404e+09, 6.105772e+09, 6.052155e+09, 5.99757e+09, 5.942029e+09, 
    5.885548e+09,
  5.937712e+09, 5.99757e+09, 6.056508e+09, 6.114508e+09, 6.171552e+09, 
    6.227619e+09, 6.282692e+09, 6.336752e+09, 6.38978e+09, 6.441759e+09, 
    6.492669e+09, 6.542493e+09, 6.591213e+09, 6.638811e+09, 6.685269e+09, 
    6.730571e+09, 6.774699e+09, 6.817636e+09, 6.859367e+09, 6.899874e+09, 
    6.939143e+09, 6.977157e+09, 7.013901e+09, 7.049361e+09, 7.083523e+09, 
    7.116371e+09, 7.147894e+09, 7.178077e+09, 7.206909e+09, 7.234377e+09, 
    7.260469e+09, 7.285175e+09, 7.308484e+09, 7.330385e+09, 7.350871e+09, 
    7.36993e+09, 7.387556e+09, 7.403741e+09, 7.418477e+09, 7.431758e+09, 
    7.443579e+09, 7.453934e+09, 7.462817e+09, 7.470226e+09, 7.476158e+09, 
    7.480609e+09, 7.483577e+09, 7.485062e+09, 7.485062e+09, 7.483577e+09, 
    7.480609e+09, 7.476158e+09, 7.470226e+09, 7.462817e+09, 7.453934e+09, 
    7.443579e+09, 7.431758e+09, 7.418477e+09, 7.403741e+09, 7.387556e+09, 
    7.36993e+09, 7.350871e+09, 7.330385e+09, 7.308484e+09, 7.285175e+09, 
    7.260469e+09, 7.234377e+09, 7.206909e+09, 7.178077e+09, 7.147894e+09, 
    7.116371e+09, 7.083523e+09, 7.049361e+09, 7.013901e+09, 6.977157e+09, 
    6.939143e+09, 6.899874e+09, 6.859367e+09, 6.817636e+09, 6.774699e+09, 
    6.730571e+09, 6.685269e+09, 6.638811e+09, 6.591213e+09, 6.542493e+09, 
    6.492669e+09, 6.441759e+09, 6.38978e+09, 6.336752e+09, 6.282692e+09, 
    6.227619e+09, 6.171552e+09, 6.114508e+09, 6.056508e+09, 5.99757e+09, 
    5.937712e+09,
  5.988909e+09, 6.052155e+09, 6.114508e+09, 6.175945e+09, 6.236442e+09, 
    6.295976e+09, 6.354524e+09, 6.412062e+09, 6.468569e+09, 6.52402e+09, 
    6.578392e+09, 6.631664e+09, 6.683811e+09, 6.734811e+09, 6.784643e+09, 
    6.833284e+09, 6.880711e+09, 6.926904e+09, 6.971842e+09, 7.015503e+09, 
    7.057866e+09, 7.098912e+09, 7.13862e+09, 7.176973e+09, 7.21395e+09, 
    7.249533e+09, 7.283705e+09, 7.316448e+09, 7.347746e+09, 7.377583e+09, 
    7.405943e+09, 7.432813e+09, 7.458176e+09, 7.482021e+09, 7.504335e+09, 
    7.525106e+09, 7.544322e+09, 7.561974e+09, 7.578052e+09, 7.592547e+09, 
    7.605452e+09, 7.616759e+09, 7.626462e+09, 7.634556e+09, 7.641037e+09, 
    7.645901e+09, 7.649145e+09, 7.650767e+09, 7.650767e+09, 7.649145e+09, 
    7.645901e+09, 7.641037e+09, 7.634556e+09, 7.626462e+09, 7.616759e+09, 
    7.605452e+09, 7.592547e+09, 7.578052e+09, 7.561974e+09, 7.544322e+09, 
    7.525106e+09, 7.504335e+09, 7.482021e+09, 7.458176e+09, 7.432813e+09, 
    7.405943e+09, 7.377583e+09, 7.347746e+09, 7.316448e+09, 7.283705e+09, 
    7.249533e+09, 7.21395e+09, 7.176973e+09, 7.13862e+09, 7.098912e+09, 
    7.057866e+09, 7.015503e+09, 6.971842e+09, 6.926904e+09, 6.880711e+09, 
    6.833284e+09, 6.784643e+09, 6.734811e+09, 6.683811e+09, 6.631664e+09, 
    6.578392e+09, 6.52402e+09, 6.468569e+09, 6.412062e+09, 6.354524e+09, 
    6.295976e+09, 6.236442e+09, 6.175945e+09, 6.114508e+09, 6.052155e+09, 
    5.988909e+09,
  6.039129e+09, 6.105772e+09, 6.171552e+09, 6.236442e+09, 6.300414e+09, 
    6.363442e+09, 6.425497e+09, 6.486551e+09, 6.546576e+09, 6.605544e+09, 
    6.663429e+09, 6.720201e+09, 6.775833e+09, 6.830297e+09, 6.883567e+09, 
    6.935614e+09, 6.986412e+09, 7.035934e+09, 7.084154e+09, 7.131045e+09, 
    7.176583e+09, 7.220742e+09, 7.263496e+09, 7.304823e+09, 7.344698e+09, 
    7.383099e+09, 7.420003e+09, 7.455388e+09, 7.489233e+09, 7.521518e+09, 
    7.552224e+09, 7.581331e+09, 7.608822e+09, 7.634681e+09, 7.65889e+09, 
    7.681435e+09, 7.702302e+09, 7.721477e+09, 7.738948e+09, 7.754704e+09, 
    7.768736e+09, 7.781033e+09, 7.791588e+09, 7.800395e+09, 7.807448e+09, 
    7.812741e+09, 7.816271e+09, 7.818037e+09, 7.818037e+09, 7.816271e+09, 
    7.812741e+09, 7.807448e+09, 7.800395e+09, 7.791588e+09, 7.781033e+09, 
    7.768736e+09, 7.754704e+09, 7.738948e+09, 7.721477e+09, 7.702302e+09, 
    7.681435e+09, 7.65889e+09, 7.634681e+09, 7.608822e+09, 7.581331e+09, 
    7.552224e+09, 7.521518e+09, 7.489233e+09, 7.455388e+09, 7.420003e+09, 
    7.383099e+09, 7.344698e+09, 7.304823e+09, 7.263496e+09, 7.220742e+09, 
    7.176583e+09, 7.131045e+09, 7.084154e+09, 7.035934e+09, 6.986412e+09, 
    6.935614e+09, 6.883567e+09, 6.830297e+09, 6.775833e+09, 6.720201e+09, 
    6.663429e+09, 6.605544e+09, 6.546576e+09, 6.486551e+09, 6.425497e+09, 
    6.363442e+09, 6.300414e+09, 6.236442e+09, 6.171552e+09, 6.105772e+09, 
    6.039129e+09,
  6.088361e+09, 6.158404e+09, 6.227619e+09, 6.295976e+09, 6.363442e+09, 
    6.429985e+09, 6.495574e+09, 6.560175e+09, 6.623755e+09, 6.686283e+09, 
    6.747724e+09, 6.808046e+09, 6.867216e+09, 6.925201e+09, 6.981969e+09, 
    7.037487e+09, 7.091722e+09, 7.144643e+09, 7.196217e+09, 7.246414e+09, 
    7.295202e+09, 7.342552e+09, 7.388432e+09, 7.432814e+09, 7.475667e+09, 
    7.516966e+09, 7.556683e+09, 7.594789e+09, 7.631261e+09, 7.666072e+09, 
    7.699199e+09, 7.73062e+09, 7.760311e+09, 7.788252e+09, 7.814423e+09, 
    7.838806e+09, 7.861382e+09, 7.882135e+09, 7.901051e+09, 7.918115e+09, 
    7.933316e+09, 7.946641e+09, 7.958081e+09, 7.967627e+09, 7.975273e+09, 
    7.981012e+09, 7.984841e+09, 7.986756e+09, 7.986756e+09, 7.984841e+09, 
    7.981012e+09, 7.975273e+09, 7.967627e+09, 7.958081e+09, 7.946641e+09, 
    7.933316e+09, 7.918115e+09, 7.901051e+09, 7.882135e+09, 7.861382e+09, 
    7.838806e+09, 7.814423e+09, 7.788252e+09, 7.760311e+09, 7.73062e+09, 
    7.699199e+09, 7.666072e+09, 7.631261e+09, 7.594789e+09, 7.556683e+09, 
    7.516966e+09, 7.475667e+09, 7.432814e+09, 7.388432e+09, 7.342552e+09, 
    7.295202e+09, 7.246414e+09, 7.196217e+09, 7.144643e+09, 7.091722e+09, 
    7.037487e+09, 6.981969e+09, 6.925201e+09, 6.867216e+09, 6.808046e+09, 
    6.747724e+09, 6.686283e+09, 6.623755e+09, 6.560175e+09, 6.495574e+09, 
    6.429985e+09, 6.363442e+09, 6.295976e+09, 6.227619e+09, 6.158404e+09, 
    6.088361e+09,
  6.136596e+09, 6.210038e+09, 6.282692e+09, 6.354524e+09, 6.425497e+09, 
    6.495574e+09, 6.564719e+09, 6.632894e+09, 6.700061e+09, 6.766183e+09, 
    6.831222e+09, 6.895139e+09, 6.957896e+09, 7.019455e+09, 7.079777e+09, 
    7.138825e+09, 7.196561e+09, 7.252946e+09, 7.307944e+09, 7.361518e+09, 
    7.41363e+09, 7.464245e+09, 7.513327e+09, 7.56084e+09, 7.606751e+09, 
    7.651027e+09, 7.693634e+09, 7.734541e+09, 7.773715e+09, 7.811129e+09, 
    7.846753e+09, 7.880559e+09, 7.912521e+09, 7.942612e+09, 7.970811e+09, 
    7.997093e+09, 8.021437e+09, 8.043825e+09, 8.064236e+09, 8.082655e+09, 
    8.099066e+09, 8.113456e+09, 8.125813e+09, 8.136126e+09, 8.144387e+09, 
    8.150589e+09, 8.154726e+09, 8.156796e+09, 8.156796e+09, 8.154726e+09, 
    8.150589e+09, 8.144387e+09, 8.136126e+09, 8.125813e+09, 8.113456e+09, 
    8.099066e+09, 8.082655e+09, 8.064236e+09, 8.043825e+09, 8.021437e+09, 
    7.997093e+09, 7.970811e+09, 7.942612e+09, 7.912521e+09, 7.880559e+09, 
    7.846753e+09, 7.811129e+09, 7.773715e+09, 7.734541e+09, 7.693634e+09, 
    7.651027e+09, 7.606751e+09, 7.56084e+09, 7.513327e+09, 7.464245e+09, 
    7.41363e+09, 7.361518e+09, 7.307944e+09, 7.252946e+09, 7.196561e+09, 
    7.138825e+09, 7.079777e+09, 7.019455e+09, 6.957896e+09, 6.895139e+09, 
    6.831222e+09, 6.766183e+09, 6.700061e+09, 6.632894e+09, 6.564719e+09, 
    6.495574e+09, 6.425497e+09, 6.354524e+09, 6.282692e+09, 6.210038e+09, 
    6.136596e+09,
  6.183825e+09, 6.260659e+09, 6.336752e+09, 6.412062e+09, 6.486551e+09, 
    6.560175e+09, 6.632894e+09, 6.704666e+09, 6.775447e+09, 6.845195e+09, 
    6.913867e+09, 6.981418e+09, 7.047806e+09, 7.112987e+09, 7.176916e+09, 
    7.23955e+09, 7.300845e+09, 7.360757e+09, 7.419243e+09, 7.47626e+09, 
    7.531766e+09, 7.585717e+09, 7.638074e+09, 7.688794e+09, 7.737838e+09, 
    7.785166e+09, 7.830739e+09, 7.874522e+09, 7.916475e+09, 7.956566e+09, 
    7.994759e+09, 8.031022e+09, 8.065324e+09, 8.097633e+09, 8.127923e+09, 
    8.156166e+09, 8.182336e+09, 8.20641e+09, 8.228367e+09, 8.248187e+09, 
    8.26585e+09, 8.281342e+09, 8.294647e+09, 8.305754e+09, 8.314652e+09, 
    8.321333e+09, 8.32579e+09, 8.32802e+09, 8.32802e+09, 8.32579e+09, 
    8.321333e+09, 8.314652e+09, 8.305754e+09, 8.294647e+09, 8.281342e+09, 
    8.26585e+09, 8.248187e+09, 8.228367e+09, 8.20641e+09, 8.182336e+09, 
    8.156166e+09, 8.127923e+09, 8.097633e+09, 8.065324e+09, 8.031022e+09, 
    7.994759e+09, 7.956566e+09, 7.916475e+09, 7.874522e+09, 7.830739e+09, 
    7.785166e+09, 7.737838e+09, 7.688794e+09, 7.638074e+09, 7.585717e+09, 
    7.531766e+09, 7.47626e+09, 7.419243e+09, 7.360757e+09, 7.300845e+09, 
    7.23955e+09, 7.176916e+09, 7.112987e+09, 7.047806e+09, 6.981418e+09, 
    6.913867e+09, 6.845195e+09, 6.775447e+09, 6.704666e+09, 6.632894e+09, 
    6.560175e+09, 6.486551e+09, 6.412062e+09, 6.336752e+09, 6.260659e+09, 
    6.183825e+09,
  6.230037e+09, 6.310255e+09, 6.38978e+09, 6.468569e+09, 6.546576e+09, 
    6.623755e+09, 6.700061e+09, 6.775447e+09, 6.849864e+09, 6.923265e+09, 
    6.9956e+09, 7.066822e+09, 7.136881e+09, 7.205726e+09, 7.273309e+09, 
    7.339579e+09, 7.404488e+09, 7.467984e+09, 7.530018e+09, 7.590542e+09, 
    7.649507e+09, 7.706863e+09, 7.762563e+09, 7.816561e+09, 7.868808e+09, 
    7.919261e+09, 7.967875e+09, 8.014606e+09, 8.059411e+09, 8.10225e+09, 
    8.143084e+09, 8.181873e+09, 8.218582e+09, 8.253174e+09, 8.285618e+09, 
    8.31588e+09, 8.343933e+09, 8.369748e+09, 8.3933e+09, 8.414565e+09, 
    8.433522e+09, 8.450151e+09, 8.464436e+09, 8.476363e+09, 8.485919e+09, 
    8.493095e+09, 8.497883e+09, 8.500278e+09, 8.500278e+09, 8.497883e+09, 
    8.493095e+09, 8.485919e+09, 8.476363e+09, 8.464436e+09, 8.450151e+09, 
    8.433522e+09, 8.414565e+09, 8.3933e+09, 8.369748e+09, 8.343933e+09, 
    8.31588e+09, 8.285618e+09, 8.253174e+09, 8.218582e+09, 8.181873e+09, 
    8.143084e+09, 8.10225e+09, 8.059411e+09, 8.014606e+09, 7.967875e+09, 
    7.919261e+09, 7.868808e+09, 7.816561e+09, 7.762563e+09, 7.706863e+09, 
    7.649507e+09, 7.590542e+09, 7.530018e+09, 7.467984e+09, 7.404488e+09, 
    7.339579e+09, 7.273309e+09, 7.205726e+09, 7.136881e+09, 7.066822e+09, 
    6.9956e+09, 6.923265e+09, 6.849864e+09, 6.775447e+09, 6.700061e+09, 
    6.623755e+09, 6.546576e+09, 6.468569e+09, 6.38978e+09, 6.310255e+09, 
    6.230037e+09,
  6.275223e+09, 6.35881e+09, 6.441759e+09, 6.52402e+09, 6.605544e+09, 
    6.686283e+09, 6.766183e+09, 6.845195e+09, 6.923265e+09, 7.000339e+09, 
    7.076365e+09, 7.151286e+09, 7.225049e+09, 7.297597e+09, 7.368877e+09, 
    7.438829e+09, 7.5074e+09, 7.574533e+09, 7.640172e+09, 7.704261e+09, 
    7.766745e+09, 7.827569e+09, 7.886679e+09, 7.94402e+09, 7.99954e+09, 
    8.053188e+09, 8.10491e+09, 8.15466e+09, 8.202386e+09, 8.248043e+09, 
    8.291585e+09, 8.332967e+09, 8.372148e+09, 8.409087e+09, 8.443745e+09, 
    8.476086e+09, 8.506077e+09, 8.533684e+09, 8.558878e+09, 8.581632e+09, 
    8.601922e+09, 8.619724e+09, 8.63502e+09, 8.647793e+09, 8.658028e+09, 
    8.665715e+09, 8.670843e+09, 8.673409e+09, 8.673409e+09, 8.670843e+09, 
    8.665715e+09, 8.658028e+09, 8.647793e+09, 8.63502e+09, 8.619724e+09, 
    8.601922e+09, 8.581632e+09, 8.558878e+09, 8.533684e+09, 8.506077e+09, 
    8.476086e+09, 8.443745e+09, 8.409087e+09, 8.372148e+09, 8.332967e+09, 
    8.291585e+09, 8.248043e+09, 8.202386e+09, 8.15466e+09, 8.10491e+09, 
    8.053188e+09, 7.99954e+09, 7.94402e+09, 7.886679e+09, 7.827569e+09, 
    7.766745e+09, 7.704261e+09, 7.640172e+09, 7.574533e+09, 7.5074e+09, 
    7.438829e+09, 7.368877e+09, 7.297597e+09, 7.225049e+09, 7.151286e+09, 
    7.076365e+09, 7.000339e+09, 6.923265e+09, 6.845195e+09, 6.766183e+09, 
    6.686283e+09, 6.605544e+09, 6.52402e+09, 6.441759e+09, 6.35881e+09, 
    6.275223e+09,
  6.319373e+09, 6.406312e+09, 6.492669e+09, 6.578392e+09, 6.663429e+09, 
    6.747724e+09, 6.831222e+09, 6.913867e+09, 6.9956e+09, 7.076365e+09, 
    7.1561e+09, 7.234745e+09, 7.312241e+09, 7.388526e+09, 7.463537e+09, 
    7.537212e+09, 7.60949e+09, 7.680307e+09, 7.749601e+09, 7.817309e+09, 
    7.883369e+09, 7.94772e+09, 8.010299e+09, 8.071048e+09, 8.129904e+09, 
    8.186811e+09, 8.241709e+09, 8.294543e+09, 8.345257e+09, 8.393798e+09, 
    8.440113e+09, 8.484152e+09, 8.525868e+09, 8.565214e+09, 8.602145e+09, 
    8.636621e+09, 8.668601e+09, 8.698051e+09, 8.724934e+09, 8.749221e+09, 
    8.770882e+09, 8.789891e+09, 8.806228e+09, 8.819871e+09, 8.830806e+09, 
    8.839017e+09, 8.844498e+09, 8.84724e+09, 8.84724e+09, 8.844498e+09, 
    8.839017e+09, 8.830806e+09, 8.819871e+09, 8.806228e+09, 8.789891e+09, 
    8.770882e+09, 8.749221e+09, 8.724934e+09, 8.698051e+09, 8.668601e+09, 
    8.636621e+09, 8.602145e+09, 8.565214e+09, 8.525868e+09, 8.484152e+09, 
    8.440113e+09, 8.393798e+09, 8.345257e+09, 8.294543e+09, 8.241709e+09, 
    8.186811e+09, 8.129904e+09, 8.071048e+09, 8.010299e+09, 7.94772e+09, 
    7.883369e+09, 7.817309e+09, 7.749601e+09, 7.680307e+09, 7.60949e+09, 
    7.537212e+09, 7.463537e+09, 7.388526e+09, 7.312241e+09, 7.234745e+09, 
    7.1561e+09, 7.076365e+09, 6.9956e+09, 6.913867e+09, 6.831222e+09, 
    6.747724e+09, 6.663429e+09, 6.578392e+09, 6.492669e+09, 6.406312e+09, 
    6.319373e+09,
  6.362479e+09, 6.452746e+09, 6.542493e+09, 6.631664e+09, 6.720201e+09, 
    6.808046e+09, 6.895139e+09, 6.981418e+09, 7.066822e+09, 7.151286e+09, 
    7.234745e+09, 7.317134e+09, 7.398386e+09, 7.478433e+09, 7.557208e+09, 
    7.634641e+09, 7.710664e+09, 7.785207e+09, 7.858201e+09, 7.929576e+09, 
    7.999264e+09, 8.067195e+09, 8.133301e+09, 8.197513e+09, 8.259766e+09, 
    8.319992e+09, 8.378128e+09, 8.434108e+09, 8.487873e+09, 8.539359e+09, 
    8.58851e+09, 8.635267e+09, 8.679578e+09, 8.721389e+09, 8.760649e+09, 
    8.797313e+09, 8.831335e+09, 8.862674e+09, 8.891291e+09, 8.917151e+09, 
    8.940219e+09, 8.96047e+09, 8.977876e+09, 8.992415e+09, 9.004068e+09, 
    9.012821e+09, 9.018663e+09, 9.021585e+09, 9.021585e+09, 9.018663e+09, 
    9.012821e+09, 9.004068e+09, 8.992415e+09, 8.977876e+09, 8.96047e+09, 
    8.940219e+09, 8.917151e+09, 8.891291e+09, 8.862674e+09, 8.831335e+09, 
    8.797313e+09, 8.760649e+09, 8.721389e+09, 8.679578e+09, 8.635267e+09, 
    8.58851e+09, 8.539359e+09, 8.487873e+09, 8.434108e+09, 8.378128e+09, 
    8.319992e+09, 8.259766e+09, 8.197513e+09, 8.133301e+09, 8.067195e+09, 
    7.999264e+09, 7.929576e+09, 7.858201e+09, 7.785207e+09, 7.710664e+09, 
    7.634641e+09, 7.557208e+09, 7.478433e+09, 7.398386e+09, 7.317134e+09, 
    7.234745e+09, 7.151286e+09, 7.066822e+09, 6.981418e+09, 6.895139e+09, 
    6.808046e+09, 6.720201e+09, 6.631664e+09, 6.542493e+09, 6.452746e+09, 
    6.362479e+09,
  6.404531e+09, 6.4981e+09, 6.591213e+09, 6.683811e+09, 6.775833e+09, 
    6.867216e+09, 6.957896e+09, 7.047806e+09, 7.136881e+09, 7.225049e+09, 
    7.312241e+09, 7.398386e+09, 7.483411e+09, 7.567242e+09, 7.649805e+09, 
    7.731025e+09, 7.810825e+09, 7.889131e+09, 7.965864e+09, 8.04095e+09, 
    8.11431e+09, 8.18587e+09, 8.255552e+09, 8.323282e+09, 8.388985e+09, 
    8.452588e+09, 8.514017e+09, 8.573202e+09, 8.630074e+09, 8.684566e+09, 
    8.736609e+09, 8.786142e+09, 8.833104e+09, 8.877434e+09, 8.919077e+09, 
    8.95798e+09, 8.994092e+09, 9.027367e+09, 9.05776e+09, 9.085231e+09, 
    9.109745e+09, 9.131267e+09, 9.14977e+09, 9.165227e+09, 9.177618e+09, 
    9.186927e+09, 9.193139e+09, 9.196247e+09, 9.196247e+09, 9.193139e+09, 
    9.186927e+09, 9.177618e+09, 9.165227e+09, 9.14977e+09, 9.131267e+09, 
    9.109745e+09, 9.085231e+09, 9.05776e+09, 9.027367e+09, 8.994092e+09, 
    8.95798e+09, 8.919077e+09, 8.877434e+09, 8.833104e+09, 8.786142e+09, 
    8.736609e+09, 8.684566e+09, 8.630074e+09, 8.573202e+09, 8.514017e+09, 
    8.452588e+09, 8.388985e+09, 8.323282e+09, 8.255552e+09, 8.18587e+09, 
    8.11431e+09, 8.04095e+09, 7.965864e+09, 7.889131e+09, 7.810825e+09, 
    7.731025e+09, 7.649805e+09, 7.567242e+09, 7.483411e+09, 7.398386e+09, 
    7.312241e+09, 7.225049e+09, 7.136881e+09, 7.047806e+09, 6.957896e+09, 
    6.867216e+09, 6.775833e+09, 6.683811e+09, 6.591213e+09, 6.4981e+09, 
    6.404531e+09,
  6.445522e+09, 6.54236e+09, 6.638811e+09, 6.734811e+09, 6.830297e+09, 
    6.925201e+09, 7.019455e+09, 7.112987e+09, 7.205726e+09, 7.297597e+09, 
    7.388526e+09, 7.478433e+09, 7.567242e+09, 7.654872e+09, 7.741242e+09, 
    7.826271e+09, 7.909876e+09, 7.991974e+09, 8.072481e+09, 8.151313e+09, 
    8.228386e+09, 8.303616e+09, 8.37692e+09, 8.448214e+09, 8.517416e+09, 
    8.584445e+09, 8.649221e+09, 8.711665e+09, 8.771699e+09, 8.829247e+09, 
    8.884238e+09, 8.936601e+09, 8.986266e+09, 9.033167e+09, 9.077242e+09, 
    9.118431e+09, 9.156679e+09, 9.191932e+09, 9.224142e+09, 9.253263e+09, 
    9.279254e+09, 9.302078e+09, 9.321703e+09, 9.338102e+09, 9.351248e+09, 
    9.361125e+09, 9.367718e+09, 9.371016e+09, 9.371016e+09, 9.367718e+09, 
    9.361125e+09, 9.351248e+09, 9.338102e+09, 9.321703e+09, 9.302078e+09, 
    9.279254e+09, 9.253263e+09, 9.224142e+09, 9.191932e+09, 9.156679e+09, 
    9.118431e+09, 9.077242e+09, 9.033167e+09, 8.986266e+09, 8.936601e+09, 
    8.884238e+09, 8.829247e+09, 8.771699e+09, 8.711665e+09, 8.649221e+09, 
    8.584445e+09, 8.517416e+09, 8.448214e+09, 8.37692e+09, 8.303616e+09, 
    8.228386e+09, 8.151313e+09, 8.072481e+09, 7.991974e+09, 7.909876e+09, 
    7.826271e+09, 7.741242e+09, 7.654872e+09, 7.567242e+09, 7.478433e+09, 
    7.388526e+09, 7.297597e+09, 7.205726e+09, 7.112987e+09, 7.019455e+09, 
    6.925201e+09, 6.830297e+09, 6.734811e+09, 6.638811e+09, 6.54236e+09, 
    6.445522e+09,
  6.485442e+09, 6.585513e+09, 6.685269e+09, 6.784643e+09, 6.883567e+09, 
    6.981969e+09, 7.079777e+09, 7.176916e+09, 7.273309e+09, 7.368877e+09, 
    7.463537e+09, 7.557208e+09, 7.649805e+09, 7.741242e+09, 7.831433e+09, 
    7.920287e+09, 8.007716e+09, 8.093629e+09, 8.177936e+09, 8.260545e+09, 
    8.341364e+09, 8.420301e+09, 8.497266e+09, 8.572165e+09, 8.64491e+09, 
    8.715411e+09, 8.78358e+09, 8.849328e+09, 8.912572e+09, 8.973229e+09, 
    9.031216e+09, 9.086456e+09, 9.138871e+09, 9.188391e+09, 9.234944e+09, 
    9.278465e+09, 9.318892e+09, 9.356163e+09, 9.390226e+09, 9.421031e+09, 
    9.448532e+09, 9.472687e+09, 9.49346e+09, 9.510819e+09, 9.524738e+09, 
    9.535196e+09, 9.542177e+09, 9.54567e+09, 9.54567e+09, 9.542177e+09, 
    9.535196e+09, 9.524738e+09, 9.510819e+09, 9.49346e+09, 9.472687e+09, 
    9.448532e+09, 9.421031e+09, 9.390226e+09, 9.356163e+09, 9.318892e+09, 
    9.278465e+09, 9.234944e+09, 9.188391e+09, 9.138871e+09, 9.086456e+09, 
    9.031216e+09, 8.973229e+09, 8.912572e+09, 8.849328e+09, 8.78358e+09, 
    8.715411e+09, 8.64491e+09, 8.572165e+09, 8.497266e+09, 8.420301e+09, 
    8.341364e+09, 8.260545e+09, 8.177936e+09, 8.093629e+09, 8.007716e+09, 
    7.920287e+09, 7.831433e+09, 7.741242e+09, 7.649805e+09, 7.557208e+09, 
    7.463537e+09, 7.368877e+09, 7.273309e+09, 7.176916e+09, 7.079777e+09, 
    6.981969e+09, 6.883567e+09, 6.784643e+09, 6.685269e+09, 6.585513e+09, 
    6.485442e+09,
  6.524282e+09, 6.627547e+09, 6.730571e+09, 6.833284e+09, 6.935614e+09, 
    7.037487e+09, 7.138825e+09, 7.23955e+09, 7.339579e+09, 7.438829e+09, 
    7.537212e+09, 7.634641e+09, 7.731025e+09, 7.826271e+09, 7.920287e+09, 
    8.012976e+09, 8.104243e+09, 8.193989e+09, 8.282116e+09, 8.368525e+09, 
    8.453116e+09, 8.53579e+09, 8.616447e+09, 8.694987e+09, 8.771312e+09, 
    8.845323e+09, 8.916924e+09, 8.986021e+09, 9.052518e+09, 9.116325e+09, 
    9.177352e+09, 9.235513e+09, 9.290724e+09, 9.342905e+09, 9.391978e+09, 
    9.437871e+09, 9.480515e+09, 9.519842e+09, 9.555794e+09, 9.588315e+09, 
    9.617354e+09, 9.642865e+09, 9.664807e+09, 9.683147e+09, 9.697854e+09, 
    9.708905e+09, 9.716282e+09, 9.719975e+09, 9.719975e+09, 9.716282e+09, 
    9.708905e+09, 9.697854e+09, 9.683147e+09, 9.664807e+09, 9.642865e+09, 
    9.617354e+09, 9.588315e+09, 9.555794e+09, 9.519842e+09, 9.480515e+09, 
    9.437871e+09, 9.391978e+09, 9.342905e+09, 9.290724e+09, 9.235513e+09, 
    9.177352e+09, 9.116325e+09, 9.052518e+09, 8.986021e+09, 8.916924e+09, 
    8.845323e+09, 8.771312e+09, 8.694987e+09, 8.616447e+09, 8.53579e+09, 
    8.453116e+09, 8.368525e+09, 8.282116e+09, 8.193989e+09, 8.104243e+09, 
    8.012976e+09, 7.920287e+09, 7.826271e+09, 7.731025e+09, 7.634641e+09, 
    7.537212e+09, 7.438829e+09, 7.339579e+09, 7.23955e+09, 7.138825e+09, 
    7.037487e+09, 6.935614e+09, 6.833284e+09, 6.730571e+09, 6.627547e+09, 
    6.524282e+09,
  6.562035e+09, 6.668449e+09, 6.774699e+09, 6.880711e+09, 6.986412e+09, 
    7.091722e+09, 7.196561e+09, 7.300845e+09, 7.404488e+09, 7.5074e+09, 
    7.60949e+09, 7.710664e+09, 7.810825e+09, 7.909876e+09, 8.007716e+09, 
    8.104243e+09, 8.199353e+09, 8.292941e+09, 8.384902e+09, 8.475127e+09, 
    8.563511e+09, 8.649944e+09, 8.734319e+09, 8.816526e+09, 8.896461e+09, 
    8.974015e+09, 9.049084e+09, 9.121564e+09, 9.191351e+09, 9.258346e+09, 
    9.322452e+09, 9.383574e+09, 9.441618e+09, 9.496498e+09, 9.548129e+09, 
    9.596429e+09, 9.641325e+09, 9.68274e+09, 9.720613e+09, 9.754878e+09, 
    9.785482e+09, 9.812372e+09, 9.835507e+09, 9.854844e+09, 9.870353e+09, 
    9.882009e+09, 9.88979e+09, 9.893683e+09, 9.893683e+09, 9.88979e+09, 
    9.882009e+09, 9.870353e+09, 9.854844e+09, 9.835507e+09, 9.812372e+09, 
    9.785482e+09, 9.754878e+09, 9.720613e+09, 9.68274e+09, 9.641325e+09, 
    9.596429e+09, 9.548129e+09, 9.496498e+09, 9.441618e+09, 9.383574e+09, 
    9.322452e+09, 9.258346e+09, 9.191351e+09, 9.121564e+09, 9.049084e+09, 
    8.974015e+09, 8.896461e+09, 8.816526e+09, 8.734319e+09, 8.649944e+09, 
    8.563511e+09, 8.475127e+09, 8.384902e+09, 8.292941e+09, 8.199353e+09, 
    8.104243e+09, 8.007716e+09, 7.909876e+09, 7.810825e+09, 7.710664e+09, 
    7.60949e+09, 7.5074e+09, 7.404488e+09, 7.300845e+09, 7.196561e+09, 
    7.091722e+09, 6.986412e+09, 6.880711e+09, 6.774699e+09, 6.668449e+09, 
    6.562035e+09,
  6.598693e+09, 6.708208e+09, 6.817636e+09, 6.926904e+09, 7.035934e+09, 
    7.144643e+09, 7.252946e+09, 7.360757e+09, 7.467984e+09, 7.574533e+09, 
    7.680307e+09, 7.785207e+09, 7.889131e+09, 7.991974e+09, 8.093629e+09, 
    8.193989e+09, 8.292941e+09, 8.390374e+09, 8.486173e+09, 8.580225e+09, 
    8.672412e+09, 8.762619e+09, 8.85073e+09, 8.936627e+09, 9.020195e+09, 
    9.101317e+09, 9.17988e+09, 9.255772e+09, 9.32888e+09, 9.399095e+09, 
    9.466312e+09, 9.530426e+09, 9.591338e+09, 9.64895e+09, 9.703171e+09, 
    9.753911e+09, 9.801088e+09, 9.844622e+09, 9.884442e+09, 9.920478e+09, 
    9.95267e+09, 9.980962e+09, 1.00053e+10, 1.002566e+10, 1.004198e+10, 
    1.005425e+10, 1.006244e+10, 1.006654e+10, 1.006654e+10, 1.006244e+10, 
    1.005425e+10, 1.004198e+10, 1.002566e+10, 1.00053e+10, 9.980962e+09, 
    9.95267e+09, 9.920478e+09, 9.884442e+09, 9.844622e+09, 9.801088e+09, 
    9.753911e+09, 9.703171e+09, 9.64895e+09, 9.591338e+09, 9.530426e+09, 
    9.466312e+09, 9.399095e+09, 9.32888e+09, 9.255772e+09, 9.17988e+09, 
    9.101317e+09, 9.020195e+09, 8.936627e+09, 8.85073e+09, 8.762619e+09, 
    8.672412e+09, 8.580225e+09, 8.486173e+09, 8.390374e+09, 8.292941e+09, 
    8.193989e+09, 8.093629e+09, 7.991974e+09, 7.889131e+09, 7.785207e+09, 
    7.680307e+09, 7.574533e+09, 7.467984e+09, 7.360757e+09, 7.252946e+09, 
    7.144643e+09, 7.035934e+09, 6.926904e+09, 6.817636e+09, 6.708208e+09, 
    6.598693e+09,
  6.634248e+09, 6.74681e+09, 6.859367e+09, 6.971842e+09, 7.084154e+09, 
    7.196217e+09, 7.307944e+09, 7.419243e+09, 7.530018e+09, 7.640172e+09, 
    7.749601e+09, 7.858201e+09, 7.965864e+09, 8.072481e+09, 8.177936e+09, 
    8.282116e+09, 8.384902e+09, 8.486173e+09, 8.585809e+09, 8.683688e+09, 
    8.779684e+09, 8.873673e+09, 8.96553e+09, 9.055129e+09, 9.142345e+09, 
    9.227054e+09, 9.309132e+09, 9.388457e+09, 9.464909e+09, 9.53837e+09, 
    9.608722e+09, 9.675857e+09, 9.739662e+09, 9.800034e+09, 9.856871e+09, 
    9.910078e+09, 9.959563e+09, 1.000524e+10, 1.004703e+10, 1.008486e+10, 
    1.011866e+10, 1.014837e+10, 1.017394e+10, 1.019532e+10, 1.021247e+10, 
    1.022536e+10, 1.023397e+10, 1.023827e+10, 1.023827e+10, 1.023397e+10, 
    1.022536e+10, 1.021247e+10, 1.019532e+10, 1.017394e+10, 1.014837e+10, 
    1.011866e+10, 1.008486e+10, 1.004703e+10, 1.000524e+10, 9.959563e+09, 
    9.910078e+09, 9.856871e+09, 9.800034e+09, 9.739662e+09, 9.675857e+09, 
    9.608722e+09, 9.53837e+09, 9.464909e+09, 9.388457e+09, 9.309132e+09, 
    9.227054e+09, 9.142345e+09, 9.055129e+09, 8.96553e+09, 8.873673e+09, 
    8.779684e+09, 8.683688e+09, 8.585809e+09, 8.486173e+09, 8.384902e+09, 
    8.282116e+09, 8.177936e+09, 8.072481e+09, 7.965864e+09, 7.858201e+09, 
    7.749601e+09, 7.640172e+09, 7.530018e+09, 7.419243e+09, 7.307944e+09, 
    7.196217e+09, 7.084154e+09, 6.971842e+09, 6.859367e+09, 6.74681e+09, 
    6.634248e+09,
  6.668692e+09, 6.784244e+09, 6.899874e+09, 7.015503e+09, 7.131045e+09, 
    7.246414e+09, 7.361518e+09, 7.47626e+09, 7.590542e+09, 7.704261e+09, 
    7.817309e+09, 7.929576e+09, 8.04095e+09, 8.151313e+09, 8.260545e+09, 
    8.368525e+09, 8.475127e+09, 8.580225e+09, 8.683688e+09, 8.785385e+09, 
    8.885187e+09, 8.982957e+09, 9.078562e+09, 9.171869e+09, 9.262742e+09, 
    9.351046e+09, 9.436652e+09, 9.519426e+09, 9.599237e+09, 9.67596e+09, 
    9.749469e+09, 9.819643e+09, 9.886363e+09, 9.949515e+09, 1.000899e+10, 
    1.006469e+10, 1.01165e+10, 1.016434e+10, 1.020812e+10, 1.024776e+10, 
    1.028319e+10, 1.031433e+10, 1.034114e+10, 1.036355e+10, 1.038154e+10, 
    1.039506e+10, 1.040409e+10, 1.040861e+10, 1.040861e+10, 1.040409e+10, 
    1.039506e+10, 1.038154e+10, 1.036355e+10, 1.034114e+10, 1.031433e+10, 
    1.028319e+10, 1.024776e+10, 1.020812e+10, 1.016434e+10, 1.01165e+10, 
    1.006469e+10, 1.000899e+10, 9.949515e+09, 9.886363e+09, 9.819643e+09, 
    9.749469e+09, 9.67596e+09, 9.599237e+09, 9.519426e+09, 9.436652e+09, 
    9.351046e+09, 9.262742e+09, 9.171869e+09, 9.078562e+09, 8.982957e+09, 
    8.885187e+09, 8.785385e+09, 8.683688e+09, 8.580225e+09, 8.475127e+09, 
    8.368525e+09, 8.260545e+09, 8.151313e+09, 8.04095e+09, 7.929576e+09, 
    7.817309e+09, 7.704261e+09, 7.590542e+09, 7.47626e+09, 7.361518e+09, 
    7.246414e+09, 7.131045e+09, 7.015503e+09, 6.899874e+09, 6.784244e+09, 
    6.668692e+09,
  6.702019e+09, 6.8205e+09, 6.939143e+09, 7.057866e+09, 7.176583e+09, 
    7.295202e+09, 7.41363e+09, 7.531766e+09, 7.649507e+09, 7.766745e+09, 
    7.883369e+09, 7.999264e+09, 8.11431e+09, 8.228386e+09, 8.341364e+09, 
    8.453116e+09, 8.563511e+09, 8.672412e+09, 8.779684e+09, 8.885187e+09, 
    8.988781e+09, 9.090322e+09, 9.18967e+09, 9.286681e+09, 9.381209e+09, 
    9.473112e+09, 9.562249e+09, 9.648477e+09, 9.731658e+09, 9.811654e+09, 
    9.88833e+09, 9.961556e+09, 1.00312e+10, 1.009715e+10, 1.015928e+10, 
    1.021748e+10, 1.027164e+10, 1.032166e+10, 1.036744e+10, 1.040891e+10, 
    1.044597e+10, 1.047856e+10, 1.050662e+10, 1.053008e+10, 1.054891e+10, 
    1.056306e+10, 1.057252e+10, 1.057725e+10, 1.057725e+10, 1.057252e+10, 
    1.056306e+10, 1.054891e+10, 1.053008e+10, 1.050662e+10, 1.047856e+10, 
    1.044597e+10, 1.040891e+10, 1.036744e+10, 1.032166e+10, 1.027164e+10, 
    1.021748e+10, 1.015928e+10, 1.009715e+10, 1.00312e+10, 9.961556e+09, 
    9.88833e+09, 9.811654e+09, 9.731658e+09, 9.648477e+09, 9.562249e+09, 
    9.473112e+09, 9.381209e+09, 9.286681e+09, 9.18967e+09, 9.090322e+09, 
    8.988781e+09, 8.885187e+09, 8.779684e+09, 8.672412e+09, 8.563511e+09, 
    8.453116e+09, 8.341364e+09, 8.228386e+09, 8.11431e+09, 7.999264e+09, 
    7.883369e+09, 7.766745e+09, 7.649507e+09, 7.531766e+09, 7.41363e+09, 
    7.295202e+09, 7.176583e+09, 7.057866e+09, 6.939143e+09, 6.8205e+09, 
    6.702019e+09,
  6.734221e+09, 6.855565e+09, 6.977157e+09, 7.098912e+09, 7.220742e+09, 
    7.342552e+09, 7.464245e+09, 7.585717e+09, 7.706863e+09, 7.827569e+09, 
    7.94772e+09, 8.067195e+09, 8.18587e+09, 8.303616e+09, 8.420301e+09, 
    8.53579e+09, 8.649944e+09, 8.762619e+09, 8.873673e+09, 8.982957e+09, 
    9.090322e+09, 9.195619e+09, 9.298694e+09, 9.399396e+09, 9.497571e+09, 
    9.593066e+09, 9.68573e+09, 9.775411e+09, 9.861961e+09, 9.945231e+09, 
    1.002508e+10, 1.010136e+10, 1.017395e+10, 1.02427e+10, 1.030749e+10, 
    1.03682e+10, 1.042471e+10, 1.047692e+10, 1.052472e+10, 1.056802e+10, 
    1.060673e+10, 1.064077e+10, 1.067009e+10, 1.06946e+10, 1.071428e+10, 
    1.072907e+10, 1.073895e+10, 1.07439e+10, 1.07439e+10, 1.073895e+10, 
    1.072907e+10, 1.071428e+10, 1.06946e+10, 1.067009e+10, 1.064077e+10, 
    1.060673e+10, 1.056802e+10, 1.052472e+10, 1.047692e+10, 1.042471e+10, 
    1.03682e+10, 1.030749e+10, 1.02427e+10, 1.017395e+10, 1.010136e+10, 
    1.002508e+10, 9.945231e+09, 9.861961e+09, 9.775411e+09, 9.68573e+09, 
    9.593066e+09, 9.497571e+09, 9.399396e+09, 9.298694e+09, 9.195619e+09, 
    9.090322e+09, 8.982957e+09, 8.873673e+09, 8.762619e+09, 8.649944e+09, 
    8.53579e+09, 8.420301e+09, 8.303616e+09, 8.18587e+09, 8.067195e+09, 
    7.94772e+09, 7.827569e+09, 7.706863e+09, 7.585717e+09, 7.464245e+09, 
    7.342552e+09, 7.220742e+09, 7.098912e+09, 6.977157e+09, 6.855565e+09, 
    6.734221e+09,
  6.76529e+09, 6.889429e+09, 7.013901e+09, 7.13862e+09, 7.263496e+09, 
    7.388432e+09, 7.513327e+09, 7.638074e+09, 7.762563e+09, 7.886679e+09, 
    8.010299e+09, 8.133301e+09, 8.255552e+09, 8.37692e+09, 8.497266e+09, 
    8.616447e+09, 8.734319e+09, 8.85073e+09, 8.96553e+09, 9.078562e+09, 
    9.18967e+09, 9.298694e+09, 9.405474e+09, 9.509846e+09, 9.61165e+09, 
    9.710721e+09, 9.806899e+09, 9.900023e+09, 9.989933e+09, 1.007647e+10, 
    1.015949e+10, 1.023883e+10, 1.031435e+10, 1.03859e+10, 1.045336e+10, 
    1.051658e+10, 1.057545e+10, 1.062985e+10, 1.067967e+10, 1.07248e+10, 
    1.076517e+10, 1.080067e+10, 1.083124e+10, 1.085682e+10, 1.087735e+10, 
    1.089278e+10, 1.090309e+10, 1.090825e+10, 1.090825e+10, 1.090309e+10, 
    1.089278e+10, 1.087735e+10, 1.085682e+10, 1.083124e+10, 1.080067e+10, 
    1.076517e+10, 1.07248e+10, 1.067967e+10, 1.062985e+10, 1.057545e+10, 
    1.051658e+10, 1.045336e+10, 1.03859e+10, 1.031435e+10, 1.023883e+10, 
    1.015949e+10, 1.007647e+10, 9.989933e+09, 9.900023e+09, 9.806899e+09, 
    9.710721e+09, 9.61165e+09, 9.509846e+09, 9.405474e+09, 9.298694e+09, 
    9.18967e+09, 9.078562e+09, 8.96553e+09, 8.85073e+09, 8.734319e+09, 
    8.616447e+09, 8.497266e+09, 8.37692e+09, 8.255552e+09, 8.133301e+09, 
    8.010299e+09, 7.886679e+09, 7.762563e+09, 7.638074e+09, 7.513327e+09, 
    7.388432e+09, 7.263496e+09, 7.13862e+09, 7.013901e+09, 6.889429e+09, 
    6.76529e+09,
  6.795221e+09, 6.922081e+09, 7.049361e+09, 7.176973e+09, 7.304823e+09, 
    7.432814e+09, 7.56084e+09, 7.688794e+09, 7.816561e+09, 7.94402e+09, 
    8.071048e+09, 8.197513e+09, 8.323282e+09, 8.448214e+09, 8.572165e+09, 
    8.694987e+09, 8.816526e+09, 8.936627e+09, 9.055129e+09, 9.171869e+09, 
    9.286681e+09, 9.399396e+09, 9.509846e+09, 9.61786e+09, 9.723264e+09, 
    9.825887e+09, 9.925557e+09, 1.00221e+10, 1.011536e+10, 1.020515e+10, 
    1.029132e+10, 1.037371e+10, 1.045215e+10, 1.05265e+10, 1.059662e+10, 
    1.066235e+10, 1.072358e+10, 1.078017e+10, 1.0832e+10, 1.087898e+10, 
    1.092099e+10, 1.095795e+10, 1.098979e+10, 1.101642e+10, 1.10378e+10, 
    1.105388e+10, 1.106461e+10, 1.106999e+10, 1.106999e+10, 1.106461e+10, 
    1.105388e+10, 1.10378e+10, 1.101642e+10, 1.098979e+10, 1.095795e+10, 
    1.092099e+10, 1.087898e+10, 1.0832e+10, 1.078017e+10, 1.072358e+10, 
    1.066235e+10, 1.059662e+10, 1.05265e+10, 1.045215e+10, 1.037371e+10, 
    1.029132e+10, 1.020515e+10, 1.011536e+10, 1.00221e+10, 9.925557e+09, 
    9.825887e+09, 9.723264e+09, 9.61786e+09, 9.509846e+09, 9.399396e+09, 
    9.286681e+09, 9.171869e+09, 9.055129e+09, 8.936627e+09, 8.816526e+09, 
    8.694987e+09, 8.572165e+09, 8.448214e+09, 8.323282e+09, 8.197513e+09, 
    8.071048e+09, 7.94402e+09, 7.816561e+09, 7.688794e+09, 7.56084e+09, 
    7.432814e+09, 7.304823e+09, 7.176973e+09, 7.049361e+09, 6.922081e+09, 
    6.795221e+09,
  6.824007e+09, 6.953512e+09, 7.083523e+09, 7.21395e+09, 7.344698e+09, 
    7.475667e+09, 7.606751e+09, 7.737838e+09, 7.868808e+09, 7.99954e+09, 
    8.129904e+09, 8.259766e+09, 8.388985e+09, 8.517416e+09, 8.64491e+09, 
    8.771312e+09, 8.896461e+09, 9.020195e+09, 9.142345e+09, 9.262742e+09, 
    9.381209e+09, 9.497571e+09, 9.61165e+09, 9.723264e+09, 9.832232e+09, 
    9.938373e+09, 1.00415e+10, 1.014144e+10, 1.023802e+10, 1.033104e+10, 
    1.042034e+10, 1.050575e+10, 1.058711e+10, 1.066424e+10, 1.0737e+10, 
    1.080523e+10, 1.08688e+10, 1.092757e+10, 1.098142e+10, 1.103023e+10, 
    1.107389e+10, 1.111231e+10, 1.11454e+10, 1.117309e+10, 1.119532e+10, 
    1.121203e+10, 1.12232e+10, 1.122879e+10, 1.122879e+10, 1.12232e+10, 
    1.121203e+10, 1.119532e+10, 1.117309e+10, 1.11454e+10, 1.111231e+10, 
    1.107389e+10, 1.103023e+10, 1.098142e+10, 1.092757e+10, 1.08688e+10, 
    1.080523e+10, 1.0737e+10, 1.066424e+10, 1.058711e+10, 1.050575e+10, 
    1.042034e+10, 1.033104e+10, 1.023802e+10, 1.014144e+10, 1.00415e+10, 
    9.938373e+09, 9.832232e+09, 9.723264e+09, 9.61165e+09, 9.497571e+09, 
    9.381209e+09, 9.262742e+09, 9.142345e+09, 9.020195e+09, 8.896461e+09, 
    8.771312e+09, 8.64491e+09, 8.517416e+09, 8.388985e+09, 8.259766e+09, 
    8.129904e+09, 7.99954e+09, 7.868808e+09, 7.737838e+09, 7.606751e+09, 
    7.475667e+09, 7.344698e+09, 7.21395e+09, 7.083523e+09, 6.953512e+09, 
    6.824007e+09,
  6.851641e+09, 6.98371e+09, 7.116371e+09, 7.249533e+09, 7.383099e+09, 
    7.516966e+09, 7.651027e+09, 7.785166e+09, 7.919261e+09, 8.053188e+09, 
    8.186811e+09, 8.319992e+09, 8.452588e+09, 8.584445e+09, 8.715411e+09, 
    8.845323e+09, 8.974015e+09, 9.101317e+09, 9.227054e+09, 9.351046e+09, 
    9.473112e+09, 9.593066e+09, 9.710721e+09, 9.825887e+09, 9.938373e+09, 
    1.004799e+10, 1.015454e+10, 1.025783e+10, 1.035769e+10, 1.045391e+10, 
    1.054631e+10, 1.063472e+10, 1.071896e+10, 1.079885e+10, 1.087423e+10, 
    1.094495e+10, 1.101085e+10, 1.107179e+10, 1.112763e+10, 1.117826e+10, 
    1.122356e+10, 1.126342e+10, 1.129776e+10, 1.13265e+10, 1.134958e+10, 
    1.136693e+10, 1.137852e+10, 1.138432e+10, 1.138432e+10, 1.137852e+10, 
    1.136693e+10, 1.134958e+10, 1.13265e+10, 1.129776e+10, 1.126342e+10, 
    1.122356e+10, 1.117826e+10, 1.112763e+10, 1.107179e+10, 1.101085e+10, 
    1.094495e+10, 1.087423e+10, 1.079885e+10, 1.071896e+10, 1.063472e+10, 
    1.054631e+10, 1.045391e+10, 1.035769e+10, 1.025783e+10, 1.015454e+10, 
    1.004799e+10, 9.938373e+09, 9.825887e+09, 9.710721e+09, 9.593066e+09, 
    9.473112e+09, 9.351046e+09, 9.227054e+09, 9.101317e+09, 8.974015e+09, 
    8.845323e+09, 8.715411e+09, 8.584445e+09, 8.452588e+09, 8.319992e+09, 
    8.186811e+09, 8.053188e+09, 7.919261e+09, 7.785166e+09, 7.651027e+09, 
    7.516966e+09, 7.383099e+09, 7.249533e+09, 7.116371e+09, 6.98371e+09, 
    6.851641e+09,
  6.878117e+09, 7.012667e+09, 7.147894e+09, 7.283705e+09, 7.420003e+09, 
    7.556683e+09, 7.693634e+09, 7.830739e+09, 7.967875e+09, 8.10491e+09, 
    8.241709e+09, 8.378128e+09, 8.514017e+09, 8.649221e+09, 8.78358e+09, 
    8.916924e+09, 9.049084e+09, 9.17988e+09, 9.309132e+09, 9.436652e+09, 
    9.562249e+09, 9.68573e+09, 9.806899e+09, 9.925557e+09, 1.00415e+10, 
    1.015454e+10, 1.026446e+10, 1.037106e+10, 1.047415e+10, 1.057352e+10, 
    1.066899e+10, 1.076036e+10, 1.084745e+10, 1.093007e+10, 1.100805e+10, 
    1.108122e+10, 1.114942e+10, 1.12125e+10, 1.127033e+10, 1.132276e+10, 
    1.136968e+10, 1.141097e+10, 1.144656e+10, 1.147634e+10, 1.150025e+10, 
    1.151823e+10, 1.153025e+10, 1.153626e+10, 1.153626e+10, 1.153025e+10, 
    1.151823e+10, 1.150025e+10, 1.147634e+10, 1.144656e+10, 1.141097e+10, 
    1.136968e+10, 1.132276e+10, 1.127033e+10, 1.12125e+10, 1.114942e+10, 
    1.108122e+10, 1.100805e+10, 1.093007e+10, 1.084745e+10, 1.076036e+10, 
    1.066899e+10, 1.057352e+10, 1.047415e+10, 1.037106e+10, 1.026446e+10, 
    1.015454e+10, 1.00415e+10, 9.925557e+09, 9.806899e+09, 9.68573e+09, 
    9.562249e+09, 9.436652e+09, 9.309132e+09, 9.17988e+09, 9.049084e+09, 
    8.916924e+09, 8.78358e+09, 8.649221e+09, 8.514017e+09, 8.378128e+09, 
    8.241709e+09, 8.10491e+09, 7.967875e+09, 7.830739e+09, 7.693634e+09, 
    7.556683e+09, 7.420003e+09, 7.283705e+09, 7.147894e+09, 7.012667e+09, 
    6.878117e+09,
  6.903431e+09, 7.040374e+09, 7.178077e+09, 7.316448e+09, 7.455388e+09, 
    7.594789e+09, 7.734541e+09, 7.874522e+09, 8.014606e+09, 8.15466e+09, 
    8.294543e+09, 8.434108e+09, 8.573202e+09, 8.711665e+09, 8.849328e+09, 
    8.986021e+09, 9.121564e+09, 9.255772e+09, 9.388457e+09, 9.519426e+09, 
    9.648477e+09, 9.775411e+09, 9.900023e+09, 1.00221e+10, 1.014144e+10, 
    1.025783e+10, 1.037106e+10, 1.048091e+10, 1.058718e+10, 1.068966e+10, 
    1.078814e+10, 1.088243e+10, 1.097232e+10, 1.105763e+10, 1.113816e+10, 
    1.121375e+10, 1.128423e+10, 1.134943e+10, 1.14092e+10, 1.146341e+10, 
    1.151193e+10, 1.155465e+10, 1.159146e+10, 1.162227e+10, 1.164701e+10, 
    1.166561e+10, 1.167804e+10, 1.168427e+10, 1.168427e+10, 1.167804e+10, 
    1.166561e+10, 1.164701e+10, 1.162227e+10, 1.159146e+10, 1.155465e+10, 
    1.151193e+10, 1.146341e+10, 1.14092e+10, 1.134943e+10, 1.128423e+10, 
    1.121375e+10, 1.113816e+10, 1.105763e+10, 1.097232e+10, 1.088243e+10, 
    1.078814e+10, 1.068966e+10, 1.058718e+10, 1.048091e+10, 1.037106e+10, 
    1.025783e+10, 1.014144e+10, 1.00221e+10, 9.900023e+09, 9.775411e+09, 
    9.648477e+09, 9.519426e+09, 9.388457e+09, 9.255772e+09, 9.121564e+09, 
    8.986021e+09, 8.849328e+09, 8.711665e+09, 8.573202e+09, 8.434108e+09, 
    8.294543e+09, 8.15466e+09, 8.014606e+09, 7.874522e+09, 7.734541e+09, 
    7.594789e+09, 7.455388e+09, 7.316448e+09, 7.178077e+09, 7.040374e+09, 
    6.903431e+09,
  6.927576e+09, 7.066821e+09, 7.206909e+09, 7.347746e+09, 7.489233e+09, 
    7.631261e+09, 7.773715e+09, 7.916475e+09, 8.059411e+09, 8.202386e+09, 
    8.345257e+09, 8.487873e+09, 8.630074e+09, 8.771699e+09, 8.912572e+09, 
    9.052518e+09, 9.191351e+09, 9.32888e+09, 9.464909e+09, 9.599237e+09, 
    9.731658e+09, 9.861961e+09, 9.989933e+09, 1.011536e+10, 1.023802e+10, 
    1.035769e+10, 1.047415e+10, 1.058718e+10, 1.069657e+10, 1.080209e+10, 
    1.090352e+10, 1.100067e+10, 1.109331e+10, 1.118125e+10, 1.12643e+10, 
    1.134227e+10, 1.141498e+10, 1.148226e+10, 1.154395e+10, 1.159992e+10, 
    1.165001e+10, 1.169412e+10, 1.173213e+10, 1.176396e+10, 1.178951e+10, 
    1.180873e+10, 1.182158e+10, 1.1828e+10, 1.1828e+10, 1.182158e+10, 
    1.180873e+10, 1.178951e+10, 1.176396e+10, 1.173213e+10, 1.169412e+10, 
    1.165001e+10, 1.159992e+10, 1.154395e+10, 1.148226e+10, 1.141498e+10, 
    1.134227e+10, 1.12643e+10, 1.118125e+10, 1.109331e+10, 1.100067e+10, 
    1.090352e+10, 1.080209e+10, 1.069657e+10, 1.058718e+10, 1.047415e+10, 
    1.035769e+10, 1.023802e+10, 1.011536e+10, 9.989933e+09, 9.861961e+09, 
    9.731658e+09, 9.599237e+09, 9.464909e+09, 9.32888e+09, 9.191351e+09, 
    9.052518e+09, 8.912572e+09, 8.771699e+09, 8.630074e+09, 8.487873e+09, 
    8.345257e+09, 8.202386e+09, 8.059411e+09, 7.916475e+09, 7.773715e+09, 
    7.631261e+09, 7.489233e+09, 7.347746e+09, 7.206909e+09, 7.066821e+09, 
    6.927576e+09,
  6.950547e+09, 7.092e+09, 7.234377e+09, 7.377583e+09, 7.521518e+09, 
    7.666072e+09, 7.811129e+09, 7.956566e+09, 8.10225e+09, 8.248043e+09, 
    8.393798e+09, 8.539359e+09, 8.684566e+09, 8.829247e+09, 8.973229e+09, 
    9.116325e+09, 9.258346e+09, 9.399095e+09, 9.53837e+09, 9.67596e+09, 
    9.811654e+09, 9.945231e+09, 1.007647e+10, 1.020515e+10, 1.033104e+10, 
    1.045391e+10, 1.057352e+10, 1.068966e+10, 1.080209e+10, 1.091057e+10, 
    1.10149e+10, 1.111483e+10, 1.121017e+10, 1.130069e+10, 1.13862e+10, 
    1.146649e+10, 1.154138e+10, 1.16107e+10, 1.167428e+10, 1.173195e+10, 
    1.17836e+10, 1.182907e+10, 1.186826e+10, 1.190108e+10, 1.192743e+10, 
    1.194726e+10, 1.19605e+10, 1.196713e+10, 1.196713e+10, 1.19605e+10, 
    1.194726e+10, 1.192743e+10, 1.190108e+10, 1.186826e+10, 1.182907e+10, 
    1.17836e+10, 1.173195e+10, 1.167428e+10, 1.16107e+10, 1.154138e+10, 
    1.146649e+10, 1.13862e+10, 1.130069e+10, 1.121017e+10, 1.111483e+10, 
    1.10149e+10, 1.091057e+10, 1.080209e+10, 1.068966e+10, 1.057352e+10, 
    1.045391e+10, 1.033104e+10, 1.020515e+10, 1.007647e+10, 9.945231e+09, 
    9.811654e+09, 9.67596e+09, 9.53837e+09, 9.399095e+09, 9.258346e+09, 
    9.116325e+09, 8.973229e+09, 8.829247e+09, 8.684566e+09, 8.539359e+09, 
    8.393798e+09, 8.248043e+09, 8.10225e+09, 7.956566e+09, 7.811129e+09, 
    7.666072e+09, 7.521518e+09, 7.377583e+09, 7.234377e+09, 7.092e+09, 
    6.950547e+09,
  6.972339e+09, 7.115902e+09, 7.260469e+09, 7.405943e+09, 7.552224e+09, 
    7.699199e+09, 7.846753e+09, 7.994759e+09, 8.143084e+09, 8.291585e+09, 
    8.440113e+09, 8.58851e+09, 8.736609e+09, 8.884238e+09, 9.031216e+09, 
    9.177352e+09, 9.322452e+09, 9.466312e+09, 9.608722e+09, 9.749469e+09, 
    9.88833e+09, 1.002508e+10, 1.015949e+10, 1.029132e+10, 1.042034e+10, 
    1.054631e+10, 1.066899e+10, 1.078814e+10, 1.090352e+10, 1.10149e+10, 
    1.112203e+10, 1.122468e+10, 1.132264e+10, 1.141567e+10, 1.150357e+10, 
    1.158613e+10, 1.166315e+10, 1.173446e+10, 1.179987e+10, 1.185922e+10, 
    1.191237e+10, 1.195917e+10, 1.199952e+10, 1.203331e+10, 1.206044e+10, 
    1.208085e+10, 1.209449e+10, 1.210132e+10, 1.210132e+10, 1.209449e+10, 
    1.208085e+10, 1.206044e+10, 1.203331e+10, 1.199952e+10, 1.195917e+10, 
    1.191237e+10, 1.185922e+10, 1.179987e+10, 1.173446e+10, 1.166315e+10, 
    1.158613e+10, 1.150357e+10, 1.141567e+10, 1.132264e+10, 1.122468e+10, 
    1.112203e+10, 1.10149e+10, 1.090352e+10, 1.078814e+10, 1.066899e+10, 
    1.054631e+10, 1.042034e+10, 1.029132e+10, 1.015949e+10, 1.002508e+10, 
    9.88833e+09, 9.749469e+09, 9.608722e+09, 9.466312e+09, 9.322452e+09, 
    9.177352e+09, 9.031216e+09, 8.884238e+09, 8.736609e+09, 8.58851e+09, 
    8.440113e+09, 8.291585e+09, 8.143084e+09, 7.994759e+09, 7.846753e+09, 
    7.699199e+09, 7.552224e+09, 7.405943e+09, 7.260469e+09, 7.115902e+09, 
    6.972339e+09,
  6.992947e+09, 7.138521e+09, 7.285175e+09, 7.432813e+09, 7.581331e+09, 
    7.73062e+09, 7.880559e+09, 8.031022e+09, 8.181873e+09, 8.332967e+09, 
    8.484152e+09, 8.635267e+09, 8.786142e+09, 8.936601e+09, 9.086456e+09, 
    9.235513e+09, 9.383574e+09, 9.530426e+09, 9.675857e+09, 9.819643e+09, 
    9.961556e+09, 1.010136e+10, 1.023883e+10, 1.037371e+10, 1.050575e+10, 
    1.063472e+10, 1.076036e+10, 1.088243e+10, 1.100067e+10, 1.111483e+10, 
    1.122468e+10, 1.132997e+10, 1.143046e+10, 1.152593e+10, 1.161615e+10, 
    1.170091e+10, 1.178001e+10, 1.185324e+10, 1.192043e+10, 1.198141e+10, 
    1.203602e+10, 1.208412e+10, 1.212559e+10, 1.216031e+10, 1.218821e+10, 
    1.220919e+10, 1.222321e+10, 1.223023e+10, 1.223023e+10, 1.222321e+10, 
    1.220919e+10, 1.218821e+10, 1.216031e+10, 1.212559e+10, 1.208412e+10, 
    1.203602e+10, 1.198141e+10, 1.192043e+10, 1.185324e+10, 1.178001e+10, 
    1.170091e+10, 1.161615e+10, 1.152593e+10, 1.143046e+10, 1.132997e+10, 
    1.122468e+10, 1.111483e+10, 1.100067e+10, 1.088243e+10, 1.076036e+10, 
    1.063472e+10, 1.050575e+10, 1.037371e+10, 1.023883e+10, 1.010136e+10, 
    9.961556e+09, 9.819643e+09, 9.675857e+09, 9.530426e+09, 9.383574e+09, 
    9.235513e+09, 9.086456e+09, 8.936601e+09, 8.786142e+09, 8.635267e+09, 
    8.484152e+09, 8.332967e+09, 8.181873e+09, 8.031022e+09, 7.880559e+09, 
    7.73062e+09, 7.581331e+09, 7.432813e+09, 7.285175e+09, 7.138521e+09, 
    6.992947e+09,
  7.012366e+09, 7.159848e+09, 7.308484e+09, 7.458176e+09, 7.608822e+09, 
    7.760311e+09, 7.912521e+09, 8.065324e+09, 8.218582e+09, 8.372148e+09, 
    8.525868e+09, 8.679578e+09, 8.833104e+09, 8.986266e+09, 9.138871e+09, 
    9.290724e+09, 9.441618e+09, 9.591338e+09, 9.739662e+09, 9.886363e+09, 
    1.00312e+10, 1.017395e+10, 1.031435e+10, 1.045215e+10, 1.058711e+10, 
    1.071896e+10, 1.084745e+10, 1.097232e+10, 1.109331e+10, 1.121017e+10, 
    1.132264e+10, 1.143046e+10, 1.153341e+10, 1.163122e+10, 1.172369e+10, 
    1.181057e+10, 1.189166e+10, 1.196675e+10, 1.203567e+10, 1.209821e+10, 
    1.215424e+10, 1.220359e+10, 1.224615e+10, 1.228178e+10, 1.231041e+10, 
    1.233195e+10, 1.234634e+10, 1.235355e+10, 1.235355e+10, 1.234634e+10, 
    1.233195e+10, 1.231041e+10, 1.228178e+10, 1.224615e+10, 1.220359e+10, 
    1.215424e+10, 1.209821e+10, 1.203567e+10, 1.196675e+10, 1.189166e+10, 
    1.181057e+10, 1.172369e+10, 1.163122e+10, 1.153341e+10, 1.143046e+10, 
    1.132264e+10, 1.121017e+10, 1.109331e+10, 1.097232e+10, 1.084745e+10, 
    1.071896e+10, 1.058711e+10, 1.045215e+10, 1.031435e+10, 1.017395e+10, 
    1.00312e+10, 9.886363e+09, 9.739662e+09, 9.591338e+09, 9.441618e+09, 
    9.290724e+09, 9.138871e+09, 8.986266e+09, 8.833104e+09, 8.679578e+09, 
    8.525868e+09, 8.372148e+09, 8.218582e+09, 8.065324e+09, 7.912521e+09, 
    7.760311e+09, 7.608822e+09, 7.458176e+09, 7.308484e+09, 7.159848e+09, 
    7.012366e+09,
  7.030593e+09, 7.179877e+09, 7.330385e+09, 7.482021e+09, 7.634681e+09, 
    7.788252e+09, 7.942612e+09, 8.097633e+09, 8.253174e+09, 8.409087e+09, 
    8.565214e+09, 8.721389e+09, 8.877434e+09, 9.033167e+09, 9.188391e+09, 
    9.342905e+09, 9.496498e+09, 9.64895e+09, 9.800034e+09, 9.949515e+09, 
    1.009715e+10, 1.02427e+10, 1.03859e+10, 1.05265e+10, 1.066424e+10, 
    1.079885e+10, 1.093007e+10, 1.105763e+10, 1.118125e+10, 1.130069e+10, 
    1.141567e+10, 1.152593e+10, 1.163122e+10, 1.17313e+10, 1.182591e+10, 
    1.191483e+10, 1.199784e+10, 1.207473e+10, 1.214529e+10, 1.220935e+10, 
    1.226673e+10, 1.231729e+10, 1.236089e+10, 1.23974e+10, 1.242673e+10, 
    1.24488e+10, 1.246355e+10, 1.247093e+10, 1.247093e+10, 1.246355e+10, 
    1.24488e+10, 1.242673e+10, 1.23974e+10, 1.236089e+10, 1.231729e+10, 
    1.226673e+10, 1.220935e+10, 1.214529e+10, 1.207473e+10, 1.199784e+10, 
    1.191483e+10, 1.182591e+10, 1.17313e+10, 1.163122e+10, 1.152593e+10, 
    1.141567e+10, 1.130069e+10, 1.118125e+10, 1.105763e+10, 1.093007e+10, 
    1.079885e+10, 1.066424e+10, 1.05265e+10, 1.03859e+10, 1.02427e+10, 
    1.009715e+10, 9.949515e+09, 9.800034e+09, 9.64895e+09, 9.496498e+09, 
    9.342905e+09, 9.188391e+09, 9.033167e+09, 8.877434e+09, 8.721389e+09, 
    8.565214e+09, 8.409087e+09, 8.253174e+09, 8.097633e+09, 7.942612e+09, 
    7.788252e+09, 7.634681e+09, 7.482021e+09, 7.330385e+09, 7.179877e+09, 
    7.030593e+09,
  7.047623e+09, 7.198601e+09, 7.350871e+09, 7.504335e+09, 7.65889e+09, 
    7.814423e+09, 7.970811e+09, 8.127923e+09, 8.285618e+09, 8.443745e+09, 
    8.602145e+09, 8.760649e+09, 8.919077e+09, 9.077242e+09, 9.234944e+09, 
    9.391978e+09, 9.548129e+09, 9.703171e+09, 9.856871e+09, 1.000899e+10, 
    1.015928e+10, 1.030749e+10, 1.045336e+10, 1.059662e+10, 1.0737e+10, 
    1.087423e+10, 1.100805e+10, 1.113816e+10, 1.12643e+10, 1.13862e+10, 
    1.150357e+10, 1.161615e+10, 1.172369e+10, 1.182591e+10, 1.192258e+10, 
    1.201345e+10, 1.209829e+10, 1.217688e+10, 1.224902e+10, 1.231452e+10, 
    1.237321e+10, 1.242492e+10, 1.246951e+10, 1.250686e+10, 1.253687e+10, 
    1.255944e+10, 1.257453e+10, 1.258209e+10, 1.258209e+10, 1.257453e+10, 
    1.255944e+10, 1.253687e+10, 1.250686e+10, 1.246951e+10, 1.242492e+10, 
    1.237321e+10, 1.231452e+10, 1.224902e+10, 1.217688e+10, 1.209829e+10, 
    1.201345e+10, 1.192258e+10, 1.182591e+10, 1.172369e+10, 1.161615e+10, 
    1.150357e+10, 1.13862e+10, 1.12643e+10, 1.113816e+10, 1.100805e+10, 
    1.087423e+10, 1.0737e+10, 1.059662e+10, 1.045336e+10, 1.030749e+10, 
    1.015928e+10, 1.000899e+10, 9.856871e+09, 9.703171e+09, 9.548129e+09, 
    9.391978e+09, 9.234944e+09, 9.077242e+09, 8.919077e+09, 8.760649e+09, 
    8.602145e+09, 8.443745e+09, 8.285618e+09, 8.127923e+09, 7.970811e+09, 
    7.814423e+09, 7.65889e+09, 7.504335e+09, 7.350871e+09, 7.198601e+09, 
    7.047623e+09,
  7.063453e+09, 7.216014e+09, 7.36993e+09, 7.525106e+09, 7.681435e+09, 
    7.838806e+09, 7.997093e+09, 8.156166e+09, 8.31588e+09, 8.476086e+09, 
    8.636621e+09, 8.797313e+09, 8.95798e+09, 9.118431e+09, 9.278465e+09, 
    9.437871e+09, 9.596429e+09, 9.753911e+09, 9.910078e+09, 1.006469e+10, 
    1.021748e+10, 1.03682e+10, 1.051658e+10, 1.066235e+10, 1.080523e+10, 
    1.094495e+10, 1.108122e+10, 1.121375e+10, 1.134227e+10, 1.146649e+10, 
    1.158613e+10, 1.170091e+10, 1.181057e+10, 1.191483e+10, 1.201345e+10, 
    1.210616e+10, 1.219274e+10, 1.227295e+10, 1.234659e+10, 1.241347e+10, 
    1.247338e+10, 1.252618e+10, 1.257172e+10, 1.260987e+10, 1.264052e+10, 
    1.266358e+10, 1.267899e+10, 1.268671e+10, 1.268671e+10, 1.267899e+10, 
    1.266358e+10, 1.264052e+10, 1.260987e+10, 1.257172e+10, 1.252618e+10, 
    1.247338e+10, 1.241347e+10, 1.234659e+10, 1.227295e+10, 1.219274e+10, 
    1.210616e+10, 1.201345e+10, 1.191483e+10, 1.181057e+10, 1.170091e+10, 
    1.158613e+10, 1.146649e+10, 1.134227e+10, 1.121375e+10, 1.108122e+10, 
    1.094495e+10, 1.080523e+10, 1.066235e+10, 1.051658e+10, 1.03682e+10, 
    1.021748e+10, 1.006469e+10, 9.910078e+09, 9.753911e+09, 9.596429e+09, 
    9.437871e+09, 9.278465e+09, 9.118431e+09, 8.95798e+09, 8.797313e+09, 
    8.636621e+09, 8.476086e+09, 8.31588e+09, 8.156166e+09, 7.997093e+09, 
    7.838806e+09, 7.681435e+09, 7.525106e+09, 7.36993e+09, 7.216014e+09, 
    7.063453e+09,
  7.078078e+09, 7.23211e+09, 7.387556e+09, 7.544322e+09, 7.702302e+09, 
    7.861382e+09, 8.021437e+09, 8.182336e+09, 8.343933e+09, 8.506077e+09, 
    8.668601e+09, 8.831335e+09, 8.994092e+09, 9.156679e+09, 9.318892e+09, 
    9.480515e+09, 9.641325e+09, 9.801088e+09, 9.959563e+09, 1.01165e+10, 
    1.027164e+10, 1.042471e+10, 1.057545e+10, 1.072358e+10, 1.08688e+10, 
    1.101085e+10, 1.114942e+10, 1.128423e+10, 1.141498e+10, 1.154138e+10, 
    1.166315e+10, 1.178001e+10, 1.189166e+10, 1.199784e+10, 1.209829e+10, 
    1.219274e+10, 1.228095e+10, 1.236269e+10, 1.243775e+10, 1.250591e+10, 
    1.256699e+10, 1.262082e+10, 1.266725e+10, 1.270614e+10, 1.273739e+10, 
    1.276091e+10, 1.277663e+10, 1.27845e+10, 1.27845e+10, 1.277663e+10, 
    1.276091e+10, 1.273739e+10, 1.270614e+10, 1.266725e+10, 1.262082e+10, 
    1.256699e+10, 1.250591e+10, 1.243775e+10, 1.236269e+10, 1.228095e+10, 
    1.219274e+10, 1.209829e+10, 1.199784e+10, 1.189166e+10, 1.178001e+10, 
    1.166315e+10, 1.154138e+10, 1.141498e+10, 1.128423e+10, 1.114942e+10, 
    1.101085e+10, 1.08688e+10, 1.072358e+10, 1.057545e+10, 1.042471e+10, 
    1.027164e+10, 1.01165e+10, 9.959563e+09, 9.801088e+09, 9.641325e+09, 
    9.480515e+09, 9.318892e+09, 9.156679e+09, 8.994092e+09, 8.831335e+09, 
    8.668601e+09, 8.506077e+09, 8.343933e+09, 8.182336e+09, 8.021437e+09, 
    7.861382e+09, 7.702302e+09, 7.544322e+09, 7.387556e+09, 7.23211e+09, 
    7.078078e+09,
  7.091497e+09, 7.246883e+09, 7.403741e+09, 7.561974e+09, 7.721477e+09, 
    7.882135e+09, 8.043825e+09, 8.20641e+09, 8.369748e+09, 8.533684e+09, 
    8.698051e+09, 8.862674e+09, 9.027367e+09, 9.191932e+09, 9.356163e+09, 
    9.519842e+09, 9.68274e+09, 9.844622e+09, 1.000524e+10, 1.016434e+10, 
    1.032166e+10, 1.047692e+10, 1.062985e+10, 1.078017e+10, 1.092757e+10, 
    1.107179e+10, 1.12125e+10, 1.134943e+10, 1.148226e+10, 1.16107e+10, 
    1.173446e+10, 1.185324e+10, 1.196675e+10, 1.207473e+10, 1.217688e+10, 
    1.227295e+10, 1.236269e+10, 1.244586e+10, 1.252223e+10, 1.25916e+10, 
    1.265377e+10, 1.270856e+10, 1.275582e+10, 1.279542e+10, 1.282723e+10, 
    1.285118e+10, 1.286718e+10, 1.287519e+10, 1.287519e+10, 1.286718e+10, 
    1.285118e+10, 1.282723e+10, 1.279542e+10, 1.275582e+10, 1.270856e+10, 
    1.265377e+10, 1.25916e+10, 1.252223e+10, 1.244586e+10, 1.236269e+10, 
    1.227295e+10, 1.217688e+10, 1.207473e+10, 1.196675e+10, 1.185324e+10, 
    1.173446e+10, 1.16107e+10, 1.148226e+10, 1.134943e+10, 1.12125e+10, 
    1.107179e+10, 1.092757e+10, 1.078017e+10, 1.062985e+10, 1.047692e+10, 
    1.032166e+10, 1.016434e+10, 1.000524e+10, 9.844622e+09, 9.68274e+09, 
    9.519842e+09, 9.356163e+09, 9.191932e+09, 9.027367e+09, 8.862674e+09, 
    8.698051e+09, 8.533684e+09, 8.369748e+09, 8.20641e+09, 8.043825e+09, 
    7.882135e+09, 7.721477e+09, 7.561974e+09, 7.403741e+09, 7.246883e+09, 
    7.091497e+09,
  7.103705e+09, 7.260329e+09, 7.418477e+09, 7.578052e+09, 7.738948e+09, 
    7.901051e+09, 8.064236e+09, 8.228367e+09, 8.3933e+09, 8.558878e+09, 
    8.724934e+09, 8.891291e+09, 9.05776e+09, 9.224142e+09, 9.390226e+09, 
    9.555794e+09, 9.720613e+09, 9.884442e+09, 1.004703e+10, 1.020812e+10, 
    1.036744e+10, 1.052472e+10, 1.067967e+10, 1.0832e+10, 1.098142e+10, 
    1.112763e+10, 1.127033e+10, 1.14092e+10, 1.154395e+10, 1.167428e+10, 
    1.179987e+10, 1.192043e+10, 1.203567e+10, 1.214529e+10, 1.224902e+10, 
    1.234659e+10, 1.243775e+10, 1.252223e+10, 1.259983e+10, 1.267031e+10, 
    1.273348e+10, 1.278916e+10, 1.283719e+10, 1.287743e+10, 1.290977e+10, 
    1.293411e+10, 1.295038e+10, 1.295852e+10, 1.295852e+10, 1.295038e+10, 
    1.293411e+10, 1.290977e+10, 1.287743e+10, 1.283719e+10, 1.278916e+10, 
    1.273348e+10, 1.267031e+10, 1.259983e+10, 1.252223e+10, 1.243775e+10, 
    1.234659e+10, 1.224902e+10, 1.214529e+10, 1.203567e+10, 1.192043e+10, 
    1.179987e+10, 1.167428e+10, 1.154395e+10, 1.14092e+10, 1.127033e+10, 
    1.112763e+10, 1.098142e+10, 1.0832e+10, 1.067967e+10, 1.052472e+10, 
    1.036744e+10, 1.020812e+10, 1.004703e+10, 9.884442e+09, 9.720613e+09, 
    9.555794e+09, 9.390226e+09, 9.224142e+09, 9.05776e+09, 8.891291e+09, 
    8.724934e+09, 8.558878e+09, 8.3933e+09, 8.228367e+09, 8.064236e+09, 
    7.901051e+09, 7.738948e+09, 7.578052e+09, 7.418477e+09, 7.260329e+09, 
    7.103705e+09,
  7.1147e+09, 7.272444e+09, 7.431758e+09, 7.592547e+09, 7.754704e+09, 
    7.918115e+09, 8.082655e+09, 8.248187e+09, 8.414565e+09, 8.581632e+09, 
    8.749221e+09, 8.917151e+09, 9.085231e+09, 9.253263e+09, 9.421031e+09, 
    9.588315e+09, 9.754878e+09, 9.920478e+09, 1.008486e+10, 1.024776e+10, 
    1.040891e+10, 1.056802e+10, 1.07248e+10, 1.087898e+10, 1.103023e+10, 
    1.117826e+10, 1.132276e+10, 1.146341e+10, 1.159992e+10, 1.173195e+10, 
    1.185922e+10, 1.198141e+10, 1.209821e+10, 1.220935e+10, 1.231452e+10, 
    1.241347e+10, 1.250591e+10, 1.25916e+10, 1.267031e+10, 1.27418e+10, 
    1.280589e+10, 1.286239e+10, 1.291113e+10, 1.295196e+10, 1.298478e+10, 
    1.300948e+10, 1.302599e+10, 1.303425e+10, 1.303425e+10, 1.302599e+10, 
    1.300948e+10, 1.298478e+10, 1.295196e+10, 1.291113e+10, 1.286239e+10, 
    1.280589e+10, 1.27418e+10, 1.267031e+10, 1.25916e+10, 1.250591e+10, 
    1.241347e+10, 1.231452e+10, 1.220935e+10, 1.209821e+10, 1.198141e+10, 
    1.185922e+10, 1.173195e+10, 1.159992e+10, 1.146341e+10, 1.132276e+10, 
    1.117826e+10, 1.103023e+10, 1.087898e+10, 1.07248e+10, 1.056802e+10, 
    1.040891e+10, 1.024776e+10, 1.008486e+10, 9.920478e+09, 9.754878e+09, 
    9.588315e+09, 9.421031e+09, 9.253263e+09, 9.085231e+09, 8.917151e+09, 
    8.749221e+09, 8.581632e+09, 8.414565e+09, 8.248187e+09, 8.082655e+09, 
    7.918115e+09, 7.754704e+09, 7.592547e+09, 7.431758e+09, 7.272444e+09, 
    7.1147e+09,
  7.124479e+09, 7.283223e+09, 7.443579e+09, 7.605452e+09, 7.768736e+09, 
    7.933316e+09, 8.099066e+09, 8.26585e+09, 8.433522e+09, 8.601922e+09, 
    8.770882e+09, 8.940219e+09, 9.109745e+09, 9.279254e+09, 9.448532e+09, 
    9.617354e+09, 9.785482e+09, 9.95267e+09, 1.011866e+10, 1.028319e+10, 
    1.044597e+10, 1.060673e+10, 1.076517e+10, 1.092099e+10, 1.107389e+10, 
    1.122356e+10, 1.136968e+10, 1.151193e+10, 1.165001e+10, 1.17836e+10, 
    1.191237e+10, 1.203602e+10, 1.215424e+10, 1.226673e+10, 1.237321e+10, 
    1.247338e+10, 1.256699e+10, 1.265377e+10, 1.273348e+10, 1.280589e+10, 
    1.287081e+10, 1.292804e+10, 1.297741e+10, 1.301878e+10, 1.305203e+10, 
    1.307706e+10, 1.309378e+10, 1.310215e+10, 1.310215e+10, 1.309378e+10, 
    1.307706e+10, 1.305203e+10, 1.301878e+10, 1.297741e+10, 1.292804e+10, 
    1.287081e+10, 1.280589e+10, 1.273348e+10, 1.265377e+10, 1.256699e+10, 
    1.247338e+10, 1.237321e+10, 1.226673e+10, 1.215424e+10, 1.203602e+10, 
    1.191237e+10, 1.17836e+10, 1.165001e+10, 1.151193e+10, 1.136968e+10, 
    1.122356e+10, 1.107389e+10, 1.092099e+10, 1.076517e+10, 1.060673e+10, 
    1.044597e+10, 1.028319e+10, 1.011866e+10, 9.95267e+09, 9.785482e+09, 
    9.617354e+09, 9.448532e+09, 9.279254e+09, 9.109745e+09, 8.940219e+09, 
    8.770882e+09, 8.601922e+09, 8.433522e+09, 8.26585e+09, 8.099066e+09, 
    7.933316e+09, 7.768736e+09, 7.605452e+09, 7.443579e+09, 7.283223e+09, 
    7.124479e+09,
  7.133041e+09, 7.292662e+09, 7.453934e+09, 7.616759e+09, 7.781033e+09, 
    7.946641e+09, 8.113456e+09, 8.281342e+09, 8.450151e+09, 8.619724e+09, 
    8.789891e+09, 8.96047e+09, 9.131267e+09, 9.302078e+09, 9.472687e+09, 
    9.642865e+09, 9.812372e+09, 9.980962e+09, 1.014837e+10, 1.031433e+10, 
    1.047856e+10, 1.064077e+10, 1.080067e+10, 1.095795e+10, 1.111231e+10, 
    1.126342e+10, 1.141097e+10, 1.155465e+10, 1.169412e+10, 1.182907e+10, 
    1.195917e+10, 1.208412e+10, 1.220359e+10, 1.231729e+10, 1.242492e+10, 
    1.252618e+10, 1.262082e+10, 1.270856e+10, 1.278916e+10, 1.286239e+10, 
    1.292804e+10, 1.298592e+10, 1.303585e+10, 1.30777e+10, 1.311133e+10, 
    1.313664e+10, 1.315356e+10, 1.316203e+10, 1.316203e+10, 1.315356e+10, 
    1.313664e+10, 1.311133e+10, 1.30777e+10, 1.303585e+10, 1.298592e+10, 
    1.292804e+10, 1.286239e+10, 1.278916e+10, 1.270856e+10, 1.262082e+10, 
    1.252618e+10, 1.242492e+10, 1.231729e+10, 1.220359e+10, 1.208412e+10, 
    1.195917e+10, 1.182907e+10, 1.169412e+10, 1.155465e+10, 1.141097e+10, 
    1.126342e+10, 1.111231e+10, 1.095795e+10, 1.080067e+10, 1.064077e+10, 
    1.047856e+10, 1.031433e+10, 1.014837e+10, 9.980962e+09, 9.812372e+09, 
    9.642865e+09, 9.472687e+09, 9.302078e+09, 9.131267e+09, 8.96047e+09, 
    8.789891e+09, 8.619724e+09, 8.450151e+09, 8.281342e+09, 8.113456e+09, 
    7.946641e+09, 7.781033e+09, 7.616759e+09, 7.453934e+09, 7.292662e+09, 
    7.133041e+09,
  7.140384e+09, 7.30076e+09, 7.462817e+09, 7.626462e+09, 7.791588e+09, 
    7.958081e+09, 8.125813e+09, 8.294647e+09, 8.464436e+09, 8.63502e+09, 
    8.806228e+09, 8.977876e+09, 9.14977e+09, 9.321703e+09, 9.49346e+09, 
    9.664807e+09, 9.835507e+09, 1.00053e+10, 1.017394e+10, 1.034114e+10, 
    1.050662e+10, 1.067009e+10, 1.083124e+10, 1.098979e+10, 1.11454e+10, 
    1.129776e+10, 1.144656e+10, 1.159146e+10, 1.173213e+10, 1.186826e+10, 
    1.199952e+10, 1.212559e+10, 1.224615e+10, 1.236089e+10, 1.246951e+10, 
    1.257172e+10, 1.266725e+10, 1.275582e+10, 1.283719e+10, 1.291113e+10, 
    1.297741e+10, 1.303585e+10, 1.308628e+10, 1.312854e+10, 1.316249e+10, 
    1.318806e+10, 1.320514e+10, 1.32137e+10, 1.32137e+10, 1.320514e+10, 
    1.318806e+10, 1.316249e+10, 1.312854e+10, 1.308628e+10, 1.303585e+10, 
    1.297741e+10, 1.291113e+10, 1.283719e+10, 1.275582e+10, 1.266725e+10, 
    1.257172e+10, 1.246951e+10, 1.236089e+10, 1.224615e+10, 1.212559e+10, 
    1.199952e+10, 1.186826e+10, 1.173213e+10, 1.159146e+10, 1.144656e+10, 
    1.129776e+10, 1.11454e+10, 1.098979e+10, 1.083124e+10, 1.067009e+10, 
    1.050662e+10, 1.034114e+10, 1.017394e+10, 1.00053e+10, 9.835507e+09, 
    9.664807e+09, 9.49346e+09, 9.321703e+09, 9.14977e+09, 8.977876e+09, 
    8.806228e+09, 8.63502e+09, 8.464436e+09, 8.294647e+09, 8.125813e+09, 
    7.958081e+09, 7.791588e+09, 7.626462e+09, 7.462817e+09, 7.30076e+09, 
    7.140384e+09,
  7.146505e+09, 7.307511e+09, 7.470226e+09, 7.634556e+09, 7.800395e+09, 
    7.967627e+09, 8.136126e+09, 8.305754e+09, 8.476363e+09, 8.647793e+09, 
    8.819871e+09, 8.992415e+09, 9.165227e+09, 9.338102e+09, 9.510819e+09, 
    9.683147e+09, 9.854844e+09, 1.002566e+10, 1.019532e+10, 1.036355e+10, 
    1.053008e+10, 1.06946e+10, 1.085682e+10, 1.101642e+10, 1.117309e+10, 
    1.13265e+10, 1.147634e+10, 1.162227e+10, 1.176396e+10, 1.190108e+10, 
    1.203331e+10, 1.216031e+10, 1.228178e+10, 1.23974e+10, 1.250686e+10, 
    1.260987e+10, 1.270614e+10, 1.279542e+10, 1.287743e+10, 1.295196e+10, 
    1.301878e+10, 1.30777e+10, 1.312854e+10, 1.317114e+10, 1.320537e+10, 
    1.323115e+10, 1.324837e+10, 1.3257e+10, 1.3257e+10, 1.324837e+10, 
    1.323115e+10, 1.320537e+10, 1.317114e+10, 1.312854e+10, 1.30777e+10, 
    1.301878e+10, 1.295196e+10, 1.287743e+10, 1.279542e+10, 1.270614e+10, 
    1.260987e+10, 1.250686e+10, 1.23974e+10, 1.228178e+10, 1.216031e+10, 
    1.203331e+10, 1.190108e+10, 1.176396e+10, 1.162227e+10, 1.147634e+10, 
    1.13265e+10, 1.117309e+10, 1.101642e+10, 1.085682e+10, 1.06946e+10, 
    1.053008e+10, 1.036355e+10, 1.019532e+10, 1.002566e+10, 9.854844e+09, 
    9.683147e+09, 9.510819e+09, 9.338102e+09, 9.165227e+09, 8.992415e+09, 
    8.819871e+09, 8.647793e+09, 8.476363e+09, 8.305754e+09, 8.136126e+09, 
    7.967627e+09, 7.800395e+09, 7.634556e+09, 7.470226e+09, 7.307511e+09, 
    7.146505e+09,
  7.151404e+09, 7.312915e+09, 7.476158e+09, 7.641037e+09, 7.807448e+09, 
    7.975273e+09, 8.144387e+09, 8.314652e+09, 8.485919e+09, 8.658028e+09, 
    8.830806e+09, 9.004068e+09, 9.177618e+09, 9.351248e+09, 9.524738e+09, 
    9.697854e+09, 9.870353e+09, 1.004198e+10, 1.021247e+10, 1.038154e+10, 
    1.054891e+10, 1.071428e+10, 1.087735e+10, 1.10378e+10, 1.119532e+10, 
    1.134958e+10, 1.150025e+10, 1.164701e+10, 1.178951e+10, 1.192743e+10, 
    1.206044e+10, 1.218821e+10, 1.231041e+10, 1.242673e+10, 1.253687e+10, 
    1.264052e+10, 1.273739e+10, 1.282723e+10, 1.290977e+10, 1.298478e+10, 
    1.305203e+10, 1.311133e+10, 1.316249e+10, 1.320537e+10, 1.323984e+10, 
    1.326578e+10, 1.328312e+10, 1.32918e+10, 1.32918e+10, 1.328312e+10, 
    1.326578e+10, 1.323984e+10, 1.320537e+10, 1.316249e+10, 1.311133e+10, 
    1.305203e+10, 1.298478e+10, 1.290977e+10, 1.282723e+10, 1.273739e+10, 
    1.264052e+10, 1.253687e+10, 1.242673e+10, 1.231041e+10, 1.218821e+10, 
    1.206044e+10, 1.192743e+10, 1.178951e+10, 1.164701e+10, 1.150025e+10, 
    1.134958e+10, 1.119532e+10, 1.10378e+10, 1.087735e+10, 1.071428e+10, 
    1.054891e+10, 1.038154e+10, 1.021247e+10, 1.004198e+10, 9.870353e+09, 
    9.697854e+09, 9.524738e+09, 9.351248e+09, 9.177618e+09, 9.004068e+09, 
    8.830806e+09, 8.658028e+09, 8.485919e+09, 8.314652e+09, 8.144387e+09, 
    7.975273e+09, 7.807448e+09, 7.641037e+09, 7.476158e+09, 7.312915e+09, 
    7.151404e+09,
  7.155078e+09, 7.316969e+09, 7.480609e+09, 7.645901e+09, 7.812741e+09, 
    7.981012e+09, 8.150589e+09, 8.321333e+09, 8.493095e+09, 8.665715e+09, 
    8.839017e+09, 9.012821e+09, 9.186927e+09, 9.361125e+09, 9.535196e+09, 
    9.708905e+09, 9.882009e+09, 1.005425e+10, 1.022536e+10, 1.039506e+10, 
    1.056306e+10, 1.072907e+10, 1.089278e+10, 1.105388e+10, 1.121203e+10, 
    1.136693e+10, 1.151823e+10, 1.166561e+10, 1.180873e+10, 1.194726e+10, 
    1.208085e+10, 1.220919e+10, 1.233195e+10, 1.24488e+10, 1.255944e+10, 
    1.266358e+10, 1.276091e+10, 1.285118e+10, 1.293411e+10, 1.300948e+10, 
    1.307706e+10, 1.313664e+10, 1.318806e+10, 1.323115e+10, 1.326578e+10, 
    1.329185e+10, 1.330927e+10, 1.3318e+10, 1.3318e+10, 1.330927e+10, 
    1.329185e+10, 1.326578e+10, 1.323115e+10, 1.318806e+10, 1.313664e+10, 
    1.307706e+10, 1.300948e+10, 1.293411e+10, 1.285118e+10, 1.276091e+10, 
    1.266358e+10, 1.255944e+10, 1.24488e+10, 1.233195e+10, 1.220919e+10, 
    1.208085e+10, 1.194726e+10, 1.180873e+10, 1.166561e+10, 1.151823e+10, 
    1.136693e+10, 1.121203e+10, 1.105388e+10, 1.089278e+10, 1.072907e+10, 
    1.056306e+10, 1.039506e+10, 1.022536e+10, 1.005425e+10, 9.882009e+09, 
    9.708905e+09, 9.535196e+09, 9.361125e+09, 9.186927e+09, 9.012821e+09, 
    8.839017e+09, 8.665715e+09, 8.493095e+09, 8.321333e+09, 8.150589e+09, 
    7.981012e+09, 7.812741e+09, 7.645901e+09, 7.480609e+09, 7.316969e+09, 
    7.155078e+09,
  7.157529e+09, 7.319673e+09, 7.483577e+09, 7.649145e+09, 7.816271e+09, 
    7.984841e+09, 8.154726e+09, 8.32579e+09, 8.497883e+09, 8.670843e+09, 
    8.844498e+09, 9.018663e+09, 9.193139e+09, 9.367718e+09, 9.542177e+09, 
    9.716282e+09, 9.88979e+09, 1.006244e+10, 1.023397e+10, 1.040409e+10, 
    1.057252e+10, 1.073895e+10, 1.090309e+10, 1.106461e+10, 1.12232e+10, 
    1.137852e+10, 1.153025e+10, 1.167804e+10, 1.182158e+10, 1.19605e+10, 
    1.209449e+10, 1.222321e+10, 1.234634e+10, 1.246355e+10, 1.257453e+10, 
    1.267899e+10, 1.277663e+10, 1.286718e+10, 1.295038e+10, 1.302599e+10, 
    1.309378e+10, 1.315356e+10, 1.320514e+10, 1.324837e+10, 1.328312e+10, 
    1.330927e+10, 1.332675e+10, 1.333551e+10, 1.333551e+10, 1.332675e+10, 
    1.330927e+10, 1.328312e+10, 1.324837e+10, 1.320514e+10, 1.315356e+10, 
    1.309378e+10, 1.302599e+10, 1.295038e+10, 1.286718e+10, 1.277663e+10, 
    1.267899e+10, 1.257453e+10, 1.246355e+10, 1.234634e+10, 1.222321e+10, 
    1.209449e+10, 1.19605e+10, 1.182158e+10, 1.167804e+10, 1.153025e+10, 
    1.137852e+10, 1.12232e+10, 1.106461e+10, 1.090309e+10, 1.073895e+10, 
    1.057252e+10, 1.040409e+10, 1.023397e+10, 1.006244e+10, 9.88979e+09, 
    9.716282e+09, 9.542177e+09, 9.367718e+09, 9.193139e+09, 9.018663e+09, 
    8.844498e+09, 8.670843e+09, 8.497883e+09, 8.32579e+09, 8.154726e+09, 
    7.984841e+09, 7.816271e+09, 7.649145e+09, 7.483577e+09, 7.319673e+09, 
    7.157529e+09,
  7.158754e+09, 7.321026e+09, 7.485062e+09, 7.650767e+09, 7.818037e+09, 
    7.986756e+09, 8.156796e+09, 8.32802e+09, 8.500278e+09, 8.673409e+09, 
    8.84724e+09, 9.021585e+09, 9.196247e+09, 9.371016e+09, 9.54567e+09, 
    9.719975e+09, 9.893683e+09, 1.006654e+10, 1.023827e+10, 1.040861e+10, 
    1.057725e+10, 1.07439e+10, 1.090825e+10, 1.106999e+10, 1.122879e+10, 
    1.138432e+10, 1.153626e+10, 1.168427e+10, 1.1828e+10, 1.196713e+10, 
    1.210132e+10, 1.223023e+10, 1.235355e+10, 1.247093e+10, 1.258209e+10, 
    1.268671e+10, 1.27845e+10, 1.287519e+10, 1.295852e+10, 1.303425e+10, 
    1.310215e+10, 1.316203e+10, 1.32137e+10, 1.3257e+10, 1.32918e+10, 
    1.3318e+10, 1.333551e+10, 1.334428e+10, 1.334428e+10, 1.333551e+10, 
    1.3318e+10, 1.32918e+10, 1.3257e+10, 1.32137e+10, 1.316203e+10, 
    1.310215e+10, 1.303425e+10, 1.295852e+10, 1.287519e+10, 1.27845e+10, 
    1.268671e+10, 1.258209e+10, 1.247093e+10, 1.235355e+10, 1.223023e+10, 
    1.210132e+10, 1.196713e+10, 1.1828e+10, 1.168427e+10, 1.153626e+10, 
    1.138432e+10, 1.122879e+10, 1.106999e+10, 1.090825e+10, 1.07439e+10, 
    1.057725e+10, 1.040861e+10, 1.023827e+10, 1.006654e+10, 9.893683e+09, 
    9.719975e+09, 9.54567e+09, 9.371016e+09, 9.196247e+09, 9.021585e+09, 
    8.84724e+09, 8.673409e+09, 8.500278e+09, 8.32802e+09, 8.156796e+09, 
    7.986756e+09, 7.818037e+09, 7.650767e+09, 7.485062e+09, 7.321026e+09, 
    7.158754e+09,
  7.158754e+09, 7.321026e+09, 7.485062e+09, 7.650767e+09, 7.818037e+09, 
    7.986756e+09, 8.156796e+09, 8.32802e+09, 8.500278e+09, 8.673409e+09, 
    8.84724e+09, 9.021585e+09, 9.196247e+09, 9.371016e+09, 9.54567e+09, 
    9.719975e+09, 9.893683e+09, 1.006654e+10, 1.023827e+10, 1.040861e+10, 
    1.057725e+10, 1.07439e+10, 1.090825e+10, 1.106999e+10, 1.122879e+10, 
    1.138432e+10, 1.153626e+10, 1.168427e+10, 1.1828e+10, 1.196713e+10, 
    1.210132e+10, 1.223023e+10, 1.235355e+10, 1.247093e+10, 1.258209e+10, 
    1.268671e+10, 1.27845e+10, 1.287519e+10, 1.295852e+10, 1.303425e+10, 
    1.310215e+10, 1.316203e+10, 1.32137e+10, 1.3257e+10, 1.32918e+10, 
    1.3318e+10, 1.333551e+10, 1.334428e+10, 1.334428e+10, 1.333551e+10, 
    1.3318e+10, 1.32918e+10, 1.3257e+10, 1.32137e+10, 1.316203e+10, 
    1.310215e+10, 1.303425e+10, 1.295852e+10, 1.287519e+10, 1.27845e+10, 
    1.268671e+10, 1.258209e+10, 1.247093e+10, 1.235355e+10, 1.223023e+10, 
    1.210132e+10, 1.196713e+10, 1.1828e+10, 1.168427e+10, 1.153626e+10, 
    1.138432e+10, 1.122879e+10, 1.106999e+10, 1.090825e+10, 1.07439e+10, 
    1.057725e+10, 1.040861e+10, 1.023827e+10, 1.006654e+10, 9.893683e+09, 
    9.719975e+09, 9.54567e+09, 9.371016e+09, 9.196247e+09, 9.021585e+09, 
    8.84724e+09, 8.673409e+09, 8.500278e+09, 8.32802e+09, 8.156796e+09, 
    7.986756e+09, 7.818037e+09, 7.650767e+09, 7.485062e+09, 7.321026e+09, 
    7.158754e+09,
  7.157529e+09, 7.319673e+09, 7.483577e+09, 7.649145e+09, 7.816271e+09, 
    7.984841e+09, 8.154726e+09, 8.32579e+09, 8.497883e+09, 8.670843e+09, 
    8.844498e+09, 9.018663e+09, 9.193139e+09, 9.367718e+09, 9.542177e+09, 
    9.716282e+09, 9.88979e+09, 1.006244e+10, 1.023397e+10, 1.040409e+10, 
    1.057252e+10, 1.073895e+10, 1.090309e+10, 1.106461e+10, 1.12232e+10, 
    1.137852e+10, 1.153025e+10, 1.167804e+10, 1.182158e+10, 1.19605e+10, 
    1.209449e+10, 1.222321e+10, 1.234634e+10, 1.246355e+10, 1.257453e+10, 
    1.267899e+10, 1.277663e+10, 1.286718e+10, 1.295038e+10, 1.302599e+10, 
    1.309378e+10, 1.315356e+10, 1.320514e+10, 1.324837e+10, 1.328312e+10, 
    1.330927e+10, 1.332675e+10, 1.333551e+10, 1.333551e+10, 1.332675e+10, 
    1.330927e+10, 1.328312e+10, 1.324837e+10, 1.320514e+10, 1.315356e+10, 
    1.309378e+10, 1.302599e+10, 1.295038e+10, 1.286718e+10, 1.277663e+10, 
    1.267899e+10, 1.257453e+10, 1.246355e+10, 1.234634e+10, 1.222321e+10, 
    1.209449e+10, 1.19605e+10, 1.182158e+10, 1.167804e+10, 1.153025e+10, 
    1.137852e+10, 1.12232e+10, 1.106461e+10, 1.090309e+10, 1.073895e+10, 
    1.057252e+10, 1.040409e+10, 1.023397e+10, 1.006244e+10, 9.88979e+09, 
    9.716282e+09, 9.542177e+09, 9.367718e+09, 9.193139e+09, 9.018663e+09, 
    8.844498e+09, 8.670843e+09, 8.497883e+09, 8.32579e+09, 8.154726e+09, 
    7.984841e+09, 7.816271e+09, 7.649145e+09, 7.483577e+09, 7.319673e+09, 
    7.157529e+09,
  7.155078e+09, 7.316969e+09, 7.480609e+09, 7.645901e+09, 7.812741e+09, 
    7.981012e+09, 8.150589e+09, 8.321333e+09, 8.493095e+09, 8.665715e+09, 
    8.839017e+09, 9.012821e+09, 9.186927e+09, 9.361125e+09, 9.535196e+09, 
    9.708905e+09, 9.882009e+09, 1.005425e+10, 1.022536e+10, 1.039506e+10, 
    1.056306e+10, 1.072907e+10, 1.089278e+10, 1.105388e+10, 1.121203e+10, 
    1.136693e+10, 1.151823e+10, 1.166561e+10, 1.180873e+10, 1.194726e+10, 
    1.208085e+10, 1.220919e+10, 1.233195e+10, 1.24488e+10, 1.255944e+10, 
    1.266358e+10, 1.276091e+10, 1.285118e+10, 1.293411e+10, 1.300948e+10, 
    1.307706e+10, 1.313664e+10, 1.318806e+10, 1.323115e+10, 1.326578e+10, 
    1.329185e+10, 1.330927e+10, 1.3318e+10, 1.3318e+10, 1.330927e+10, 
    1.329185e+10, 1.326578e+10, 1.323115e+10, 1.318806e+10, 1.313664e+10, 
    1.307706e+10, 1.300948e+10, 1.293411e+10, 1.285118e+10, 1.276091e+10, 
    1.266358e+10, 1.255944e+10, 1.24488e+10, 1.233195e+10, 1.220919e+10, 
    1.208085e+10, 1.194726e+10, 1.180873e+10, 1.166561e+10, 1.151823e+10, 
    1.136693e+10, 1.121203e+10, 1.105388e+10, 1.089278e+10, 1.072907e+10, 
    1.056306e+10, 1.039506e+10, 1.022536e+10, 1.005425e+10, 9.882009e+09, 
    9.708905e+09, 9.535196e+09, 9.361125e+09, 9.186927e+09, 9.012821e+09, 
    8.839017e+09, 8.665715e+09, 8.493095e+09, 8.321333e+09, 8.150589e+09, 
    7.981012e+09, 7.812741e+09, 7.645901e+09, 7.480609e+09, 7.316969e+09, 
    7.155078e+09,
  7.151404e+09, 7.312915e+09, 7.476158e+09, 7.641037e+09, 7.807448e+09, 
    7.975273e+09, 8.144387e+09, 8.314652e+09, 8.485919e+09, 8.658028e+09, 
    8.830806e+09, 9.004068e+09, 9.177618e+09, 9.351248e+09, 9.524738e+09, 
    9.697854e+09, 9.870353e+09, 1.004198e+10, 1.021247e+10, 1.038154e+10, 
    1.054891e+10, 1.071428e+10, 1.087735e+10, 1.10378e+10, 1.119532e+10, 
    1.134958e+10, 1.150025e+10, 1.164701e+10, 1.178951e+10, 1.192743e+10, 
    1.206044e+10, 1.218821e+10, 1.231041e+10, 1.242673e+10, 1.253687e+10, 
    1.264052e+10, 1.273739e+10, 1.282723e+10, 1.290977e+10, 1.298478e+10, 
    1.305203e+10, 1.311133e+10, 1.316249e+10, 1.320537e+10, 1.323984e+10, 
    1.326578e+10, 1.328312e+10, 1.32918e+10, 1.32918e+10, 1.328312e+10, 
    1.326578e+10, 1.323984e+10, 1.320537e+10, 1.316249e+10, 1.311133e+10, 
    1.305203e+10, 1.298478e+10, 1.290977e+10, 1.282723e+10, 1.273739e+10, 
    1.264052e+10, 1.253687e+10, 1.242673e+10, 1.231041e+10, 1.218821e+10, 
    1.206044e+10, 1.192743e+10, 1.178951e+10, 1.164701e+10, 1.150025e+10, 
    1.134958e+10, 1.119532e+10, 1.10378e+10, 1.087735e+10, 1.071428e+10, 
    1.054891e+10, 1.038154e+10, 1.021247e+10, 1.004198e+10, 9.870353e+09, 
    9.697854e+09, 9.524738e+09, 9.351248e+09, 9.177618e+09, 9.004068e+09, 
    8.830806e+09, 8.658028e+09, 8.485919e+09, 8.314652e+09, 8.144387e+09, 
    7.975273e+09, 7.807448e+09, 7.641037e+09, 7.476158e+09, 7.312915e+09, 
    7.151404e+09,
  7.146505e+09, 7.307511e+09, 7.470226e+09, 7.634556e+09, 7.800395e+09, 
    7.967627e+09, 8.136126e+09, 8.305754e+09, 8.476363e+09, 8.647793e+09, 
    8.819871e+09, 8.992415e+09, 9.165227e+09, 9.338102e+09, 9.510819e+09, 
    9.683147e+09, 9.854844e+09, 1.002566e+10, 1.019532e+10, 1.036355e+10, 
    1.053008e+10, 1.06946e+10, 1.085682e+10, 1.101642e+10, 1.117309e+10, 
    1.13265e+10, 1.147634e+10, 1.162227e+10, 1.176396e+10, 1.190108e+10, 
    1.203331e+10, 1.216031e+10, 1.228178e+10, 1.23974e+10, 1.250686e+10, 
    1.260987e+10, 1.270614e+10, 1.279542e+10, 1.287743e+10, 1.295196e+10, 
    1.301878e+10, 1.30777e+10, 1.312854e+10, 1.317114e+10, 1.320537e+10, 
    1.323115e+10, 1.324837e+10, 1.3257e+10, 1.3257e+10, 1.324837e+10, 
    1.323115e+10, 1.320537e+10, 1.317114e+10, 1.312854e+10, 1.30777e+10, 
    1.301878e+10, 1.295196e+10, 1.287743e+10, 1.279542e+10, 1.270614e+10, 
    1.260987e+10, 1.250686e+10, 1.23974e+10, 1.228178e+10, 1.216031e+10, 
    1.203331e+10, 1.190108e+10, 1.176396e+10, 1.162227e+10, 1.147634e+10, 
    1.13265e+10, 1.117309e+10, 1.101642e+10, 1.085682e+10, 1.06946e+10, 
    1.053008e+10, 1.036355e+10, 1.019532e+10, 1.002566e+10, 9.854844e+09, 
    9.683147e+09, 9.510819e+09, 9.338102e+09, 9.165227e+09, 8.992415e+09, 
    8.819871e+09, 8.647793e+09, 8.476363e+09, 8.305754e+09, 8.136126e+09, 
    7.967627e+09, 7.800395e+09, 7.634556e+09, 7.470226e+09, 7.307511e+09, 
    7.146505e+09,
  7.140384e+09, 7.30076e+09, 7.462817e+09, 7.626462e+09, 7.791588e+09, 
    7.958081e+09, 8.125813e+09, 8.294647e+09, 8.464436e+09, 8.63502e+09, 
    8.806228e+09, 8.977876e+09, 9.14977e+09, 9.321703e+09, 9.49346e+09, 
    9.664807e+09, 9.835507e+09, 1.00053e+10, 1.017394e+10, 1.034114e+10, 
    1.050662e+10, 1.067009e+10, 1.083124e+10, 1.098979e+10, 1.11454e+10, 
    1.129776e+10, 1.144656e+10, 1.159146e+10, 1.173213e+10, 1.186826e+10, 
    1.199952e+10, 1.212559e+10, 1.224615e+10, 1.236089e+10, 1.246951e+10, 
    1.257172e+10, 1.266725e+10, 1.275582e+10, 1.283719e+10, 1.291113e+10, 
    1.297741e+10, 1.303585e+10, 1.308628e+10, 1.312854e+10, 1.316249e+10, 
    1.318806e+10, 1.320514e+10, 1.32137e+10, 1.32137e+10, 1.320514e+10, 
    1.318806e+10, 1.316249e+10, 1.312854e+10, 1.308628e+10, 1.303585e+10, 
    1.297741e+10, 1.291113e+10, 1.283719e+10, 1.275582e+10, 1.266725e+10, 
    1.257172e+10, 1.246951e+10, 1.236089e+10, 1.224615e+10, 1.212559e+10, 
    1.199952e+10, 1.186826e+10, 1.173213e+10, 1.159146e+10, 1.144656e+10, 
    1.129776e+10, 1.11454e+10, 1.098979e+10, 1.083124e+10, 1.067009e+10, 
    1.050662e+10, 1.034114e+10, 1.017394e+10, 1.00053e+10, 9.835507e+09, 
    9.664807e+09, 9.49346e+09, 9.321703e+09, 9.14977e+09, 8.977876e+09, 
    8.806228e+09, 8.63502e+09, 8.464436e+09, 8.294647e+09, 8.125813e+09, 
    7.958081e+09, 7.791588e+09, 7.626462e+09, 7.462817e+09, 7.30076e+09, 
    7.140384e+09,
  7.133041e+09, 7.292662e+09, 7.453934e+09, 7.616759e+09, 7.781033e+09, 
    7.946641e+09, 8.113456e+09, 8.281342e+09, 8.450151e+09, 8.619724e+09, 
    8.789891e+09, 8.96047e+09, 9.131267e+09, 9.302078e+09, 9.472687e+09, 
    9.642865e+09, 9.812372e+09, 9.980962e+09, 1.014837e+10, 1.031433e+10, 
    1.047856e+10, 1.064077e+10, 1.080067e+10, 1.095795e+10, 1.111231e+10, 
    1.126342e+10, 1.141097e+10, 1.155465e+10, 1.169412e+10, 1.182907e+10, 
    1.195917e+10, 1.208412e+10, 1.220359e+10, 1.231729e+10, 1.242492e+10, 
    1.252618e+10, 1.262082e+10, 1.270856e+10, 1.278916e+10, 1.286239e+10, 
    1.292804e+10, 1.298592e+10, 1.303585e+10, 1.30777e+10, 1.311133e+10, 
    1.313664e+10, 1.315356e+10, 1.316203e+10, 1.316203e+10, 1.315356e+10, 
    1.313664e+10, 1.311133e+10, 1.30777e+10, 1.303585e+10, 1.298592e+10, 
    1.292804e+10, 1.286239e+10, 1.278916e+10, 1.270856e+10, 1.262082e+10, 
    1.252618e+10, 1.242492e+10, 1.231729e+10, 1.220359e+10, 1.208412e+10, 
    1.195917e+10, 1.182907e+10, 1.169412e+10, 1.155465e+10, 1.141097e+10, 
    1.126342e+10, 1.111231e+10, 1.095795e+10, 1.080067e+10, 1.064077e+10, 
    1.047856e+10, 1.031433e+10, 1.014837e+10, 9.980962e+09, 9.812372e+09, 
    9.642865e+09, 9.472687e+09, 9.302078e+09, 9.131267e+09, 8.96047e+09, 
    8.789891e+09, 8.619724e+09, 8.450151e+09, 8.281342e+09, 8.113456e+09, 
    7.946641e+09, 7.781033e+09, 7.616759e+09, 7.453934e+09, 7.292662e+09, 
    7.133041e+09,
  7.124479e+09, 7.283223e+09, 7.443579e+09, 7.605452e+09, 7.768736e+09, 
    7.933316e+09, 8.099066e+09, 8.26585e+09, 8.433522e+09, 8.601922e+09, 
    8.770882e+09, 8.940219e+09, 9.109745e+09, 9.279254e+09, 9.448532e+09, 
    9.617354e+09, 9.785482e+09, 9.95267e+09, 1.011866e+10, 1.028319e+10, 
    1.044597e+10, 1.060673e+10, 1.076517e+10, 1.092099e+10, 1.107389e+10, 
    1.122356e+10, 1.136968e+10, 1.151193e+10, 1.165001e+10, 1.17836e+10, 
    1.191237e+10, 1.203602e+10, 1.215424e+10, 1.226673e+10, 1.237321e+10, 
    1.247338e+10, 1.256699e+10, 1.265377e+10, 1.273348e+10, 1.280589e+10, 
    1.287081e+10, 1.292804e+10, 1.297741e+10, 1.301878e+10, 1.305203e+10, 
    1.307706e+10, 1.309378e+10, 1.310215e+10, 1.310215e+10, 1.309378e+10, 
    1.307706e+10, 1.305203e+10, 1.301878e+10, 1.297741e+10, 1.292804e+10, 
    1.287081e+10, 1.280589e+10, 1.273348e+10, 1.265377e+10, 1.256699e+10, 
    1.247338e+10, 1.237321e+10, 1.226673e+10, 1.215424e+10, 1.203602e+10, 
    1.191237e+10, 1.17836e+10, 1.165001e+10, 1.151193e+10, 1.136968e+10, 
    1.122356e+10, 1.107389e+10, 1.092099e+10, 1.076517e+10, 1.060673e+10, 
    1.044597e+10, 1.028319e+10, 1.011866e+10, 9.95267e+09, 9.785482e+09, 
    9.617354e+09, 9.448532e+09, 9.279254e+09, 9.109745e+09, 8.940219e+09, 
    8.770882e+09, 8.601922e+09, 8.433522e+09, 8.26585e+09, 8.099066e+09, 
    7.933316e+09, 7.768736e+09, 7.605452e+09, 7.443579e+09, 7.283223e+09, 
    7.124479e+09,
  7.1147e+09, 7.272444e+09, 7.431758e+09, 7.592547e+09, 7.754704e+09, 
    7.918115e+09, 8.082655e+09, 8.248187e+09, 8.414565e+09, 8.581632e+09, 
    8.749221e+09, 8.917151e+09, 9.085231e+09, 9.253263e+09, 9.421031e+09, 
    9.588315e+09, 9.754878e+09, 9.920478e+09, 1.008486e+10, 1.024776e+10, 
    1.040891e+10, 1.056802e+10, 1.07248e+10, 1.087898e+10, 1.103023e+10, 
    1.117826e+10, 1.132276e+10, 1.146341e+10, 1.159992e+10, 1.173195e+10, 
    1.185922e+10, 1.198141e+10, 1.209821e+10, 1.220935e+10, 1.231452e+10, 
    1.241347e+10, 1.250591e+10, 1.25916e+10, 1.267031e+10, 1.27418e+10, 
    1.280589e+10, 1.286239e+10, 1.291113e+10, 1.295196e+10, 1.298478e+10, 
    1.300948e+10, 1.302599e+10, 1.303425e+10, 1.303425e+10, 1.302599e+10, 
    1.300948e+10, 1.298478e+10, 1.295196e+10, 1.291113e+10, 1.286239e+10, 
    1.280589e+10, 1.27418e+10, 1.267031e+10, 1.25916e+10, 1.250591e+10, 
    1.241347e+10, 1.231452e+10, 1.220935e+10, 1.209821e+10, 1.198141e+10, 
    1.185922e+10, 1.173195e+10, 1.159992e+10, 1.146341e+10, 1.132276e+10, 
    1.117826e+10, 1.103023e+10, 1.087898e+10, 1.07248e+10, 1.056802e+10, 
    1.040891e+10, 1.024776e+10, 1.008486e+10, 9.920478e+09, 9.754878e+09, 
    9.588315e+09, 9.421031e+09, 9.253263e+09, 9.085231e+09, 8.917151e+09, 
    8.749221e+09, 8.581632e+09, 8.414565e+09, 8.248187e+09, 8.082655e+09, 
    7.918115e+09, 7.754704e+09, 7.592547e+09, 7.431758e+09, 7.272444e+09, 
    7.1147e+09,
  7.103705e+09, 7.260329e+09, 7.418477e+09, 7.578052e+09, 7.738948e+09, 
    7.901051e+09, 8.064236e+09, 8.228367e+09, 8.3933e+09, 8.558878e+09, 
    8.724934e+09, 8.891291e+09, 9.05776e+09, 9.224142e+09, 9.390226e+09, 
    9.555794e+09, 9.720613e+09, 9.884442e+09, 1.004703e+10, 1.020812e+10, 
    1.036744e+10, 1.052472e+10, 1.067967e+10, 1.0832e+10, 1.098142e+10, 
    1.112763e+10, 1.127033e+10, 1.14092e+10, 1.154395e+10, 1.167428e+10, 
    1.179987e+10, 1.192043e+10, 1.203567e+10, 1.214529e+10, 1.224902e+10, 
    1.234659e+10, 1.243775e+10, 1.252223e+10, 1.259983e+10, 1.267031e+10, 
    1.273348e+10, 1.278916e+10, 1.283719e+10, 1.287743e+10, 1.290977e+10, 
    1.293411e+10, 1.295038e+10, 1.295852e+10, 1.295852e+10, 1.295038e+10, 
    1.293411e+10, 1.290977e+10, 1.287743e+10, 1.283719e+10, 1.278916e+10, 
    1.273348e+10, 1.267031e+10, 1.259983e+10, 1.252223e+10, 1.243775e+10, 
    1.234659e+10, 1.224902e+10, 1.214529e+10, 1.203567e+10, 1.192043e+10, 
    1.179987e+10, 1.167428e+10, 1.154395e+10, 1.14092e+10, 1.127033e+10, 
    1.112763e+10, 1.098142e+10, 1.0832e+10, 1.067967e+10, 1.052472e+10, 
    1.036744e+10, 1.020812e+10, 1.004703e+10, 9.884442e+09, 9.720613e+09, 
    9.555794e+09, 9.390226e+09, 9.224142e+09, 9.05776e+09, 8.891291e+09, 
    8.724934e+09, 8.558878e+09, 8.3933e+09, 8.228367e+09, 8.064236e+09, 
    7.901051e+09, 7.738948e+09, 7.578052e+09, 7.418477e+09, 7.260329e+09, 
    7.103705e+09,
  7.091497e+09, 7.246883e+09, 7.403741e+09, 7.561974e+09, 7.721477e+09, 
    7.882135e+09, 8.043825e+09, 8.20641e+09, 8.369748e+09, 8.533684e+09, 
    8.698051e+09, 8.862674e+09, 9.027367e+09, 9.191932e+09, 9.356163e+09, 
    9.519842e+09, 9.68274e+09, 9.844622e+09, 1.000524e+10, 1.016434e+10, 
    1.032166e+10, 1.047692e+10, 1.062985e+10, 1.078017e+10, 1.092757e+10, 
    1.107179e+10, 1.12125e+10, 1.134943e+10, 1.148226e+10, 1.16107e+10, 
    1.173446e+10, 1.185324e+10, 1.196675e+10, 1.207473e+10, 1.217688e+10, 
    1.227295e+10, 1.236269e+10, 1.244586e+10, 1.252223e+10, 1.25916e+10, 
    1.265377e+10, 1.270856e+10, 1.275582e+10, 1.279542e+10, 1.282723e+10, 
    1.285118e+10, 1.286718e+10, 1.287519e+10, 1.287519e+10, 1.286718e+10, 
    1.285118e+10, 1.282723e+10, 1.279542e+10, 1.275582e+10, 1.270856e+10, 
    1.265377e+10, 1.25916e+10, 1.252223e+10, 1.244586e+10, 1.236269e+10, 
    1.227295e+10, 1.217688e+10, 1.207473e+10, 1.196675e+10, 1.185324e+10, 
    1.173446e+10, 1.16107e+10, 1.148226e+10, 1.134943e+10, 1.12125e+10, 
    1.107179e+10, 1.092757e+10, 1.078017e+10, 1.062985e+10, 1.047692e+10, 
    1.032166e+10, 1.016434e+10, 1.000524e+10, 9.844622e+09, 9.68274e+09, 
    9.519842e+09, 9.356163e+09, 9.191932e+09, 9.027367e+09, 8.862674e+09, 
    8.698051e+09, 8.533684e+09, 8.369748e+09, 8.20641e+09, 8.043825e+09, 
    7.882135e+09, 7.721477e+09, 7.561974e+09, 7.403741e+09, 7.246883e+09, 
    7.091497e+09,
  7.078078e+09, 7.23211e+09, 7.387556e+09, 7.544322e+09, 7.702302e+09, 
    7.861382e+09, 8.021437e+09, 8.182336e+09, 8.343933e+09, 8.506077e+09, 
    8.668601e+09, 8.831335e+09, 8.994092e+09, 9.156679e+09, 9.318892e+09, 
    9.480515e+09, 9.641325e+09, 9.801088e+09, 9.959563e+09, 1.01165e+10, 
    1.027164e+10, 1.042471e+10, 1.057545e+10, 1.072358e+10, 1.08688e+10, 
    1.101085e+10, 1.114942e+10, 1.128423e+10, 1.141498e+10, 1.154138e+10, 
    1.166315e+10, 1.178001e+10, 1.189166e+10, 1.199784e+10, 1.209829e+10, 
    1.219274e+10, 1.228095e+10, 1.236269e+10, 1.243775e+10, 1.250591e+10, 
    1.256699e+10, 1.262082e+10, 1.266725e+10, 1.270614e+10, 1.273739e+10, 
    1.276091e+10, 1.277663e+10, 1.27845e+10, 1.27845e+10, 1.277663e+10, 
    1.276091e+10, 1.273739e+10, 1.270614e+10, 1.266725e+10, 1.262082e+10, 
    1.256699e+10, 1.250591e+10, 1.243775e+10, 1.236269e+10, 1.228095e+10, 
    1.219274e+10, 1.209829e+10, 1.199784e+10, 1.189166e+10, 1.178001e+10, 
    1.166315e+10, 1.154138e+10, 1.141498e+10, 1.128423e+10, 1.114942e+10, 
    1.101085e+10, 1.08688e+10, 1.072358e+10, 1.057545e+10, 1.042471e+10, 
    1.027164e+10, 1.01165e+10, 9.959563e+09, 9.801088e+09, 9.641325e+09, 
    9.480515e+09, 9.318892e+09, 9.156679e+09, 8.994092e+09, 8.831335e+09, 
    8.668601e+09, 8.506077e+09, 8.343933e+09, 8.182336e+09, 8.021437e+09, 
    7.861382e+09, 7.702302e+09, 7.544322e+09, 7.387556e+09, 7.23211e+09, 
    7.078078e+09,
  7.063453e+09, 7.216014e+09, 7.36993e+09, 7.525106e+09, 7.681435e+09, 
    7.838806e+09, 7.997093e+09, 8.156166e+09, 8.31588e+09, 8.476086e+09, 
    8.636621e+09, 8.797313e+09, 8.95798e+09, 9.118431e+09, 9.278465e+09, 
    9.437871e+09, 9.596429e+09, 9.753911e+09, 9.910078e+09, 1.006469e+10, 
    1.021748e+10, 1.03682e+10, 1.051658e+10, 1.066235e+10, 1.080523e+10, 
    1.094495e+10, 1.108122e+10, 1.121375e+10, 1.134227e+10, 1.146649e+10, 
    1.158613e+10, 1.170091e+10, 1.181057e+10, 1.191483e+10, 1.201345e+10, 
    1.210616e+10, 1.219274e+10, 1.227295e+10, 1.234659e+10, 1.241347e+10, 
    1.247338e+10, 1.252618e+10, 1.257172e+10, 1.260987e+10, 1.264052e+10, 
    1.266358e+10, 1.267899e+10, 1.268671e+10, 1.268671e+10, 1.267899e+10, 
    1.266358e+10, 1.264052e+10, 1.260987e+10, 1.257172e+10, 1.252618e+10, 
    1.247338e+10, 1.241347e+10, 1.234659e+10, 1.227295e+10, 1.219274e+10, 
    1.210616e+10, 1.201345e+10, 1.191483e+10, 1.181057e+10, 1.170091e+10, 
    1.158613e+10, 1.146649e+10, 1.134227e+10, 1.121375e+10, 1.108122e+10, 
    1.094495e+10, 1.080523e+10, 1.066235e+10, 1.051658e+10, 1.03682e+10, 
    1.021748e+10, 1.006469e+10, 9.910078e+09, 9.753911e+09, 9.596429e+09, 
    9.437871e+09, 9.278465e+09, 9.118431e+09, 8.95798e+09, 8.797313e+09, 
    8.636621e+09, 8.476086e+09, 8.31588e+09, 8.156166e+09, 7.997093e+09, 
    7.838806e+09, 7.681435e+09, 7.525106e+09, 7.36993e+09, 7.216014e+09, 
    7.063453e+09,
  7.047623e+09, 7.198601e+09, 7.350871e+09, 7.504335e+09, 7.65889e+09, 
    7.814423e+09, 7.970811e+09, 8.127923e+09, 8.285618e+09, 8.443745e+09, 
    8.602145e+09, 8.760649e+09, 8.919077e+09, 9.077242e+09, 9.234944e+09, 
    9.391978e+09, 9.548129e+09, 9.703171e+09, 9.856871e+09, 1.000899e+10, 
    1.015928e+10, 1.030749e+10, 1.045336e+10, 1.059662e+10, 1.0737e+10, 
    1.087423e+10, 1.100805e+10, 1.113816e+10, 1.12643e+10, 1.13862e+10, 
    1.150357e+10, 1.161615e+10, 1.172369e+10, 1.182591e+10, 1.192258e+10, 
    1.201345e+10, 1.209829e+10, 1.217688e+10, 1.224902e+10, 1.231452e+10, 
    1.237321e+10, 1.242492e+10, 1.246951e+10, 1.250686e+10, 1.253687e+10, 
    1.255944e+10, 1.257453e+10, 1.258209e+10, 1.258209e+10, 1.257453e+10, 
    1.255944e+10, 1.253687e+10, 1.250686e+10, 1.246951e+10, 1.242492e+10, 
    1.237321e+10, 1.231452e+10, 1.224902e+10, 1.217688e+10, 1.209829e+10, 
    1.201345e+10, 1.192258e+10, 1.182591e+10, 1.172369e+10, 1.161615e+10, 
    1.150357e+10, 1.13862e+10, 1.12643e+10, 1.113816e+10, 1.100805e+10, 
    1.087423e+10, 1.0737e+10, 1.059662e+10, 1.045336e+10, 1.030749e+10, 
    1.015928e+10, 1.000899e+10, 9.856871e+09, 9.703171e+09, 9.548129e+09, 
    9.391978e+09, 9.234944e+09, 9.077242e+09, 8.919077e+09, 8.760649e+09, 
    8.602145e+09, 8.443745e+09, 8.285618e+09, 8.127923e+09, 7.970811e+09, 
    7.814423e+09, 7.65889e+09, 7.504335e+09, 7.350871e+09, 7.198601e+09, 
    7.047623e+09,
  7.030593e+09, 7.179877e+09, 7.330385e+09, 7.482021e+09, 7.634681e+09, 
    7.788252e+09, 7.942612e+09, 8.097633e+09, 8.253174e+09, 8.409087e+09, 
    8.565214e+09, 8.721389e+09, 8.877434e+09, 9.033167e+09, 9.188391e+09, 
    9.342905e+09, 9.496498e+09, 9.64895e+09, 9.800034e+09, 9.949515e+09, 
    1.009715e+10, 1.02427e+10, 1.03859e+10, 1.05265e+10, 1.066424e+10, 
    1.079885e+10, 1.093007e+10, 1.105763e+10, 1.118125e+10, 1.130069e+10, 
    1.141567e+10, 1.152593e+10, 1.163122e+10, 1.17313e+10, 1.182591e+10, 
    1.191483e+10, 1.199784e+10, 1.207473e+10, 1.214529e+10, 1.220935e+10, 
    1.226673e+10, 1.231729e+10, 1.236089e+10, 1.23974e+10, 1.242673e+10, 
    1.24488e+10, 1.246355e+10, 1.247093e+10, 1.247093e+10, 1.246355e+10, 
    1.24488e+10, 1.242673e+10, 1.23974e+10, 1.236089e+10, 1.231729e+10, 
    1.226673e+10, 1.220935e+10, 1.214529e+10, 1.207473e+10, 1.199784e+10, 
    1.191483e+10, 1.182591e+10, 1.17313e+10, 1.163122e+10, 1.152593e+10, 
    1.141567e+10, 1.130069e+10, 1.118125e+10, 1.105763e+10, 1.093007e+10, 
    1.079885e+10, 1.066424e+10, 1.05265e+10, 1.03859e+10, 1.02427e+10, 
    1.009715e+10, 9.949515e+09, 9.800034e+09, 9.64895e+09, 9.496498e+09, 
    9.342905e+09, 9.188391e+09, 9.033167e+09, 8.877434e+09, 8.721389e+09, 
    8.565214e+09, 8.409087e+09, 8.253174e+09, 8.097633e+09, 7.942612e+09, 
    7.788252e+09, 7.634681e+09, 7.482021e+09, 7.330385e+09, 7.179877e+09, 
    7.030593e+09,
  7.012366e+09, 7.159848e+09, 7.308484e+09, 7.458176e+09, 7.608822e+09, 
    7.760311e+09, 7.912521e+09, 8.065324e+09, 8.218582e+09, 8.372148e+09, 
    8.525868e+09, 8.679578e+09, 8.833104e+09, 8.986266e+09, 9.138871e+09, 
    9.290724e+09, 9.441618e+09, 9.591338e+09, 9.739662e+09, 9.886363e+09, 
    1.00312e+10, 1.017395e+10, 1.031435e+10, 1.045215e+10, 1.058711e+10, 
    1.071896e+10, 1.084745e+10, 1.097232e+10, 1.109331e+10, 1.121017e+10, 
    1.132264e+10, 1.143046e+10, 1.153341e+10, 1.163122e+10, 1.172369e+10, 
    1.181057e+10, 1.189166e+10, 1.196675e+10, 1.203567e+10, 1.209821e+10, 
    1.215424e+10, 1.220359e+10, 1.224615e+10, 1.228178e+10, 1.231041e+10, 
    1.233195e+10, 1.234634e+10, 1.235355e+10, 1.235355e+10, 1.234634e+10, 
    1.233195e+10, 1.231041e+10, 1.228178e+10, 1.224615e+10, 1.220359e+10, 
    1.215424e+10, 1.209821e+10, 1.203567e+10, 1.196675e+10, 1.189166e+10, 
    1.181057e+10, 1.172369e+10, 1.163122e+10, 1.153341e+10, 1.143046e+10, 
    1.132264e+10, 1.121017e+10, 1.109331e+10, 1.097232e+10, 1.084745e+10, 
    1.071896e+10, 1.058711e+10, 1.045215e+10, 1.031435e+10, 1.017395e+10, 
    1.00312e+10, 9.886363e+09, 9.739662e+09, 9.591338e+09, 9.441618e+09, 
    9.290724e+09, 9.138871e+09, 8.986266e+09, 8.833104e+09, 8.679578e+09, 
    8.525868e+09, 8.372148e+09, 8.218582e+09, 8.065324e+09, 7.912521e+09, 
    7.760311e+09, 7.608822e+09, 7.458176e+09, 7.308484e+09, 7.159848e+09, 
    7.012366e+09,
  6.992947e+09, 7.138521e+09, 7.285175e+09, 7.432813e+09, 7.581331e+09, 
    7.73062e+09, 7.880559e+09, 8.031022e+09, 8.181873e+09, 8.332967e+09, 
    8.484152e+09, 8.635267e+09, 8.786142e+09, 8.936601e+09, 9.086456e+09, 
    9.235513e+09, 9.383574e+09, 9.530426e+09, 9.675857e+09, 9.819643e+09, 
    9.961556e+09, 1.010136e+10, 1.023883e+10, 1.037371e+10, 1.050575e+10, 
    1.063472e+10, 1.076036e+10, 1.088243e+10, 1.100067e+10, 1.111483e+10, 
    1.122468e+10, 1.132997e+10, 1.143046e+10, 1.152593e+10, 1.161615e+10, 
    1.170091e+10, 1.178001e+10, 1.185324e+10, 1.192043e+10, 1.198141e+10, 
    1.203602e+10, 1.208412e+10, 1.212559e+10, 1.216031e+10, 1.218821e+10, 
    1.220919e+10, 1.222321e+10, 1.223023e+10, 1.223023e+10, 1.222321e+10, 
    1.220919e+10, 1.218821e+10, 1.216031e+10, 1.212559e+10, 1.208412e+10, 
    1.203602e+10, 1.198141e+10, 1.192043e+10, 1.185324e+10, 1.178001e+10, 
    1.170091e+10, 1.161615e+10, 1.152593e+10, 1.143046e+10, 1.132997e+10, 
    1.122468e+10, 1.111483e+10, 1.100067e+10, 1.088243e+10, 1.076036e+10, 
    1.063472e+10, 1.050575e+10, 1.037371e+10, 1.023883e+10, 1.010136e+10, 
    9.961556e+09, 9.819643e+09, 9.675857e+09, 9.530426e+09, 9.383574e+09, 
    9.235513e+09, 9.086456e+09, 8.936601e+09, 8.786142e+09, 8.635267e+09, 
    8.484152e+09, 8.332967e+09, 8.181873e+09, 8.031022e+09, 7.880559e+09, 
    7.73062e+09, 7.581331e+09, 7.432813e+09, 7.285175e+09, 7.138521e+09, 
    6.992947e+09,
  6.972339e+09, 7.115902e+09, 7.260469e+09, 7.405943e+09, 7.552224e+09, 
    7.699199e+09, 7.846753e+09, 7.994759e+09, 8.143084e+09, 8.291585e+09, 
    8.440113e+09, 8.58851e+09, 8.736609e+09, 8.884238e+09, 9.031216e+09, 
    9.177352e+09, 9.322452e+09, 9.466312e+09, 9.608722e+09, 9.749469e+09, 
    9.88833e+09, 1.002508e+10, 1.015949e+10, 1.029132e+10, 1.042034e+10, 
    1.054631e+10, 1.066899e+10, 1.078814e+10, 1.090352e+10, 1.10149e+10, 
    1.112203e+10, 1.122468e+10, 1.132264e+10, 1.141567e+10, 1.150357e+10, 
    1.158613e+10, 1.166315e+10, 1.173446e+10, 1.179987e+10, 1.185922e+10, 
    1.191237e+10, 1.195917e+10, 1.199952e+10, 1.203331e+10, 1.206044e+10, 
    1.208085e+10, 1.209449e+10, 1.210132e+10, 1.210132e+10, 1.209449e+10, 
    1.208085e+10, 1.206044e+10, 1.203331e+10, 1.199952e+10, 1.195917e+10, 
    1.191237e+10, 1.185922e+10, 1.179987e+10, 1.173446e+10, 1.166315e+10, 
    1.158613e+10, 1.150357e+10, 1.141567e+10, 1.132264e+10, 1.122468e+10, 
    1.112203e+10, 1.10149e+10, 1.090352e+10, 1.078814e+10, 1.066899e+10, 
    1.054631e+10, 1.042034e+10, 1.029132e+10, 1.015949e+10, 1.002508e+10, 
    9.88833e+09, 9.749469e+09, 9.608722e+09, 9.466312e+09, 9.322452e+09, 
    9.177352e+09, 9.031216e+09, 8.884238e+09, 8.736609e+09, 8.58851e+09, 
    8.440113e+09, 8.291585e+09, 8.143084e+09, 7.994759e+09, 7.846753e+09, 
    7.699199e+09, 7.552224e+09, 7.405943e+09, 7.260469e+09, 7.115902e+09, 
    6.972339e+09,
  6.950547e+09, 7.092e+09, 7.234377e+09, 7.377583e+09, 7.521518e+09, 
    7.666072e+09, 7.811129e+09, 7.956566e+09, 8.10225e+09, 8.248043e+09, 
    8.393798e+09, 8.539359e+09, 8.684566e+09, 8.829247e+09, 8.973229e+09, 
    9.116325e+09, 9.258346e+09, 9.399095e+09, 9.53837e+09, 9.67596e+09, 
    9.811654e+09, 9.945231e+09, 1.007647e+10, 1.020515e+10, 1.033104e+10, 
    1.045391e+10, 1.057352e+10, 1.068966e+10, 1.080209e+10, 1.091057e+10, 
    1.10149e+10, 1.111483e+10, 1.121017e+10, 1.130069e+10, 1.13862e+10, 
    1.146649e+10, 1.154138e+10, 1.16107e+10, 1.167428e+10, 1.173195e+10, 
    1.17836e+10, 1.182907e+10, 1.186826e+10, 1.190108e+10, 1.192743e+10, 
    1.194726e+10, 1.19605e+10, 1.196713e+10, 1.196713e+10, 1.19605e+10, 
    1.194726e+10, 1.192743e+10, 1.190108e+10, 1.186826e+10, 1.182907e+10, 
    1.17836e+10, 1.173195e+10, 1.167428e+10, 1.16107e+10, 1.154138e+10, 
    1.146649e+10, 1.13862e+10, 1.130069e+10, 1.121017e+10, 1.111483e+10, 
    1.10149e+10, 1.091057e+10, 1.080209e+10, 1.068966e+10, 1.057352e+10, 
    1.045391e+10, 1.033104e+10, 1.020515e+10, 1.007647e+10, 9.945231e+09, 
    9.811654e+09, 9.67596e+09, 9.53837e+09, 9.399095e+09, 9.258346e+09, 
    9.116325e+09, 8.973229e+09, 8.829247e+09, 8.684566e+09, 8.539359e+09, 
    8.393798e+09, 8.248043e+09, 8.10225e+09, 7.956566e+09, 7.811129e+09, 
    7.666072e+09, 7.521518e+09, 7.377583e+09, 7.234377e+09, 7.092e+09, 
    6.950547e+09,
  6.927576e+09, 7.066821e+09, 7.206909e+09, 7.347746e+09, 7.489233e+09, 
    7.631261e+09, 7.773715e+09, 7.916475e+09, 8.059411e+09, 8.202386e+09, 
    8.345257e+09, 8.487873e+09, 8.630074e+09, 8.771699e+09, 8.912572e+09, 
    9.052518e+09, 9.191351e+09, 9.32888e+09, 9.464909e+09, 9.599237e+09, 
    9.731658e+09, 9.861961e+09, 9.989933e+09, 1.011536e+10, 1.023802e+10, 
    1.035769e+10, 1.047415e+10, 1.058718e+10, 1.069657e+10, 1.080209e+10, 
    1.090352e+10, 1.100067e+10, 1.109331e+10, 1.118125e+10, 1.12643e+10, 
    1.134227e+10, 1.141498e+10, 1.148226e+10, 1.154395e+10, 1.159992e+10, 
    1.165001e+10, 1.169412e+10, 1.173213e+10, 1.176396e+10, 1.178951e+10, 
    1.180873e+10, 1.182158e+10, 1.1828e+10, 1.1828e+10, 1.182158e+10, 
    1.180873e+10, 1.178951e+10, 1.176396e+10, 1.173213e+10, 1.169412e+10, 
    1.165001e+10, 1.159992e+10, 1.154395e+10, 1.148226e+10, 1.141498e+10, 
    1.134227e+10, 1.12643e+10, 1.118125e+10, 1.109331e+10, 1.100067e+10, 
    1.090352e+10, 1.080209e+10, 1.069657e+10, 1.058718e+10, 1.047415e+10, 
    1.035769e+10, 1.023802e+10, 1.011536e+10, 9.989933e+09, 9.861961e+09, 
    9.731658e+09, 9.599237e+09, 9.464909e+09, 9.32888e+09, 9.191351e+09, 
    9.052518e+09, 8.912572e+09, 8.771699e+09, 8.630074e+09, 8.487873e+09, 
    8.345257e+09, 8.202386e+09, 8.059411e+09, 7.916475e+09, 7.773715e+09, 
    7.631261e+09, 7.489233e+09, 7.347746e+09, 7.206909e+09, 7.066821e+09, 
    6.927576e+09,
  6.903431e+09, 7.040374e+09, 7.178077e+09, 7.316448e+09, 7.455388e+09, 
    7.594789e+09, 7.734541e+09, 7.874522e+09, 8.014606e+09, 8.15466e+09, 
    8.294543e+09, 8.434108e+09, 8.573202e+09, 8.711665e+09, 8.849328e+09, 
    8.986021e+09, 9.121564e+09, 9.255772e+09, 9.388457e+09, 9.519426e+09, 
    9.648477e+09, 9.775411e+09, 9.900023e+09, 1.00221e+10, 1.014144e+10, 
    1.025783e+10, 1.037106e+10, 1.048091e+10, 1.058718e+10, 1.068966e+10, 
    1.078814e+10, 1.088243e+10, 1.097232e+10, 1.105763e+10, 1.113816e+10, 
    1.121375e+10, 1.128423e+10, 1.134943e+10, 1.14092e+10, 1.146341e+10, 
    1.151193e+10, 1.155465e+10, 1.159146e+10, 1.162227e+10, 1.164701e+10, 
    1.166561e+10, 1.167804e+10, 1.168427e+10, 1.168427e+10, 1.167804e+10, 
    1.166561e+10, 1.164701e+10, 1.162227e+10, 1.159146e+10, 1.155465e+10, 
    1.151193e+10, 1.146341e+10, 1.14092e+10, 1.134943e+10, 1.128423e+10, 
    1.121375e+10, 1.113816e+10, 1.105763e+10, 1.097232e+10, 1.088243e+10, 
    1.078814e+10, 1.068966e+10, 1.058718e+10, 1.048091e+10, 1.037106e+10, 
    1.025783e+10, 1.014144e+10, 1.00221e+10, 9.900023e+09, 9.775411e+09, 
    9.648477e+09, 9.519426e+09, 9.388457e+09, 9.255772e+09, 9.121564e+09, 
    8.986021e+09, 8.849328e+09, 8.711665e+09, 8.573202e+09, 8.434108e+09, 
    8.294543e+09, 8.15466e+09, 8.014606e+09, 7.874522e+09, 7.734541e+09, 
    7.594789e+09, 7.455388e+09, 7.316448e+09, 7.178077e+09, 7.040374e+09, 
    6.903431e+09,
  6.878117e+09, 7.012667e+09, 7.147894e+09, 7.283705e+09, 7.420003e+09, 
    7.556683e+09, 7.693634e+09, 7.830739e+09, 7.967875e+09, 8.10491e+09, 
    8.241709e+09, 8.378128e+09, 8.514017e+09, 8.649221e+09, 8.78358e+09, 
    8.916924e+09, 9.049084e+09, 9.17988e+09, 9.309132e+09, 9.436652e+09, 
    9.562249e+09, 9.68573e+09, 9.806899e+09, 9.925557e+09, 1.00415e+10, 
    1.015454e+10, 1.026446e+10, 1.037106e+10, 1.047415e+10, 1.057352e+10, 
    1.066899e+10, 1.076036e+10, 1.084745e+10, 1.093007e+10, 1.100805e+10, 
    1.108122e+10, 1.114942e+10, 1.12125e+10, 1.127033e+10, 1.132276e+10, 
    1.136968e+10, 1.141097e+10, 1.144656e+10, 1.147634e+10, 1.150025e+10, 
    1.151823e+10, 1.153025e+10, 1.153626e+10, 1.153626e+10, 1.153025e+10, 
    1.151823e+10, 1.150025e+10, 1.147634e+10, 1.144656e+10, 1.141097e+10, 
    1.136968e+10, 1.132276e+10, 1.127033e+10, 1.12125e+10, 1.114942e+10, 
    1.108122e+10, 1.100805e+10, 1.093007e+10, 1.084745e+10, 1.076036e+10, 
    1.066899e+10, 1.057352e+10, 1.047415e+10, 1.037106e+10, 1.026446e+10, 
    1.015454e+10, 1.00415e+10, 9.925557e+09, 9.806899e+09, 9.68573e+09, 
    9.562249e+09, 9.436652e+09, 9.309132e+09, 9.17988e+09, 9.049084e+09, 
    8.916924e+09, 8.78358e+09, 8.649221e+09, 8.514017e+09, 8.378128e+09, 
    8.241709e+09, 8.10491e+09, 7.967875e+09, 7.830739e+09, 7.693634e+09, 
    7.556683e+09, 7.420003e+09, 7.283705e+09, 7.147894e+09, 7.012667e+09, 
    6.878117e+09,
  6.851641e+09, 6.98371e+09, 7.116371e+09, 7.249533e+09, 7.383099e+09, 
    7.516966e+09, 7.651027e+09, 7.785166e+09, 7.919261e+09, 8.053188e+09, 
    8.186811e+09, 8.319992e+09, 8.452588e+09, 8.584445e+09, 8.715411e+09, 
    8.845323e+09, 8.974015e+09, 9.101317e+09, 9.227054e+09, 9.351046e+09, 
    9.473112e+09, 9.593066e+09, 9.710721e+09, 9.825887e+09, 9.938373e+09, 
    1.004799e+10, 1.015454e+10, 1.025783e+10, 1.035769e+10, 1.045391e+10, 
    1.054631e+10, 1.063472e+10, 1.071896e+10, 1.079885e+10, 1.087423e+10, 
    1.094495e+10, 1.101085e+10, 1.107179e+10, 1.112763e+10, 1.117826e+10, 
    1.122356e+10, 1.126342e+10, 1.129776e+10, 1.13265e+10, 1.134958e+10, 
    1.136693e+10, 1.137852e+10, 1.138432e+10, 1.138432e+10, 1.137852e+10, 
    1.136693e+10, 1.134958e+10, 1.13265e+10, 1.129776e+10, 1.126342e+10, 
    1.122356e+10, 1.117826e+10, 1.112763e+10, 1.107179e+10, 1.101085e+10, 
    1.094495e+10, 1.087423e+10, 1.079885e+10, 1.071896e+10, 1.063472e+10, 
    1.054631e+10, 1.045391e+10, 1.035769e+10, 1.025783e+10, 1.015454e+10, 
    1.004799e+10, 9.938373e+09, 9.825887e+09, 9.710721e+09, 9.593066e+09, 
    9.473112e+09, 9.351046e+09, 9.227054e+09, 9.101317e+09, 8.974015e+09, 
    8.845323e+09, 8.715411e+09, 8.584445e+09, 8.452588e+09, 8.319992e+09, 
    8.186811e+09, 8.053188e+09, 7.919261e+09, 7.785166e+09, 7.651027e+09, 
    7.516966e+09, 7.383099e+09, 7.249533e+09, 7.116371e+09, 6.98371e+09, 
    6.851641e+09,
  6.824007e+09, 6.953512e+09, 7.083523e+09, 7.21395e+09, 7.344698e+09, 
    7.475667e+09, 7.606751e+09, 7.737838e+09, 7.868808e+09, 7.99954e+09, 
    8.129904e+09, 8.259766e+09, 8.388985e+09, 8.517416e+09, 8.64491e+09, 
    8.771312e+09, 8.896461e+09, 9.020195e+09, 9.142345e+09, 9.262742e+09, 
    9.381209e+09, 9.497571e+09, 9.61165e+09, 9.723264e+09, 9.832232e+09, 
    9.938373e+09, 1.00415e+10, 1.014144e+10, 1.023802e+10, 1.033104e+10, 
    1.042034e+10, 1.050575e+10, 1.058711e+10, 1.066424e+10, 1.0737e+10, 
    1.080523e+10, 1.08688e+10, 1.092757e+10, 1.098142e+10, 1.103023e+10, 
    1.107389e+10, 1.111231e+10, 1.11454e+10, 1.117309e+10, 1.119532e+10, 
    1.121203e+10, 1.12232e+10, 1.122879e+10, 1.122879e+10, 1.12232e+10, 
    1.121203e+10, 1.119532e+10, 1.117309e+10, 1.11454e+10, 1.111231e+10, 
    1.107389e+10, 1.103023e+10, 1.098142e+10, 1.092757e+10, 1.08688e+10, 
    1.080523e+10, 1.0737e+10, 1.066424e+10, 1.058711e+10, 1.050575e+10, 
    1.042034e+10, 1.033104e+10, 1.023802e+10, 1.014144e+10, 1.00415e+10, 
    9.938373e+09, 9.832232e+09, 9.723264e+09, 9.61165e+09, 9.497571e+09, 
    9.381209e+09, 9.262742e+09, 9.142345e+09, 9.020195e+09, 8.896461e+09, 
    8.771312e+09, 8.64491e+09, 8.517416e+09, 8.388985e+09, 8.259766e+09, 
    8.129904e+09, 7.99954e+09, 7.868808e+09, 7.737838e+09, 7.606751e+09, 
    7.475667e+09, 7.344698e+09, 7.21395e+09, 7.083523e+09, 6.953512e+09, 
    6.824007e+09,
  6.795221e+09, 6.922081e+09, 7.049361e+09, 7.176973e+09, 7.304823e+09, 
    7.432814e+09, 7.56084e+09, 7.688794e+09, 7.816561e+09, 7.94402e+09, 
    8.071048e+09, 8.197513e+09, 8.323282e+09, 8.448214e+09, 8.572165e+09, 
    8.694987e+09, 8.816526e+09, 8.936627e+09, 9.055129e+09, 9.171869e+09, 
    9.286681e+09, 9.399396e+09, 9.509846e+09, 9.61786e+09, 9.723264e+09, 
    9.825887e+09, 9.925557e+09, 1.00221e+10, 1.011536e+10, 1.020515e+10, 
    1.029132e+10, 1.037371e+10, 1.045215e+10, 1.05265e+10, 1.059662e+10, 
    1.066235e+10, 1.072358e+10, 1.078017e+10, 1.0832e+10, 1.087898e+10, 
    1.092099e+10, 1.095795e+10, 1.098979e+10, 1.101642e+10, 1.10378e+10, 
    1.105388e+10, 1.106461e+10, 1.106999e+10, 1.106999e+10, 1.106461e+10, 
    1.105388e+10, 1.10378e+10, 1.101642e+10, 1.098979e+10, 1.095795e+10, 
    1.092099e+10, 1.087898e+10, 1.0832e+10, 1.078017e+10, 1.072358e+10, 
    1.066235e+10, 1.059662e+10, 1.05265e+10, 1.045215e+10, 1.037371e+10, 
    1.029132e+10, 1.020515e+10, 1.011536e+10, 1.00221e+10, 9.925557e+09, 
    9.825887e+09, 9.723264e+09, 9.61786e+09, 9.509846e+09, 9.399396e+09, 
    9.286681e+09, 9.171869e+09, 9.055129e+09, 8.936627e+09, 8.816526e+09, 
    8.694987e+09, 8.572165e+09, 8.448214e+09, 8.323282e+09, 8.197513e+09, 
    8.071048e+09, 7.94402e+09, 7.816561e+09, 7.688794e+09, 7.56084e+09, 
    7.432814e+09, 7.304823e+09, 7.176973e+09, 7.049361e+09, 6.922081e+09, 
    6.795221e+09,
  6.76529e+09, 6.889429e+09, 7.013901e+09, 7.13862e+09, 7.263496e+09, 
    7.388432e+09, 7.513327e+09, 7.638074e+09, 7.762563e+09, 7.886679e+09, 
    8.010299e+09, 8.133301e+09, 8.255552e+09, 8.37692e+09, 8.497266e+09, 
    8.616447e+09, 8.734319e+09, 8.85073e+09, 8.96553e+09, 9.078562e+09, 
    9.18967e+09, 9.298694e+09, 9.405474e+09, 9.509846e+09, 9.61165e+09, 
    9.710721e+09, 9.806899e+09, 9.900023e+09, 9.989933e+09, 1.007647e+10, 
    1.015949e+10, 1.023883e+10, 1.031435e+10, 1.03859e+10, 1.045336e+10, 
    1.051658e+10, 1.057545e+10, 1.062985e+10, 1.067967e+10, 1.07248e+10, 
    1.076517e+10, 1.080067e+10, 1.083124e+10, 1.085682e+10, 1.087735e+10, 
    1.089278e+10, 1.090309e+10, 1.090825e+10, 1.090825e+10, 1.090309e+10, 
    1.089278e+10, 1.087735e+10, 1.085682e+10, 1.083124e+10, 1.080067e+10, 
    1.076517e+10, 1.07248e+10, 1.067967e+10, 1.062985e+10, 1.057545e+10, 
    1.051658e+10, 1.045336e+10, 1.03859e+10, 1.031435e+10, 1.023883e+10, 
    1.015949e+10, 1.007647e+10, 9.989933e+09, 9.900023e+09, 9.806899e+09, 
    9.710721e+09, 9.61165e+09, 9.509846e+09, 9.405474e+09, 9.298694e+09, 
    9.18967e+09, 9.078562e+09, 8.96553e+09, 8.85073e+09, 8.734319e+09, 
    8.616447e+09, 8.497266e+09, 8.37692e+09, 8.255552e+09, 8.133301e+09, 
    8.010299e+09, 7.886679e+09, 7.762563e+09, 7.638074e+09, 7.513327e+09, 
    7.388432e+09, 7.263496e+09, 7.13862e+09, 7.013901e+09, 6.889429e+09, 
    6.76529e+09,
  6.734221e+09, 6.855565e+09, 6.977157e+09, 7.098912e+09, 7.220742e+09, 
    7.342552e+09, 7.464245e+09, 7.585717e+09, 7.706863e+09, 7.827569e+09, 
    7.94772e+09, 8.067195e+09, 8.18587e+09, 8.303616e+09, 8.420301e+09, 
    8.53579e+09, 8.649944e+09, 8.762619e+09, 8.873673e+09, 8.982957e+09, 
    9.090322e+09, 9.195619e+09, 9.298694e+09, 9.399396e+09, 9.497571e+09, 
    9.593066e+09, 9.68573e+09, 9.775411e+09, 9.861961e+09, 9.945231e+09, 
    1.002508e+10, 1.010136e+10, 1.017395e+10, 1.02427e+10, 1.030749e+10, 
    1.03682e+10, 1.042471e+10, 1.047692e+10, 1.052472e+10, 1.056802e+10, 
    1.060673e+10, 1.064077e+10, 1.067009e+10, 1.06946e+10, 1.071428e+10, 
    1.072907e+10, 1.073895e+10, 1.07439e+10, 1.07439e+10, 1.073895e+10, 
    1.072907e+10, 1.071428e+10, 1.06946e+10, 1.067009e+10, 1.064077e+10, 
    1.060673e+10, 1.056802e+10, 1.052472e+10, 1.047692e+10, 1.042471e+10, 
    1.03682e+10, 1.030749e+10, 1.02427e+10, 1.017395e+10, 1.010136e+10, 
    1.002508e+10, 9.945231e+09, 9.861961e+09, 9.775411e+09, 9.68573e+09, 
    9.593066e+09, 9.497571e+09, 9.399396e+09, 9.298694e+09, 9.195619e+09, 
    9.090322e+09, 8.982957e+09, 8.873673e+09, 8.762619e+09, 8.649944e+09, 
    8.53579e+09, 8.420301e+09, 8.303616e+09, 8.18587e+09, 8.067195e+09, 
    7.94772e+09, 7.827569e+09, 7.706863e+09, 7.585717e+09, 7.464245e+09, 
    7.342552e+09, 7.220742e+09, 7.098912e+09, 6.977157e+09, 6.855565e+09, 
    6.734221e+09,
  6.702019e+09, 6.8205e+09, 6.939143e+09, 7.057866e+09, 7.176583e+09, 
    7.295202e+09, 7.41363e+09, 7.531766e+09, 7.649507e+09, 7.766745e+09, 
    7.883369e+09, 7.999264e+09, 8.11431e+09, 8.228386e+09, 8.341364e+09, 
    8.453116e+09, 8.563511e+09, 8.672412e+09, 8.779684e+09, 8.885187e+09, 
    8.988781e+09, 9.090322e+09, 9.18967e+09, 9.286681e+09, 9.381209e+09, 
    9.473112e+09, 9.562249e+09, 9.648477e+09, 9.731658e+09, 9.811654e+09, 
    9.88833e+09, 9.961556e+09, 1.00312e+10, 1.009715e+10, 1.015928e+10, 
    1.021748e+10, 1.027164e+10, 1.032166e+10, 1.036744e+10, 1.040891e+10, 
    1.044597e+10, 1.047856e+10, 1.050662e+10, 1.053008e+10, 1.054891e+10, 
    1.056306e+10, 1.057252e+10, 1.057725e+10, 1.057725e+10, 1.057252e+10, 
    1.056306e+10, 1.054891e+10, 1.053008e+10, 1.050662e+10, 1.047856e+10, 
    1.044597e+10, 1.040891e+10, 1.036744e+10, 1.032166e+10, 1.027164e+10, 
    1.021748e+10, 1.015928e+10, 1.009715e+10, 1.00312e+10, 9.961556e+09, 
    9.88833e+09, 9.811654e+09, 9.731658e+09, 9.648477e+09, 9.562249e+09, 
    9.473112e+09, 9.381209e+09, 9.286681e+09, 9.18967e+09, 9.090322e+09, 
    8.988781e+09, 8.885187e+09, 8.779684e+09, 8.672412e+09, 8.563511e+09, 
    8.453116e+09, 8.341364e+09, 8.228386e+09, 8.11431e+09, 7.999264e+09, 
    7.883369e+09, 7.766745e+09, 7.649507e+09, 7.531766e+09, 7.41363e+09, 
    7.295202e+09, 7.176583e+09, 7.057866e+09, 6.939143e+09, 6.8205e+09, 
    6.702019e+09,
  6.668692e+09, 6.784244e+09, 6.899874e+09, 7.015503e+09, 7.131045e+09, 
    7.246414e+09, 7.361518e+09, 7.47626e+09, 7.590542e+09, 7.704261e+09, 
    7.817309e+09, 7.929576e+09, 8.04095e+09, 8.151313e+09, 8.260545e+09, 
    8.368525e+09, 8.475127e+09, 8.580225e+09, 8.683688e+09, 8.785385e+09, 
    8.885187e+09, 8.982957e+09, 9.078562e+09, 9.171869e+09, 9.262742e+09, 
    9.351046e+09, 9.436652e+09, 9.519426e+09, 9.599237e+09, 9.67596e+09, 
    9.749469e+09, 9.819643e+09, 9.886363e+09, 9.949515e+09, 1.000899e+10, 
    1.006469e+10, 1.01165e+10, 1.016434e+10, 1.020812e+10, 1.024776e+10, 
    1.028319e+10, 1.031433e+10, 1.034114e+10, 1.036355e+10, 1.038154e+10, 
    1.039506e+10, 1.040409e+10, 1.040861e+10, 1.040861e+10, 1.040409e+10, 
    1.039506e+10, 1.038154e+10, 1.036355e+10, 1.034114e+10, 1.031433e+10, 
    1.028319e+10, 1.024776e+10, 1.020812e+10, 1.016434e+10, 1.01165e+10, 
    1.006469e+10, 1.000899e+10, 9.949515e+09, 9.886363e+09, 9.819643e+09, 
    9.749469e+09, 9.67596e+09, 9.599237e+09, 9.519426e+09, 9.436652e+09, 
    9.351046e+09, 9.262742e+09, 9.171869e+09, 9.078562e+09, 8.982957e+09, 
    8.885187e+09, 8.785385e+09, 8.683688e+09, 8.580225e+09, 8.475127e+09, 
    8.368525e+09, 8.260545e+09, 8.151313e+09, 8.04095e+09, 7.929576e+09, 
    7.817309e+09, 7.704261e+09, 7.590542e+09, 7.47626e+09, 7.361518e+09, 
    7.246414e+09, 7.131045e+09, 7.015503e+09, 6.899874e+09, 6.784244e+09, 
    6.668692e+09,
  6.634248e+09, 6.74681e+09, 6.859367e+09, 6.971842e+09, 7.084154e+09, 
    7.196217e+09, 7.307944e+09, 7.419243e+09, 7.530018e+09, 7.640172e+09, 
    7.749601e+09, 7.858201e+09, 7.965864e+09, 8.072481e+09, 8.177936e+09, 
    8.282116e+09, 8.384902e+09, 8.486173e+09, 8.585809e+09, 8.683688e+09, 
    8.779684e+09, 8.873673e+09, 8.96553e+09, 9.055129e+09, 9.142345e+09, 
    9.227054e+09, 9.309132e+09, 9.388457e+09, 9.464909e+09, 9.53837e+09, 
    9.608722e+09, 9.675857e+09, 9.739662e+09, 9.800034e+09, 9.856871e+09, 
    9.910078e+09, 9.959563e+09, 1.000524e+10, 1.004703e+10, 1.008486e+10, 
    1.011866e+10, 1.014837e+10, 1.017394e+10, 1.019532e+10, 1.021247e+10, 
    1.022536e+10, 1.023397e+10, 1.023827e+10, 1.023827e+10, 1.023397e+10, 
    1.022536e+10, 1.021247e+10, 1.019532e+10, 1.017394e+10, 1.014837e+10, 
    1.011866e+10, 1.008486e+10, 1.004703e+10, 1.000524e+10, 9.959563e+09, 
    9.910078e+09, 9.856871e+09, 9.800034e+09, 9.739662e+09, 9.675857e+09, 
    9.608722e+09, 9.53837e+09, 9.464909e+09, 9.388457e+09, 9.309132e+09, 
    9.227054e+09, 9.142345e+09, 9.055129e+09, 8.96553e+09, 8.873673e+09, 
    8.779684e+09, 8.683688e+09, 8.585809e+09, 8.486173e+09, 8.384902e+09, 
    8.282116e+09, 8.177936e+09, 8.072481e+09, 7.965864e+09, 7.858201e+09, 
    7.749601e+09, 7.640172e+09, 7.530018e+09, 7.419243e+09, 7.307944e+09, 
    7.196217e+09, 7.084154e+09, 6.971842e+09, 6.859367e+09, 6.74681e+09, 
    6.634248e+09,
  6.598693e+09, 6.708208e+09, 6.817636e+09, 6.926904e+09, 7.035934e+09, 
    7.144643e+09, 7.252946e+09, 7.360757e+09, 7.467984e+09, 7.574533e+09, 
    7.680307e+09, 7.785207e+09, 7.889131e+09, 7.991974e+09, 8.093629e+09, 
    8.193989e+09, 8.292941e+09, 8.390374e+09, 8.486173e+09, 8.580225e+09, 
    8.672412e+09, 8.762619e+09, 8.85073e+09, 8.936627e+09, 9.020195e+09, 
    9.101317e+09, 9.17988e+09, 9.255772e+09, 9.32888e+09, 9.399095e+09, 
    9.466312e+09, 9.530426e+09, 9.591338e+09, 9.64895e+09, 9.703171e+09, 
    9.753911e+09, 9.801088e+09, 9.844622e+09, 9.884442e+09, 9.920478e+09, 
    9.95267e+09, 9.980962e+09, 1.00053e+10, 1.002566e+10, 1.004198e+10, 
    1.005425e+10, 1.006244e+10, 1.006654e+10, 1.006654e+10, 1.006244e+10, 
    1.005425e+10, 1.004198e+10, 1.002566e+10, 1.00053e+10, 9.980962e+09, 
    9.95267e+09, 9.920478e+09, 9.884442e+09, 9.844622e+09, 9.801088e+09, 
    9.753911e+09, 9.703171e+09, 9.64895e+09, 9.591338e+09, 9.530426e+09, 
    9.466312e+09, 9.399095e+09, 9.32888e+09, 9.255772e+09, 9.17988e+09, 
    9.101317e+09, 9.020195e+09, 8.936627e+09, 8.85073e+09, 8.762619e+09, 
    8.672412e+09, 8.580225e+09, 8.486173e+09, 8.390374e+09, 8.292941e+09, 
    8.193989e+09, 8.093629e+09, 7.991974e+09, 7.889131e+09, 7.785207e+09, 
    7.680307e+09, 7.574533e+09, 7.467984e+09, 7.360757e+09, 7.252946e+09, 
    7.144643e+09, 7.035934e+09, 6.926904e+09, 6.817636e+09, 6.708208e+09, 
    6.598693e+09,
  6.562035e+09, 6.668449e+09, 6.774699e+09, 6.880711e+09, 6.986412e+09, 
    7.091722e+09, 7.196561e+09, 7.300845e+09, 7.404488e+09, 7.5074e+09, 
    7.60949e+09, 7.710664e+09, 7.810825e+09, 7.909876e+09, 8.007716e+09, 
    8.104243e+09, 8.199353e+09, 8.292941e+09, 8.384902e+09, 8.475127e+09, 
    8.563511e+09, 8.649944e+09, 8.734319e+09, 8.816526e+09, 8.896461e+09, 
    8.974015e+09, 9.049084e+09, 9.121564e+09, 9.191351e+09, 9.258346e+09, 
    9.322452e+09, 9.383574e+09, 9.441618e+09, 9.496498e+09, 9.548129e+09, 
    9.596429e+09, 9.641325e+09, 9.68274e+09, 9.720613e+09, 9.754878e+09, 
    9.785482e+09, 9.812372e+09, 9.835507e+09, 9.854844e+09, 9.870353e+09, 
    9.882009e+09, 9.88979e+09, 9.893683e+09, 9.893683e+09, 9.88979e+09, 
    9.882009e+09, 9.870353e+09, 9.854844e+09, 9.835507e+09, 9.812372e+09, 
    9.785482e+09, 9.754878e+09, 9.720613e+09, 9.68274e+09, 9.641325e+09, 
    9.596429e+09, 9.548129e+09, 9.496498e+09, 9.441618e+09, 9.383574e+09, 
    9.322452e+09, 9.258346e+09, 9.191351e+09, 9.121564e+09, 9.049084e+09, 
    8.974015e+09, 8.896461e+09, 8.816526e+09, 8.734319e+09, 8.649944e+09, 
    8.563511e+09, 8.475127e+09, 8.384902e+09, 8.292941e+09, 8.199353e+09, 
    8.104243e+09, 8.007716e+09, 7.909876e+09, 7.810825e+09, 7.710664e+09, 
    7.60949e+09, 7.5074e+09, 7.404488e+09, 7.300845e+09, 7.196561e+09, 
    7.091722e+09, 6.986412e+09, 6.880711e+09, 6.774699e+09, 6.668449e+09, 
    6.562035e+09,
  6.524282e+09, 6.627547e+09, 6.730571e+09, 6.833284e+09, 6.935614e+09, 
    7.037487e+09, 7.138825e+09, 7.23955e+09, 7.339579e+09, 7.438829e+09, 
    7.537212e+09, 7.634641e+09, 7.731025e+09, 7.826271e+09, 7.920287e+09, 
    8.012976e+09, 8.104243e+09, 8.193989e+09, 8.282116e+09, 8.368525e+09, 
    8.453116e+09, 8.53579e+09, 8.616447e+09, 8.694987e+09, 8.771312e+09, 
    8.845323e+09, 8.916924e+09, 8.986021e+09, 9.052518e+09, 9.116325e+09, 
    9.177352e+09, 9.235513e+09, 9.290724e+09, 9.342905e+09, 9.391978e+09, 
    9.437871e+09, 9.480515e+09, 9.519842e+09, 9.555794e+09, 9.588315e+09, 
    9.617354e+09, 9.642865e+09, 9.664807e+09, 9.683147e+09, 9.697854e+09, 
    9.708905e+09, 9.716282e+09, 9.719975e+09, 9.719975e+09, 9.716282e+09, 
    9.708905e+09, 9.697854e+09, 9.683147e+09, 9.664807e+09, 9.642865e+09, 
    9.617354e+09, 9.588315e+09, 9.555794e+09, 9.519842e+09, 9.480515e+09, 
    9.437871e+09, 9.391978e+09, 9.342905e+09, 9.290724e+09, 9.235513e+09, 
    9.177352e+09, 9.116325e+09, 9.052518e+09, 8.986021e+09, 8.916924e+09, 
    8.845323e+09, 8.771312e+09, 8.694987e+09, 8.616447e+09, 8.53579e+09, 
    8.453116e+09, 8.368525e+09, 8.282116e+09, 8.193989e+09, 8.104243e+09, 
    8.012976e+09, 7.920287e+09, 7.826271e+09, 7.731025e+09, 7.634641e+09, 
    7.537212e+09, 7.438829e+09, 7.339579e+09, 7.23955e+09, 7.138825e+09, 
    7.037487e+09, 6.935614e+09, 6.833284e+09, 6.730571e+09, 6.627547e+09, 
    6.524282e+09,
  6.485442e+09, 6.585513e+09, 6.685269e+09, 6.784643e+09, 6.883567e+09, 
    6.981969e+09, 7.079777e+09, 7.176916e+09, 7.273309e+09, 7.368877e+09, 
    7.463537e+09, 7.557208e+09, 7.649805e+09, 7.741242e+09, 7.831433e+09, 
    7.920287e+09, 8.007716e+09, 8.093629e+09, 8.177936e+09, 8.260545e+09, 
    8.341364e+09, 8.420301e+09, 8.497266e+09, 8.572165e+09, 8.64491e+09, 
    8.715411e+09, 8.78358e+09, 8.849328e+09, 8.912572e+09, 8.973229e+09, 
    9.031216e+09, 9.086456e+09, 9.138871e+09, 9.188391e+09, 9.234944e+09, 
    9.278465e+09, 9.318892e+09, 9.356163e+09, 9.390226e+09, 9.421031e+09, 
    9.448532e+09, 9.472687e+09, 9.49346e+09, 9.510819e+09, 9.524738e+09, 
    9.535196e+09, 9.542177e+09, 9.54567e+09, 9.54567e+09, 9.542177e+09, 
    9.535196e+09, 9.524738e+09, 9.510819e+09, 9.49346e+09, 9.472687e+09, 
    9.448532e+09, 9.421031e+09, 9.390226e+09, 9.356163e+09, 9.318892e+09, 
    9.278465e+09, 9.234944e+09, 9.188391e+09, 9.138871e+09, 9.086456e+09, 
    9.031216e+09, 8.973229e+09, 8.912572e+09, 8.849328e+09, 8.78358e+09, 
    8.715411e+09, 8.64491e+09, 8.572165e+09, 8.497266e+09, 8.420301e+09, 
    8.341364e+09, 8.260545e+09, 8.177936e+09, 8.093629e+09, 8.007716e+09, 
    7.920287e+09, 7.831433e+09, 7.741242e+09, 7.649805e+09, 7.557208e+09, 
    7.463537e+09, 7.368877e+09, 7.273309e+09, 7.176916e+09, 7.079777e+09, 
    6.981969e+09, 6.883567e+09, 6.784643e+09, 6.685269e+09, 6.585513e+09, 
    6.485442e+09,
  6.445522e+09, 6.54236e+09, 6.638811e+09, 6.734811e+09, 6.830297e+09, 
    6.925201e+09, 7.019455e+09, 7.112987e+09, 7.205726e+09, 7.297597e+09, 
    7.388526e+09, 7.478433e+09, 7.567242e+09, 7.654872e+09, 7.741242e+09, 
    7.826271e+09, 7.909876e+09, 7.991974e+09, 8.072481e+09, 8.151313e+09, 
    8.228386e+09, 8.303616e+09, 8.37692e+09, 8.448214e+09, 8.517416e+09, 
    8.584445e+09, 8.649221e+09, 8.711665e+09, 8.771699e+09, 8.829247e+09, 
    8.884238e+09, 8.936601e+09, 8.986266e+09, 9.033167e+09, 9.077242e+09, 
    9.118431e+09, 9.156679e+09, 9.191932e+09, 9.224142e+09, 9.253263e+09, 
    9.279254e+09, 9.302078e+09, 9.321703e+09, 9.338102e+09, 9.351248e+09, 
    9.361125e+09, 9.367718e+09, 9.371016e+09, 9.371016e+09, 9.367718e+09, 
    9.361125e+09, 9.351248e+09, 9.338102e+09, 9.321703e+09, 9.302078e+09, 
    9.279254e+09, 9.253263e+09, 9.224142e+09, 9.191932e+09, 9.156679e+09, 
    9.118431e+09, 9.077242e+09, 9.033167e+09, 8.986266e+09, 8.936601e+09, 
    8.884238e+09, 8.829247e+09, 8.771699e+09, 8.711665e+09, 8.649221e+09, 
    8.584445e+09, 8.517416e+09, 8.448214e+09, 8.37692e+09, 8.303616e+09, 
    8.228386e+09, 8.151313e+09, 8.072481e+09, 7.991974e+09, 7.909876e+09, 
    7.826271e+09, 7.741242e+09, 7.654872e+09, 7.567242e+09, 7.478433e+09, 
    7.388526e+09, 7.297597e+09, 7.205726e+09, 7.112987e+09, 7.019455e+09, 
    6.925201e+09, 6.830297e+09, 6.734811e+09, 6.638811e+09, 6.54236e+09, 
    6.445522e+09,
  6.404531e+09, 6.4981e+09, 6.591213e+09, 6.683811e+09, 6.775833e+09, 
    6.867216e+09, 6.957896e+09, 7.047806e+09, 7.136881e+09, 7.225049e+09, 
    7.312241e+09, 7.398386e+09, 7.483411e+09, 7.567242e+09, 7.649805e+09, 
    7.731025e+09, 7.810825e+09, 7.889131e+09, 7.965864e+09, 8.04095e+09, 
    8.11431e+09, 8.18587e+09, 8.255552e+09, 8.323282e+09, 8.388985e+09, 
    8.452588e+09, 8.514017e+09, 8.573202e+09, 8.630074e+09, 8.684566e+09, 
    8.736609e+09, 8.786142e+09, 8.833104e+09, 8.877434e+09, 8.919077e+09, 
    8.95798e+09, 8.994092e+09, 9.027367e+09, 9.05776e+09, 9.085231e+09, 
    9.109745e+09, 9.131267e+09, 9.14977e+09, 9.165227e+09, 9.177618e+09, 
    9.186927e+09, 9.193139e+09, 9.196247e+09, 9.196247e+09, 9.193139e+09, 
    9.186927e+09, 9.177618e+09, 9.165227e+09, 9.14977e+09, 9.131267e+09, 
    9.109745e+09, 9.085231e+09, 9.05776e+09, 9.027367e+09, 8.994092e+09, 
    8.95798e+09, 8.919077e+09, 8.877434e+09, 8.833104e+09, 8.786142e+09, 
    8.736609e+09, 8.684566e+09, 8.630074e+09, 8.573202e+09, 8.514017e+09, 
    8.452588e+09, 8.388985e+09, 8.323282e+09, 8.255552e+09, 8.18587e+09, 
    8.11431e+09, 8.04095e+09, 7.965864e+09, 7.889131e+09, 7.810825e+09, 
    7.731025e+09, 7.649805e+09, 7.567242e+09, 7.483411e+09, 7.398386e+09, 
    7.312241e+09, 7.225049e+09, 7.136881e+09, 7.047806e+09, 6.957896e+09, 
    6.867216e+09, 6.775833e+09, 6.683811e+09, 6.591213e+09, 6.4981e+09, 
    6.404531e+09,
  6.362479e+09, 6.452746e+09, 6.542493e+09, 6.631664e+09, 6.720201e+09, 
    6.808046e+09, 6.895139e+09, 6.981418e+09, 7.066822e+09, 7.151286e+09, 
    7.234745e+09, 7.317134e+09, 7.398386e+09, 7.478433e+09, 7.557208e+09, 
    7.634641e+09, 7.710664e+09, 7.785207e+09, 7.858201e+09, 7.929576e+09, 
    7.999264e+09, 8.067195e+09, 8.133301e+09, 8.197513e+09, 8.259766e+09, 
    8.319992e+09, 8.378128e+09, 8.434108e+09, 8.487873e+09, 8.539359e+09, 
    8.58851e+09, 8.635267e+09, 8.679578e+09, 8.721389e+09, 8.760649e+09, 
    8.797313e+09, 8.831335e+09, 8.862674e+09, 8.891291e+09, 8.917151e+09, 
    8.940219e+09, 8.96047e+09, 8.977876e+09, 8.992415e+09, 9.004068e+09, 
    9.012821e+09, 9.018663e+09, 9.021585e+09, 9.021585e+09, 9.018663e+09, 
    9.012821e+09, 9.004068e+09, 8.992415e+09, 8.977876e+09, 8.96047e+09, 
    8.940219e+09, 8.917151e+09, 8.891291e+09, 8.862674e+09, 8.831335e+09, 
    8.797313e+09, 8.760649e+09, 8.721389e+09, 8.679578e+09, 8.635267e+09, 
    8.58851e+09, 8.539359e+09, 8.487873e+09, 8.434108e+09, 8.378128e+09, 
    8.319992e+09, 8.259766e+09, 8.197513e+09, 8.133301e+09, 8.067195e+09, 
    7.999264e+09, 7.929576e+09, 7.858201e+09, 7.785207e+09, 7.710664e+09, 
    7.634641e+09, 7.557208e+09, 7.478433e+09, 7.398386e+09, 7.317134e+09, 
    7.234745e+09, 7.151286e+09, 7.066822e+09, 6.981418e+09, 6.895139e+09, 
    6.808046e+09, 6.720201e+09, 6.631664e+09, 6.542493e+09, 6.452746e+09, 
    6.362479e+09,
  6.319373e+09, 6.406312e+09, 6.492669e+09, 6.578392e+09, 6.663429e+09, 
    6.747724e+09, 6.831222e+09, 6.913867e+09, 6.9956e+09, 7.076365e+09, 
    7.1561e+09, 7.234745e+09, 7.312241e+09, 7.388526e+09, 7.463537e+09, 
    7.537212e+09, 7.60949e+09, 7.680307e+09, 7.749601e+09, 7.817309e+09, 
    7.883369e+09, 7.94772e+09, 8.010299e+09, 8.071048e+09, 8.129904e+09, 
    8.186811e+09, 8.241709e+09, 8.294543e+09, 8.345257e+09, 8.393798e+09, 
    8.440113e+09, 8.484152e+09, 8.525868e+09, 8.565214e+09, 8.602145e+09, 
    8.636621e+09, 8.668601e+09, 8.698051e+09, 8.724934e+09, 8.749221e+09, 
    8.770882e+09, 8.789891e+09, 8.806228e+09, 8.819871e+09, 8.830806e+09, 
    8.839017e+09, 8.844498e+09, 8.84724e+09, 8.84724e+09, 8.844498e+09, 
    8.839017e+09, 8.830806e+09, 8.819871e+09, 8.806228e+09, 8.789891e+09, 
    8.770882e+09, 8.749221e+09, 8.724934e+09, 8.698051e+09, 8.668601e+09, 
    8.636621e+09, 8.602145e+09, 8.565214e+09, 8.525868e+09, 8.484152e+09, 
    8.440113e+09, 8.393798e+09, 8.345257e+09, 8.294543e+09, 8.241709e+09, 
    8.186811e+09, 8.129904e+09, 8.071048e+09, 8.010299e+09, 7.94772e+09, 
    7.883369e+09, 7.817309e+09, 7.749601e+09, 7.680307e+09, 7.60949e+09, 
    7.537212e+09, 7.463537e+09, 7.388526e+09, 7.312241e+09, 7.234745e+09, 
    7.1561e+09, 7.076365e+09, 6.9956e+09, 6.913867e+09, 6.831222e+09, 
    6.747724e+09, 6.663429e+09, 6.578392e+09, 6.492669e+09, 6.406312e+09, 
    6.319373e+09,
  6.275223e+09, 6.35881e+09, 6.441759e+09, 6.52402e+09, 6.605544e+09, 
    6.686283e+09, 6.766183e+09, 6.845195e+09, 6.923265e+09, 7.000339e+09, 
    7.076365e+09, 7.151286e+09, 7.225049e+09, 7.297597e+09, 7.368877e+09, 
    7.438829e+09, 7.5074e+09, 7.574533e+09, 7.640172e+09, 7.704261e+09, 
    7.766745e+09, 7.827569e+09, 7.886679e+09, 7.94402e+09, 7.99954e+09, 
    8.053188e+09, 8.10491e+09, 8.15466e+09, 8.202386e+09, 8.248043e+09, 
    8.291585e+09, 8.332967e+09, 8.372148e+09, 8.409087e+09, 8.443745e+09, 
    8.476086e+09, 8.506077e+09, 8.533684e+09, 8.558878e+09, 8.581632e+09, 
    8.601922e+09, 8.619724e+09, 8.63502e+09, 8.647793e+09, 8.658028e+09, 
    8.665715e+09, 8.670843e+09, 8.673409e+09, 8.673409e+09, 8.670843e+09, 
    8.665715e+09, 8.658028e+09, 8.647793e+09, 8.63502e+09, 8.619724e+09, 
    8.601922e+09, 8.581632e+09, 8.558878e+09, 8.533684e+09, 8.506077e+09, 
    8.476086e+09, 8.443745e+09, 8.409087e+09, 8.372148e+09, 8.332967e+09, 
    8.291585e+09, 8.248043e+09, 8.202386e+09, 8.15466e+09, 8.10491e+09, 
    8.053188e+09, 7.99954e+09, 7.94402e+09, 7.886679e+09, 7.827569e+09, 
    7.766745e+09, 7.704261e+09, 7.640172e+09, 7.574533e+09, 7.5074e+09, 
    7.438829e+09, 7.368877e+09, 7.297597e+09, 7.225049e+09, 7.151286e+09, 
    7.076365e+09, 7.000339e+09, 6.923265e+09, 6.845195e+09, 6.766183e+09, 
    6.686283e+09, 6.605544e+09, 6.52402e+09, 6.441759e+09, 6.35881e+09, 
    6.275223e+09,
  6.230037e+09, 6.310255e+09, 6.38978e+09, 6.468569e+09, 6.546576e+09, 
    6.623755e+09, 6.700061e+09, 6.775447e+09, 6.849864e+09, 6.923265e+09, 
    6.9956e+09, 7.066822e+09, 7.136881e+09, 7.205726e+09, 7.273309e+09, 
    7.339579e+09, 7.404488e+09, 7.467984e+09, 7.530018e+09, 7.590542e+09, 
    7.649507e+09, 7.706863e+09, 7.762563e+09, 7.816561e+09, 7.868808e+09, 
    7.919261e+09, 7.967875e+09, 8.014606e+09, 8.059411e+09, 8.10225e+09, 
    8.143084e+09, 8.181873e+09, 8.218582e+09, 8.253174e+09, 8.285618e+09, 
    8.31588e+09, 8.343933e+09, 8.369748e+09, 8.3933e+09, 8.414565e+09, 
    8.433522e+09, 8.450151e+09, 8.464436e+09, 8.476363e+09, 8.485919e+09, 
    8.493095e+09, 8.497883e+09, 8.500278e+09, 8.500278e+09, 8.497883e+09, 
    8.493095e+09, 8.485919e+09, 8.476363e+09, 8.464436e+09, 8.450151e+09, 
    8.433522e+09, 8.414565e+09, 8.3933e+09, 8.369748e+09, 8.343933e+09, 
    8.31588e+09, 8.285618e+09, 8.253174e+09, 8.218582e+09, 8.181873e+09, 
    8.143084e+09, 8.10225e+09, 8.059411e+09, 8.014606e+09, 7.967875e+09, 
    7.919261e+09, 7.868808e+09, 7.816561e+09, 7.762563e+09, 7.706863e+09, 
    7.649507e+09, 7.590542e+09, 7.530018e+09, 7.467984e+09, 7.404488e+09, 
    7.339579e+09, 7.273309e+09, 7.205726e+09, 7.136881e+09, 7.066822e+09, 
    6.9956e+09, 6.923265e+09, 6.849864e+09, 6.775447e+09, 6.700061e+09, 
    6.623755e+09, 6.546576e+09, 6.468569e+09, 6.38978e+09, 6.310255e+09, 
    6.230037e+09,
  6.183825e+09, 6.260659e+09, 6.336752e+09, 6.412062e+09, 6.486551e+09, 
    6.560175e+09, 6.632894e+09, 6.704666e+09, 6.775447e+09, 6.845195e+09, 
    6.913867e+09, 6.981418e+09, 7.047806e+09, 7.112987e+09, 7.176916e+09, 
    7.23955e+09, 7.300845e+09, 7.360757e+09, 7.419243e+09, 7.47626e+09, 
    7.531766e+09, 7.585717e+09, 7.638074e+09, 7.688794e+09, 7.737838e+09, 
    7.785166e+09, 7.830739e+09, 7.874522e+09, 7.916475e+09, 7.956566e+09, 
    7.994759e+09, 8.031022e+09, 8.065324e+09, 8.097633e+09, 8.127923e+09, 
    8.156166e+09, 8.182336e+09, 8.20641e+09, 8.228367e+09, 8.248187e+09, 
    8.26585e+09, 8.281342e+09, 8.294647e+09, 8.305754e+09, 8.314652e+09, 
    8.321333e+09, 8.32579e+09, 8.32802e+09, 8.32802e+09, 8.32579e+09, 
    8.321333e+09, 8.314652e+09, 8.305754e+09, 8.294647e+09, 8.281342e+09, 
    8.26585e+09, 8.248187e+09, 8.228367e+09, 8.20641e+09, 8.182336e+09, 
    8.156166e+09, 8.127923e+09, 8.097633e+09, 8.065324e+09, 8.031022e+09, 
    7.994759e+09, 7.956566e+09, 7.916475e+09, 7.874522e+09, 7.830739e+09, 
    7.785166e+09, 7.737838e+09, 7.688794e+09, 7.638074e+09, 7.585717e+09, 
    7.531766e+09, 7.47626e+09, 7.419243e+09, 7.360757e+09, 7.300845e+09, 
    7.23955e+09, 7.176916e+09, 7.112987e+09, 7.047806e+09, 6.981418e+09, 
    6.913867e+09, 6.845195e+09, 6.775447e+09, 6.704666e+09, 6.632894e+09, 
    6.560175e+09, 6.486551e+09, 6.412062e+09, 6.336752e+09, 6.260659e+09, 
    6.183825e+09,
  6.136596e+09, 6.210038e+09, 6.282692e+09, 6.354524e+09, 6.425497e+09, 
    6.495574e+09, 6.564719e+09, 6.632894e+09, 6.700061e+09, 6.766183e+09, 
    6.831222e+09, 6.895139e+09, 6.957896e+09, 7.019455e+09, 7.079777e+09, 
    7.138825e+09, 7.196561e+09, 7.252946e+09, 7.307944e+09, 7.361518e+09, 
    7.41363e+09, 7.464245e+09, 7.513327e+09, 7.56084e+09, 7.606751e+09, 
    7.651027e+09, 7.693634e+09, 7.734541e+09, 7.773715e+09, 7.811129e+09, 
    7.846753e+09, 7.880559e+09, 7.912521e+09, 7.942612e+09, 7.970811e+09, 
    7.997093e+09, 8.021437e+09, 8.043825e+09, 8.064236e+09, 8.082655e+09, 
    8.099066e+09, 8.113456e+09, 8.125813e+09, 8.136126e+09, 8.144387e+09, 
    8.150589e+09, 8.154726e+09, 8.156796e+09, 8.156796e+09, 8.154726e+09, 
    8.150589e+09, 8.144387e+09, 8.136126e+09, 8.125813e+09, 8.113456e+09, 
    8.099066e+09, 8.082655e+09, 8.064236e+09, 8.043825e+09, 8.021437e+09, 
    7.997093e+09, 7.970811e+09, 7.942612e+09, 7.912521e+09, 7.880559e+09, 
    7.846753e+09, 7.811129e+09, 7.773715e+09, 7.734541e+09, 7.693634e+09, 
    7.651027e+09, 7.606751e+09, 7.56084e+09, 7.513327e+09, 7.464245e+09, 
    7.41363e+09, 7.361518e+09, 7.307944e+09, 7.252946e+09, 7.196561e+09, 
    7.138825e+09, 7.079777e+09, 7.019455e+09, 6.957896e+09, 6.895139e+09, 
    6.831222e+09, 6.766183e+09, 6.700061e+09, 6.632894e+09, 6.564719e+09, 
    6.495574e+09, 6.425497e+09, 6.354524e+09, 6.282692e+09, 6.210038e+09, 
    6.136596e+09,
  6.088361e+09, 6.158404e+09, 6.227619e+09, 6.295976e+09, 6.363442e+09, 
    6.429985e+09, 6.495574e+09, 6.560175e+09, 6.623755e+09, 6.686283e+09, 
    6.747724e+09, 6.808046e+09, 6.867216e+09, 6.925201e+09, 6.981969e+09, 
    7.037487e+09, 7.091722e+09, 7.144643e+09, 7.196217e+09, 7.246414e+09, 
    7.295202e+09, 7.342552e+09, 7.388432e+09, 7.432814e+09, 7.475667e+09, 
    7.516966e+09, 7.556683e+09, 7.594789e+09, 7.631261e+09, 7.666072e+09, 
    7.699199e+09, 7.73062e+09, 7.760311e+09, 7.788252e+09, 7.814423e+09, 
    7.838806e+09, 7.861382e+09, 7.882135e+09, 7.901051e+09, 7.918115e+09, 
    7.933316e+09, 7.946641e+09, 7.958081e+09, 7.967627e+09, 7.975273e+09, 
    7.981012e+09, 7.984841e+09, 7.986756e+09, 7.986756e+09, 7.984841e+09, 
    7.981012e+09, 7.975273e+09, 7.967627e+09, 7.958081e+09, 7.946641e+09, 
    7.933316e+09, 7.918115e+09, 7.901051e+09, 7.882135e+09, 7.861382e+09, 
    7.838806e+09, 7.814423e+09, 7.788252e+09, 7.760311e+09, 7.73062e+09, 
    7.699199e+09, 7.666072e+09, 7.631261e+09, 7.594789e+09, 7.556683e+09, 
    7.516966e+09, 7.475667e+09, 7.432814e+09, 7.388432e+09, 7.342552e+09, 
    7.295202e+09, 7.246414e+09, 7.196217e+09, 7.144643e+09, 7.091722e+09, 
    7.037487e+09, 6.981969e+09, 6.925201e+09, 6.867216e+09, 6.808046e+09, 
    6.747724e+09, 6.686283e+09, 6.623755e+09, 6.560175e+09, 6.495574e+09, 
    6.429985e+09, 6.363442e+09, 6.295976e+09, 6.227619e+09, 6.158404e+09, 
    6.088361e+09,
  6.039129e+09, 6.105772e+09, 6.171552e+09, 6.236442e+09, 6.300414e+09, 
    6.363442e+09, 6.425497e+09, 6.486551e+09, 6.546576e+09, 6.605544e+09, 
    6.663429e+09, 6.720201e+09, 6.775833e+09, 6.830297e+09, 6.883567e+09, 
    6.935614e+09, 6.986412e+09, 7.035934e+09, 7.084154e+09, 7.131045e+09, 
    7.176583e+09, 7.220742e+09, 7.263496e+09, 7.304823e+09, 7.344698e+09, 
    7.383099e+09, 7.420003e+09, 7.455388e+09, 7.489233e+09, 7.521518e+09, 
    7.552224e+09, 7.581331e+09, 7.608822e+09, 7.634681e+09, 7.65889e+09, 
    7.681435e+09, 7.702302e+09, 7.721477e+09, 7.738948e+09, 7.754704e+09, 
    7.768736e+09, 7.781033e+09, 7.791588e+09, 7.800395e+09, 7.807448e+09, 
    7.812741e+09, 7.816271e+09, 7.818037e+09, 7.818037e+09, 7.816271e+09, 
    7.812741e+09, 7.807448e+09, 7.800395e+09, 7.791588e+09, 7.781033e+09, 
    7.768736e+09, 7.754704e+09, 7.738948e+09, 7.721477e+09, 7.702302e+09, 
    7.681435e+09, 7.65889e+09, 7.634681e+09, 7.608822e+09, 7.581331e+09, 
    7.552224e+09, 7.521518e+09, 7.489233e+09, 7.455388e+09, 7.420003e+09, 
    7.383099e+09, 7.344698e+09, 7.304823e+09, 7.263496e+09, 7.220742e+09, 
    7.176583e+09, 7.131045e+09, 7.084154e+09, 7.035934e+09, 6.986412e+09, 
    6.935614e+09, 6.883567e+09, 6.830297e+09, 6.775833e+09, 6.720201e+09, 
    6.663429e+09, 6.605544e+09, 6.546576e+09, 6.486551e+09, 6.425497e+09, 
    6.363442e+09, 6.300414e+09, 6.236442e+09, 6.171552e+09, 6.105772e+09, 
    6.039129e+09,
  5.988909e+09, 6.052155e+09, 6.114508e+09, 6.175945e+09, 6.236442e+09, 
    6.295976e+09, 6.354524e+09, 6.412062e+09, 6.468569e+09, 6.52402e+09, 
    6.578392e+09, 6.631664e+09, 6.683811e+09, 6.734811e+09, 6.784643e+09, 
    6.833284e+09, 6.880711e+09, 6.926904e+09, 6.971842e+09, 7.015503e+09, 
    7.057866e+09, 7.098912e+09, 7.13862e+09, 7.176973e+09, 7.21395e+09, 
    7.249533e+09, 7.283705e+09, 7.316448e+09, 7.347746e+09, 7.377583e+09, 
    7.405943e+09, 7.432813e+09, 7.458176e+09, 7.482021e+09, 7.504335e+09, 
    7.525106e+09, 7.544322e+09, 7.561974e+09, 7.578052e+09, 7.592547e+09, 
    7.605452e+09, 7.616759e+09, 7.626462e+09, 7.634556e+09, 7.641037e+09, 
    7.645901e+09, 7.649145e+09, 7.650767e+09, 7.650767e+09, 7.649145e+09, 
    7.645901e+09, 7.641037e+09, 7.634556e+09, 7.626462e+09, 7.616759e+09, 
    7.605452e+09, 7.592547e+09, 7.578052e+09, 7.561974e+09, 7.544322e+09, 
    7.525106e+09, 7.504335e+09, 7.482021e+09, 7.458176e+09, 7.432813e+09, 
    7.405943e+09, 7.377583e+09, 7.347746e+09, 7.316448e+09, 7.283705e+09, 
    7.249533e+09, 7.21395e+09, 7.176973e+09, 7.13862e+09, 7.098912e+09, 
    7.057866e+09, 7.015503e+09, 6.971842e+09, 6.926904e+09, 6.880711e+09, 
    6.833284e+09, 6.784643e+09, 6.734811e+09, 6.683811e+09, 6.631664e+09, 
    6.578392e+09, 6.52402e+09, 6.468569e+09, 6.412062e+09, 6.354524e+09, 
    6.295976e+09, 6.236442e+09, 6.175945e+09, 6.114508e+09, 6.052155e+09, 
    5.988909e+09,
  5.937712e+09, 5.99757e+09, 6.056508e+09, 6.114508e+09, 6.171552e+09, 
    6.227619e+09, 6.282692e+09, 6.336752e+09, 6.38978e+09, 6.441759e+09, 
    6.492669e+09, 6.542493e+09, 6.591213e+09, 6.638811e+09, 6.685269e+09, 
    6.730571e+09, 6.774699e+09, 6.817636e+09, 6.859367e+09, 6.899874e+09, 
    6.939143e+09, 6.977157e+09, 7.013901e+09, 7.049361e+09, 7.083523e+09, 
    7.116371e+09, 7.147894e+09, 7.178077e+09, 7.206909e+09, 7.234377e+09, 
    7.260469e+09, 7.285175e+09, 7.308484e+09, 7.330385e+09, 7.350871e+09, 
    7.36993e+09, 7.387556e+09, 7.403741e+09, 7.418477e+09, 7.431758e+09, 
    7.443579e+09, 7.453934e+09, 7.462817e+09, 7.470226e+09, 7.476158e+09, 
    7.480609e+09, 7.483577e+09, 7.485062e+09, 7.485062e+09, 7.483577e+09, 
    7.480609e+09, 7.476158e+09, 7.470226e+09, 7.462817e+09, 7.453934e+09, 
    7.443579e+09, 7.431758e+09, 7.418477e+09, 7.403741e+09, 7.387556e+09, 
    7.36993e+09, 7.350871e+09, 7.330385e+09, 7.308484e+09, 7.285175e+09, 
    7.260469e+09, 7.234377e+09, 7.206909e+09, 7.178077e+09, 7.147894e+09, 
    7.116371e+09, 7.083523e+09, 7.049361e+09, 7.013901e+09, 6.977157e+09, 
    6.939143e+09, 6.899874e+09, 6.859367e+09, 6.817636e+09, 6.774699e+09, 
    6.730571e+09, 6.685269e+09, 6.638811e+09, 6.591213e+09, 6.542493e+09, 
    6.492669e+09, 6.441759e+09, 6.38978e+09, 6.336752e+09, 6.282692e+09, 
    6.227619e+09, 6.171552e+09, 6.114508e+09, 6.056508e+09, 5.99757e+09, 
    5.937712e+09,
  5.885548e+09, 5.942029e+09, 5.99757e+09, 6.052155e+09, 6.105772e+09, 
    6.158404e+09, 6.210038e+09, 6.260659e+09, 6.310255e+09, 6.35881e+09, 
    6.406312e+09, 6.452746e+09, 6.4981e+09, 6.54236e+09, 6.585513e+09, 
    6.627547e+09, 6.668449e+09, 6.708208e+09, 6.74681e+09, 6.784244e+09, 
    6.8205e+09, 6.855565e+09, 6.889429e+09, 6.922081e+09, 6.953512e+09, 
    6.98371e+09, 7.012667e+09, 7.040374e+09, 7.066821e+09, 7.092e+09, 
    7.115902e+09, 7.138521e+09, 7.159848e+09, 7.179877e+09, 7.198601e+09, 
    7.216014e+09, 7.23211e+09, 7.246883e+09, 7.260329e+09, 7.272444e+09, 
    7.283223e+09, 7.292662e+09, 7.30076e+09, 7.307511e+09, 7.312915e+09, 
    7.316969e+09, 7.319673e+09, 7.321026e+09, 7.321026e+09, 7.319673e+09, 
    7.316969e+09, 7.312915e+09, 7.307511e+09, 7.30076e+09, 7.292662e+09, 
    7.283223e+09, 7.272444e+09, 7.260329e+09, 7.246883e+09, 7.23211e+09, 
    7.216014e+09, 7.198601e+09, 7.179877e+09, 7.159848e+09, 7.138521e+09, 
    7.115902e+09, 7.092e+09, 7.066821e+09, 7.040374e+09, 7.012667e+09, 
    6.98371e+09, 6.953512e+09, 6.922081e+09, 6.889429e+09, 6.855565e+09, 
    6.8205e+09, 6.784244e+09, 6.74681e+09, 6.708208e+09, 6.668449e+09, 
    6.627547e+09, 6.585513e+09, 6.54236e+09, 6.4981e+09, 6.452746e+09, 
    6.406312e+09, 6.35881e+09, 6.310255e+09, 6.260659e+09, 6.210038e+09, 
    6.158404e+09, 6.105772e+09, 6.052155e+09, 5.99757e+09, 5.942029e+09, 
    5.885548e+09,
  5.832426e+09, 5.885548e+09, 5.937712e+09, 5.988909e+09, 6.039129e+09, 
    6.088361e+09, 6.136596e+09, 6.183825e+09, 6.230037e+09, 6.275223e+09, 
    6.319373e+09, 6.362479e+09, 6.404531e+09, 6.445522e+09, 6.485442e+09, 
    6.524282e+09, 6.562035e+09, 6.598693e+09, 6.634248e+09, 6.668692e+09, 
    6.702019e+09, 6.734221e+09, 6.76529e+09, 6.795221e+09, 6.824007e+09, 
    6.851641e+09, 6.878117e+09, 6.903431e+09, 6.927576e+09, 6.950547e+09, 
    6.972339e+09, 6.992947e+09, 7.012366e+09, 7.030593e+09, 7.047623e+09, 
    7.063453e+09, 7.078078e+09, 7.091497e+09, 7.103705e+09, 7.1147e+09, 
    7.124479e+09, 7.133041e+09, 7.140384e+09, 7.146505e+09, 7.151404e+09, 
    7.155078e+09, 7.157529e+09, 7.158754e+09, 7.158754e+09, 7.157529e+09, 
    7.155078e+09, 7.151404e+09, 7.146505e+09, 7.140384e+09, 7.133041e+09, 
    7.124479e+09, 7.1147e+09, 7.103705e+09, 7.091497e+09, 7.078078e+09, 
    7.063453e+09, 7.047623e+09, 7.030593e+09, 7.012366e+09, 6.992947e+09, 
    6.972339e+09, 6.950547e+09, 6.927576e+09, 6.903431e+09, 6.878117e+09, 
    6.851641e+09, 6.824007e+09, 6.795221e+09, 6.76529e+09, 6.734221e+09, 
    6.702019e+09, 6.668692e+09, 6.634248e+09, 6.598693e+09, 6.562035e+09, 
    6.524282e+09, 6.485442e+09, 6.445522e+09, 6.404531e+09, 6.362479e+09, 
    6.319373e+09, 6.275223e+09, 6.230037e+09, 6.183825e+09, 6.136596e+09, 
    6.088361e+09, 6.039129e+09, 5.988909e+09, 5.937712e+09, 5.885548e+09, 
    5.832426e+09 ;

 bk = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.01253, 0.04887, 0.10724, 0.18455, 0.27461, 0.36914, 
    0.46103, 0.54623, 0.62305, 0.69099, 0.75016, 0.8011, 0.84453, 0.88125, 
    0.9121, 0.93766, 0.95849, 0.97495, 0.98743, 0.9958, 1 ;

 pk = 1, 2.69722, 5.17136, 8.89455, 14.2479, 22.07157, 33.61283, 50.48096, 
    74.79993, 109.4006, 158.0046, 225.4411, 317.8956, 443.1935, 611.1156, 
    833.7439, 1125.834, 1505.208, 1993.158, 2614.863, 3399.784, 4382.062, 
    5600.87, 7100.731, 8931.782, 11149.97, 13817.17, 17001.21, 20775.82, 
    23967.34, 25527.65, 25671.22, 24609.3, 22640.51, 20147.13, 17477.63, 
    14859.86, 12414.93, 10201.44, 8241.503, 6534.432, 5066.179, 3815.607, 
    2758.603, 1880.646, 1169.339, 618.4799, 225, 10, 0 ;

 sftlf =
  0, 0.2884085, 0.9991118, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9922887, 0.3335225, 
    0.004607826, 0.003236954, 0.508559, 0.9850757, 0.9911836, 0.1925444, 0, 
    0, 0,
  0.02305815, 0.1375988, 0.944828, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.8519247, 
    0.1034592, 0, 0, 0.02152651, 0.1580271, 0.214971, 0, 0, 0, 0.004275662,
  0.6877087, 0.944828, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.7618825, 
    4.015537e-05, 0.2204578, 0.0836201, 0, 0, 0, 0, 0.006251427, 0.5966954,
  0.9875305, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.6890369, 0.02053772, 
    0.7023288, 0.225828, 0, 0, 0.2833943, 0.1682406, 0.614427, 1,
  0.9998894, 1, 1, 1, 1, 1, 1, 1, 1, 0.982605, 0.4463286, 0.2774308, 
    0.6133593, 0.9973181, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 0.5015463, 0.3794187, 0.9844274, 0.1219514, 0, 0.5, 
    1, 0.9917114, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 0.9341351, 0.2591562, 0, 0, 0, 0.778241, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.7423904, 
    0.641713, 1, 0.7179503, 0.7577073, 1, 1, 1, 0.9345905, 0.7734837,
  1, 1, 1, 1, 1, 1, 1, 1, 0.6711941, 0, 0, 0, 0, 0.7003056, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.7377394, 0.5135806, 0.05480789, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 0.5039137, 0, 0, 0, 0.02591443, 0.9401757, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 0.7924682, 0.0008498987, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 0.3537756, 0, 0, 0, 0, 0.8171846, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.8385026, 0.01230605, 0, 0, 0,
  0.9900191, 1, 1, 1, 0.982605, 0.8792336, 0.6995067, 0.5093474, 0.0169677, 
    0, 0, 0, 0, 0.7583464, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.5511215, 0, 0, 0, 0,
  0.6112348, 1, 0.995035, 0.7029089, 0.810859, 0.09081139, 0, 0, 0, 0, 0, 0, 
    0.01839714, 0.9189041, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.7265073, 0.04310679, 0, 0, 0, 0,
  0.4115516, 0.9695646, 0.32083, 0.3587675, 0.2985553, 0, 0, 0, 0, 0, 
    0.1353143, 0.3167184, 0.5955938, 0.2275586, 0.3671458, 0.9835829, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.3382995, 0, 0, 0, 0, 0,
  0, 0.1277016, 0.7127959, 0.9866941, 0.6133593, 0, 0, 0, 0, 0, 0.2077407, 
    0.931155, 0.5506355, 0.03697443, 0.1507062, 0.5356609, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9921315, 
    0.147725, 0, 0, 0, 0, 0,
  0.01037147, 0.1938587, 0.8625931, 1, 0.9973181, 0.4946559, 0.0311923, 0, 0, 
    0, 0.00735819, 0.5864723, 0.9627873, 0.8827814, 0.9648471, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9980701, 
    0.1807344, 0, 0, 0, 0, 0,
  0.7028435, 0.9317848, 1, 1, 1, 1, 0.9336721, 0.3483783, 0.07686493, 0, 0, 
    0.3183673, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 0.6919137, 0.0003099618, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 0.888535, 0.5828943, 0.380111, 0.6304355, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 0.983552, 0.1295606, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.8518441, 0.01128992, 
    0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.999961, 0.276726, 0, 0, 
    0, 0, 0.01621984,
  0.6853452, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.8485698, 
    0.009902901, 0, 0, 0, 0.1625293, 0.2812916,
  0.1046904, 0.9492866, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.5342661, 
    0, 0, 0, 0.2437459, 0.5925891, 0.1728241,
  0, 0.6909669, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9896021, 0.19564, 
    0, 0, 1.512684e-05, 0.6681376, 0.5249494, 0.001406433,
  0.104618, 0.3731309, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.516663, 0, 
    0, 0, 0.179388, 0.9754534, 0.9489582, 0.4696769,
  0.1094959, 0.1844557, 0.9892092, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.8602238, 0.005510823, 0, 0.005748244, 0.4703873, 0.9732017, 1, 
    0.8608779, 0.03971616,
  0.04849377, 0.01244223, 0.9232286, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.3732215, 0, 0, 0.02369886, 0.5267625, 0.6938574, 0.9234961, 0.9547111, 
    0.04446942,
  0.5122615, 0.02757481, 0.5740731, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.840474, 
    0.01930639, 0.0865661, 0.5162175, 0.1518759, 0, 0, 0.2306587, 0.5255683, 0,
  1, 0.5190924, 0.05039959, 0.9774919, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9979244, 
    0.6173158, 0.06360614, 0.3239541, 0.6181117, 0.3434, 0.08735604, 0, 0, 0, 
    0, 0,
  1, 0.6923935, 2.081939e-06, 0.6747068, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9996232, 1, 1, 1, 1, 
    0.3280995, 0.1371462, 0.7053908, 0.4147068, 0, 0, 0, 0, 0, 0, 0, 0,
  0.9767516, 0.9616271, 0.1639549, 0.271809, 0.9999644, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 0.79072, 0.9954807, 0.6932396, 0.992215, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 0.9982526, 0.7430784, 0.3342112, 0.9753816, 1, 1, 0.5895154, 
    0.4768312, 0.9639986, 0.7426976, 0.1318247, 0, 0, 0, 0, 0, 0, 0, 0,
  0.3953824, 1, 0.9443728, 0.9979815, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.8859383, 0.6344793, 0.8400888, 1, 0.6961708, 0.6793767, 1, 0.9887459, 
    0.4841065, 0.8715914, 1, 1, 1, 1, 0.9284868, 0.7849948, 0.7127485, 1, 
    0.9687542, 0.9541373, 0.7891752, 1, 1, 0.9629303, 0.8951254, 0.6504759, 
    0.8937041, 0.7830405, 0.342161, 1, 0.6261792, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.8566951, 0.02276905, 0.002447544, 0.514191, 0.722188, 0.6127455, 
    0.7949336, 0.7562089, 0.5650142, 0.06637619, 0.01120179, 0, 0, 0, 0, 0, 
    0, 0, 0,
  0.05505988, 0.888244, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.5507722, 
    0.0006194019, 0.116053, 0.619944, 0.742622, 0.1034394, 0.9146509, 
    0.4991146, 0.2116089, 0.9242266, 1, 1, 1, 1, 0.8386455, 0.4342496, 
    0.06022686, 0.5132908, 0.3214224, 0.5160704, 0.224035, 0.4073008, 
    0.5465707, 0.3329684, 0, 0.07634896, 0.5107231, 0.03671252, 0.2859505, 1, 
    0.6545428, 0.9156184, 0.97225, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.3421438, 0, 0, 0, 
    0.2840079, 0.6098053, 0.106933, 0.001375207, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  0.4128869, 0.9714226, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9036868, 
    0.3452899, 0, 0, 0, 0.0115361, 0.1913566, 0.1288761, 0.5540914, 
    0.9598167, 1, 1, 1, 1, 1, 1, 0.3918472, 0.3429512, 1, 0.8047241, 
    0.02029391, 0.7208738, 0.03791168, 0.4779267, 0, 0.01079109, 0.2673898, 
    0.04183982, 0, 0.1123773, 0.8191687, 0.7129377, 0.5516703, 0.9328146, 
    0.75521, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 0.9617294, 0.06184853, 0, 0, 0.000967195, 0.1277687, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0.9957435, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.8395773, 0.1179296, 
    0.01795836, 0.02010509, 0.007536734, 0.2286892, 0.04640759, 0, 0, 
    0.6564662, 1, 1, 1, 1, 1, 1, 1, 0.834378, 0.7319705, 1, 0.9198699, 
    0.01201014, 0.04465218, 0, 0, 0, 0.3684395, 0.5827318, 0, 0, 0, 
    0.2186891, 0.6873481, 0.1364655, 0.186791, 0.7450449, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.5434414, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.889401, 0.122736, 0.3139295, 
    0.7522845, 0.8038401, 0.3664241, 0.24319, 0.52267, 0.1478724, 0.09243008, 
    0.6729867, 0.9999971, 1, 1, 1, 1, 1, 0.9871168, 0.9992952, 1, 0.8422172, 
    0, 0, 0, 0, 0, 0.3275236, 0.8442517, 0.08887865, 0, 0, 0, 0.156116, 
    0.02045131, 3.470624e-05, 0.2521144, 0.6287342, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9975308, 0.149125, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.4399916, 0.4513926, 0.6248305, 1, 
    1, 1, 1, 1, 0.5065262, 0, 0, 0.4453909, 0.5339093, 0.4254689, 0.5834806, 
    1, 1, 1, 1, 1, 0.5982459, 0, 0, 0, 0, 0, 0, 0.3391043, 0.852947, 
    0.1592709, 0, 0, 0, 0, 0, 0.03027248, 0.4168469, 0.9877434, 1, 1, 1, 1, 
    0.8619069, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.9664218, 0.08247031, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.8920162, 0.5407821, 0.4654229, 
    0.2409135, 0.3909343, 0.988422, 1, 1, 1, 0.8909804, 0.531373, 0.2580832, 
    0.3792476, 0.7087116, 0.4061886, 0.4193644, 1, 1, 1, 1, 1, 0.2638651, 0, 
    0, 0, 0, 0, 0, 0, 0.2239696, 0.9176144, 0.4488631, 0.1449512, 
    0.001410662, 0, 0, 0.03603189, 0, 0.3868065, 0.9493498, 1, 1, 1, 
    0.7200027, 0.8212039, 0.990998, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 0.4792888, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.7146486, 0.118375, 0.4868317, 0.9180648, 
    0.8884519, 0.3578016, 0.3644181, 0.9821022, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 0.9876617, 0.3491453, 0, 0, 0, 0, 0, 0, 0, 0, 0.08260295, 
    0.4333614, 0.5040144, 0.3614931, 0, 0, 0, 0.005346482, 0.01236961, 
    0.2922967, 0.7454089, 1, 1, 0.8454538, 0.1922676, 0.3820402, 0.5675731, 
    0.9620153, 1, 1, 0.9772007, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.8661066, 0.00407539, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 0.7854356, 0.5305065, 0.2314634, 0, 0, 
    0.2847562, 0.6988515, 0.3205059, 0.001980788, 0.5282913, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 0.9088889, 0.3662374, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.002319489, 0.003097083, 0.006384837, 0.4009853, 
    0.9520847, 0.9565648, 0.7851307, 0.003207061, 0, 0.03928687, 0.8853757, 
    0.9915587, 0.4154324, 0.5028495, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.9239731, 0.04490227, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1532502, 0, 0, 0, 
    0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 0.6720341, 0.02851992, 0.0008780628, 0, 0, 0, 0, 0, 
    0.08552671, 0.7316995, 0.9995651, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.7766737, 0.4137197, 0.01565327, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.00839087, 0.179177, 0.3358206, 0.1938771, 0.08693577, 
    0.01849443, 0, 0, 0, 0.04255971, 0.1354656, 0, 0.2326064, 0.9961697, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9906443, 0.6093469, 0.08272952, 0, 0, 
    0, 0, 0, 0, 0.003714734, 0.04793612, 0.195166, 0.1305265, 0, 0, 0, 0, 0, 
    0, 0,
  1, 1, 1, 1, 1, 1, 0.997851, 0.8851513, 0.2218852, 0, 0, 0, 0, 0, 0, 0, 
    0.01474294, 0.9223265, 0.9997482, 1, 1, 1, 1, 0.8567648, 0.7138887, 
    0.7556022, 0.7419234, 0.5976552, 0.7780174, 0.7167592, 0.4319452, 
    0.02324593, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.02652722, 0.7279592, 0.6135988, 0.341273, 0.007845606, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.01614682, 0.6782818, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.9998435, 0.2067607, 0, 0, 0.091288, 0.5062699, 0.6916178, 0.7767209, 
    0.8624772, 0.9701989, 0.364688, 0, 0, 0, 0, 0, 0, 0, 0,
  0.4190771, 0.6497226, 0.9545459, 1, 1, 1, 0.6781163, 0.06010642, 0.5008612, 
    0.4229959, 0.1875891, 0, 0, 0, 0, 0, 0, 0.0595316, 0.5124435, 0.9682307, 
    1, 0.9258996, 0.5065909, 0.04083258, 0, 0, 0, 0.03120807, 0.1286479, 
    0.006753318, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1067706, 0.3340207, 
    0.2393772, 0, 0.002743472, 0.01939562, 0.08303384, 0.6292495, 0.01828023, 
    0, 0, 0, 0, 0, 0, 0, 0, 0.03133215, 0.007111566, 0.2436219, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9708926, 0.4725524, 0.1960722, 0, 0.1848622, 
    0.8739176, 1, 1, 1, 0.9030244, 0.3938256, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0.6705055, 1, 1, 0.9502218, 0.107991, 0.4462324, 1, 1, 0.7277706, 
    0.004069345, 0, 0, 0, 0, 0, 0, 0, 0.05657173, 0.3351253, 0.1607299, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.03699553, 
    0.2052931, 0.1163417, 0.04926136, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.3625355, 0.506983, 0.2779973, 0.5109867, 0.7485809, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 0.5927411, 0, 0, 0.1106688, 0.9105396, 1, 1, 1, 
    0.9959307, 0.4352124, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0.01193915, 0.7290006, 0.9996663, 0.09786085, 0.1382244, 0.5658905, 
    1, 1, 1, 0.8744788, 0.08482047, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1665618, 0.3248779, 0.0230974, 
    0.01594665, 0.02927415, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.2599293, 0.8565587, 0.00678506, 0, 0.0779523, 0.699297, 0.9691742, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 0.8166098, 0.03916229, 0, 0.005817841, 
    0.692153, 1, 1, 1, 0.9411603, 0.2435686, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0.2993191, 0.9495773, 0, 0.01423644, 0.7039637, 1, 1, 1, 1, 
    0.7995175, 0.254755, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.2888699, 0.705927, 0.7486029, 0.6040528, 0.3449149, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1760819, 
    0.4655593, 0, 0, 0, 0.1594579, 0.9752054, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.8951882, 0.2522649, 0.004452626, 0.5549645, 1, 1, 1, 0.8623571, 
    0.6075783, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0.07980675, 0.2809722, 0, 0.1385953, 0.7865735, 0.7880519, 
    0.968846, 0.5791082, 0.4798856, 0.9172074, 0.927383, 0.83219, 0.3994447, 
    0.04030702, 0, 0.07399552, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.0004920398, 0.3404756, 0.9613062, 0.4522832, 0.03017027, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01749192, 0.01128817, 
    0.1379025, 0, 0, 0, 0.04587796, 0.9871097, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.6999564, 0.3755875, 0.9989443, 0.6214731, 0.5969585, 0.5454745, 
    0.1750769, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0.1596749, 0.01195103, 0.1571471, 0.02306698, 0.028618, 
    0.3427889, 0.721784, 1, 1, 0.8513392, 0.3177238, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.02060047, 0.2733825, 0.02397867, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.4457313, 0.7043854, 1, 1, 1, 1, 1, 1, 1, 1, 0.6029556, 0.9542752, 
    0.4643725, 0.2527745, 0.02328439, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0.007150483, 0.7961679, 0.8434761, 0.9726763, 
    0.4238593, 0.5026287, 0.622201, 0.4973026, 0.0772241, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.2232726, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 0.9596362, 0.2153704, 0.02692382, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0.5481955, 1, 1, 0.9846066, 0.5166809, 0, 0, 
    0.0605782, 0, 0, 0, 0.02565648, 0.2292144, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.002742995, 0.9592576, 1, 1, 1, 1, 
    1, 1, 1, 1, 0.8386291, 0.06731934, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0.7911306, 0.744423, 0.9958476, 0.3917643, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.1602756, 0.7774471, 1, 1, 1, 1, 1, 1, 1, 1, 0.7282078, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0.2763341, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.02465551, 0.5389555, 
    0.09023141, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.3491064, 0.7970511, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.7709398, 0.05621546, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.02616456, 0.4072716, 0.02764438, 0, 0, 0, 0, 0, 0, 0, 0, 0.007946228, 
    0.0215098, 0.1481985, 0.1512895, 0.2826785, 0.7654743, 0.9869945, 
    0.5499371, 0.567008, 0.05657073, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.3411054, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.7214631, 0.1254226, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.5718764, 1, 0.617721, 0, 0, 0, 0, 0, 0, 0, 0.148285, 0.6013126, 
    0.7386797, 0.8317872, 0.9721572, 0.9878897, 1, 1, 1, 1, 0.5187135, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.04601588, 0.1928452, 0.9953901, 1, 1, 1, 1, 1, 1, 0.9362985, 0.1519071, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.02308159, 
    0.9368013, 1, 0.5605719, 0, 0, 0, 0, 0.0994027, 0.1519942, 0.4023046, 
    0.8973336, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.6283081, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.2124189, 0.437899, 0, 
    0.7649915, 1, 1, 1, 0.9788436, 0.7998188, 1, 0.4011095, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1528232, 
    0.9851291, 1, 0.5690181, 0.007882722, 0, 0, 0.3224736, 0.4599625, 
    0.9042956, 0.999677, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.4572058, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.006458772, 
    0.0237647, 0, 0.227326, 0.9942815, 1, 0.6645961, 0.4432212, 0.03989381, 
    0.5392244, 0.2095875, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.430079, 
    0.7312796, 0.8450026, 0.1614028, 0, 0.04361914, 0.8531964, 0.8497482, 
    0.9997948, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.8977383, 0.3332031, 
    0.3655361, 0.04765641, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.7132292, 1, 0.816526, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.05260738, 0.07836438, 0, 0, 0.2491814, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 0.9207466, 0.7041428, 1, 0.7042463, 0.01935159, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1916869, 0.997572, 
    0.9664844, 0.2796616, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.3168469, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.8713294, 
    0.7350758, 1, 0.9985892, 0.5351546, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1795665, 0.9986884, 0.8846707, 0.5677841, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.3550282, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.279303, 
    0.6442038, 1, 0.6813606, 0.6184936, 0.1960024, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0251202, 0.260837, 0, 0.0004929128, 
    0.3365258, 0.0114776, 0.03985736, 0.1344334, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.1158035, 0.890343, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.7351844, 0.5533677, 1, 0.7738451, 0.9701509, 0.3894742, 0.001606799, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.005773118, 0.3039451, 0.7407112, 
    0.7999177, 0.9048856, 0.0141415, 0.1831883, 0.4115106, 0, 0.1069227, 
    0.2025667, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1092487, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.5193717, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.994473, 0.5692437, 
    0.4542774, 0.9261664, 0.8238658, 0.2153217, 0.5868801, 1, 0.7394806, 
    0.8058553, 0.1632256, 0.547113, 0.06057538, 0.09398247, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.7215818, 1, 1, 1, 1, 0.4168746, 0.8358276, 0.9664901, 
    0.1808136, 0.01235209, 0.0244422, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.02900386, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.6050302, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.8627397, 0.2401952, 0, 0, 
    0.121907, 0.1521004, 0, 0.644744, 0.9510419, 0.301559, 0.2032923, 
    0.2832184, 0.1715124, 0.0642454, 0.3894436, 0.355457, 0.1890444, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.07950651, 0.9975182, 1, 1, 1, 1, 0.8763351, 
    0.9740863, 0.9582601, 0.05713792, 0.006239007, 0.08203404, 0.03931703, 
    0.00247307, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.06966187, 0.06613558, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.003755757, 0.5864659, 1, 1, 1, 1, 1, 0.9925512, 0.8724307, 0.6710725, 
    0.7534792, 0.07587746, 0, 0, 0, 0, 0, 0, 0.3674421, 0.5488101, 0.6089712, 
    0.5379397, 0.2472398, 0.1861075, 0.1012413, 0.1267425, 0.4983214, 
    0.6058319, 0.03750185, 0, 0, 0, 0, 0, 0, 0, 0, 0.5366537, 1, 1, 1, 1, 1, 
    1, 1, 0.6697894, 0.2345046, 0.8237509, 0.9863058, 0.4740853, 0.4750053, 
    0.1235425, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.4309661, 0.9817041, 1, 1, 1, 1, 1, 0.571421, 0.7863377, 0.1386277, 
    0.02245102, 0, 0, 0, 0, 0, 0, 0.05556273, 0.9789172, 0.7375769, 
    0.8189688, 0.3559348, 0.6307323, 0.6821151, 0.5123709, 0.6651374, 
    0.8837627, 0.1572086, 0.05174712, 0.09259965, 0, 0, 0, 0, 0, 0, 
    0.06662905, 0.9413299, 1, 1, 1, 1, 1, 1, 1, 0.9999163, 0.9697776, 1, 1, 
    1, 0.4300958, 0.003663761, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.1867139, 0.9595957, 1, 1, 1, 1, 1, 1, 0.284351, 0.2819466, 0, 0, 0, 0, 
    0, 0, 0, 0.221816, 0.234015, 0.1498427, 0.4379888, 0.4701115, 0.3815823, 
    0.202223, 0.06689857, 0.1760091, 0.348862, 0.2906938, 0.3599098, 
    0.8773224, 0.6843942, 1.096974e-05, 0, 0, 0, 0, 0, 0.729326, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 0.9291328, 0.1750867, 0, 0, 0, 0, 0, 0, 0, 
    0.1284918, 0.03147244, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.2094367, 0.9369895, 1, 1, 1, 1, 1, 1, 0.8089225, 0.05077393, 0, 0, 0, 
    0, 0, 0, 0.1286864, 0.5131698, 0.9357795, 0.9835859, 0.6595818, 
    0.6586512, 0.5519477, 0.6267641, 0.5283211, 0.1642075, 0.2885776, 
    0.04336228, 0.04232852, 0.7210842, 0.8761302, 1, 0.4428093, 0, 0, 0, 0, 
    0.2362406, 0.9876587, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.8892759, 
    0.2210028, 0, 0, 0, 0, 0.01768243, 0.2350183, 0.2126607, 0.007313905, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.09397414, 0.9518533, 1, 1, 1, 1, 1, 0.9310701, 0.6551082, 0.02464128, 
    0, 0, 0, 0, 0.001893531, 0.428525, 0.660005, 0.9646558, 0.9979754, 1, 1, 
    0.7802781, 0.8504569, 0.2165388, 0.643451, 0.9057896, 0.4174795, 
    0.5542305, 0.6763288, 0.8081042, 0.988646, 0.6779991, 0.7144226, 
    0.3391109, 0.03010433, 0.1083374, 0.3236497, 0.4993806, 0.6720286, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.7566548, 0.09032444, 0, 0, 0, 
    0.1800638, 0.2171838, 0.04050701, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.5591969, 0.9228026, 1, 1, 1, 0.9221501, 0.5172973, 0.05100384, 0, 0, 0, 
    0.0007068556, 0.01091526, 0.0301949, 0.2755317, 0.965713, 1, 1, 
    0.9936191, 1, 1, 0.9859811, 0.619966, 0.1089375, 0.4886177, 0.6999307, 
    0.07001494, 0.6258047, 0.9147264, 1, 1, 0.6264263, 0, 0, 0.1941441, 
    0.9471765, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.5419797, 
    0, 0.015395, 0.2036542, 0.6540743, 0.4381296, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.006838025, 0.01351406, 0.4722523, 0.538614, 0.2337886, 0.001982945, 0, 
    0, 0, 0, 0, 0.7464898, 0.9450542, 0.9789113, 0.99442, 1, 0.9895004, 
    0.7432182, 0.2929687, 0.8314089, 0.8995512, 0.7964581, 0.1749706, 
    0.6521643, 0.7756425, 0.008177926, 0.1344325, 0.8013356, 1, 0.9843748, 
    0.6497664, 0.5200529, 0.04047306, 0.6355119, 0.8531175, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 0.8961154, 0.9560985, 0.9943568, 1, 0.9338681, 
    0.5818689, 0.7449133, 0.7265122, 0.293891, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.0579614, 0.9415749, 0.8603365, 0.9990121, 1, 
    0.803029, 0.3949734, 0.1770097, 0.005452511, 0.510583, 0.7336312, 
    0.001113111, 0.1646328, 0.8604911, 0.5931268, 0.1902591, 0.5364736, 
    0.9966938, 0.956994, 1, 0.9285627, 0.4400202, 0.722735, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9410389, 0.5555537, 0.3014219, 0.601414, 
    0.4825325, 0.2935872, 0.08583173, 0.004107873, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.03901332, 0.3728116, 0.4575627, 1, 1, 0.3147727, 
    0.3332067, 0.2217817, 0.05301935, 0.7761925, 0.6799878, 0.399193, 
    0.7055106, 0.8377438, 0.6134337, 0.4755627, 0.2565599, 0.4595538, 
    0.6566908, 0.4802974, 0.3227839, 0.6104215, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 0.9089081, 0.5222241, 0.4558146, 0.1927821, 0.1057313, 
    0.7160483, 0.6894037, 0.0001066323, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.001781516, 0.5839874, 0.9946612, 1, 1, 0.9786469, 
    0.2361013, 0, 0, 0.2998931, 1, 0.8093447, 0.6758854, 0.9936388, 
    0.9348447, 0.6461143, 0.534321, 0.2699139, 0.8118511, 0.9714402, 
    0.7283285, 0.8378774, 0.9670031, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 0.8234991, 0.08674643, 0.0131576, 0, 0, 0.02502642, 0.01614379, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.1014065, 0.7311866, 0.7506915, 1, 1, 0.9619322, 
    0.6062644, 0.1703102, 0, 0.04583564, 0.6992308, 0.8417487, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9660713, 
    0.2967638, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.01285044, 0.1548295, 0.6499813, 0.889262, 0.9474576, 
    0.3051719, 0.1076564, 0.5899696, 0.2210208, 0, 0.1423286, 0.6488663, 
    0.7522198, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 0.9999971, 0.4893933, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.1127665, 0.1135007, 0, 6.399585e-05, 0.0003775573, 
    0.03852168, 0.05766925, 0, 0.171762, 0.01750567, 0.4126715, 0.8537696, 
    0.8530025, 0.672665, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 0.9984903, 0.1519116, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.0262549, 0.4324569, 0.9188194, 0.03891509, 0.07369219, 0.2784357, 
    0.439794, 0.9090685, 0.8842618, 0.613674, 0.169175, 0.0007593664, 
    0.05496632, 0.3555141, 0.4366377, 0.1746797, 0.660701, 0.9513029, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9929273, 
    0.1262638, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0152431, 0.3903114, 0.8834387, 1, 0.809934, 0, 0.08427224, 0.9253466, 
    1, 1, 1, 0.7736004, 0.162165, 0.0586152, 0.3602923, 0.03943993, 
    0.001398534, 0, 0.2553839, 0.8987577, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9784375, 0.07446165, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.006909454, 
    0.02203574, 0.2018838, 0.2004992, 0.2420584, 0.6730793, 0.9998235, 1, 1, 
    0.9541899, 0.6909702, 0.8539598, 1, 1, 1, 0.9992172, 0.3129094, 0, 0, 0, 
    0, 0, 0, 0, 0.5284762, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 0.9821761, 0.7433433, 0.2581827, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.004164889, 
    0.598833, 0.912891, 0.9848074, 1, 0.9949051, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 0.8401424, 0, 0, 0, 0, 0, 0, 0, 0, 0.1808639, 0.9999599, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9998994, 0.5513852, 
    0.3237998, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.6889238, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.7519505, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.8577955, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 0.9713004, 0.1253456, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.03594787, 0, 0.0008203032, 
    0.4332399, 0.5592608, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9933216, 
    0.4570104, 0.01265947, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.8118156, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.942905, 0.6050133, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0007849386, 0.06672296, 0.6196942, 
    0.3867162, 0.3914538, 0.7130988, 0.1269462, 0.9995891, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 0.6703829, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.06998937, 
    0.5995811, 0.9730762, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 0.4093178, 0.145072, 0.09990545, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.003637707, 0.559929, 0.9073727, 1, 
    0.9975478, 0.999097, 0.3226125, 0.1728628, 0.996939, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 0.618335, 0.03839462, 0.163095, 0, 0, 0, 0, 0, 0.00750303, 
    0.003358266, 0.3714445, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 0.8540727, 0.2479777, 0.566503, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1012027, 0.4235917, 0.7059572, 
    0.9331499, 1, 0.8808568, 0.05236256, 0, 0.6189646, 0.9339727, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 0.8560801, 0.09653471, 0, 0, 0, 0, 0.001193712, 
    0.3857171, 0.8091468, 0.9605917, 0.8586759, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9887962, 0.08099455, 0.4007379, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0009469227, 0.2329264, 0.444853, 
    0.8093558, 0.5496757, 0, 0.002437673, 0.227669, 0.2634807, 0.7164366, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9659117, 0.3167773, 0, 0.4677332, 0.5943365, 
    0.5637257, 0.8562685, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.8810632, 0.004721967, 0.05446313, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.2208384, 0.1411825, 0, 
    0.01509914, 0.3049383, 0.1022427, 0.001643809, 0.7302889, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 0.5155249, 0, 0.2220955, 0.925254, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9658247, 
    0.04132003, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.03023492, 0.1040698, 0, 
    0, 0.2589638, 0.8127933, 0.4118724, 0.5901706, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.6797279, 0.03147244, 0.148788, 0.8013205, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9649417, 
    0.2472448, 0.0001925075, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.2116711, 0.7594843, 
    0.04181511, 0, 0, 0.2791559, 0.9919224, 0.9871036, 0.5026899, 1, 1, 1, 1, 
    1, 1, 1, 1, 0.6875119, 0.1673929, 0.6100693, 0.9931602, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 0.9986221, 0.9031882, 0.02072693, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1597966, 0.6263976, 
    0.3037237, 0.3064115, 0.3001947, 0.9453359, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 0.9858415, 0.9203051, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9886171, 0.999054, 
    0.7919562, 0.001658652, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.106327, 0.9335366, 
    0.7329312, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 0.5367375, 0.8222567, 0.3355962, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.002422816, 0.6366513, 
    0.9978582, 0.7376231, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 0.998466, 0.4211002, 0.5821907, 0.06182952, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.2501551, 0.9984199, 
    0.2726648, 0.9098034, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 0.657743, 0.8075415, 0.4442849, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.221493, 0.713844, 
    0.009902901, 0.6008854, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 0.9938447, 0.7752694, 0.610476, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.006310866, 0, 
    0.1160645, 0.9701369, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 0.9781886, 0.1501769, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.5544846, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.7063521, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.5219765, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.9999979, 0.291099, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0005927939, 0.3538766, 
    0.271129, 0.9385704, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 0.8661439, 0.2963106, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.03236142, 0.5147032, 
    0.9229311, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 0.9242505, 0.07807732, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 orog =
  1.957085, 182.3516, 345.853, 566.5532, 583.9197, 703.0031, 841.8619, 
    930.701, 1327.418, 1866.999, 2029.211, 1998.469, 1606.435, 2058.914, 
    894.809, 267.2261, 1038.635, 95.99315, -29, -29, -14.74468, 50.54665, 
    131.9456, 149.8255, 180.3951, 144.0376, 117.0449, 65.4011, 47.57902, 
    52.56764, 62.57636, 88.29622, 103.0397, 116.2788, 146.1452, 149.0459, 
    260.9405, 209.8252, 240.3782, 305.7633, 380.0433, 410.2039, 401.1645, 
    344.6812, 350.6726, 420.6497, 639.9168, 1359.416, 1773.189, 1596.877, 
    1193.995, 945.0976, 478.8944, 313.0052, 364.5321, 544.9355, 728.1349, 
    913.1708, 1094.162, 1205.655, 1103.695, 1186.761, 1181.66, 1198.702, 
    1409.169, 1265.896, 1273.084, 1305.134, 1441.755, 1591.454, 1519.917, 
    1441.886, 1330.869, 1070.649, 1189.587, 1315.408, 1415.29, 1531.97, 
    1529.214, 1473.449, 1430.014, 1306.896, 1270.828, 872.1915, 165.6583, 
    2.112291, 1.155395, 0.02070807, 0.08559992, 13.39372, 105.9956, 72.41502, 
    2.817191, 0, 0, 0.04834903,
  0.02893994, 4.580082, 170.3799, 581.9701, 947.2767, 1071.069, 1146.666, 
    1154.808, 1640.017, 1900.844, 1998.073, 1884.909, 1641.079, 1859.79, 
    780.6656, 620.8061, 1727.327, 225.5852, -29, -29, -29, 38.14354, 
    126.9196, 155.8592, 184.8903, 179.1412, 129.6505, 97.10344, 37.13656, 
    33.23013, 51.04347, 71.70508, 91.74311, 103.1298, 126.9913, 145.6968, 
    179.7494, 230.5837, 298.0778, 375.3928, 434.7722, 459.8557, 350.7677, 
    343.3709, 347.6726, 356.1186, 381.6495, 446.8376, 603.9845, 758.576, 
    881.1244, 1095.882, 904.9011, 568.9519, 433.0408, 654.4484, 862.9261, 
    1147.874, 1391.479, 1546.497, 1694.146, 1655.956, 1846.877, 1863.535, 
    1773.414, 1861.801, 1658.115, 1432.014, 1446.591, 1505.779, 1598.366, 
    1639.378, 1501.092, 1183.134, 1002.323, 1205.448, 1280.397, 1347.836, 
    1565.089, 1583.707, 1551.659, 1326.685, 1098.686, 688.5358, 124.0418, 
    3.131963, 2.67241, 0, 0, 0.3741298, 0, 14.65283, 0, 0, 0, 0.08931515,
  735.5396, 867.0506, 660.6748, 924.9462, 1301.789, 1480.976, 1317.01, 
    1341.343, 1806.828, 2025.722, 2183.452, 2051.318, 1930.586, 1732.126, 
    665.5182, 1034.291, 2036.85, 544.5954, -29, -29, -28.76467, 38.63471, 
    172.218, 155.2569, 183.3024, 142.7022, 156.3304, 131.9387, 71.52921, 
    29.83442, 38.42982, 63.1153, 82.10826, 123.0225, 117.6491, 159.6424, 
    210.2419, 265.2799, 324.6303, 429.2385, 526.7354, 552.8436, 445.1412, 
    408.4677, 410.2799, 482.5757, 457.1882, 425.4275, 467.3434, 724.1971, 
    978.342, 1341.993, 1428.619, 1158.37, 714.2965, 634.1248, 1100.511, 
    1729.557, 2079.457, 2205.601, 2096.228, 1923.082, 2023.244, 2032.364, 
    2087.194, 1819.859, 1741.359, 1652.907, 1411.046, 1353.822, 1332.2, 
    1373.966, 1373.264, 1169.126, 951.4221, 1059.032, 1129.511, 1144.062, 
    1270.443, 1435.999, 1450.52, 1447.836, 1236.854, 758.832, 350.9756, 
    181.3987, 25.64147, 0, 7.676435, 3.285792, 0, 0, 0, 0, 4.333813, 55.45658,
  1304.387, 1437.602, 1376.26, 1494.452, 1659.236, 1723.898, 1639.994, 
    1657.578, 1850.001, 2092.416, 1922.954, 1856.68, 1913.263, 1612.252, 
    1244.188, 1688.415, 1823.349, 597.8655, -28.95335, -29, -29, 36.93167, 
    126.3385, 56.37119, 89.7822, 66.37797, 91.53525, 123.4684, 92.97884, 
    64.8284, 57.79882, 59.7579, 86.7978, 105.0893, 148.6383, 195.5772, 
    329.0817, 307.0089, 342.0926, 436.9752, 591.1713, 694.5746, 679.3177, 
    636.2111, 632.0756, 646.1209, 669.288, 648.6287, 782.5434, 883.3128, 
    793.3741, 676.8798, 926.3399, 801.6874, 746.4554, 1202.792, 1920.346, 
    2443.33, 2322.053, 1982.287, 1837.848, 1673.851, 1988.25, 2200.716, 
    1986.238, 1899.81, 1884.782, 1790.649, 1548.873, 1296.591, 1256.828, 
    1255.077, 1205.229, 1093.803, 927.5923, 972.8065, 1059.568, 1028.104, 
    1103.09, 1202.041, 1344.654, 1430.761, 1304.095, 857.4107, 614.5168, 
    408.0826, 142.5798, 1.184603, 40.65562, 3.480806, 0, 1.402507, 22.73934, 
    1.869505, 22.95708, 208.0578,
  1176.996, 1274.15, 1167.862, 1260.973, 1305.267, 1444.57, 1547.88, 
    1561.639, 1724.48, 1392.404, 542.0779, 297.3251, 709.7617, 908.8043, 
    1689.685, 1619.551, 990.7944, 115.7064, -24.46063, -28.99723, -29, 11.77, 
    -18.20284, -18.30782, -26.05886, -15.76914, 55.73129, 98.28559, 125.4715, 
    138.3384, 126.8703, 111.3977, 77.0961, 90.02938, 117.3675, 253.6755, 
    387.6956, 435.0849, 377.246, 411.8622, 531.7675, 673.597, 770.8846, 
    853.8765, 854.3976, 850.265, 792.6041, 745.4413, 733.783, 735.1926, 
    603.2223, 591.2675, 993.4567, 1367.18, 1860.522, 2238.518, 2511.91, 
    2284.058, 1663.224, 1322.216, 1438.35, 1776.375, 2169.013, 2455.426, 
    2488.388, 2387.191, 2351.167, 2100.744, 1704.273, 1439.597, 1375.393, 
    1281.368, 1147.538, 1084.584, 931.0007, 951.1368, 1033.676, 1018.033, 
    1023.891, 1108.402, 1268.471, 1365.725, 1364.301, 974.9635, 739.7955, 
    399.5302, 73.64684, 12.84806, 147.529, 5.471954, 0, 24.00544, 116.3721, 
    114.7116, 240.0056, 341.1817,
  1120.788, 1306.315, 1094.511, 1054.712, 1080.561, 1158.717, 1213.522, 
    1205.066, 948.7064, 166.4328, 0, 0, 7.011492, 766.0705, 1910.302, 
    1318.522, 220.8738, 20.13437, -22.87948, -28.96292, -28.99967, -28.96005, 
    -28.95333, -28.95845, -28.27328, -19.16533, 25.35257, 78.57539, 126.1784, 
    178.1593, 206.8317, 152.6626, 97.64114, 76.05511, 110.28, 209.1862, 
    385.8008, 487.759, 490.3545, 435.6064, 477.5195, 573.1337, 679.9717, 
    815.3858, 863.851, 795.056, 638.4842, 521.1765, 490.9408, 599.1897, 
    654.6764, 994.7811, 1491.828, 2086.955, 2473.281, 2589.081, 2203.682, 
    1937.777, 1327.908, 1322.338, 1643.389, 1980.04, 2347.152, 2586.005, 
    2474.671, 2249.25, 1973.765, 1742.107, 1577.967, 1488.696, 1454.051, 
    1334.462, 1222.04, 1055.741, 975.7679, 973.0269, 1098.012, 1137.429, 
    1093.573, 1125.746, 1300.224, 1360.541, 1194.296, 881.052, 581.177, 
    281.8254, 19.61534, 84.07046, 212.6468, 69.3125, 29.19267, 158.5775, 
    304.7471, 402.8232, 454.9509, 428.1056,
  1187.477, 1316.139, 1129.726, 991.171, 1030.374, 1016.187, 1020.988, 
    818.59, 381.7968, 0, 0, 0, 0, 1129.767, 1979.666, 998.5098, 264.3186, 
    59.78041, -4.723167, -24.42554, -28.50731, -28.65225, -28.92911, -29, 
    -28.607, -24.37205, 20.2152, 104.2612, 164.2149, 231.1236, 260.2584, 
    221.0597, 141.5681, 105.8174, 115.9729, 151.8276, 274.3087, 439.8468, 
    448.8825, 399.3673, 408.2239, 453.6656, 569.141, 609.5902, 626.4427, 
    521.6019, 365.9188, 284.7949, 285.1086, 423.1974, 846.5926, 1237.006, 
    1726.326, 2102.346, 2434.645, 2372.822, 2198.263, 1666.205, 1424.405, 
    1409.403, 1744.127, 2013.176, 2073.452, 2140.749, 2030.338, 1827.267, 
    1580.342, 1325.149, 1298.67, 1349.97, 1428.83, 1395.826, 1250.978, 
    1179.868, 1037.025, 1015.187, 1152.761, 1271.608, 1141.957, 1128.437, 
    1250.247, 1118.777, 820.3528, 513.1799, 459.0807, 201.0253, 50.98212, 
    173.3005, 353.3956, 272.952, 377.204, 340.7662, 338.8821, 282.7307, 
    42.52118, 0,
  911.2604, 1162.884, 1137.084, 979.4952, 1010.004, 1126.895, 1059.642, 
    869.5664, 252.7621, 0, 0, 0, 0, 1150.678, 1275, 595.7617, 273.573, 
    133.9935, 32.51972, -16.08583, -22.48619, -23.88273, -23.75681, 
    -24.06026, -24.22806, -20.21073, 10.21312, 100.5829, 164.7874, 248.1127, 
    306.6323, 287.0247, 220.7695, 169.7234, 135.2546, 137.2507, 172.6728, 
    311.0542, 341.0001, 327.2497, 348.4995, 425.6412, 463.1763, 447.4398, 
    353.7435, 252.8357, 186.9208, 193.5265, 269.0485, 416.4105, 833.4974, 
    1255.776, 1478.953, 1658.504, 2096.166, 2288.637, 1723.026, 1429.502, 
    949.519, 1162.872, 1667.993, 1924.058, 2051.646, 1868.885, 1679.083, 
    1502.363, 1410.3, 1248.582, 1158.49, 1393.645, 1598.457, 1420.972, 
    1293.249, 1159.699, 1133.274, 1037.51, 1155.602, 1250.937, 1090.242, 
    1007.832, 1146.141, 923.0365, 519.2554, 340.7791, 297.567, 152.0113, 
    84.55415, 319.1597, 474.4228, 619.5093, 846.3072, 366.6542, 0.09596219, 
    0, 0, 0,
  612.0165, 1024.829, 1129.861, 947.5595, 1080.557, 1194.547, 1150.219, 
    904.1955, 156.9333, 0, 0, 0, 0, 583.678, 439.6959, 309.7408, 232.4993, 
    133.5744, 75.71014, -1.082752, -7.73104, -16.27212, -16.11549, -15.90899, 
    -15.91451, -10.86247, 4.381418, 61.24113, 156.1658, 234.102, 316.4874, 
    335.1181, 275.5302, 255.234, 212.9649, 181.6552, 180.8939, 256.1131, 
    302.8167, 311.314, 343.6282, 353.8376, 353.0165, 257.5091, 195.26, 
    136.4342, 132.6939, 165.401, 204.5192, 263.7407, 417.9625, 651.0251, 
    757.1484, 1176.346, 1630.802, 1775.998, 1641.073, 1216.329, 1179.213, 
    1361.391, 1647.038, 1987.515, 2015.377, 1927.813, 1564.168, 1375.637, 
    1276.543, 1056.094, 1081.178, 1433.004, 1697.667, 1528.249, 1249.511, 
    1163.054, 1084.624, 1005.993, 992.0644, 1018.707, 950.4731, 940.6085, 
    1033.09, 798.034, 387.972, 229.6093, 197.4241, 132.7397, 211.0327, 
    408.1602, 644.9759, 902.4259, 1280.562, 421.0834, 0, 0, 0, 0,
  358.6493, 740.4105, 851.3992, 682.4423, 613.3671, 561.9201, 439.3097, 
    284.2988, 0, 0, 0, 0, 0, 164.7004, 99.19429, 101.628, 107.9559, 74.77886, 
    89.1244, 63.77163, 1.608809, -6.549558, -9.00685, -8.677175, -9.026371, 
    -3.706912, 1.230656, 51.11661, 139.9139, 209.1897, 282.7745, 328.7339, 
    305.7128, 303.4295, 269.2504, 220.6103, 194.5171, 252.9004, 301.2274, 
    362.1626, 362.2566, 319.3198, 217.928, 137.8181, 105.979, 105.6061, 
    114.0887, 135.0031, 185.067, 190.351, 191.2327, 234.4863, 323.938, 
    543.4288, 1060.478, 1268.447, 1192.681, 1328.727, 1228.022, 1216.701, 
    1586.167, 1872.411, 2054.413, 1874.194, 1613.623, 1458.215, 1250.402, 
    935.8388, 937.23, 1296.085, 1562.618, 1421.365, 1164.499, 1045.977, 
    969.0322, 885.1325, 801.2127, 811.7344, 891.5575, 953.3035, 938.8203, 
    644.8547, 285.5817, 157.9158, 154.0628, 172.5158, 282.7875, 469.8745, 
    706.7769, 1102.511, 1230.183, 277.3174, 0, 0, 0, 0,
  132.9001, 385.4105, 339.2654, 181.7644, 142.398, 0.8909621, 0, 0, 0, 0, 0, 
    0, 4.920471, 45.10483, 8.741613, 47.47253, 68.29308, 52.40722, 93.38539, 
    77.34655, 43.84061, 4.212869, 4.007848, 10.19131, 4.169814, 0.9422171, 
    9.296235, 56.39237, 118.7264, 170.1291, 210.7619, 320.4744, 331.2771, 
    318.584, 273.9849, 219.1942, 178.2944, 198.5368, 260.3773, 310.2903, 
    314.4893, 238.4738, 144.5557, 99.9539, 97.97208, 100.8626, 114.6869, 
    130.8342, 169.4516, 185.3304, 185.0731, 235.592, 278.8924, 478.6136, 
    764.5692, 685.5565, 811.843, 974.8875, 1184.866, 1309.973, 1492.49, 
    1975.901, 2111.276, 1920.701, 1584.152, 1393.754, 1227.47, 867.7672, 
    863.7648, 1180.989, 1434.811, 1408.729, 1119.982, 937.4036, 832.1047, 
    725.7586, 654.3876, 681.5729, 879.4352, 1001.297, 813.8375, 472.1414, 
    186.7852, 145.5977, 173.9421, 209.2027, 326.0379, 476.7007, 804.9005, 
    1109.927, 922.321, 75.55848, 0, 0, 0, 0,
  55.06753, 268.7123, 117.1969, 34.0993, 31.63307, 0, 0, 0, 0, 0, 75.30566, 
    123.2075, 25.73137, 4.677011, 0.4355646, 21.74989, 39.51146, 59.60038, 
    56.39664, 83.5396, 72.77475, 42.05199, 25.05266, 18.50826, 21.90979, 
    18.97606, 32.88521, 52.70894, 108.0705, 133.6327, 212.1806, 346.0227, 
    454.2986, 381.998, 286.2616, 211.4252, 172.9534, 157.5838, 173.7746, 
    195.4111, 173.0165, 139.0157, 104.9335, 99.12243, 103.3306, 100.5489, 
    103.4557, 134.8257, 162.8266, 185.8695, 232.4137, 269.2041, 308.7599, 
    614.8231, 747.6427, 544.698, 422.7588, 738.6674, 1183.856, 1471.337, 
    1606.683, 1839.523, 1757.208, 1367.475, 928.4243, 840.8771, 759.8136, 
    793.3425, 873.0726, 1079.337, 1313.67, 1351.702, 1047.42, 866.4039, 
    745.4284, 686.4276, 600.6986, 676.6058, 942.1893, 1006.475, 678.2116, 
    313.3897, 146.0503, 136.1638, 173.3874, 203.2215, 423.4491, 556.2217, 
    687.7593, 707.8784, 130.9646, 0, 0, 0, 0, 0,
  7.121133, 32.15426, 84.65013, 100.6684, 128.3299, 0, 0, 0, 0, 0, 37.53299, 
    141.1044, 20.04803, 0.0226125, 4.211974, 29.80108, 80.3756, 118.8334, 
    109.4529, 114.3332, 124.4319, 101.2349, 79.91515, 62.1116, 42.87167, 
    62.06577, 74.78121, 105.4743, 125.4183, 177.7379, 223.2901, 362.0724, 
    497.8951, 520.5967, 347.3084, 218.1198, 160.7832, 142.836, 141.2242, 
    142.3133, 130.3157, 119.2133, 114.2978, 107.0357, 102.9367, 104.6058, 
    110.6453, 123.0354, 142.3407, 155.8816, 175.0349, 218.0002, 336.6488, 
    481.0204, 622.3756, 464.2339, 567.8765, 821.3962, 1203.486, 1431.367, 
    1332.833, 1153.785, 908.6243, 652.9219, 598.5366, 569.8493, 665.6304, 
    778.8425, 895.4351, 980.2097, 1137.299, 1139.964, 917.5201, 727.8011, 
    697.3036, 645.4094, 611.8453, 750.6511, 997.3835, 898.4934, 452.9046, 
    187.9874, 131.9667, 132.1604, 162.3042, 257.2846, 519.6144, 578.7543, 
    534.0048, 299.177, 10.42934, 0, 0, 0, 0, 0,
  29.01102, 22.0339, 235.5383, 205.7878, 202.3339, 34.00895, 0, 0, 0, 0, 
    0.7499724, 39.96126, 8.142411, 27.61915, 77.46246, 141.4588, 165.7684, 
    167.3914, 132.9326, 131.5184, 138.1546, 130.3924, 147.073, 128.6659, 
    88.82133, 71.90593, 79.99207, 93.95091, 122.2475, 174.1009, 224.5994, 
    264.6025, 432.1731, 552.0823, 489.6333, 281.8752, 171.4949, 136.2069, 
    133.1193, 125.4225, 126.965, 120.7626, 111.4299, 101.8144, 99.97607, 
    113.2573, 118.6737, 130.7982, 136.456, 127.7007, 138.2258, 178.1324, 
    196.5107, 345.3022, 326.9236, 389.049, 456.8989, 544.9363, 644.9791, 
    795.9853, 714.1006, 626.2784, 512.6625, 545.9469, 686.3776, 774.8943, 
    722.8535, 808.6535, 999.6533, 978.3033, 988.0608, 965.1602, 774.5897, 
    743.5015, 720.1992, 658.6784, 645.7189, 780.3297, 934.1503, 668.8269, 
    269.4187, 138.0441, 142.1439, 151.7155, 169.5889, 303.9595, 540.4365, 
    608.5374, 528.3405, 294.674, 2.237589, 0, 0, 0, 0, 0,
  111.4144, 193.5326, 681.5145, 360.9993, 352.8302, 226.3572, 174.55, 
    37.86699, 0.2644904, 0.002788612, 0, 3.079878, 23.88782, 46.11481, 
    80.04777, 123.263, 147.1195, 144.2522, 130.5605, 152.2023, 141.6269, 
    132.931, 157.0246, 184.9375, 164.1916, 154.953, 124.2921, 92.66442, 
    103.1418, 164.1006, 233.3318, 178.8902, 210.3269, 409.1046, 418.7644, 
    336.8872, 189.2744, 130.1919, 111.7867, 105.783, 110.7427, 102.534, 
    94.83035, 91.60812, 107.021, 117.6856, 130.0774, 128.3777, 127.6499, 
    111.2988, 106.9357, 137.1521, 166.8579, 176.284, 241.0266, 287.8779, 
    322.1338, 316.6681, 333.3232, 405.2602, 465.2554, 453.8713, 526.2246, 
    631.4445, 775.7401, 794.0515, 706.1703, 873.7288, 1141.089, 1067.214, 
    1009.558, 878.1597, 765.5309, 814.0995, 825.5641, 682.4036, 688.0043, 
    821.9866, 793.0577, 482.589, 210.6379, 172.7338, 171.0665, 163.2869, 
    239.3744, 290.9917, 518.2194, 476.0343, 344.188, 253.0163, 199.3618, 
    0.09988576, 0, 0, 0, 0,
  396.4076, 461.4612, 931.6284, 727.4689, 459.6009, 316.0923, 161.0612, 
    61.08897, 39.84538, 14.21865, 16.21696, 14.69456, 42.59837, 83.79881, 
    96.42057, 106.7112, 127.726, 139.3746, 149.1176, 158.2953, 146.0142, 
    133.0698, 149.0564, 185.547, 219.5478, 236.7041, 204.2428, 142.1788, 
    111.0571, 152.1457, 197.096, 162.3448, 145.3164, 257.3849, 359.7718, 
    344.883, 231.0725, 134.1741, 96.72655, 77.17216, 67.97431, 71.95205, 
    78.97033, 92.42341, 106.5057, 121.7666, 113.3711, 112.7681, 100.1774, 
    90.3449, 93.89151, 126.1822, 144.4522, 167.8977, 184.3656, 222.1504, 
    216.4159, 276.5192, 273.3236, 330.4809, 405.03, 466.5895, 519.9902, 
    669.0401, 778.4682, 755.4747, 760.0569, 995.1483, 1292.865, 1133.658, 
    1035.321, 891.3419, 745.2759, 794.439, 820.8765, 731.4034, 825.5676, 
    816.8707, 654.7597, 365.2853, 254.1914, 241.2478, 251.6084, 300.0577, 
    283.1929, 314.035, 356.0846, 297.13, 224.8416, 403.2619, 439.1473, 
    0.3467962, 0, 0, 0, 0,
  855.1598, 709.2625, 1002.592, 837.1132, 519.1252, 130.5939, 71.12158, 
    81.11422, 142.1018, 51.00807, 96.93317, 79.51467, 95.48483, 129.0423, 
    140.4562, 103.5044, 126.4621, 151.7047, 177.8282, 174.2761, 156.9096, 
    144.2187, 154.5808, 180.015, 203.6465, 223.6183, 210.2678, 151.1036, 
    112.8854, 117.9561, 134.9364, 127.8695, 129.1225, 218.7797, 270.9187, 
    350.6521, 238.6366, 134.1218, 93.92628, 66.70253, 59.81225, 64.58974, 
    83.67481, 91.74277, 99.39961, 97.78426, 98.12943, 79.38904, 76.33865, 
    79.66943, 96.24992, 117.7307, 139.8467, 146.7351, 147.0995, 206.1468, 
    254.7715, 275.4333, 300.4858, 331.8605, 412.4602, 458.4528, 508.2016, 
    647.9883, 697.1085, 851.0264, 924.2222, 1209.887, 1389.744, 1105.53, 
    981.9774, 946.9201, 772.724, 746.0531, 774.8968, 822.0195, 896.6089, 
    762.1265, 469.3407, 356.1171, 319.8726, 356.8423, 393.546, 402.3568, 
    300.6212, 214.0752, 218.7073, 138.1364, 184.7563, 493.152, 362.86, 0, 0, 
    0, 0, 0,
  886.0403, 899.0963, 842.0179, 772.5779, 432.9344, 92.04449, 177.5087, 
    546.1584, 477.8832, 337.027, 119.8037, 133.9722, 151.3862, 176.6996, 
    157.914, 107.5661, 123.6268, 163.6318, 191.2482, 207.9477, 183.4089, 
    166.7186, 150.5348, 152.3792, 164.6893, 178.3489, 177.4384, 146.3247, 
    116.5272, 132.4336, 138.0589, 139.9558, 167.7014, 180.2253, 221.528, 
    303.055, 258.0195, 122.0804, 91.42705, 76.97997, 52.65008, 55.3461, 
    72.29636, 81.25592, 81.83448, 87.9664, 75.1608, 69.10935, 76.35617, 
    101.0703, 128.3883, 140.7466, 138.2242, 132.6284, 251.6389, 360.3346, 
    363.8312, 345.4504, 282.5562, 300.7509, 352.1882, 428.2724, 480.032, 
    508.1172, 638.3249, 969.0288, 1175.973, 1303.747, 1379.587, 1075.456, 
    939.7833, 971.2458, 876.7556, 679.537, 703.0974, 840.0677, 888.4769, 
    685.1582, 465.5422, 392.8445, 362.4918, 364.3657, 413.9269, 386.9064, 
    151.63, 102.4381, 140.1844, 97.34532, 357.6024, 508.7825, 100.0093, 0, 0, 
    0, 0.4358488, 0,
  377.0912, 777.9293, 847.1389, 613.7839, 347.3856, 183.928, 503.8705, 
    767.5604, 736.3063, 591.572, 261.3434, 142.1519, 203.053, 216.3297, 
    177.3449, 117.8392, 131.8621, 155.6192, 186.6643, 210.5387, 213.1024, 
    198.3484, 171.8902, 133.9252, 133.7206, 147.76, 149.0784, 123.2078, 
    117.5802, 128.9419, 142.8373, 162.3329, 190.3584, 196.8235, 191.6556, 
    277.8559, 336.0329, 136.4615, 78.44816, 67.13183, 57.19013, 45.63347, 
    56.64672, 62.35668, 62.41399, 58.50655, 64.08222, 61.68793, 82.98176, 
    109.022, 132.2926, 141.4133, 130.0148, 202.6298, 352.5894, 478.8041, 
    483.1053, 383.9174, 324.0171, 288.2619, 333.3291, 429.6476, 498.3948, 
    476.5586, 511.4784, 972.3265, 1117.176, 1333.446, 1231.988, 1100.885, 
    955.795, 961.8926, 865.2928, 707.8149, 605.3251, 700.6523, 739.4321, 
    558.5131, 402.4283, 297.584, 211.9652, 189.1523, 300.2366, 262.1036, 
    80.62009, 63.98812, 122.1838, 218.2967, 512.9334, 462.9636, 1.060671, 0, 
    0, 0, 37.38868, 81.3967,
  0, 594.21, 1018.811, 745.1058, 412.2401, 385.4236, 638.6064, 788.1194, 
    668.9521, 749.03, 562.7498, 197.1136, 243.5414, 257.3966, 197.9897, 
    130.8538, 123.876, 145.1576, 174.6566, 198.9581, 214.8165, 215.6441, 
    189.8338, 139.6603, 120.3094, 124.8503, 116.1674, 109.7017, 110.3707, 
    135.235, 142.0241, 170.4792, 213.9434, 209.5347, 167.4813, 264.8561, 
    348.0725, 240.3373, 75.87767, 79.91491, 71.83314, 45.36616, 48.33675, 
    52.77137, 49.97958, 59.72789, 63.37616, 71.72295, 88.81493, 109.8572, 
    136.8765, 144.6113, 151.7365, 193.6578, 319.4838, 403.0927, 398.4877, 
    411.3876, 349.0669, 324.9615, 351.6237, 448.8545, 494.1817, 457.7076, 
    444.8627, 679.2474, 972.8405, 1012.391, 1150.945, 1145.6, 1127.534, 
    944.8821, 822.8835, 703.0647, 531.0294, 464.5009, 428.4065, 363.7079, 
    263.4396, 211.7635, 198.9796, 267.8853, 350.3128, 264.7803, 65.758, 
    59.44502, 199.1785, 430.2982, 657.9562, 212.0221, 0, 0, 0, 97.63541, 
    113.3308, 41.61473,
  0, 399.1143, 1120.441, 820.4569, 297.3376, 195.9688, 434.3469, 519.7678, 
    533.1642, 758.1817, 711.3763, 342.4791, 278.5041, 278.4136, 214.2995, 
    149.314, 124.3232, 138.1995, 163.2455, 188.7315, 200.2267, 205.1242, 
    191.2654, 153.1303, 140.5527, 120.2366, 117.1466, 119.59, 127.6191, 
    134.2686, 149.6515, 164.0252, 186.4469, 196.4661, 161.6761, 177.2666, 
    334.9556, 307.35, 143.2057, 109.0354, 87.71973, 79.37965, 65.37148, 
    76.016, 76.0844, 78.8138, 85.20406, 92.65923, 120.6024, 124.1407, 
    141.3281, 120.2449, 152.1772, 252.603, 380.783, 423.7603, 464.9473, 
    420.7524, 383.9003, 365.9595, 382.3451, 404.967, 427.5276, 426.6728, 
    395.3827, 540.5605, 755.1957, 952.8699, 1084.376, 1365.629, 1383.233, 
    963.2598, 743.7776, 748.3361, 583.3853, 439.8699, 330.5274, 274.6473, 
    239.082, 218.2501, 375.178, 416.6259, 488.4598, 300.3638, 65.87481, 
    54.1222, 354.7472, 673.2607, 622.6516, 29.62266, 0, 0, 0, 206.3307, 
    149.5761, 0,
  0.003310259, 133.1911, 940.6332, 781.675, 248.0849, 90.08338, 116.6424, 
    220.5476, 304.2039, 419.5131, 703.8474, 411.9249, 301.6213, 267.3719, 
    209.3017, 160.7548, 131.8181, 134.4422, 157.0661, 185.6122, 207.0094, 
    210.453, 201.0542, 179.5661, 159.3497, 148.5723, 124.2159, 138.4398, 
    148.6608, 162.3591, 173.3146, 175.035, 184.1364, 181.5239, 173.0168, 
    157.8075, 250.5602, 304.8704, 179.2655, 67.08978, 85.99716, 73.47701, 
    103.1553, 107.7299, 100.9882, 96.31065, 80.26945, 83.55797, 94.24591, 
    113.5028, 87.01515, 83.67673, 216.3896, 356.1998, 462.2934, 496.7366, 
    464.9568, 424.9034, 395.8524, 405.8656, 396.2522, 369.3352, 362.0952, 
    392.2811, 403.4277, 532.8717, 897.1837, 937.3101, 997.2128, 1238.674, 
    1234.297, 916.9507, 798.6755, 785.5186, 683.3135, 527.7955, 404.3859, 
    329.3802, 251.766, 331.9852, 519.2047, 603.6315, 693.9681, 306.4999, 
    50.3644, 206.1701, 627.575, 741.8391, 292.8152, 0, 0, 0.002287545, 
    47.08162, 366.3271, 345.8133, 140.5091,
  0.1355318, 54.76622, 752.4495, 779.2272, 233.4452, 90.45777, 81.94717, 
    83.38457, 113.8429, 180.5548, 517.6541, 398.6514, 294.062, 222.6104, 
    177.3117, 146.8111, 135.3791, 142.748, 161.5963, 189.4258, 213.6966, 
    218.6755, 216.248, 169.9221, 153.2071, 133.3895, 136.4664, 149.2455, 
    169.6985, 177.9319, 169.0834, 158.8819, 153.8374, 154.3419, 155.6863, 
    159.3348, 168.2593, 263.9666, 210.4024, 63.44218, 42.57559, 53.28033, 
    74.75113, 94.46678, 84.90047, 77.8112, 56.29344, 41.15648, 64.81905, 
    77.03599, 86.15321, 102.1669, 314.0604, 390.679, 394.7146, 406.8066, 
    419.1735, 403.4146, 401.5237, 394.1876, 379.7701, 337.2509, 349.9233, 
    401.1396, 396.1155, 511.2408, 755.8575, 709.9775, 686.9054, 793.6512, 
    1004.453, 980.0493, 971.1741, 917.5543, 726.7474, 512.3557, 394.0262, 
    441.8013, 404.3204, 456.4452, 727.2965, 845.9907, 812.4409, 408.3134, 
    83.84931, 448.7415, 730.8319, 467.4902, 0.9863583, 0, 1.720724, 35.83591, 
    297.3234, 472.4654, 318.6473, 2.667824,
  2.786609, 2.644013, 504.1062, 684.3657, 243.8393, 124.4904, 120.2434, 
    118.8162, 136.5323, 274.2844, 459.7988, 323.3001, 252.3182, 197.7955, 
    158.2456, 143.8349, 155.14, 171.036, 179.7861, 181.361, 194.9534, 
    211.9559, 228.9097, 199.0386, 153.3901, 145.1039, 136.1797, 149.812, 
    166.3282, 157.6181, 154.2063, 126.907, 146.2792, 140.0006, 147.5358, 
    162.919, 152.3721, 222.5984, 246.1506, 256.06, 62.73549, 34.49001, 
    46.63019, 67.38826, 49.56528, 57.15746, 51.01564, 36.49106, 33.8912, 
    64.45266, 63.10199, 144.3528, 351.2276, 400.1565, 401.1474, 439.6917, 
    469.2003, 431.5126, 411.8654, 369.9917, 321.8169, 323.1301, 326.4559, 
    382.4082, 378.7637, 344.4705, 461.5488, 414.4735, 376.186, 542.0886, 
    713.6682, 832.4791, 967.1309, 1007.369, 852.7335, 704.9957, 550.9443, 
    581.854, 539.4864, 852.6191, 1003.918, 778.0033, 665.1097, 266.5093, 
    311.5761, 683.8643, 705.9689, 96.01817, 0, 1.189999, 8.842051, 47.33828, 
    140.6496, 324.6157, 137.269, 0,
  276.4731, 0, 179.3712, 525.0765, 251.7486, 132.691, 157.0414, 154.7416, 
    302.1239, 580.2548, 583.1707, 323.0918, 206.9382, 174.8136, 156.9467, 
    158.7047, 172.3876, 199.9602, 184.0974, 164.6234, 165.0962, 185.8372, 
    203.0004, 193.7835, 175.1679, 146.9807, 142.3714, 150.1652, 157.6037, 
    163.3478, 129.6109, 129.2951, 159.414, 161.3647, 162.9705, 181.9612, 
    128.0042, 147.4346, 353.2044, 345.6928, 272.2606, 81.65241, 31.30544, 
    29.65827, 24.55814, 44.82172, 50.73238, 36.99446, 29.24441, 45.64774, 
    56.69508, 147.8097, 350.2406, 446.015, 517.4972, 568.1435, 509.0543, 
    480.6918, 464.3664, 407.0969, 359.9652, 325.3537, 336.1723, 338.7549, 
    334.156, 299.1234, 313.2734, 332.2038, 383.9116, 472.8965, 632.2615, 
    813.0618, 1026.41, 1103.619, 1136.821, 1031.338, 975.8419, 689.2612, 
    568.7227, 943.745, 852.9982, 485.5357, 236.3455, 271.7433, 463.5656, 
    614.2126, 345.1251, 0, 16.48282, 105.6186, 7.521848, 0, 0, 87.10019, 
    40.73374, 0,
  508.8716, 70.13601, 6.784113, 372.3694, 322.6259, 293.2125, 242.353, 
    173.0082, 268.3181, 591.1161, 536.0643, 296.8539, 202.5906, 164.5604, 
    144.654, 150.5097, 161.7568, 165.6213, 170.2032, 147.5072, 145.3487, 
    118.8593, 111.2818, 111.6931, 136.4204, 155.4414, 171.5328, 140.8391, 
    169.3844, 138.0114, 124.348, 104.4207, 145.8794, 164.8125, 186.8414, 
    188.481, 126.0499, 90.26923, 110.4248, 252.1565, 185.2361, 152.9825, 
    177.3863, 27.33101, 14.74302, 22.59383, 32.78283, 24.52886, 36.56748, 
    50.80676, 80.63863, 201.0317, 398.6272, 570.3611, 631.2753, 643.4182, 
    537.705, 514.1293, 540.4216, 502.6988, 444.1647, 409.5107, 358.6469, 
    313.3456, 229.5331, 227.212, 262.0572, 326.5652, 403.6352, 469.1498, 
    543.0381, 673.6775, 820.8776, 1047.744, 949.5495, 1148.552, 1111.228, 
    855.2848, 484.6896, 661.6188, 513.8441, 249.184, 299.0674, 415.421, 
    493.6745, 252.4404, 5.99207, 59.10885, 97.5045, 79.21317, 10.46941, 0, 0, 
    43.29576, 3.355622, 0,
  443.5912, 255.1915, 0.09644534, 195.873, 487.8073, 735.0255, 695.2324, 
    348.3268, 280.6532, 412.6371, 385.954, 220.2776, 204.6375, 127.3774, 
    125.8829, 139.0522, 124.0497, 124.0424, 125.5306, 122.1397, 132.0455, 
    96.83639, 60.97416, 63.26183, 70.19158, 96.56532, 138.9745, 127.6716, 
    134.1593, 150.0386, 90.46266, 84.52273, 112.2292, 121.4295, 151.5019, 
    166.1176, 108.1869, 79.91405, 92.42285, 97.96801, 124.7679, 221.8664, 
    228.2843, 115.3288, 24.56494, 14.8802, 20.65261, 31.73664, 49.24442, 
    60.99174, 105.08, 244.0706, 521.9723, 723.241, 767.3787, 664.4177, 
    487.5122, 513.0247, 515.0753, 538.3448, 511.0675, 463.2043, 376.3399, 
    264.3518, 201.9225, 193.3568, 293.2623, 334.261, 373.6343, 439.8721, 
    490.5887, 493.9969, 600.4854, 755.9476, 924.3199, 950.3077, 1052.388, 
    779.1483, 183.5563, 265.7245, 179.8311, 213.6126, 282.3783, 202.5462, 
    128.2361, 30.74742, 219.925, 102.526, 0, 0, 0, 0, 0, 16.26684, 0.6956787, 0,
  260.7036, 393.7766, 11.27141, 23.8249, 678.2915, 1205.305, 983.3217, 
    600.5497, 405.7943, 426.7081, 384.4165, 217.486, 141.1087, 113.0105, 
    118.703, 126.1676, 90.83533, 74.9175, 85.22266, 86.1847, 108.5499, 
    97.74491, 85.57736, 64.07814, 40.13272, 24.09916, 78.24743, 80.76043, 
    124.5104, 132.6886, 90.25305, 50.69267, 81.38572, 64.80839, 89.60198, 
    115.1036, 102.3747, 89.09599, 91.98434, 106.8285, 90.62163, 137.0851, 
    183.7695, 40.38134, 27.67106, 11.31515, 23.2658, 37.70986, 46.24703, 
    62.2045, 86.09678, 336.5412, 717.0566, 919.0491, 854.2428, 596.1452, 
    380.2888, 384.9098, 468.5178, 498.7417, 522.8006, 451.6152, 351.5222, 
    233.9609, 161.0052, 184.1114, 234.4022, 294.4582, 302.137, 342.4128, 
    411.9693, 392.7577, 351.6703, 590.9839, 653.2507, 725.2677, 801.4582, 
    656.3619, 55.66471, 28.70166, 97.66091, 137.6178, 146.7572, 75.24693, 
    99.51981, 291.1764, 193.6622, 6.543282, 0, 0, 0, 0, 10.53877, 52.14492, 
    0, 0,
  43.77597, 464.1584, 56.89383, 468.3003, 1272.138, 1580.384, 1018.172, 
    560.8243, 492.4376, 414.2195, 387.2528, 175.9947, 96.38813, 88.09875, 
    109.2793, 71.96533, 25.01822, 58.2986, 73.01802, 38.57325, 49.70271, 
    62.90857, 57.06133, 27.90662, 27.32676, 23.32841, 78.08787, 112.5397, 
    118.9064, 113.533, 66.1688, 38.50869, 78.81353, 50.76294, 38.3057, 
    62.43602, 80.58298, 45.74772, 40.23263, 38.5184, 22.24349, 97.94888, 
    42.41491, 12.44253, 28.08678, 14.85801, 30.86785, 37.11079, 35.73439, 
    33.91776, 124.3871, 381.5867, 780.6381, 921.0138, 807.3401, 514.1893, 
    283.6758, 323.1736, 314.6895, 374.642, 395.0815, 392.9985, 310.7736, 
    226.0156, 184.2313, 147.4343, 164.883, 202.6225, 252.7558, 260.424, 
    307.9431, 309.5395, 311.4832, 401.2553, 517.3415, 550.1964, 679.3637, 
    525.896, 1.616105, 2.896513, 88.79086, 59.5556, 70.75466, 69.71838, 
    122.3319, 154.2911, 15.59744, 0, 0, 0, 0, 0, 27.71455, 6.569491, 0, 0,
  0, 439.4178, 195.6855, 907.5368, 1805.264, 1501.639, 712.643, 483.2295, 
    497.7593, 420.5321, 315.0768, 136.8431, 80.70911, 102.5947, 110.8975, 
    56.06786, 0.2648131, 3.387826, 36.63493, 22.48626, 4.213938, 32.13628, 
    34.12004, 9.394886, 55.34244, 71.22887, 124.1325, 164.2337, 141.1722, 
    73.3173, 29.08077, 2.917876, 50.12897, 16.72008, 8.767165, 20.09276, 
    6.12492, 9.995467, 2.303684, 0.02967453, 7.202766, 15.59999, 0, 4.923676, 
    28.76822, 14.64493, 19.81721, 22.2378, 29.72172, 55.51414, 46.22926, 
    135.3196, 311.9851, 389.0701, 426.3514, 394.7778, 346.0056, 381.4013, 
    311.8159, 286.077, 316.2218, 321.0644, 306.4557, 227.0812, 163.6294, 
    111.7403, 127.4932, 171.2171, 128.8476, 186.4454, 234.3389, 277.8444, 
    263.8623, 387.7439, 507.9923, 593.5289, 671.5868, 151.9244, 0, 0, 
    0.1526855, 11.12141, 27.27045, 5.642293, 0, 0, 0, 0, 0, 0, 0, 0, 
    29.69389, 0, 0, 0,
  336.1212, 283.2744, 280.2505, 1349.746, 1791.143, 1240.253, 581.5303, 
    454.5894, 529.9597, 451.9621, 271.3024, 88.98106, 65.69213, 79.26176, 
    83.76402, 15.86282, 0, 0, 0, 0.01159282, 3.559813, 3.361201, 26.5549, 
    78.995, 104.8708, 111.296, 123.7502, 183.7094, 170.4765, 96.75568, 
    18.82452, 36.92904, 173.0009, 147.0736, 0.6561724, 40.09827, 1.400087, 
    18.67419, 0, 4.921213, 17.68606, 0.02064603, 0, 0.5728964, 18.75198, 
    13.3812, 8.656983, 8.488718, 38.44683, 61.09453, 51.83106, 52.62397, 
    58.6014, 59.39347, 165.6035, 290.221, 454.3603, 531.7468, 356.0366, 
    250.5548, 230.6507, 267.4886, 263.0035, 170.9993, 101.3395, 226.0812, 
    405.6003, 438.8228, 243.4076, 140.5213, 194.1314, 222.0123, 325.5292, 
    476.0626, 621.8958, 708.6229, 614.3857, 5.007009, 0, 0, 0.5131387, 
    10.68596, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 30.96639, 0, 0, 0,
  1014.961, 1059.676, 999.4585, 1486.217, 1353.48, 822.1008, 483.4728, 
    423.429, 432.9811, 400.1913, 184.7545, 59.76541, 51.08024, 32.45238, 
    3.397727, 1.339373, 0.5192116, 1.949396, 6.878533, 0.8359628, 0, 
    0.4469217, 32.46057, 94.17204, 138.7826, 139.0123, 142.075, 170.2651, 
    199.8437, 156.3874, 66.95568, 99.59976, 214.9215, 163.2938, 0, 
    0.00557197, 0, 0, 0, 37.75103, 85.04147, 0, 0, 0, 2.593199, 6.704577, 
    0.9132928, 2.0938, 109.5198, 89.66087, 71.78169, 61.52934, 55.7276, 
    50.0367, 66.96713, 204.8958, 385.6734, 415.6871, 273.868, 163.4537, 
    185.3572, 235.6016, 183.325, 121.5506, 331.4378, 656.7086, 973.7778, 
    936.9366, 698.6102, 315.4651, 158.0312, 304.8352, 599.1711, 767.9793, 
    739.1931, 587.2299, 272.567, 0, 0, 0.0005063568, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.3449626, 0.8638448, 0, 0, 0,
  1276.519, 1596.647, 1710.525, 1532.737, 942.0485, 525.4172, 468.8974, 
    340.8898, 335.7376, 367.5742, 202.7082, 87.97628, 47.15509, 23.6611, 
    2.109894, 16.11546, 63.89506, 99.67946, 35.14595, 6.804534, 11.33926, 
    3.489694, 4.426375, 51.48684, 116.296, 132.7959, 119.1194, 141.0041, 
    206.496, 213.7981, 189.8233, 189.694, 225.2005, 137.5171, 0, 0, 0, 0, 0, 
    51.36637, 209.3645, 35.64569, 0, 0, 0, 0.1678525, 0, 0, 2.154153, 
    17.08876, 89.85088, 131.7713, 127.0772, 66.14963, 54.64122, 98.0938, 
    154.5197, 216.6144, 122.0288, 144.2869, 194.6717, 195.0684, 113.4059, 
    305.1859, 773.1769, 944.6837, 944.9396, 1041.262, 1010.897, 714.8572, 
    441.2517, 615.52, 994.8956, 1017.131, 735.3895, 398.553, 39.48136, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16.48005, 0, 0, 0, 0,
  576.1854, 931.6247, 906.6362, 782.9591, 492.1016, 465.3861, 284.8566, 
    247.166, 278.3712, 328.5902, 197.9191, 70.77742, 37.59184, 12.53315, 
    7.181137, 43.26176, 121.2297, 201.0618, 133.2232, 65.32127, 50.51119, 
    18.33489, 0, 0.11232, 20.32129, 27.82987, 23.76683, 29.30825, 141.2721, 
    243.3896, 253.101, 230.2507, 183.3705, 51.35647, 0, 0, 0, 0, 0, 0, 
    70.44017, 221.9524, 66.5798, 0, 0, 0, 0, 0, 0.3017679, 8.757327, 
    127.2703, 222.3685, 176.8489, 129.8425, 56.31729, 30.53881, 53.13721, 
    56.63842, 85.90793, 110.0528, 170.028, 155.7422, 181.1576, 658.582, 
    891.925, 765.0097, 566.7166, 683.1484, 938.3599, 946.0663, 950.6962, 
    1152.784, 1400.864, 1190.112, 699.8245, 303.8513, 1.38781, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 4.373055, 0.3063857, 0, 0, 0, 0,
  645.5978, 651.4741, 348.0461, 338.1821, 333.729, 297.324, 274.5483, 
    329.6071, 320.4292, 242.4523, 142.7768, 33.2918, 19.17206, 13.50416, 
    14.204, 8.873847, 37.03663, 147.5774, 138.1909, 116.1385, 174.9569, 
    163.6211, 73.71962, 29.18241, 51.88186, 92.01063, 38.92251, 26.84706, 
    114.0117, 203.6541, 270.5715, 215.7726, 151.7382, 14.68677, 0, 0, 0, 0, 
    0, 0, 0, 40.54074, 369.3293, 317.3165, 114.3371, 3.862887, 0, 0, 0.11153, 
    0.006048144, 19.55387, 142.5781, 154.5665, 123.9076, 179.1985, 79.16, 
    14.5393, 34.07465, 42.74265, 97.64807, 169.0159, 219.1613, 396.9012, 
    642.2534, 732.5916, 397.1309, 377.0508, 643.4995, 985.1297, 1109.908, 
    1146.201, 1363.316, 1434.265, 1369.427, 928.765, 436.3409, 111.6556, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5.772016, 0.006933623, 0, 0, 0, 0, 0,
  832.0802, 796.4195, 452.5931, 305.7719, 293.3802, 263.662, 251.0075, 
    350.6158, 214.3606, 118.4772, 23.99523, 9.823727, 0.9374197, 9.133391, 
    30.28316, 31.31364, 7.673902, 30.12636, 73.6406, 163.2412, 282.5515, 
    383.3724, 343.9316, 270.9898, 269.3295, 315.7319, 274.4701, 208.2753, 
    218.7913, 263.5744, 306.8953, 271.2532, 182.3894, 67.36945, 0, 0, 0, 0, 
    0, 0, 0, 0, 5.676641, 71.09753, 100.5261, 93.03223, 0, 0, 0, 0.029983, 
    0.2834589, 5.7791, 29.0103, 202.0174, 299.2979, 245.8783, 10.45641, 
    3.441845, 9.227307, 65.13091, 143.5608, 212.5292, 258.0329, 406.613, 
    314.3367, 276.2676, 445.5888, 781.3271, 1096.255, 1218.235, 1079.923, 
    998.8617, 1214.761, 1232.076, 1011.277, 597.6057, 136.1366, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 2.308824, 17.42456, 0, 0, 0, 0, 0, 0,
  522.8505, 646.8199, 434.2559, 254.1983, 198.1381, 141.3106, 157.4017, 
    202.436, 98.83956, 4.720938, 5.80146, 1.222248, 0.002537446, 0, 6.751021, 
    16.09051, 4.110047, 0, 67.87675, 217.9813, 406.6455, 577.1392, 615.5616, 
    464.1506, 415.4912, 491.5859, 515.1653, 499.5445, 526.2872, 472.2782, 
    484.1233, 346.7195, 209.6823, 28.12877, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.04541712, 0.1208085, 35.22072, 93.14128, 169.8435, 
    92.35309, 0, 0, 0.01013316, 4.865694, 16.84927, 23.22182, 27.02969, 
    119.0616, 246.3213, 518.4421, 657.4585, 736.8021, 1052.213, 1052.852, 
    1112.684, 1157.132, 1119.51, 1128.288, 975.9925, 711.0227, 271.4639, 
    11.86194, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10.20065, 51.1852, 0, 0, 0, 0, 0, 0, 0,
  189.5987, 372.6584, 272.8972, 153.0684, 129.0797, 107.2802, 101.2548, 
    98.52764, 13.1368, 0.6186931, -0.0932398, 0.01887309, 0, 0, 0, 0, 
    5.934471, 249.3546, 496.3241, 641.0406, 712.6684, 883.3423, 769.7581, 
    568.9565, 546.6921, 654.5696, 742.6288, 773.7735, 770.8872, 664.8349, 
    517.9086, 240.3035, 48.13427, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 25.80465, 75.88532, 127.7064, 5.597481, 0.01321575, 0.01744381, 
    0, 0, 0, 0.008600875, 0.2463465, 0, 3.196367, 26.82889, 218.4336, 
    438.3653, 500.2625, 445.5697, 536.2654, 907.6587, 1133.265, 1245.885, 
    1148.132, 918.5613, 905.1179, 873.1757, 565.6349, 139.6936, 9.307497, 0, 
    0, 0, 0, 0, 0, 0, 5.973339, 51.01183, 18.53154, 0, 0, 0, 0, 0, 0, 0,
  66.53913, 126.0707, 158.3924, 101.3495, 129.9872, 153.1423, 111.0585, 
    69.88337, 5.909921, 0, 0, 0, 0, 0, 0, 0, 6.110831, 443.8941, 822.0618, 
    1065.257, 1147.54, 1026.579, 615.9289, 217.0476, 161.5421, 240.8548, 
    308.3307, 226.1226, 224.5132, 167.3122, 91.86687, 2.702835, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 1.687579, 0, 0, 0, 0, 2.009178, 150.2296, 
    137.6718, 53.3191, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01111945, 8.059679, 
    76.88058, 223.2468, 192.0626, 54.48991, 351.7439, 523.5924, 854.4131, 
    841.848, 774.7855, 709.6036, 701.8489, 900.449, 776.0449, 283.2952, 
    20.40456, 0, 0, 3.21502, 41.93052, 145.8842, 257.1946, 238.5102, 
    233.1759, 92.08567, 0, 0, 0, 0, 0, 0, 0, 0,
  10.54719, 38.52236, 89.41316, 88.45621, 129.8748, 140.0378, 1.758609, 
    3.622372, 20.79722, 16.84281, 3.764497, 0, 0, 0, 0, 0, 0, 9.974582, 
    203.0671, 552.9215, 723.358, 628.1764, 114.8102, 1.827135, 0, 0, 
    0.02597354, 4.145141, 11.91014, 1.813728, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 2.070437, 19.12915, 65.26246, 40.89855, 0, 1.946335, 0.4316256, 
    4.962647, 138.3129, 0, 0, 0, 0, 0, 0, 0, 0, 0.7391827, 0.9985219, 
    0.398542, 4.360011, 16.71775, 12.17988, 71.93053, 79.30731, 98.12679, 
    133.4162, 234.3277, 244.6326, 294.9109, 406.4966, 458.4559, 607.9581, 
    806.5295, 651.6235, 97.59635, 26.42796, 0, 11.91634, 142.9294, 523.1003, 
    623.8453, 728.3721, 414.541, 179.0205, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0.2375568, 35.22453, 45.78533, 100.8335, 98.73385, 0, 19.24257, 
    69.95895, 49.19936, 14.10529, 0.5963095, 0, 0, 0, 0, 0, 0, 0, 14.52876, 
    100.917, 29.60974, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.002305, 0, 0, 
    0.049075, 0, 0, 0, 0, 10.97873, 31.62269, 20.17602, 8.189528, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 24.33025, 35.88162, 3.392136, 8.202249, 
    9.667623, 4.784458, 29.97687, 95.48793, 70.86581, 107.1511, 47.01993, 
    186.0479, 250.5408, 327.3635, 495.9941, 663.1337, 707.337, 343.3452, 0, 
    0, 12.89661, 177.2778, 526.8167, 650.3031, 730.8545, 475.256, 140.5307, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0.1563355, 32.96153, 93.6973, 8.055909, 7.271522, 46.84789, 107.1797, 
    96.87433, 65.0823, 5.47474, 1.638984, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 46.7029, 45.70561, 2.701415, 
    1.950268, 1.063997, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1.490511, 10.38847, 0.8451264, 0, 0.1427283, 5.747555, 26.19526, 
    79.84738, 54.79946, 32.89713, 97.37908, 252.4611, 375.3538, 398.1776, 
    596.9442, 749.3185, 517.8513, 3.130794, 0, 0, 92.81933, 348.3482, 
    500.1969, 715.4668, 515.3165, 78.95136, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 23.82193, 117.2348, 1.692671, 2.966081, 75.61375, 119.2401, 
    156.9432, 150.2247, 187.7098, 168.4926, 20.22646, 0, 0, 0, 0, 
    0.008525716, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 112.4393, 
    187.7537, 277.7043, 196.2434, 63.29765, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0.6239529, 13.39494, 0, 0, 0, 1.266546, 41.70436, 
    25.22967, 28.20456, 109.732, 279.7055, 394.6047, 507.9118, 776.3243, 
    775.1523, 364.5099, 50.67634, 5.433064, 185.3506, 421.2495, 414.1049, 
    393.2517, 297.5771, 294.7875, 7.586363, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 2.931184, 22.6025, 0, 26.93795, 109.4093, 139.878, 177.1416, 
    88.31774, 86.30247, 174.0245, 163.1162, 240.8645, 75.69065, 3.21588, 
    0.5801046, 6.936382, 0.1045908, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 1.200257, 139.026, 418.142, 149.2554, 1.2402, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.164914, 0.7948571, 0, 0, 0, 
    0.001168255, 16.67364, 19.89136, 43.50631, 130.2915, 266.5667, 415.8081, 
    554.9022, 713.0673, 638.9822, 273.1252, 216.0703, 123.0732, 400.6276, 
    240.1565, 113.1827, 94.77327, 41.31813, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 12.43825, 0.1656403, 16.24762, 3.12718, 2.06611, 
    13.84467, 122.0781, 227.2487, 363.1719, 217.4649, 58.97001, 0.598401, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4.693333, 86.21237, 
    0.054159, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    9.497975e-05, 0, 0, 0, 0, 0, 4.237197, 6.721555, 63.53002, 114.1027, 
    265.6567, 554.0557, 724.3539, 712.1773, 539.7785, 160.6944, 68.24227, 
    103.9293, 73.31152, 28.09826, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0.03340246, 0, 4.537661, 95.45872, 73.8838, 90.62366, 
    59.25259, 54.20035, 152.8858, 94.76863, 8.248804, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1057689, 19.82886, 
    233.0814, 269.9969, 373.4673, 617.0306, 770.7498, 660.8774, 426.0227, 
    199.58, 211.4468, 198.4001, 14.72842, 0, 0, 0, 0, 15.84741, 3.091941, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 68.96684, 105.0802, 102.1657, 102.4648, 46.12123, 
    0.1862036, 4.137225, 14.37615, 0, 0, 0, 5.570907, 19.88484, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1777319, 
    320.2881, 508.4323, 575.6027, 669.407, 672.3879, 490.291, 289.8031, 
    238.265, 313.8378, 200.7386, 9.265935, 0, 0, 0, 0, 0.1091187, 4.402359, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0.1957944, 113.7033, 75.3949, 52.71202, 37.44812, 
    0.2004635, 0, 0, 0.123569, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    13.78675, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5.807943, 138.4678, 
    425.4565, 693.1362, 582.7962, 419.3349, 270.5754, 275.724, 489.4667, 
    545.7513, 206.3423, 1.7709, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 20.8598, 0.006193054, 2.341495, 0.4137827, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.4644903, 19.146, 0.3230906, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 76.46013, 93.74072, 366.0079, 
    496.2035, 424.2791, 175.4117, 154.8367, 347.1221, 670.9517, 666.6006, 
    261.9197, 13.65668, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6.259748, 
    120.2423, 2.125335, 0, 0, 0, 0, 0, 0, 0, 0, 0.5916959, 0, 2.078349, 
    11.29419, 52.72276, 269.5899, 324.7525, 54.04507, 40.68792, 0.01734185, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    27.23831, 326.5949, 448.5767, 470.8265, 265.0998, 97.36693, 175.0721, 
    356.4594, 464.9758, 296.394, 24.18855, 0, 0, 0, 0, 0, 0, 0, 0, 6.498864, 
    0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 434.9876, 
    549.625, 194.8289, 0, 0, 0, 0, 0, 0, 0, 49.79148, 229.9053, 270.3666, 
    218.3152, 435.0714, 763.8671, 711.7297, 577.2573, 432.7135, 282.8728, 
    35.13057, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 9.57939, 23.93509, 458.746, 758.4965, 540.113, 253.5558, 102.6653, 
    138.8913, 305.0443, 234.599, 15.73475, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    26.66078, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7.860931, 
    705.9603, 764.272, 264.1802, 0.009830754, 0, 0, 0, 26.49382, 30.51307, 
    107.7551, 497.813, 1169.735, 1488.845, 1487.634, 1470.97, 1528.288, 
    1292.458, 1079.739, 876.5819, 425.0653, 38.33871, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9.993676, 78.49228, 0, 
    302.9012, 626.1432, 557.4089, 253.4888, 65.42033, 56.02234, 195.751, 
    71.06109, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.04533782, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 39.38756, 
    486.9271, 529.4836, 132.7024, 0, 0, 0, 188.4812, 192.5964, 498.543, 
    708.6475, 1124.227, 1743.003, 2079.127, 2174.609, 2030.333, 2037.837, 
    1968.742, 1794.981, 1306.613, 536.4325, 38.71229, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.2987449, 0.9965169, 0, 
    24.91258, 299.2193, 349.5217, 135.9241, 25.71449, 1.858234, 83.3325, 
    37.25776, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.5446421, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.008149051, 
    79.37028, 181.9968, 190.1527, 16.7675, 0, 13.55061, 980.6506, 768.5872, 
    1105.977, 1530.174, 1995.253, 2289.703, 2406.146, 2417.229, 2295.283, 
    2278.623, 2349.081, 2062.894, 1572.461, 794.2656, 199.4317, 65.12003, 
    90.86436, 1.968355, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 58.45197, 215.2836, 156.8912, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 1.912825, 3.799026, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    10.55764, 11.55569, 0, 0, 140.3663, 1585.396, 1665.679, 1860.954, 
    2327.909, 2685.942, 2719.711, 2651.773, 2599.41, 2509.09, 2444.553, 
    2411.1, 2231.088, 1777.786, 1073.075, 389.2512, 394.257, 742.5377, 
    431.4628, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 6.323763, 161.9636, 163.3663, 42.97362, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.2813061, 5.751188, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 162.3825, 1830.881, 2420.234, 2799.512, 2933.921, 3054.115, 
    3021.108, 2897.282, 2813.163, 2631.317, 2454.22, 2377.28, 2253.893, 
    1763.675, 967.3515, 294.468, 567.5514, 896.8688, 723.8139, 165.1352, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22.55821, 
    205.1908, 176.4454, 100.5338, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5.576109, 1.351869, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 224.3244, 1715.302, 2661.883, 3042.112, 3078.042, 3083.966, 
    3056.699, 2966.114, 2775.983, 2461.252, 2203.078, 2069.804, 2055.312, 
    1617.411, 858.8635, 63.53865, 565.2546, 820.6309, 464.1451, 208.9816, 
    21.89472, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.308722, 
    41.45142, 0, 0, 39.56498, 1.861557, 0.9454954, 8.430882, 0, 0, 0.2580895, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 15.21186, 1.925179, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 69.28409, 1442.782, 2432.051, 3022.305, 3064.017, 2982.046, 2920.952, 
    2867.871, 2768.787, 2520.354, 2211.113, 1641.312, 1364.499, 1291.194, 
    1387.434, 845.2209, 244.3112, 296.0118, 614.2589, 358.0775, 523.442, 
    111.5307, 0.1241507, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6.110101, 52.63713, 243.9889, 184.6683, 0.4007951, 7.643325, 46.26271, 
    0.01746987, 11.53573, 9.214417, 0, 0, 2.880076, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 20.27884, 0.2822629, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 388.4866, 1897.231, 2823.74, 3016.014, 2869.568, 2752.483, 2647.189, 
    2529.865, 2443.268, 2159.798, 1604.969, 955.6561, 423.3286, 422.3328, 
    778.8141, 553.3457, 156.9905, 464.2124, 635.9963, 351.1034, 437.6381, 
    20.91868, 26.49133, 1.27366, 1.299142, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 3.944896, 32.97338, 270.1112, 460.1797, 328.6203, 29.76436, 98.42758, 
    162.2669, 21.47914, 0.01439463, 0.09217066, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.01224168, 16.85926, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 220.2471, 1591.738, 2466.678, 2747.279, 2660.819, 2426.795, 2163.563, 
    1904.25, 1726.834, 1309.499, 717.4695, 72.1908, 0.01969476, 0, 139.6303, 
    56.38565, 0.01733694, 280.8316, 373.5753, 88.71832, 60.37281, 22.64031, 
    35.58979, 1.627476, 11.44019, 3.820878, 2.149208, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.01889744, 6.854713, 95.4062, 415.7192, 609.9531, 237.4828, 87.95111, 
    174.6365, 179.5905, 1.821839, 0.4608677, 1.038414, 1.955436, 0, 0, 0, 0, 
    0.4032466, 0, 0, 0, 0, 0, 23.75265, 6.992056, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 344.95, 1579.479, 2305.747, 2500.39, 2205.512, 1810.193, 1200.209, 
    851.3199, 495.871, 307.6716, 18.7188, 0, 0, 0, 0, 0, 0.007190464, 
    328.6132, 334.6894, 151.1666, 47.72522, 19.96992, 2.669097, 2.000999, 
    5.087904, 39.56742, 29.48166, 1.290598, 0, 0, 0, 0, 0, 0, 0, 0, 7.210662, 
    34.74933, 341.6028, 763.1323, 677.7067, 334.8472, 120.0849, 233.7542, 
    94.9697, 21.47264, 47.76735, 13.35156, 8.629306, 32.41949, 2.232151, 0, 
    0, 0, 1.06906, 0, 0, 0, 0, 12.63473, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    220.6236, 1349.775, 2132.709, 2395.235, 2048.53, 1480.806, 855.7775, 
    314.9611, 477.5641, 130.0667, 3.648897, 0, 0, 0, 0, 0, 0, 10.08162, 
    642.4855, 281.7012, 101.1102, 60.59174, 61.11189, 54.33709, 36.61767, 
    64.51082, 191.8937, 50.27359, 0.1158935, 0.7644691, 0, 0, 0, 0, 0, 0, 0, 
    127.1192, 404.733, 737.6123, 874.3842, 641.8504, 235.5844, 192.8914, 
    214.4153, 206.9348, 198.1494, 125.9625, 26.56938, 2.941694, 5.601278, 0, 
    0, 0, 0, 0, 0, 0, 0, 4.25005, 1.223589, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    123.0767, 1440.606, 2345.219, 2595.379, 2201.878, 1579.878, 765.6243, 
    263.2791, 17.18813, 95.84882, 0, 0, 0, 0, 0, 0, 0, 18.90151, 14.24182, 
    240.224, 244.171, 170.7711, 72.88946, 36.88171, 3.688538, 30.90802, 
    42.64079, 82.76118, 41.20324, 110.692, 64.07503, 0, 0, 0, 0, 0, 0, 
    116.6442, 851.2905, 1040.522, 1011.616, 761.973, 391.5457, 285.8691, 
    222.6031, 231.2289, 132.9321, 127.5657, 79.20253, 79.93398, 60.85431, 
    7.069205, 0, 0, 0, 0, 0, 0, 0.002840273, 31.90177, 12.23519, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    113.4006, 1133.138, 2195.308, 2608.468, 2239.793, 1572.94, 1003.211, 
    518.9925, 189.4889, 0.6126093, 0, 0, 0, 0, 0, 0, 0.1651795, 133.9569, 
    417.8274, 384.9297, 215.625, 141.7358, 90.05803, 79.19399, 29.33371, 
    2.240706, 12.30619, 0.2534847, 0, 94.7438, 162.481, 149.9046, 37.89026, 
    0, 0, 0, 0, 5.356696, 552.9598, 964.9863, 891.923, 640.1644, 439.5914, 
    361.2435, 278.5941, 283.0451, 244.8269, 280.0539, 219.772, 241.4119, 
    332.4167, 319.8716, 147.7597, 7.835948, 0, 0, 0, 0, 0.3774112, 84.49905, 
    37.25802, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 30.39107, 
    914.6385, 1832.73, 2461.096, 2238.884, 1490.557, 718.7988, 432.395, 
    372.0842, 0.9015442, 0, 0, 0, 0, 0, 105.8306, 357.3896, 523.8076, 
    521.7178, 440.9008, 328.9724, 202.1082, 166.6164, 82.55063, 126.2423, 
    70.6189, 12.28226, 42.67114, 60.72597, 91.16128, 142.8304, 148.7395, 
    152.2123, 97.86357, 0, 0.3341298, 0.6432131, 4.719822, 37.05452, 468.78, 
    599.9188, 399.7013, 211.5083, 353.3973, 316.7687, 280.8083, 341.3538, 
    511.3751, 442.6859, 504.624, 253.1497, 250.1017, 213.2764, 67.04365, 
    3.304585, 0, 0, 0.1683532, 53.87643, 48.47186, 10.75609, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 89.8662, 
    469.3024, 1154.713, 1449.781, 1272.478, 681.3491, 128.84, 4.544834, 0, 0, 
    0, 0, 0, 5.419511, 61.07015, 489.1122, 578.3217, 527.3911, 395.0327, 
    218.0269, 167.6713, 137.974, 115.5373, 0.6435879, 88.33016, 45.21404, 
    6.509036, 44.30594, 115.2863, 242.208, 245.5465, 151.2771, 0.4254271, 
    11.1162, 1.786039, 48.14689, 37.55202, 70.14665, 156.7791, 498.9786, 
    523.2408, 473.1295, 354.968, 545.134, 489.5596, 703.8699, 925.6036, 
    986.3214, 886.7418, 869.757, 604.8533, 197.4831, 113.1076, 12.6825, 0, 
    0.02486209, 6.962315, 96.1065, 54.04581, 0.01545697, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.1216824, 0.9288862, 134.0087, 201.5549, 60.90172, 0.3555474, 0, 0, 0, 
    0, 0, 355.5598, 602.0829, 651.0312, 450.9958, 386.381, 256.653, 158.6886, 
    43.34907, 61.85168, 159.5036, 113.3953, 25.31179, 87.31884, 165.2257, 
    4.966446, 0.1061549, 45.43877, 108.6841, 188.0823, 174.495, 113.4314, 
    0.01686891, 145.4191, 132.487, 172.8789, 193.6581, 150.9564, 166.1918, 
    400.6677, 583.3967, 722.2389, 745.6167, 800.6808, 849.4872, 1009.411, 
    1053.753, 947.8483, 415.5219, 584.1187, 491.2827, 259.1023, 215.041, 
    112.3413, 76.86075, 134.8813, 221.4578, 45.61331, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 3.875198, 477.9095, 533.1882, 461.8639, 235.7978, 
    111.7738, 22.34331, 6.797899, 1.574463, 51.39446, 134.1712, 4.203103, 
    6.980784, 108.1984, 118.4102, 3.881124, 11.86376, 72.39351, 102.465, 
    159.5778, 156.6727, 107.9339, 109.4576, 488.6499, 418.6319, 300.2693, 
    237.9754, 185.1014, 104.7926, 403.3925, 659.502, 1010.157, 881.0416, 
    936.1367, 774.4136, 1186.745, 1002.815, 1015.139, 535.5046, 386.2178, 
    179.3871, 69.36623, 267.0681, 111.3501, 67.82533, 6.994944, 1.526611, 
    3.172025, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 5.725166, 102.8057, 111.4602, 125.5778, 65.69091, 
    11.31183, 6.297175, 5.844241, 2.358717, 171.9062, 167.7866, 43.11033, 
    79.99084, 74.58493, 27.5016, 14.16823, 6.523846, 31.63298, 63.06898, 
    67.15324, 85.22324, 67.61577, 224.0022, 476.0859, 396.943, 309.3507, 
    246.142, 132.8316, 335.7784, 784.7097, 1053.235, 1127.867, 967.6097, 
    771.317, 924.9985, 1333.487, 1034.066, 789.8601, 234.963, 249.6979, 
    81.2932, 14.26598, 163.186, 164.9658, 5.164979, 1.026154, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.19746, 170.4447, 463.7712, 416.7452, 239.2617, 
    79.01589, 6.674962, 0, 0, 49.56345, 226.9828, 192.8199, 164.6065, 
    182.8128, 118.2701, 17.30331, 8.986745, 3.3333, 23.55511, 61.35153, 
    53.04255, 132.2586, 229.133, 315.2996, 329.1717, 262.2387, 250.0072, 
    217.4491, 311.0166, 854.7855, 1325.855, 1237.892, 1063.641, 815.3153, 
    855.515, 1043.939, 1759.73, 1143.116, 371.2457, 14.33288, 2.286062, 0, 0, 
    0.1220521, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 13.13908, 199.9922, 369.35, 332.041, 183.8263, 
    84.41653, 28.31347, 5.11356, 0, 3.346521, 94.1303, 145.3444, 260.3771, 
    308.1046, 216.5467, 65.93798, 66.89045, 91.82342, 129.8517, 169.2161, 
    212.0327, 380.3462, 430.9281, 398.8634, 271.8267, 213.1764, 198.3177, 
    260.7658, 507.0705, 1261.594, 1556.329, 1201.677, 977.4053, 903.3651, 
    1023.128, 1437.7, 2083.172, 1221.35, 86.26831, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 1.492808, 28.12763, 241.1122, 312.6933, 227.4316, 
    40.73929, 3.901017, 60.77868, 29.63254, 0, 37.46666, 47.92201, 90.67201, 
    252.6916, 297.8447, 250.6762, 146.2321, 137.6703, 164.451, 210.1363, 
    267.7924, 336.6427, 471.1196, 486.8597, 425.3645, 315.1228, 279.0462, 
    273.7747, 290.0505, 636.9206, 1410.759, 1544.152, 1250.766, 1127.925, 
    1065.812, 1110.734, 1416.591, 1600.496, 408.8422, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 8.41072, 11.77269, 0, 0, 1.62508, 8.022939, 6.219764, 0, 
    20.28673, 0.6057806, 40.99087, 150.5031, 84.34249, 84.26646, 195.8636, 
    227.4629, 190.5297, 136.6387, 154.2375, 176.6017, 216.4878, 304.6136, 
    374.8836, 462.7287, 472.5354, 402.6108, 307.9417, 327.0253, 306.5867, 
    373.0538, 668.3615, 1415.796, 1557.029, 1306.125, 1279.073, 1162.341, 
    1153.206, 1149.406, 1078.977, 41.16324, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 4.901734, 217.5294, 284.0266, 9.755486, 12.21576, 30.38478, 
    126.8581, 295.4576, 261.4576, 148.2994, 19.41799, 0.001383794, 4.122153, 
    25.35506, 13.69719, 14.41783, 64.17224, 71.70509, 82.17438, 88.62575, 
    143.002, 168.497, 227.1901, 295.2106, 377.9786, 424.9349, 434.2556, 
    359.2029, 243.9208, 256.3825, 320.5891, 276.9689, 544.5539, 1255.969, 
    1424.041, 1287.706, 1179.742, 1196.443, 1053.201, 1167.506, 829.4473, 
    18.81178, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.3367717, 55.36858, 332.4312, 482.9248, 279.4982, 0, 4.759403, 138.2639, 
    246.2088, 336.8652, 256.5343, 116.4693, 7.490035, 1.586183, 5.608893, 
    0.125523, 0.02205558, 0, 18.84512, 43.35651, 73.8119, 134.7575, 190.767, 
    245.426, 262.851, 321.6095, 350.954, 368.8531, 361.5361, 275.9557, 
    193.2714, 264.4291, 287.2755, 295.1925, 454.3226, 894.5059, 1154.717, 
    973.0314, 1099.105, 1148.796, 1120.024, 862.0306, 375.9889, 12.88452, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.2140546, 
    0.1701733, 26.3982, 16.54789, 11.51096, 64.69183, 320.2927, 487.4863, 
    486.2169, 178.1183, 52.80968, 111.4205, 188.5571, 226.6747, 194.1454, 
    121.9309, 19.68636, 0, 0, 0, 0, 0, 0, 0.08443239, 12.21449, 77.40128, 
    139.2317, 232.2935, 274.8673, 306.887, 328.7855, 366.2649, 352.3075, 
    297.598, 212.2141, 162.9654, 161.8156, 294.4319, 331.9783, 424.2078, 
    668.4012, 775.5222, 991.9241, 1072.528, 1282.538, 1139.612, 931.2537, 
    216.4193, 62.45685, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3.731169, 
    99.69241, 145.8221, 164.5461, 190.2277, 222.6298, 352.1655, 453.9755, 
    483.7257, 366.7473, 201.0961, 195.8921, 224.278, 247.8174, 199.336, 
    145.5127, 58.51702, 0.01620398, 1.724691, 0, 0, 0, 0, 0, 0, 3.441099, 
    66.59528, 167.6643, 266.4513, 312.1495, 332.5176, 373.2896, 422.7214, 
    417.7817, 331.4211, 227.7531, 191.2091, 276.8271, 346.7453, 491.9813, 
    515.8571, 477.7105, 837.2191, 1215.665, 1373.787, 1364.735, 1284.096, 
    957.2903, 218.0976, 83.97918, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7.299129, 134.0267, 
    294.2319, 344.9782, 270.6827, 318.7709, 384.5544, 494.1917, 494.657, 
    473.3284, 365.3275, 308.8357, 293.0063, 310.0292, 272.0663, 223.5598, 
    135.7657, 49.15474, 0.05388123, 0.2981069, 0, 0, 0, 0, 0, 0, 0.2216611, 
    69.87698, 190.6432, 286.7062, 330.1897, 367.8758, 406.1044, 450.1877, 
    427.9415, 330.3656, 250.8139, 289.5048, 447.8335, 462.0058, 478.6495, 
    494.2013, 530.5643, 958.8607, 1535.851, 1566.941, 1493.999, 1267.836, 
    1004.899, 187.0762, 37.84942, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.2778322, 1.216981, 0.320554, 
    82.15788, 124.0773, 328.814, 414.2038, 370.9027, 408.5572, 474.0244, 
    515.583, 504.9358, 517.7888, 478.3085, 405.8519, 390.0446, 340.6481, 
    284.1749, 193.1102, 63.77376, 0.2711483, 0.001171568, 0, 0, 0, 0, 0, 0, 
    0, 0.01659026, 97.79198, 225.3099, 301.7682, 358.1664, 393.5924, 
    409.4816, 387.7672, 372.0033, 279.7969, 234.8109, 369.993, 486.2102, 
    487.3097, 453.6224, 565.4487, 638.8194, 1025.565, 1495.267, 1465.116, 
    1353.271, 1132.2, 829.127, 232.6918, 86.18745, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.03872748, 20.11839, 53.78059, 
    33.44499, 88.68514, 177.8256, 19.69762, 253.2851, 404.7767, 437.9373, 
    469.3643, 499.6412, 501.7674, 551.6224, 574.769, 536.6869, 488.521, 
    416.7465, 350.7989, 264.6436, 127.1555, 0.415809, 0.4254224, 0, 0, 0, 0, 
    0, 0, 0, 0.6914847, 19.04652, 131.946, 247.1787, 306.9858, 363.0714, 
    397.9942, 400.0674, 409.7594, 398.0919, 355.8009, 291.4016, 333.1392, 
    498.2859, 440.002, 539.7181, 723.6176, 765.5291, 965.6453, 1312.768, 
    1339.947, 1188.61, 996.9376, 753.3426, 184.1582, 17.82256, 30.13374, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.789168, 70.13921, 107.3934, 180.0283, 
    234.5805, 241.1893, 107.9595, 15.09211, 188.5137, 368.2224, 514.8614, 
    566.2856, 554.1669, 566.897, 608.2187, 604.4344, 543.1758, 479.5136, 
    420.2968, 358.7137, 272.7408, 113.1928, 4.518106, 5.010964, 0, 0, 0, 0, 
    0, 0, 0.7098004, 13.29282, 97.01318, 193.7101, 286.6924, 317.051, 
    366.6038, 397.0652, 432.3381, 481.5545, 519.4891, 467.0329, 436.6177, 
    526.4904, 556.9227, 596.2275, 609.3391, 692.4142, 720.394, 862.9467, 
    1120.028, 1117.907, 1092.196, 985.4866, 917.553, 349.6905, 24.9056, 
    102.5677, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18.45255, 45.57545, 90.12004, 208.861, 
    326.2532, 247.4885, 3.031927, 0.8162752, 62.72859, 240.1284, 478.4014, 
    642.7585, 624.4623, 612.9011, 633.5761, 635.511, 540.0829, 464.6622, 
    389.1842, 327.2373, 250.5822, 128.0566, 4.151914, 0.01724564, 0, 0, 0, 
    0.06221788, 16.14303, 56.51927, 60.10637, 63.71621, 129.8515, 214.7995, 
    265.7689, 302.5134, 336.1973, 365.2288, 442.3849, 504.6011, 502.0141, 
    480.3363, 467.8888, 553.1976, 593.0986, 637.1354, 629.6438, 659.4634, 
    735.4026, 1028.44, 1056.044, 946.681, 926.314, 1064.744, 949.1011, 
    392.1784, 18.68724, 70.3578, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18.13205, 81.59405, 283.5952, 
    99.12554, 0, 2.600603, 22.27865, 40.11892, 259.8885, 493.662, 624.6654, 
    578.1021, 631.7147, 627.2502, 560.2089, 436.4544, 359.2498, 263.4945, 
    198.2276, 96.85187, 8.224985, 0.006419148, 10.41262, 28.47488, 33.42284, 
    63.55798, 89.37606, 117.4287, 123.5775, 113.715, 153.6499, 198.5007, 
    238.3534, 277.4305, 321.2411, 352.9605, 414.103, 455.9593, 452.3423, 
    458.7655, 565.2747, 608.5494, 639.5411, 687.265, 764.0191, 736.5245, 
    987.5319, 1266.858, 1113.241, 848.986, 966.5779, 1123.773, 1059.529, 
    375.9788, 5.606318, 11.23915, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 50.03308, 18.7767, 0, 
    1.26797, 38.3414, 37.16248, 6.458248, 236.8902, 463.1305, 562.8348, 
    578.8032, 630.9438, 520.6262, 426.2543, 325.3188, 244.9647, 138.4487, 
    36.07342, 0.5078325, 2.94648, 57.33051, 95.80891, 105.8, 111.6879, 
    121.1859, 142.7138, 152.8308, 160.8624, 182.531, 201.2338, 222.661, 
    264.4805, 303.7233, 333.4624, 371.3336, 438.1491, 455.2211, 496.9004, 
    597.2755, 643.8214, 617.1034, 691.8447, 823.0101, 988.5286, 1358.407, 
    1648.078, 1373.022, 979.8769, 1118.349, 1293.235, 1281.518, 524.8214, 
    12.07863, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18.53168, 7.44618, 
    0.2774768, 0, 35.85915, 285.9109, 179.5872, 150.5524, 421.4404, 514.148, 
    569.3135, 533.7565, 453.5545, 348.8341, 297.6014, 196.2376, 72.14723, 
    1.141348, 3.445107, 14.83014, 68.87897, 118.991, 129.5745, 158.0152, 
    182.8073, 209.6761, 221.1556, 222.757, 222.7252, 225.1968, 215.3978, 
    252.5812, 274.6012, 313.8231, 378.8444, 483.5266, 526.6315, 559.9622, 
    581.9632, 617.732, 638.4788, 691.2427, 829.9338, 1126.817, 1687.072, 
    1798.549, 1466.908, 1100.552, 1091.336, 1508.885, 1401.512, 703.5411, 
    81.51077, 0.2449444, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15.97898, 137.8128, 2.629696, 
    0.1815157, 0, 28.15523, 299.744, 311.1771, 79.97313, 377.6644, 488.9033, 
    461.6871, 486.7418, 409.492, 350.8954, 279.0941, 180.3749, 25.7736, 
    3.397881, 18.72686, 43.95182, 103.1606, 144.6976, 190.1044, 222.457, 
    259.2217, 285.7209, 287.2361, 281.1645, 272.6286, 249.3425, 225.9028, 
    238.7993, 272.0008, 332.6962, 384.1511, 468.3911, 546.1947, 577.4488, 
    627.5869, 635.5259, 700.1279, 776.9152, 929.8552, 1510.917, 1895.887, 
    1799.537, 1355.943, 1119.573, 1392.253, 1618.039, 1311.142, 575.1276, 
    257.3511, 0.8315546, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8.894205, 72.59029, 14.85453, 
    7.508962, 13.51235, 142.9096, 296.0406, 327.9227, 156.2393, 437.1971, 
    388.5025, 385.3842, 401.033, 394.5582, 335.838, 280.1766, 193.5683, 
    96.386, 35.52516, 58.84515, 86.79417, 122.0659, 181.4595, 237.5804, 
    289.2039, 326.9966, 354.348, 356.1935, 336.6149, 307.5397, 253.4356, 
    225.7552, 236.1096, 334.7573, 444.7771, 494.1808, 514.2294, 524.8425, 
    587.1181, 631.0831, 694.0496, 751.4611, 825.4266, 1097.83, 1658.775, 
    2006.745, 1602.702, 1223.444, 1127.629, 1333.478, 1458.12, 871.0525, 
    466.6771, 267.9041, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01038057, 0, 6.643703, 101.4879, 
    82.98901, 51.23274, 85.14922, 210.2779, 283.6747, 309.324, 233.2301, 
    492.1425, 371.6667, 362.65, 444.5501, 397.6977, 330.4786, 280.92, 
    273.9966, 219.3448, 153.7401, 126.073, 117.5657, 150.8828, 219.6838, 
    283.4588, 333.4008, 374.8239, 400.1253, 395.6437, 375.5026, 312.2456, 
    243.2001, 227.2077, 279.3844, 409.5839, 514.515, 561.0614, 561.6627, 
    541.6973, 592.7158, 646.3815, 705.6855, 755.9585, 820.3306, 1077.465, 
    1725.695, 1795.541, 1577.446, 1249.411, 1148.976, 1319.127, 995.0981, 
    382.848, 349.3625, 65.2517, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 49.50258, 104.9451, 82.473, 
    92.12851, 176.1149, 268.6027, 316.0862, 341.2645, 486.9077, 443.9214, 
    441.7123, 453.1961, 411.6028, 339.4975, 305.282, 294.3625, 287.3364, 
    230.1652, 207.584, 207.6316, 229.0633, 299.8941, 320.3898, 366.2971, 
    403.0446, 399.9144, 400.9593, 372.4525, 306.9135, 239.632, 240.6821, 
    343.6025, 474.4823, 553.2586, 592.0007, 575.3657, 602.5383, 624.6992, 
    700.6254, 727.1317, 764.283, 781.6901, 1065.684, 1631.907, 1692.728, 
    1571.499, 1298.507, 1313.886, 1286.554, 934.9397, 106.3758, 289.6695, 
    15.00103, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11.55675, 115.867, 
    22.48811, 65.3556, 149.1486, 286.7424, 407.3988, 236.5376, 274.9689, 
    357.7444, 443.3862, 421.6057, 401.2734, 343.1813, 298.683, 307.432, 
    300.7722, 291.2484, 308.8382, 334.8492, 323.8983, 337.6805, 341.7525, 
    399.8321, 429.9846, 410.5637, 382.6377, 354.2699, 306.8083, 234.6121, 
    282.1734, 378.2628, 513.45, 570.4268, 609.7987, 630.7244, 657.3438, 
    763.2346, 822.8828, 897.2252, 876.2137, 902.7307, 1085.887, 1506.075, 
    1453.561, 1306.629, 1103.886, 1026.492, 1225.022, 985.5616, 402.682, 
    411.0314, 92.16769, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8.036347, 62.52849, 
    3.547037, 32.43497, 104.1824, 329.8143, 462.2404, 251.2797, 109.8259, 
    300.0777, 382.1133, 340.6129, 357.1865, 326.0741, 305.6071, 339.9389, 
    372.1312, 391.5172, 407.5522, 352.1345, 293.8417, 268.1846, 292.7089, 
    444.7627, 466.584, 417.2143, 374.3411, 349.6299, 313.55, 266.888, 
    336.9229, 432.6651, 484.9139, 546.2026, 630.8204, 650.4514, 755.9393, 
    824.0303, 861.4523, 911.7997, 958.1385, 976.4166, 1254.706, 1563.365, 
    1293.88, 1170.993, 864.0294, 700.7004, 757.6398, 917.2304, 682.3601, 
    402.354, 43.28111, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.05915249, 0.08011421, 0, 
    6.02283, 76.62966, 347.7174, 469.9626, 235.3439, 100.1177, 160.2919, 
    227.011, 263.368, 336.6925, 322.0186, 290.6877, 363.0302, 432.0052, 
    448.0348, 357.6713, 268.9411, 179.2584, 179, 233.9073, 359.2671, 
    464.7566, 411.7307, 372.834, 358.2526, 326.1168, 293.7316, 402.5888, 
    470.521, 497.5835, 578.8224, 635.5013, 674.5109, 734.5461, 763.5286, 
    810.0879, 885.3263, 939.2901, 1104.282, 1317.147, 1582.151, 1373.822, 
    1213.066, 873.9077, 635.079, 382.4486, 656.3605, 884.5526, 664.905, 
    217.4573, 32.62277, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.014362, 
    61.41228, 327.5756, 417.7493, 328.8751, 249.4016, 131.7789, 157.5266, 
    287.179, 367.0403, 311.7421, 237.5124, 263.4082, 315.4411, 318.5938, 
    269.0101, 179.5965, 192.4013, 228.7823, 193.9452, 278.2494, 363.2266, 
    430.6738, 408.0237, 404.8087, 350.7692, 302.6519, 419.8691, 508.0556, 
    530.116, 605.4689, 677.9661, 698.0052, 724.3315, 784.8451, 801.787, 
    928.4433, 1166.382, 1351.242, 1463.7, 1691.588, 1541.213, 1399.71, 
    1026.168, 717.6241, 512.4301, 377.8375, 697.6708, 594.645, 397.4904, 
    142.8448, 0.532489, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.2053152, 
    67.53915, 303.6299, 379.2345, 436.3914, 423.1708, 180.6438, 155.2336, 
    276.7622, 326.9408, 266.7624, 175.7495, 176.1388, 195.9187, 226.1668, 
    186.327, 215.0712, 291.8131, 416.8516, 394.0894, 300.8634, 340.7516, 
    360.322, 408.5583, 425.7607, 360.9985, 326.2549, 435.8652, 544.7354, 
    572.8199, 653.0318, 746.2729, 793.1929, 824.189, 828.2086, 914.1102, 
    1028.284, 1346.432, 1671.313, 1678.606, 1814.529, 1881.197, 1709.896, 
    1406.109, 1219.147, 1059.282, 948.7432, 834.345, 919.3475, 724.296, 
    356.6761, 76.5276, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.8787696, 13.35174, 
    137.5124, 287.6332, 345.7241, 417.4199, 379.3897, 131.3522, 106.2649, 
    169.0464, 272.2558, 288.1475, 201.0602, 176.5896, 223.6827, 266.1863, 
    218.2081, 176.9505, 269.0522, 436.2097, 486.094, 402.9827, 347.54, 
    334.3905, 365.894, 393.4282, 347.4721, 379.8949, 443.5723, 566.2279, 
    602.1741, 676.5858, 812.3363, 900.5889, 908.915, 931.9954, 944.5102, 
    1117.414, 1304.28, 1882.296, 1832.433, 1976.871, 2069.233, 2070.061, 
    1899.477, 1551.457, 1340.278, 1386.592, 1314.673, 1244.868, 1230.34, 
    806.1844, 287.225, 40.42369, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2.817714, 35.69061, 
    138.5443, 281.9023, 361.2498, 453.4521, 359.1906, 222.1722, 156.6933, 
    136.975, 236.7071, 325.3279, 228.1469, 196.3775, 242.6227, 329.216, 
    249.9151, 180.1256, 229.7955, 351.343, 390.6742, 362.7199, 313.2054, 
    299.3227, 315.3665, 337.3273, 403.3815, 440.4469, 459.0341, 544.0665, 
    574.6163, 685.2004, 805.9506, 978.1014, 1079.502, 1060.385, 1335.979, 
    1386.026, 1736.179, 2369.993, 2377.097, 2108.683, 2192.729, 2248.685, 
    2160.981, 1428.064, 1097.215, 1308.715, 1435.482, 1437.344, 1562.363, 
    1290.539, 805.3401, 441.8997, 16.92101, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 land_mask =
  0, 0.2884085, 0.9991118, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9922887, 0.3335225, 
    0.004607826, 0.003236954, 0.508559, 0.9850757, 0.9911836, 0.1925444, 0, 
    0, 0,
  0.02305815, 0.1375988, 0.944828, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.8519247, 
    0.1034592, 0, 0, 0.02152651, 0.1580271, 0.214971, 0, 0, 0, 0.004275662,
  0.6877087, 0.944828, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.7618825, 
    4.015537e-05, 0.2204578, 0.0836201, 0, 0, 0, 0, 0.006251427, 0.5966954,
  0.9875305, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.6890369, 0.02053772, 
    0.7023288, 0.225828, 0, 0, 0.2833943, 0.1682406, 0.614427, 1,
  0.9998894, 1, 1, 1, 1, 1, 1, 1, 1, 0.982605, 0.4463286, 0.2774308, 
    0.6133593, 0.9973181, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 0.5015463, 0.3794187, 0.9844274, 0.1219514, 0, 0.5, 
    1, 0.9917114, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 0.9341351, 0.2591562, 0, 0, 0, 0.778241, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.7423904, 
    0.641713, 1, 0.7179503, 0.7577073, 1, 1, 1, 0.9345905, 0.7734837,
  1, 1, 1, 1, 1, 1, 1, 1, 0.6711941, 0, 0, 0, 0, 0.7003056, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.7377394, 0.5135806, 0.05480789, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 0.5039137, 0, 0, 0, 0.02591443, 0.9401757, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 0.7924682, 0.0008498987, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 0.3537756, 0, 0, 0, 0, 0.8171846, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.8385026, 0.01230605, 0, 0, 0,
  0.9900191, 1, 1, 1, 0.982605, 0.8792336, 0.6995067, 0.5093474, 0.0169677, 
    0, 0, 0, 0, 0.7583464, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.5511215, 0, 0, 0, 0,
  0.6112348, 1, 0.995035, 0.7029089, 0.810859, 0.09081139, 0, 0, 0, 0, 0, 0, 
    0.01839714, 0.9189041, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.7265073, 0.04310679, 0, 0, 0, 0,
  0.4115516, 0.9695646, 0.32083, 0.3587675, 0.2985553, 0, 0, 0, 0, 0, 
    0.1353143, 0.3167184, 0.5955938, 0.2275586, 0.3671458, 0.9835829, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.3382995, 0, 0, 0, 0, 0,
  0, 0.1277016, 0.7127959, 0.9866941, 0.6133593, 0, 0, 0, 0, 0, 0.2077407, 
    0.931155, 0.5506355, 0.03697443, 0.1507062, 0.5356609, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9921315, 
    0.147725, 0, 0, 0, 0, 0,
  0.01037147, 0.1938587, 0.8625931, 1, 0.9973181, 0.4946559, 0.0311923, 0, 0, 
    0, 0.00735819, 0.5864723, 0.9627873, 0.8827814, 0.9648471, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9980701, 
    0.1807344, 0, 0, 0, 0, 0,
  0.7028435, 0.9317848, 1, 1, 1, 1, 0.9336721, 0.3483783, 0.07686493, 0, 0, 
    0.3183673, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 0.6919137, 0.0003099618, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 0.888535, 0.5828943, 0.380111, 0.6304355, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 0.983552, 0.1295606, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.8518441, 0.01128992, 
    0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.999961, 0.276726, 0, 0, 
    0, 0, 0.01621984,
  0.6853452, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.8485698, 
    0.009902901, 0, 0, 0, 0.1625293, 0.2812916,
  0.1046904, 0.9492866, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.5342661, 
    0, 0, 0, 0.2437459, 0.5925891, 0.1728241,
  0, 0.6909669, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9896021, 0.19564, 
    0, 0, 1.512684e-05, 0.6681376, 0.5249494, 0.001406433,
  0.104618, 0.3731309, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.516663, 0, 
    0, 0, 0.179388, 0.9754534, 0.9489582, 0.4696769,
  0.1094959, 0.1844557, 0.9892092, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.8602238, 0.005510823, 0, 0.005748244, 0.4703873, 0.9732017, 1, 
    0.8608779, 0.03971616,
  0.04849377, 0.01244223, 0.9232286, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.3732215, 0, 0, 0.02369886, 0.5267625, 0.6938574, 0.9234961, 0.9547111, 
    0.04446942,
  0.5122615, 0.02757481, 0.5740731, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.840474, 
    0.01930639, 0.0865661, 0.5162175, 0.1518759, 0, 0, 0.2306587, 0.5255683, 0,
  1, 0.5190924, 0.05039959, 0.9774919, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9979244, 
    0.6173158, 0.06360614, 0.3239541, 0.6181117, 0.3434, 0.08735604, 0, 0, 0, 
    0, 0,
  1, 0.6923935, 2.081939e-06, 0.6747068, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9996232, 1, 1, 1, 1, 
    0.3280995, 0.1371462, 0.7053908, 0.4147068, 0, 0, 0, 0, 0, 0, 0, 0,
  0.9767516, 0.9616271, 0.1639549, 0.271809, 0.9999644, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 0.79072, 0.9954807, 0.6932396, 0.992215, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 0.9982526, 0.7430784, 0.3342112, 0.9753816, 1, 1, 0.5895154, 
    0.4768312, 0.9639986, 0.7426976, 0.1318247, 0, 0, 0, 0, 0, 0, 0, 0,
  0.3953824, 1, 0.9443728, 0.9979815, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.8859383, 0.6344793, 0.8400888, 1, 0.6961708, 0.6793767, 1, 0.9887459, 
    0.4841065, 0.8715914, 1, 1, 1, 1, 0.9284868, 0.7849948, 0.7127485, 1, 
    0.9687542, 0.9541373, 0.7891752, 1, 1, 0.9629303, 0.8951254, 0.6504759, 
    0.8937041, 0.7830405, 0.342161, 1, 0.6261792, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.8566951, 0.02276905, 0.002447544, 0.514191, 0.722188, 0.6127455, 
    0.7949336, 0.7562089, 0.5650142, 0.06637619, 0.01120179, 0, 0, 0, 0, 0, 
    0, 0, 0,
  0.05505988, 0.888244, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.5507722, 
    0.0006194019, 0.116053, 0.619944, 0.742622, 0.1034394, 0.9146509, 
    0.4991146, 0.2116089, 0.9242266, 1, 1, 1, 1, 0.8386455, 0.4342496, 
    0.06022686, 0.5132908, 0.3214224, 0.5160704, 0.224035, 0.4073008, 
    0.5465707, 0.3329684, 0, 0.07634896, 0.5107231, 0.03671252, 0.2859505, 1, 
    0.6545428, 0.9156184, 0.97225, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.3421438, 0, 0, 0, 
    0.2840079, 0.6098053, 0.106933, 0.001375207, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  0.4128869, 0.9714226, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9036868, 
    0.3452899, 0, 0, 0, 0.0115361, 0.1913566, 0.1288761, 0.5540914, 
    0.9598167, 1, 1, 1, 1, 1, 1, 0.3918472, 0.3429512, 1, 0.8047241, 
    0.02029391, 0.7208738, 0.03791168, 0.4779267, 0, 0.01079109, 0.2673898, 
    0.04183982, 0, 0.1123773, 0.8191687, 0.7129377, 0.5516703, 0.9328146, 
    0.75521, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 0.9617294, 0.06184853, 0, 0, 0.000967195, 0.1277687, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0.9957435, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.8395773, 0.1179296, 
    0.01795836, 0.02010509, 0.007536734, 0.2286892, 0.04640759, 0, 0, 
    0.6564662, 1, 1, 1, 1, 1, 1, 1, 0.834378, 0.7319705, 1, 0.9198699, 
    0.01201014, 0.04465218, 0, 0, 0, 0.3684395, 0.5827318, 0, 0, 0, 
    0.2186891, 0.6873481, 0.1364655, 0.186791, 0.7450449, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.5434414, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.889401, 0.122736, 0.3139295, 
    0.7522845, 0.8038401, 0.3664241, 0.24319, 0.52267, 0.1478724, 0.09243008, 
    0.6729867, 0.9999971, 1, 1, 1, 1, 1, 0.9871168, 0.9992952, 1, 0.8422172, 
    0, 0, 0, 0, 0, 0.3275236, 0.8442517, 0.08887865, 0, 0, 0, 0.156116, 
    0.02045131, 3.470624e-05, 0.2521144, 0.6287342, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9975308, 0.149125, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.4399916, 0.4513926, 0.6248305, 1, 
    1, 1, 1, 1, 0.5065262, 0, 0, 0.4453909, 0.5339093, 0.4254689, 0.5834806, 
    1, 1, 1, 1, 1, 0.5982459, 0, 0, 0, 0, 0, 0, 0.3391043, 0.852947, 
    0.1592709, 0, 0, 0, 0, 0, 0.03027248, 0.4168469, 0.9877434, 1, 1, 1, 1, 
    0.8619069, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.9664218, 0.08247031, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.8920162, 0.5407821, 0.4654229, 
    0.2409135, 0.3909343, 0.988422, 1, 1, 1, 0.8909804, 0.531373, 0.2580832, 
    0.3792476, 0.7087116, 0.4061886, 0.4193644, 1, 1, 1, 1, 1, 0.2638651, 0, 
    0, 0, 0, 0, 0, 0, 0.2239696, 0.9176144, 0.4488631, 0.1449512, 
    0.001410662, 0, 0, 0.03603189, 0, 0.3868065, 0.9493498, 1, 1, 1, 
    0.7200027, 0.8212039, 0.990998, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 0.4792888, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.7146486, 0.118375, 0.4868317, 0.9180648, 
    0.8884519, 0.3578016, 0.3644181, 0.9821022, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 0.9876617, 0.3491453, 0, 0, 0, 0, 0, 0, 0, 0, 0.08260295, 
    0.4333614, 0.5040144, 0.3614931, 0, 0, 0, 0.005346482, 0.01236961, 
    0.2922967, 0.7454089, 1, 1, 0.8454538, 0.1922676, 0.3820402, 0.5675731, 
    0.9620153, 1, 1, 0.9772007, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.8661066, 0.00407539, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 0.7854356, 0.5305065, 0.2314634, 0, 0, 
    0.2847562, 0.6988515, 0.3205059, 0.001980788, 0.5282913, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 0.9088889, 0.3662374, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.002319489, 0.003097083, 0.006384837, 0.4009853, 
    0.9520847, 0.9565648, 0.7851307, 0.003207061, 0, 0.03928687, 0.8853757, 
    0.9915587, 0.4154324, 0.5028495, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.9239731, 0.04490227, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1532502, 0, 0, 0, 
    0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 0.6720341, 0.02851992, 0.0008780628, 0, 0, 0, 0, 0, 
    0.08552671, 0.7316995, 0.9995651, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.7766737, 0.4137197, 0.01565327, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.00839087, 0.179177, 0.3358206, 0.1938771, 0.08693577, 
    0.01849443, 0, 0, 0, 0.04255971, 0.1354656, 0, 0.2326064, 0.9961697, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9906443, 0.6093469, 0.08272952, 0, 0, 
    0, 0, 0, 0, 0.003714734, 0.04793612, 0.195166, 0.1305265, 0, 0, 0, 0, 0, 
    0, 0,
  1, 1, 1, 1, 1, 1, 0.997851, 0.8851513, 0.2218852, 0, 0, 0, 0, 0, 0, 0, 
    0.01474294, 0.9223265, 0.9997482, 1, 1, 1, 1, 0.8567648, 0.7138887, 
    0.7556022, 0.7419234, 0.5976552, 0.7780174, 0.7167592, 0.4319452, 
    0.02324593, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.02652722, 0.7279592, 0.6135988, 0.341273, 0.007845606, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.01614682, 0.6782818, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.9998435, 0.2067607, 0, 0, 0.091288, 0.5062699, 0.6916178, 0.7767209, 
    0.8624772, 0.9701989, 0.364688, 0, 0, 0, 0, 0, 0, 0, 0,
  0.4190771, 0.6497226, 0.9545459, 1, 1, 1, 0.6781163, 0.06010642, 0.5008612, 
    0.4229959, 0.1875891, 0, 0, 0, 0, 0, 0, 0.0595316, 0.5124435, 0.9682307, 
    1, 0.9258996, 0.5065909, 0.04083258, 0, 0, 0, 0.03120807, 0.1286479, 
    0.006753318, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1067706, 0.3340207, 
    0.2393772, 0, 0.002743472, 0.01939562, 0.08303384, 0.6292495, 0.01828023, 
    0, 0, 0, 0, 0, 0, 0, 0, 0.03133215, 0.007111566, 0.2436219, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9708926, 0.4725524, 0.1960722, 0, 0.1848622, 
    0.8739176, 1, 1, 1, 0.9030244, 0.3938256, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0.6705055, 1, 1, 0.9502218, 0.107991, 0.4462324, 1, 1, 0.7277706, 
    0.004069345, 0, 0, 0, 0, 0, 0, 0, 0.05657173, 0.3351253, 0.1607299, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.03699553, 
    0.2052931, 0.1163417, 0.04926136, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.3625355, 0.506983, 0.2779973, 0.5109867, 0.7485809, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 0.5927411, 0, 0, 0.1106688, 0.9105396, 1, 1, 1, 
    0.9959307, 0.4352124, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0.01193915, 0.7290006, 0.9996663, 0.09786085, 0.1382244, 0.5658905, 
    1, 1, 1, 0.8744788, 0.08482047, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1665618, 0.3248779, 0.0230974, 
    0.01594665, 0.02927415, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.2599293, 0.8565587, 0.00678506, 0, 0.0779523, 0.699297, 0.9691742, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 0.8166098, 0.03916229, 0, 0.005817841, 
    0.692153, 1, 1, 1, 0.9411603, 0.2435686, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0.2993191, 0.9495773, 0, 0.01423644, 0.7039637, 1, 1, 1, 1, 
    0.7995175, 0.254755, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.2888699, 0.705927, 0.7486029, 0.6040528, 0.3449149, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1760819, 
    0.4655593, 0, 0, 0, 0.1594579, 0.9752054, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.8951882, 0.2522649, 0.004452626, 0.5549645, 1, 1, 1, 0.8623571, 
    0.6075783, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0.07980675, 0.2809722, 0, 0.1385953, 0.7865735, 0.7880519, 
    0.968846, 0.5791082, 0.4798856, 0.9172074, 0.927383, 0.83219, 0.3994447, 
    0.04030702, 0, 0.07399552, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.0004920398, 0.3404756, 0.9613062, 0.4522832, 0.03017027, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01749192, 0.01128817, 
    0.1379025, 0, 0, 0, 0.04587796, 0.9871097, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.6999564, 0.3755875, 0.9989443, 0.6214731, 0.5969585, 0.5454745, 
    0.1750769, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0.1596749, 0.01195103, 0.1571471, 0.02306698, 0.028618, 
    0.3427889, 0.721784, 1, 1, 0.8513392, 0.3177238, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.02060047, 0.2733825, 0.02397867, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.4457313, 0.7043854, 1, 1, 1, 1, 1, 1, 1, 1, 0.6029556, 0.9542752, 
    0.4643725, 0.2527745, 0.02328439, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0.007150483, 0.7961679, 0.8434761, 0.9726763, 
    0.4238593, 0.5026287, 0.622201, 0.4973026, 0.0772241, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.2232726, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 0.9596362, 0.2153704, 0.02692382, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0.5481955, 1, 1, 0.9846066, 0.5166809, 0, 0, 
    0.0605782, 0, 0, 0, 0.02565648, 0.2292144, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.002742995, 0.9592576, 1, 1, 1, 1, 
    1, 1, 1, 1, 0.8386291, 0.06731934, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0.7911306, 0.744423, 0.9958476, 0.3917643, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.1602756, 0.7774471, 1, 1, 1, 1, 1, 1, 1, 1, 0.7282078, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0.2763341, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.02465551, 0.5389555, 
    0.09023141, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.3491064, 0.7970511, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.7709398, 0.05621546, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.02616456, 0.4072716, 0.02764438, 0, 0, 0, 0, 0, 0, 0, 0, 0.007946228, 
    0.0215098, 0.1481985, 0.1512895, 0.2826785, 0.7654743, 0.9869945, 
    0.5499371, 0.567008, 0.05657073, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.3411054, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.7214631, 0.1254226, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.5718764, 1, 0.617721, 0, 0, 0, 0, 0, 0, 0, 0.148285, 0.6013126, 
    0.7386797, 0.8317872, 0.9721572, 0.9878897, 1, 1, 1, 1, 0.5187135, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.04601588, 0.1928452, 0.9953901, 1, 1, 1, 1, 1, 1, 0.9362985, 0.1519071, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.02308159, 
    0.9368013, 1, 0.5605719, 0, 0, 0, 0, 0.0994027, 0.1519942, 0.4023046, 
    0.8973336, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.6283081, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.2124189, 0.437899, 0, 
    0.7649915, 1, 1, 1, 0.9788436, 0.7998188, 1, 0.4011095, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1528232, 
    0.9851291, 1, 0.5690181, 0.007882722, 0, 0, 0.3224736, 0.4599625, 
    0.9042956, 0.999677, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.4572058, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.006458772, 
    0.0237647, 0, 0.227326, 0.9942815, 1, 0.6645961, 0.4432212, 0.03989381, 
    0.5392244, 0.2095875, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.430079, 
    0.7312796, 0.8450026, 0.1614028, 0, 0.04361914, 0.8531964, 0.8497482, 
    0.9997948, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.8977383, 0.3332031, 
    0.3655361, 0.04765641, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.7132292, 1, 0.816526, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.05260738, 0.07836438, 0, 0, 0.2491814, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 0.9207466, 0.7041428, 1, 0.7042463, 0.01935159, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1916869, 0.997572, 
    0.9664844, 0.2796616, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.3168469, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.8713294, 
    0.7350758, 1, 0.9985892, 0.5351546, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1795665, 0.9986884, 0.8846707, 0.5677841, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.3550282, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.279303, 
    0.6442038, 1, 0.6813606, 0.6184936, 0.1960024, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0251202, 0.260837, 0, 0.0004929128, 
    0.3365258, 0.0114776, 0.03985736, 0.1344334, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.1158035, 0.890343, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.7351844, 0.5533677, 1, 0.7738451, 0.9701509, 0.3894742, 0.001606799, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.005773118, 0.3039451, 0.7407112, 
    0.7999177, 0.9048856, 0.0141415, 0.1831883, 0.4115106, 0, 0.1069227, 
    0.2025667, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1092487, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.5193717, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.994473, 0.5692437, 
    0.4542774, 0.9261664, 0.8238658, 0.2153217, 0.5868801, 1, 0.7394806, 
    0.8058553, 0.1632256, 0.547113, 0.06057538, 0.09398247, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.7215818, 1, 1, 1, 1, 0.4168746, 0.8358276, 0.9664901, 
    0.1808136, 0.01235209, 0.0244422, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.02900386, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.6050302, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.8627397, 0.2401952, 0, 0, 
    0.121907, 0.1521004, 0, 0.644744, 0.9510419, 0.301559, 0.2032923, 
    0.2832184, 0.1715124, 0.0642454, 0.3894436, 0.355457, 0.1890444, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.07950651, 0.9975182, 1, 1, 1, 1, 0.8763351, 
    0.9740863, 0.9582601, 0.05713792, 0.006239007, 0.08203404, 0.03931703, 
    0.00247307, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.06966187, 0.06613558, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.003755757, 0.5864659, 1, 1, 1, 1, 1, 0.9925512, 0.8724307, 0.6710725, 
    0.7534792, 0.07587746, 0, 0, 0, 0, 0, 0, 0.3674421, 0.5488101, 0.6089712, 
    0.5379397, 0.2472398, 0.1861075, 0.1012413, 0.1267425, 0.4983214, 
    0.6058319, 0.03750185, 0, 0, 0, 0, 0, 0, 0, 0, 0.5366537, 1, 1, 1, 1, 1, 
    1, 1, 0.6697894, 0.2345046, 0.8237509, 0.9863058, 0.4740853, 0.4750053, 
    0.1235425, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.4309661, 0.9817041, 1, 1, 1, 1, 1, 0.571421, 0.7863377, 0.1386277, 
    0.02245102, 0, 0, 0, 0, 0, 0, 0.05556273, 0.9789172, 0.7375769, 
    0.8189688, 0.3559348, 0.6307323, 0.6821151, 0.5123709, 0.6651374, 
    0.8837627, 0.1572086, 0.05174712, 0.09259965, 0, 0, 0, 0, 0, 0, 
    0.06662905, 0.9413299, 1, 1, 1, 1, 1, 1, 1, 0.9999163, 0.9697776, 1, 1, 
    1, 0.4300958, 0.003663761, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.1867139, 0.9595957, 1, 1, 1, 1, 1, 1, 0.284351, 0.2819466, 0, 0, 0, 0, 
    0, 0, 0, 0.221816, 0.234015, 0.1498427, 0.4379888, 0.4701115, 0.3815823, 
    0.202223, 0.06689857, 0.1760091, 0.348862, 0.2906938, 0.3599098, 
    0.8773224, 0.6843942, 1.096974e-05, 0, 0, 0, 0, 0, 0.729326, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 0.9291328, 0.1750867, 0, 0, 0, 0, 0, 0, 0, 
    0.1284918, 0.03147244, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.2094367, 0.9369895, 1, 1, 1, 1, 1, 1, 0.8089225, 0.05077393, 0, 0, 0, 
    0, 0, 0, 0.1286864, 0.5131698, 0.9357795, 0.9835859, 0.6595818, 
    0.6586512, 0.5519477, 0.6267641, 0.5283211, 0.1642075, 0.2885776, 
    0.04336228, 0.04232852, 0.7210842, 0.8761302, 1, 0.4428093, 0, 0, 0, 0, 
    0.2362406, 0.9876587, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.8892759, 
    0.2210028, 0, 0, 0, 0, 0.01768243, 0.2350183, 0.2126607, 0.007313905, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.09397414, 0.9518533, 1, 1, 1, 1, 1, 0.9310701, 0.6551082, 0.02464128, 
    0, 0, 0, 0, 0.001893531, 0.428525, 0.660005, 0.9646558, 0.9979754, 1, 1, 
    0.7802781, 0.8504569, 0.2165388, 0.643451, 0.9057896, 0.4174795, 
    0.5542305, 0.6763288, 0.8081042, 0.988646, 0.6779991, 0.7144226, 
    0.3391109, 0.03010433, 0.1083374, 0.3236497, 0.4993806, 0.6720286, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.7566548, 0.09032444, 0, 0, 0, 
    0.1800638, 0.2171838, 0.04050701, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.5591969, 0.9228026, 1, 1, 1, 0.9221501, 0.5172973, 0.05100384, 0, 0, 0, 
    0.0007068556, 0.01091526, 0.0301949, 0.2755317, 0.965713, 1, 1, 
    0.9936191, 1, 1, 0.9859811, 0.619966, 0.1089375, 0.4886177, 0.6999307, 
    0.07001494, 0.6258047, 0.9147264, 1, 1, 0.6264263, 0, 0, 0.1941441, 
    0.9471765, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.5419797, 
    0, 0.015395, 0.2036542, 0.6540743, 0.4381296, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.006838025, 0.01351406, 0.4722523, 0.538614, 0.2337886, 0.001982945, 0, 
    0, 0, 0, 0, 0.7464898, 0.9450542, 0.9789113, 0.99442, 1, 0.9895004, 
    0.7432182, 0.2929687, 0.8314089, 0.8995512, 0.7964581, 0.1749706, 
    0.6521643, 0.7756425, 0.008177926, 0.1344325, 0.8013356, 1, 0.9843748, 
    0.6497664, 0.5200529, 0.04047306, 0.6355119, 0.8531175, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 0.8961154, 0.9560985, 0.9943568, 1, 0.9338681, 
    0.5818689, 0.7449133, 0.7265122, 0.293891, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.0579614, 0.9415749, 0.8603365, 0.9990121, 1, 
    0.803029, 0.3949734, 0.1770097, 0.005452511, 0.510583, 0.7336312, 
    0.001113111, 0.1646328, 0.8604911, 0.5931268, 0.1902591, 0.5364736, 
    0.9966938, 0.956994, 1, 0.9285627, 0.4400202, 0.722735, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9410389, 0.5555537, 0.3014219, 0.601414, 
    0.4825325, 0.2935872, 0.08583173, 0.004107873, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.03901332, 0.3728116, 0.4575627, 1, 1, 0.3147727, 
    0.3332067, 0.2217817, 0.05301935, 0.7761925, 0.6799878, 0.399193, 
    0.7055106, 0.8377438, 0.6134337, 0.4755627, 0.2565599, 0.4595538, 
    0.6566908, 0.4802974, 0.3227839, 0.6104215, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 0.9089081, 0.5222241, 0.4558146, 0.1927821, 0.1057313, 
    0.7160483, 0.6894037, 0.0001066323, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.001781516, 0.5839874, 0.9946612, 1, 1, 0.9786469, 
    0.2361013, 0, 0, 0.2998931, 1, 0.8093447, 0.6758854, 0.9936388, 
    0.9348447, 0.6461143, 0.534321, 0.2699139, 0.8118511, 0.9714402, 
    0.7283285, 0.8378774, 0.9670031, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 0.8234991, 0.08674643, 0.0131576, 0, 0, 0.02502642, 0.01614379, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.1014065, 0.7311866, 0.7506915, 1, 1, 0.9619322, 
    0.6062644, 0.1703102, 0, 0.04583564, 0.6992308, 0.8417487, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9660713, 
    0.2967638, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.01285044, 0.1548295, 0.6499813, 0.889262, 0.9474576, 
    0.3051719, 0.1076564, 0.5899696, 0.2210208, 0, 0.1423286, 0.6488663, 
    0.7522198, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 0.9999971, 0.4893933, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.1127665, 0.1135007, 0, 6.399585e-05, 0.0003775573, 
    0.03852168, 0.05766925, 0, 0.171762, 0.01750567, 0.4126715, 0.8537696, 
    0.8530025, 0.672665, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 0.9984903, 0.1519116, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.0262549, 0.4324569, 0.9188194, 0.03891509, 0.07369219, 0.2784357, 
    0.439794, 0.9090685, 0.8842618, 0.613674, 0.169175, 0.0007593664, 
    0.05496632, 0.3555141, 0.4366377, 0.1746797, 0.660701, 0.9513029, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9929273, 
    0.1262638, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0152431, 0.3903114, 0.8834387, 1, 0.809934, 0, 0.08427224, 0.9253466, 
    1, 1, 1, 0.7736004, 0.162165, 0.0586152, 0.3602923, 0.03943993, 
    0.001398534, 0, 0.2553839, 0.8987577, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9784375, 0.07446165, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.006909454, 
    0.02203574, 0.2018838, 0.2004992, 0.2420584, 0.6730793, 0.9998235, 1, 1, 
    0.9541899, 0.6909702, 0.8539598, 1, 1, 1, 0.9992172, 0.3129094, 0, 0, 0, 
    0, 0, 0, 0, 0.5284762, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 0.9821761, 0.7433433, 0.2581827, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.004164889, 
    0.598833, 0.912891, 0.9848074, 1, 0.9949051, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 0.8401424, 0, 0, 0, 0, 0, 0, 0, 0, 0.1808639, 0.9999599, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9998994, 0.5513852, 
    0.3237998, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.6889238, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.7519505, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.8577955, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 0.9713004, 0.1253456, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.03594787, 0, 0.0008203032, 
    0.4332399, 0.5592608, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9933216, 
    0.4570104, 0.01265947, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.8118156, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.942905, 0.6050133, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0007849386, 0.06672296, 0.6196942, 
    0.3867162, 0.3914538, 0.7130988, 0.1269462, 0.9995891, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 0.6703829, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.06998937, 
    0.5995811, 0.9730762, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 0.4093178, 0.145072, 0.09990545, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.003637707, 0.559929, 0.9073727, 1, 
    0.9975478, 0.999097, 0.3226125, 0.1728628, 0.996939, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 0.618335, 0.03839462, 0.163095, 0, 0, 0, 0, 0, 0.00750303, 
    0.003358266, 0.3714445, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 0.8540727, 0.2479777, 0.566503, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1012027, 0.4235917, 0.7059572, 
    0.9331499, 1, 0.8808568, 0.05236256, 0, 0.6189646, 0.9339727, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 0.8560801, 0.09653471, 0, 0, 0, 0, 0.001193712, 
    0.3857171, 0.8091468, 0.9605917, 0.8586759, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9887962, 0.08099455, 0.4007379, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0009469227, 0.2329264, 0.444853, 
    0.8093558, 0.5496757, 0, 0.002437673, 0.227669, 0.2634807, 0.7164366, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9659117, 0.3167773, 0, 0.4677332, 0.5943365, 
    0.5637257, 0.8562685, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.8810632, 0.004721967, 0.05446313, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.2208384, 0.1411825, 0, 
    0.01509914, 0.3049383, 0.1022427, 0.001643809, 0.7302889, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 0.5155249, 0, 0.2220955, 0.925254, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9658247, 
    0.04132003, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.03023492, 0.1040698, 0, 
    0, 0.2589638, 0.8127933, 0.4118724, 0.5901706, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.6797279, 0.03147244, 0.148788, 0.8013205, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9649417, 
    0.2472448, 0.0001925075, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.2116711, 0.7594843, 
    0.04181511, 0, 0, 0.2791559, 0.9919224, 0.9871036, 0.5026899, 1, 1, 1, 1, 
    1, 1, 1, 1, 0.6875119, 0.1673929, 0.6100693, 0.9931602, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 0.9986221, 0.9031882, 0.02072693, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1597966, 0.6263976, 
    0.3037237, 0.3064115, 0.3001947, 0.9453359, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 0.9858415, 0.9203051, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9886171, 0.999054, 
    0.7919562, 0.001658652, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.106327, 0.9335366, 
    0.7329312, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 0.5367375, 0.8222567, 0.3355962, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.002422816, 0.6366513, 
    0.9978582, 0.7376231, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 0.998466, 0.4211002, 0.5821907, 0.06182952, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.2501551, 0.9984199, 
    0.2726648, 0.9098034, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 0.657743, 0.8075415, 0.4442849, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.221493, 0.713844, 
    0.009902901, 0.6008854, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 0.9938447, 0.7752694, 0.610476, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.006310866, 0, 
    0.1160645, 0.9701369, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 0.9781886, 0.1501769, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.5544846, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.7063521, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.5219765, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.9999979, 0.291099, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0005927939, 0.3538766, 
    0.271129, 0.9385704, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 0.8661439, 0.2963106, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.03236142, 0.5147032, 
    0.9229311, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 0.9242505, 0.07807732, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 zsurf =
  1.957085, 182.3516, 345.853, 566.5532, 583.9197, 703.0031, 841.8619, 
    930.701, 1327.418, 1866.999, 2029.211, 1998.469, 1606.435, 2058.914, 
    894.809, 267.2261, 1038.635, 95.99315, -29, -29, -14.74468, 50.54665, 
    131.9456, 149.8255, 180.3951, 144.0376, 117.0449, 65.4011, 47.57902, 
    52.56764, 62.57636, 88.29622, 103.0397, 116.2788, 146.1452, 149.0459, 
    260.9405, 209.8252, 240.3782, 305.7633, 380.0433, 410.2039, 401.1645, 
    344.6812, 350.6726, 420.6497, 639.9168, 1359.416, 1773.189, 1596.877, 
    1193.995, 945.0976, 478.8944, 313.0052, 364.5321, 544.9355, 728.1349, 
    913.1708, 1094.162, 1205.655, 1103.695, 1186.761, 1181.66, 1198.702, 
    1409.169, 1265.896, 1273.084, 1305.134, 1441.755, 1591.454, 1519.917, 
    1441.886, 1330.869, 1070.649, 1189.587, 1315.408, 1415.29, 1531.97, 
    1529.214, 1473.449, 1430.014, 1306.896, 1270.828, 872.1915, 165.6583, 
    2.112291, 1.155395, 0.02070807, 0.08559992, 13.39372, 105.9956, 72.41502, 
    2.817191, 0, 0, 0.04834903,
  0.02893994, 4.580082, 170.3799, 581.9701, 947.2767, 1071.069, 1146.666, 
    1154.808, 1640.017, 1900.844, 1998.073, 1884.909, 1641.079, 1859.79, 
    780.6656, 620.8061, 1727.327, 225.5852, -29, -29, -29, 38.14354, 
    126.9196, 155.8592, 184.8903, 179.1412, 129.6505, 97.10344, 37.13656, 
    33.23013, 51.04347, 71.70508, 91.74311, 103.1298, 126.9913, 145.6968, 
    179.7494, 230.5837, 298.0778, 375.3928, 434.7722, 459.8557, 350.7677, 
    343.3709, 347.6726, 356.1186, 381.6495, 446.8376, 603.9845, 758.576, 
    881.1244, 1095.882, 904.9011, 568.9519, 433.0408, 654.4484, 862.9261, 
    1147.874, 1391.479, 1546.497, 1694.146, 1655.956, 1846.877, 1863.535, 
    1773.414, 1861.801, 1658.115, 1432.014, 1446.591, 1505.779, 1598.366, 
    1639.378, 1501.092, 1183.134, 1002.323, 1205.448, 1280.397, 1347.836, 
    1565.089, 1583.707, 1551.659, 1326.685, 1098.686, 688.5358, 124.0418, 
    3.131963, 2.67241, 0, 0, 0.3741298, 0, 14.65283, 0, 0, 0, 0.08931515,
  735.5396, 867.0506, 660.6748, 924.9462, 1301.789, 1480.976, 1317.01, 
    1341.343, 1806.828, 2025.722, 2183.452, 2051.318, 1930.586, 1732.126, 
    665.5182, 1034.291, 2036.85, 544.5954, -29, -29, -28.76467, 38.63471, 
    172.218, 155.2569, 183.3024, 142.7022, 156.3304, 131.9387, 71.52921, 
    29.83442, 38.42982, 63.1153, 82.10826, 123.0225, 117.6491, 159.6424, 
    210.2419, 265.2799, 324.6303, 429.2385, 526.7354, 552.8436, 445.1412, 
    408.4677, 410.2799, 482.5757, 457.1882, 425.4275, 467.3434, 724.1971, 
    978.342, 1341.993, 1428.619, 1158.37, 714.2965, 634.1248, 1100.511, 
    1729.557, 2079.457, 2205.601, 2096.228, 1923.082, 2023.244, 2032.364, 
    2087.194, 1819.859, 1741.359, 1652.907, 1411.046, 1353.822, 1332.2, 
    1373.966, 1373.264, 1169.126, 951.4221, 1059.032, 1129.511, 1144.062, 
    1270.443, 1435.999, 1450.52, 1447.836, 1236.854, 758.832, 350.9756, 
    181.3987, 25.64147, 0, 7.676435, 3.285792, 0, 0, 0, 0, 4.333813, 55.45658,
  1304.387, 1437.602, 1376.26, 1494.452, 1659.236, 1723.898, 1639.994, 
    1657.578, 1850.001, 2092.416, 1922.954, 1856.68, 1913.263, 1612.252, 
    1244.188, 1688.415, 1823.349, 597.8655, -28.95335, -29, -29, 36.93167, 
    126.3385, 56.37119, 89.7822, 66.37797, 91.53525, 123.4684, 92.97884, 
    64.8284, 57.79882, 59.7579, 86.7978, 105.0893, 148.6383, 195.5772, 
    329.0817, 307.0089, 342.0926, 436.9752, 591.1713, 694.5746, 679.3177, 
    636.2111, 632.0756, 646.1209, 669.288, 648.6287, 782.5434, 883.3128, 
    793.3741, 676.8798, 926.3399, 801.6874, 746.4554, 1202.792, 1920.346, 
    2443.33, 2322.053, 1982.287, 1837.848, 1673.851, 1988.25, 2200.716, 
    1986.238, 1899.81, 1884.782, 1790.649, 1548.873, 1296.591, 1256.828, 
    1255.077, 1205.229, 1093.803, 927.5923, 972.8065, 1059.568, 1028.104, 
    1103.09, 1202.041, 1344.654, 1430.761, 1304.095, 857.4107, 614.5168, 
    408.0826, 142.5798, 1.184603, 40.65562, 3.480806, 0, 1.402507, 22.73934, 
    1.869505, 22.95708, 208.0578,
  1176.996, 1274.15, 1167.862, 1260.973, 1305.267, 1444.57, 1547.88, 
    1561.639, 1724.48, 1392.404, 542.0779, 297.3251, 709.7617, 908.8043, 
    1689.685, 1619.551, 990.7944, 115.7064, -24.46063, -28.99723, -29, 11.77, 
    -18.20284, -18.30782, -26.05886, -15.76914, 55.73129, 98.28559, 125.4715, 
    138.3384, 126.8703, 111.3977, 77.0961, 90.02938, 117.3675, 253.6755, 
    387.6956, 435.0849, 377.246, 411.8622, 531.7675, 673.597, 770.8846, 
    853.8765, 854.3976, 850.265, 792.6041, 745.4413, 733.783, 735.1926, 
    603.2223, 591.2675, 993.4567, 1367.18, 1860.522, 2238.518, 2511.91, 
    2284.058, 1663.224, 1322.216, 1438.35, 1776.375, 2169.013, 2455.426, 
    2488.388, 2387.191, 2351.167, 2100.744, 1704.273, 1439.597, 1375.393, 
    1281.368, 1147.538, 1084.584, 931.0007, 951.1368, 1033.676, 1018.033, 
    1023.891, 1108.402, 1268.471, 1365.725, 1364.301, 974.9635, 739.7955, 
    399.5302, 73.64684, 12.84806, 147.529, 5.471954, 0, 24.00544, 116.3721, 
    114.7116, 240.0056, 341.1817,
  1120.788, 1306.315, 1094.511, 1054.712, 1080.561, 1158.717, 1213.522, 
    1205.066, 948.7064, 166.4328, 0, 0, 7.011492, 766.0705, 1910.302, 
    1318.522, 220.8738, 20.13437, -22.87948, -28.96292, -28.99967, -28.96005, 
    -28.95333, -28.95845, -28.27328, -19.16533, 25.35257, 78.57539, 126.1784, 
    178.1593, 206.8317, 152.6626, 97.64114, 76.05511, 110.28, 209.1862, 
    385.8008, 487.759, 490.3545, 435.6064, 477.5195, 573.1337, 679.9717, 
    815.3858, 863.851, 795.056, 638.4842, 521.1765, 490.9408, 599.1897, 
    654.6764, 994.7811, 1491.828, 2086.955, 2473.281, 2589.081, 2203.682, 
    1937.777, 1327.908, 1322.338, 1643.389, 1980.04, 2347.152, 2586.005, 
    2474.671, 2249.25, 1973.765, 1742.107, 1577.967, 1488.696, 1454.051, 
    1334.462, 1222.04, 1055.741, 975.7679, 973.0269, 1098.012, 1137.429, 
    1093.573, 1125.746, 1300.224, 1360.541, 1194.296, 881.052, 581.177, 
    281.8254, 19.61534, 84.07046, 212.6468, 69.3125, 29.19267, 158.5775, 
    304.7471, 402.8232, 454.9509, 428.1056,
  1187.477, 1316.139, 1129.726, 991.171, 1030.374, 1016.187, 1020.988, 
    818.59, 381.7968, 0, 0, 0, 0, 1129.767, 1979.666, 998.5098, 264.3186, 
    59.78041, -4.723167, -24.42554, -28.50731, -28.65225, -28.92911, -29, 
    -28.607, -24.37205, 20.2152, 104.2612, 164.2149, 231.1236, 260.2584, 
    221.0597, 141.5681, 105.8174, 115.9729, 151.8276, 274.3087, 439.8468, 
    448.8825, 399.3673, 408.2239, 453.6656, 569.141, 609.5902, 626.4427, 
    521.6019, 365.9188, 284.7949, 285.1086, 423.1974, 846.5926, 1237.006, 
    1726.326, 2102.346, 2434.645, 2372.822, 2198.263, 1666.205, 1424.405, 
    1409.403, 1744.127, 2013.176, 2073.452, 2140.749, 2030.338, 1827.267, 
    1580.342, 1325.149, 1298.67, 1349.97, 1428.83, 1395.826, 1250.978, 
    1179.868, 1037.025, 1015.187, 1152.761, 1271.608, 1141.957, 1128.437, 
    1250.247, 1118.777, 820.3528, 513.1799, 459.0807, 201.0253, 50.98212, 
    173.3005, 353.3956, 272.952, 377.204, 340.7662, 338.8821, 282.7307, 
    42.52118, 0,
  911.2604, 1162.884, 1137.084, 979.4952, 1010.004, 1126.895, 1059.642, 
    869.5664, 252.7621, 0, 0, 0, 0, 1150.678, 1275, 595.7617, 273.573, 
    133.9935, 32.51972, -16.08583, -22.48619, -23.88273, -23.75681, 
    -24.06026, -24.22806, -20.21073, 10.21312, 100.5829, 164.7874, 248.1127, 
    306.6323, 287.0247, 220.7695, 169.7234, 135.2546, 137.2507, 172.6728, 
    311.0542, 341.0001, 327.2497, 348.4995, 425.6412, 463.1763, 447.4398, 
    353.7435, 252.8357, 186.9208, 193.5265, 269.0485, 416.4105, 833.4974, 
    1255.776, 1478.953, 1658.504, 2096.166, 2288.637, 1723.026, 1429.502, 
    949.519, 1162.872, 1667.993, 1924.058, 2051.646, 1868.885, 1679.083, 
    1502.363, 1410.3, 1248.582, 1158.49, 1393.645, 1598.457, 1420.972, 
    1293.249, 1159.699, 1133.274, 1037.51, 1155.602, 1250.937, 1090.242, 
    1007.832, 1146.141, 923.0365, 519.2554, 340.7791, 297.567, 152.0113, 
    84.55415, 319.1597, 474.4228, 619.5093, 846.3072, 366.6542, 0.09596219, 
    0, 0, 0,
  612.0165, 1024.829, 1129.861, 947.5595, 1080.557, 1194.547, 1150.219, 
    904.1955, 156.9333, 0, 0, 0, 0, 583.678, 439.6959, 309.7408, 232.4993, 
    133.5744, 75.71014, -1.082752, -7.73104, -16.27212, -16.11549, -15.90899, 
    -15.91451, -10.86247, 4.381418, 61.24113, 156.1658, 234.102, 316.4874, 
    335.1181, 275.5302, 255.234, 212.9649, 181.6552, 180.8939, 256.1131, 
    302.8167, 311.314, 343.6282, 353.8376, 353.0165, 257.5091, 195.26, 
    136.4342, 132.6939, 165.401, 204.5192, 263.7407, 417.9625, 651.0251, 
    757.1484, 1176.346, 1630.802, 1775.998, 1641.073, 1216.329, 1179.213, 
    1361.391, 1647.038, 1987.515, 2015.377, 1927.813, 1564.168, 1375.637, 
    1276.543, 1056.094, 1081.178, 1433.004, 1697.667, 1528.249, 1249.511, 
    1163.054, 1084.624, 1005.993, 992.0644, 1018.707, 950.4731, 940.6085, 
    1033.09, 798.034, 387.972, 229.6093, 197.4241, 132.7397, 211.0327, 
    408.1602, 644.9759, 902.4259, 1280.562, 421.0834, 0, 0, 0, 0,
  358.6493, 740.4105, 851.3992, 682.4423, 613.3671, 561.9201, 439.3097, 
    284.2988, 0, 0, 0, 0, 0, 164.7004, 99.19429, 101.628, 107.9559, 74.77886, 
    89.1244, 63.77163, 1.608809, -6.549558, -9.00685, -8.677175, -9.026371, 
    -3.706912, 1.230656, 51.11661, 139.9139, 209.1897, 282.7745, 328.7339, 
    305.7128, 303.4295, 269.2504, 220.6103, 194.5171, 252.9004, 301.2274, 
    362.1626, 362.2566, 319.3198, 217.928, 137.8181, 105.979, 105.6061, 
    114.0887, 135.0031, 185.067, 190.351, 191.2327, 234.4863, 323.938, 
    543.4288, 1060.478, 1268.447, 1192.681, 1328.727, 1228.022, 1216.701, 
    1586.167, 1872.411, 2054.413, 1874.194, 1613.623, 1458.215, 1250.402, 
    935.8388, 937.23, 1296.085, 1562.618, 1421.365, 1164.499, 1045.977, 
    969.0322, 885.1325, 801.2127, 811.7344, 891.5575, 953.3035, 938.8203, 
    644.8547, 285.5817, 157.9158, 154.0628, 172.5158, 282.7875, 469.8745, 
    706.7769, 1102.511, 1230.183, 277.3174, 0, 0, 0, 0,
  132.9001, 385.4105, 339.2654, 181.7644, 142.398, 0.8909621, 0, 0, 0, 0, 0, 
    0, 4.920471, 45.10483, 8.741613, 47.47253, 68.29308, 52.40722, 93.38539, 
    77.34655, 43.84061, 4.212869, 4.007848, 10.19131, 4.169814, 0.9422171, 
    9.296235, 56.39237, 118.7264, 170.1291, 210.7619, 320.4744, 331.2771, 
    318.584, 273.9849, 219.1942, 178.2944, 198.5368, 260.3773, 310.2903, 
    314.4893, 238.4738, 144.5557, 99.9539, 97.97208, 100.8626, 114.6869, 
    130.8342, 169.4516, 185.3304, 185.0731, 235.592, 278.8924, 478.6136, 
    764.5692, 685.5565, 811.843, 974.8875, 1184.866, 1309.973, 1492.49, 
    1975.901, 2111.276, 1920.701, 1584.152, 1393.754, 1227.47, 867.7672, 
    863.7648, 1180.989, 1434.811, 1408.729, 1119.982, 937.4036, 832.1047, 
    725.7586, 654.3876, 681.5729, 879.4352, 1001.297, 813.8375, 472.1414, 
    186.7852, 145.5977, 173.9421, 209.2027, 326.0379, 476.7007, 804.9005, 
    1109.927, 922.321, 75.55848, 0, 0, 0, 0,
  55.06753, 268.7123, 117.1969, 34.0993, 31.63307, 0, 0, 0, 0, 0, 75.30566, 
    123.2075, 25.73137, 4.677011, 0.4355646, 21.74989, 39.51146, 59.60038, 
    56.39664, 83.5396, 72.77475, 42.05199, 25.05266, 18.50826, 21.90979, 
    18.97606, 32.88521, 52.70894, 108.0705, 133.6327, 212.1806, 346.0227, 
    454.2986, 381.998, 286.2616, 211.4252, 172.9534, 157.5838, 173.7746, 
    195.4111, 173.0165, 139.0157, 104.9335, 99.12243, 103.3306, 100.5489, 
    103.4557, 134.8257, 162.8266, 185.8695, 232.4137, 269.2041, 308.7599, 
    614.8231, 747.6427, 544.698, 422.7588, 738.6674, 1183.856, 1471.337, 
    1606.683, 1839.523, 1757.208, 1367.475, 928.4243, 840.8771, 759.8136, 
    793.3425, 873.0726, 1079.337, 1313.67, 1351.702, 1047.42, 866.4039, 
    745.4284, 686.4276, 600.6986, 676.6058, 942.1893, 1006.475, 678.2116, 
    313.3897, 146.0503, 136.1638, 173.3874, 203.2215, 423.4491, 556.2217, 
    687.7593, 707.8784, 130.9646, 0, 0, 0, 0, 0,
  7.121133, 32.15426, 84.65013, 100.6684, 128.3299, 0, 0, 0, 0, 0, 37.53299, 
    141.1044, 20.04803, 0.0226125, 4.211974, 29.80108, 80.3756, 118.8334, 
    109.4529, 114.3332, 124.4319, 101.2349, 79.91515, 62.1116, 42.87167, 
    62.06577, 74.78121, 105.4743, 125.4183, 177.7379, 223.2901, 362.0724, 
    497.8951, 520.5967, 347.3084, 218.1198, 160.7832, 142.836, 141.2242, 
    142.3133, 130.3157, 119.2133, 114.2978, 107.0357, 102.9367, 104.6058, 
    110.6453, 123.0354, 142.3407, 155.8816, 175.0349, 218.0002, 336.6488, 
    481.0204, 622.3756, 464.2339, 567.8765, 821.3962, 1203.486, 1431.367, 
    1332.833, 1153.785, 908.6243, 652.9219, 598.5366, 569.8493, 665.6304, 
    778.8425, 895.4351, 980.2097, 1137.299, 1139.964, 917.5201, 727.8011, 
    697.3036, 645.4094, 611.8453, 750.6511, 997.3835, 898.4934, 452.9046, 
    187.9874, 131.9667, 132.1604, 162.3042, 257.2846, 519.6144, 578.7543, 
    534.0048, 299.177, 10.42934, 0, 0, 0, 0, 0,
  29.01102, 22.0339, 235.5383, 205.7878, 202.3339, 34.00895, 0, 0, 0, 0, 
    0.7499724, 39.96126, 8.142411, 27.61915, 77.46246, 141.4588, 165.7684, 
    167.3914, 132.9326, 131.5184, 138.1546, 130.3924, 147.073, 128.6659, 
    88.82133, 71.90593, 79.99207, 93.95091, 122.2475, 174.1009, 224.5994, 
    264.6025, 432.1731, 552.0823, 489.6333, 281.8752, 171.4949, 136.2069, 
    133.1193, 125.4225, 126.965, 120.7626, 111.4299, 101.8144, 99.97607, 
    113.2573, 118.6737, 130.7982, 136.456, 127.7007, 138.2258, 178.1324, 
    196.5107, 345.3022, 326.9236, 389.049, 456.8989, 544.9363, 644.9791, 
    795.9853, 714.1006, 626.2784, 512.6625, 545.9469, 686.3776, 774.8943, 
    722.8535, 808.6535, 999.6533, 978.3033, 988.0608, 965.1602, 774.5897, 
    743.5015, 720.1992, 658.6784, 645.7189, 780.3297, 934.1503, 668.8269, 
    269.4187, 138.0441, 142.1439, 151.7155, 169.5889, 303.9595, 540.4365, 
    608.5374, 528.3405, 294.674, 2.237589, 0, 0, 0, 0, 0,
  111.4144, 193.5326, 681.5145, 360.9993, 352.8302, 226.3572, 174.55, 
    37.86699, 0.2644904, 0.002788612, 0, 3.079878, 23.88782, 46.11481, 
    80.04777, 123.263, 147.1195, 144.2522, 130.5605, 152.2023, 141.6269, 
    132.931, 157.0246, 184.9375, 164.1916, 154.953, 124.2921, 92.66442, 
    103.1418, 164.1006, 233.3318, 178.8902, 210.3269, 409.1046, 418.7644, 
    336.8872, 189.2744, 130.1919, 111.7867, 105.783, 110.7427, 102.534, 
    94.83035, 91.60812, 107.021, 117.6856, 130.0774, 128.3777, 127.6499, 
    111.2988, 106.9357, 137.1521, 166.8579, 176.284, 241.0266, 287.8779, 
    322.1338, 316.6681, 333.3232, 405.2602, 465.2554, 453.8713, 526.2246, 
    631.4445, 775.7401, 794.0515, 706.1703, 873.7288, 1141.089, 1067.214, 
    1009.558, 878.1597, 765.5309, 814.0995, 825.5641, 682.4036, 688.0043, 
    821.9866, 793.0577, 482.589, 210.6379, 172.7338, 171.0665, 163.2869, 
    239.3744, 290.9917, 518.2194, 476.0343, 344.188, 253.0163, 199.3618, 
    0.09988576, 0, 0, 0, 0,
  396.4076, 461.4612, 931.6284, 727.4689, 459.6009, 316.0923, 161.0612, 
    61.08897, 39.84538, 14.21865, 16.21696, 14.69456, 42.59837, 83.79881, 
    96.42057, 106.7112, 127.726, 139.3746, 149.1176, 158.2953, 146.0142, 
    133.0698, 149.0564, 185.547, 219.5478, 236.7041, 204.2428, 142.1788, 
    111.0571, 152.1457, 197.096, 162.3448, 145.3164, 257.3849, 359.7718, 
    344.883, 231.0725, 134.1741, 96.72655, 77.17216, 67.97431, 71.95205, 
    78.97033, 92.42341, 106.5057, 121.7666, 113.3711, 112.7681, 100.1774, 
    90.3449, 93.89151, 126.1822, 144.4522, 167.8977, 184.3656, 222.1504, 
    216.4159, 276.5192, 273.3236, 330.4809, 405.03, 466.5895, 519.9902, 
    669.0401, 778.4682, 755.4747, 760.0569, 995.1483, 1292.865, 1133.658, 
    1035.321, 891.3419, 745.2759, 794.439, 820.8765, 731.4034, 825.5676, 
    816.8707, 654.7597, 365.2853, 254.1914, 241.2478, 251.6084, 300.0577, 
    283.1929, 314.035, 356.0846, 297.13, 224.8416, 403.2619, 439.1473, 
    0.3467962, 0, 0, 0, 0,
  855.1598, 709.2625, 1002.592, 837.1132, 519.1252, 130.5939, 71.12158, 
    81.11422, 142.1018, 51.00807, 96.93317, 79.51467, 95.48483, 129.0423, 
    140.4562, 103.5044, 126.4621, 151.7047, 177.8282, 174.2761, 156.9096, 
    144.2187, 154.5808, 180.015, 203.6465, 223.6183, 210.2678, 151.1036, 
    112.8854, 117.9561, 134.9364, 127.8695, 129.1225, 218.7797, 270.9187, 
    350.6521, 238.6366, 134.1218, 93.92628, 66.70253, 59.81225, 64.58974, 
    83.67481, 91.74277, 99.39961, 97.78426, 98.12943, 79.38904, 76.33865, 
    79.66943, 96.24992, 117.7307, 139.8467, 146.7351, 147.0995, 206.1468, 
    254.7715, 275.4333, 300.4858, 331.8605, 412.4602, 458.4528, 508.2016, 
    647.9883, 697.1085, 851.0264, 924.2222, 1209.887, 1389.744, 1105.53, 
    981.9774, 946.9201, 772.724, 746.0531, 774.8968, 822.0195, 896.6089, 
    762.1265, 469.3407, 356.1171, 319.8726, 356.8423, 393.546, 402.3568, 
    300.6212, 214.0752, 218.7073, 138.1364, 184.7563, 493.152, 362.86, 0, 0, 
    0, 0, 0,
  886.0403, 899.0963, 842.0179, 772.5779, 432.9344, 92.04449, 177.5087, 
    546.1584, 477.8832, 337.027, 119.8037, 133.9722, 151.3862, 176.6996, 
    157.914, 107.5661, 123.6268, 163.6318, 191.2482, 207.9477, 183.4089, 
    166.7186, 150.5348, 152.3792, 164.6893, 178.3489, 177.4384, 146.3247, 
    116.5272, 132.4336, 138.0589, 139.9558, 167.7014, 180.2253, 221.528, 
    303.055, 258.0195, 122.0804, 91.42705, 76.97997, 52.65008, 55.3461, 
    72.29636, 81.25592, 81.83448, 87.9664, 75.1608, 69.10935, 76.35617, 
    101.0703, 128.3883, 140.7466, 138.2242, 132.6284, 251.6389, 360.3346, 
    363.8312, 345.4504, 282.5562, 300.7509, 352.1882, 428.2724, 480.032, 
    508.1172, 638.3249, 969.0288, 1175.973, 1303.747, 1379.587, 1075.456, 
    939.7833, 971.2458, 876.7556, 679.537, 703.0974, 840.0677, 888.4769, 
    685.1582, 465.5422, 392.8445, 362.4918, 364.3657, 413.9269, 386.9064, 
    151.63, 102.4381, 140.1844, 97.34532, 357.6024, 508.7825, 100.0093, 0, 0, 
    0, 0.4358488, 0,
  377.0912, 777.9293, 847.1389, 613.7839, 347.3856, 183.928, 503.8705, 
    767.5604, 736.3063, 591.572, 261.3434, 142.1519, 203.053, 216.3297, 
    177.3449, 117.8392, 131.8621, 155.6192, 186.6643, 210.5387, 213.1024, 
    198.3484, 171.8902, 133.9252, 133.7206, 147.76, 149.0784, 123.2078, 
    117.5802, 128.9419, 142.8373, 162.3329, 190.3584, 196.8235, 191.6556, 
    277.8559, 336.0329, 136.4615, 78.44816, 67.13183, 57.19013, 45.63347, 
    56.64672, 62.35668, 62.41399, 58.50655, 64.08222, 61.68793, 82.98176, 
    109.022, 132.2926, 141.4133, 130.0148, 202.6298, 352.5894, 478.8041, 
    483.1053, 383.9174, 324.0171, 288.2619, 333.3291, 429.6476, 498.3948, 
    476.5586, 511.4784, 972.3265, 1117.176, 1333.446, 1231.988, 1100.885, 
    955.795, 961.8926, 865.2928, 707.8149, 605.3251, 700.6523, 739.4321, 
    558.5131, 402.4283, 297.584, 211.9652, 189.1523, 300.2366, 262.1036, 
    80.62009, 63.98812, 122.1838, 218.2967, 512.9334, 462.9636, 1.060671, 0, 
    0, 0, 37.38868, 81.3967,
  0, 594.21, 1018.811, 745.1058, 412.2401, 385.4236, 638.6064, 788.1194, 
    668.9521, 749.03, 562.7498, 197.1136, 243.5414, 257.3966, 197.9897, 
    130.8538, 123.876, 145.1576, 174.6566, 198.9581, 214.8165, 215.6441, 
    189.8338, 139.6603, 120.3094, 124.8503, 116.1674, 109.7017, 110.3707, 
    135.235, 142.0241, 170.4792, 213.9434, 209.5347, 167.4813, 264.8561, 
    348.0725, 240.3373, 75.87767, 79.91491, 71.83314, 45.36616, 48.33675, 
    52.77137, 49.97958, 59.72789, 63.37616, 71.72295, 88.81493, 109.8572, 
    136.8765, 144.6113, 151.7365, 193.6578, 319.4838, 403.0927, 398.4877, 
    411.3876, 349.0669, 324.9615, 351.6237, 448.8545, 494.1817, 457.7076, 
    444.8627, 679.2474, 972.8405, 1012.391, 1150.945, 1145.6, 1127.534, 
    944.8821, 822.8835, 703.0647, 531.0294, 464.5009, 428.4065, 363.7079, 
    263.4396, 211.7635, 198.9796, 267.8853, 350.3128, 264.7803, 65.758, 
    59.44502, 199.1785, 430.2982, 657.9562, 212.0221, 0, 0, 0, 97.63541, 
    113.3308, 41.61473,
  0, 399.1143, 1120.441, 820.4569, 297.3376, 195.9688, 434.3469, 519.7678, 
    533.1642, 758.1817, 711.3763, 342.4791, 278.5041, 278.4136, 214.2995, 
    149.314, 124.3232, 138.1995, 163.2455, 188.7315, 200.2267, 205.1242, 
    191.2654, 153.1303, 140.5527, 120.2366, 117.1466, 119.59, 127.6191, 
    134.2686, 149.6515, 164.0252, 186.4469, 196.4661, 161.6761, 177.2666, 
    334.9556, 307.35, 143.2057, 109.0354, 87.71973, 79.37965, 65.37148, 
    76.016, 76.0844, 78.8138, 85.20406, 92.65923, 120.6024, 124.1407, 
    141.3281, 120.2449, 152.1772, 252.603, 380.783, 423.7603, 464.9473, 
    420.7524, 383.9003, 365.9595, 382.3451, 404.967, 427.5276, 426.6728, 
    395.3827, 540.5605, 755.1957, 952.8699, 1084.376, 1365.629, 1383.233, 
    963.2598, 743.7776, 748.3361, 583.3853, 439.8699, 330.5274, 274.6473, 
    239.082, 218.2501, 375.178, 416.6259, 488.4598, 300.3638, 65.87481, 
    54.1222, 354.7472, 673.2607, 622.6516, 29.62266, 0, 0, 0, 206.3307, 
    149.5761, 0,
  0.003310259, 133.1911, 940.6332, 781.675, 248.0849, 90.08338, 116.6424, 
    220.5476, 304.2039, 419.5131, 703.8474, 411.9249, 301.6213, 267.3719, 
    209.3017, 160.7548, 131.8181, 134.4422, 157.0661, 185.6122, 207.0094, 
    210.453, 201.0542, 179.5661, 159.3497, 148.5723, 124.2159, 138.4398, 
    148.6608, 162.3591, 173.3146, 175.035, 184.1364, 181.5239, 173.0168, 
    157.8075, 250.5602, 304.8704, 179.2655, 67.08978, 85.99716, 73.47701, 
    103.1553, 107.7299, 100.9882, 96.31065, 80.26945, 83.55797, 94.24591, 
    113.5028, 87.01515, 83.67673, 216.3896, 356.1998, 462.2934, 496.7366, 
    464.9568, 424.9034, 395.8524, 405.8656, 396.2522, 369.3352, 362.0952, 
    392.2811, 403.4277, 532.8717, 897.1837, 937.3101, 997.2128, 1238.674, 
    1234.297, 916.9507, 798.6755, 785.5186, 683.3135, 527.7955, 404.3859, 
    329.3802, 251.766, 331.9852, 519.2047, 603.6315, 693.9681, 306.4999, 
    50.3644, 206.1701, 627.575, 741.8391, 292.8152, 0, 0, 0.002287545, 
    47.08162, 366.3271, 345.8133, 140.5091,
  0.1355318, 54.76622, 752.4495, 779.2272, 233.4452, 90.45777, 81.94717, 
    83.38457, 113.8429, 180.5548, 517.6541, 398.6514, 294.062, 222.6104, 
    177.3117, 146.8111, 135.3791, 142.748, 161.5963, 189.4258, 213.6966, 
    218.6755, 216.248, 169.9221, 153.2071, 133.3895, 136.4664, 149.2455, 
    169.6985, 177.9319, 169.0834, 158.8819, 153.8374, 154.3419, 155.6863, 
    159.3348, 168.2593, 263.9666, 210.4024, 63.44218, 42.57559, 53.28033, 
    74.75113, 94.46678, 84.90047, 77.8112, 56.29344, 41.15648, 64.81905, 
    77.03599, 86.15321, 102.1669, 314.0604, 390.679, 394.7146, 406.8066, 
    419.1735, 403.4146, 401.5237, 394.1876, 379.7701, 337.2509, 349.9233, 
    401.1396, 396.1155, 511.2408, 755.8575, 709.9775, 686.9054, 793.6512, 
    1004.453, 980.0493, 971.1741, 917.5543, 726.7474, 512.3557, 394.0262, 
    441.8013, 404.3204, 456.4452, 727.2965, 845.9907, 812.4409, 408.3134, 
    83.84931, 448.7415, 730.8319, 467.4902, 0.9863583, 0, 1.720724, 35.83591, 
    297.3234, 472.4654, 318.6473, 2.667824,
  2.786609, 2.644013, 504.1062, 684.3657, 243.8393, 124.4904, 120.2434, 
    118.8162, 136.5323, 274.2844, 459.7988, 323.3001, 252.3182, 197.7955, 
    158.2456, 143.8349, 155.14, 171.036, 179.7861, 181.361, 194.9534, 
    211.9559, 228.9097, 199.0386, 153.3901, 145.1039, 136.1797, 149.812, 
    166.3282, 157.6181, 154.2063, 126.907, 146.2792, 140.0006, 147.5358, 
    162.919, 152.3721, 222.5984, 246.1506, 256.06, 62.73549, 34.49001, 
    46.63019, 67.38826, 49.56528, 57.15746, 51.01564, 36.49106, 33.8912, 
    64.45266, 63.10199, 144.3528, 351.2276, 400.1565, 401.1474, 439.6917, 
    469.2003, 431.5126, 411.8654, 369.9917, 321.8169, 323.1301, 326.4559, 
    382.4082, 378.7637, 344.4705, 461.5488, 414.4735, 376.186, 542.0886, 
    713.6682, 832.4791, 967.1309, 1007.369, 852.7335, 704.9957, 550.9443, 
    581.854, 539.4864, 852.6191, 1003.918, 778.0033, 665.1097, 266.5093, 
    311.5761, 683.8643, 705.9689, 96.01817, 0, 1.189999, 8.842051, 47.33828, 
    140.6496, 324.6157, 137.269, 0,
  276.4731, 0, 179.3712, 525.0765, 251.7486, 132.691, 157.0414, 154.7416, 
    302.1239, 580.2548, 583.1707, 323.0918, 206.9382, 174.8136, 156.9467, 
    158.7047, 172.3876, 199.9602, 184.0974, 164.6234, 165.0962, 185.8372, 
    203.0004, 193.7835, 175.1679, 146.9807, 142.3714, 150.1652, 157.6037, 
    163.3478, 129.6109, 129.2951, 159.414, 161.3647, 162.9705, 181.9612, 
    128.0042, 147.4346, 353.2044, 345.6928, 272.2606, 81.65241, 31.30544, 
    29.65827, 24.55814, 44.82172, 50.73238, 36.99446, 29.24441, 45.64774, 
    56.69508, 147.8097, 350.2406, 446.015, 517.4972, 568.1435, 509.0543, 
    480.6918, 464.3664, 407.0969, 359.9652, 325.3537, 336.1723, 338.7549, 
    334.156, 299.1234, 313.2734, 332.2038, 383.9116, 472.8965, 632.2615, 
    813.0618, 1026.41, 1103.619, 1136.821, 1031.338, 975.8419, 689.2612, 
    568.7227, 943.745, 852.9982, 485.5357, 236.3455, 271.7433, 463.5656, 
    614.2126, 345.1251, 0, 16.48282, 105.6186, 7.521848, 0, 0, 87.10019, 
    40.73374, 0,
  508.8716, 70.13601, 6.784113, 372.3694, 322.6259, 293.2125, 242.353, 
    173.0082, 268.3181, 591.1161, 536.0643, 296.8539, 202.5906, 164.5604, 
    144.654, 150.5097, 161.7568, 165.6213, 170.2032, 147.5072, 145.3487, 
    118.8593, 111.2818, 111.6931, 136.4204, 155.4414, 171.5328, 140.8391, 
    169.3844, 138.0114, 124.348, 104.4207, 145.8794, 164.8125, 186.8414, 
    188.481, 126.0499, 90.26923, 110.4248, 252.1565, 185.2361, 152.9825, 
    177.3863, 27.33101, 14.74302, 22.59383, 32.78283, 24.52886, 36.56748, 
    50.80676, 80.63863, 201.0317, 398.6272, 570.3611, 631.2753, 643.4182, 
    537.705, 514.1293, 540.4216, 502.6988, 444.1647, 409.5107, 358.6469, 
    313.3456, 229.5331, 227.212, 262.0572, 326.5652, 403.6352, 469.1498, 
    543.0381, 673.6775, 820.8776, 1047.744, 949.5495, 1148.552, 1111.228, 
    855.2848, 484.6896, 661.6188, 513.8441, 249.184, 299.0674, 415.421, 
    493.6745, 252.4404, 5.99207, 59.10885, 97.5045, 79.21317, 10.46941, 0, 0, 
    43.29576, 3.355622, 0,
  443.5912, 255.1915, 0.09644534, 195.873, 487.8073, 735.0255, 695.2324, 
    348.3268, 280.6532, 412.6371, 385.954, 220.2776, 204.6375, 127.3774, 
    125.8829, 139.0522, 124.0497, 124.0424, 125.5306, 122.1397, 132.0455, 
    96.83639, 60.97416, 63.26183, 70.19158, 96.56532, 138.9745, 127.6716, 
    134.1593, 150.0386, 90.46266, 84.52273, 112.2292, 121.4295, 151.5019, 
    166.1176, 108.1869, 79.91405, 92.42285, 97.96801, 124.7679, 221.8664, 
    228.2843, 115.3288, 24.56494, 14.8802, 20.65261, 31.73664, 49.24442, 
    60.99174, 105.08, 244.0706, 521.9723, 723.241, 767.3787, 664.4177, 
    487.5122, 513.0247, 515.0753, 538.3448, 511.0675, 463.2043, 376.3399, 
    264.3518, 201.9225, 193.3568, 293.2623, 334.261, 373.6343, 439.8721, 
    490.5887, 493.9969, 600.4854, 755.9476, 924.3199, 950.3077, 1052.388, 
    779.1483, 183.5563, 265.7245, 179.8311, 213.6126, 282.3783, 202.5462, 
    128.2361, 30.74742, 219.925, 102.526, 0, 0, 0, 0, 0, 16.26684, 0.6956787, 0,
  260.7036, 393.7766, 11.27141, 23.8249, 678.2915, 1205.305, 983.3217, 
    600.5497, 405.7943, 426.7081, 384.4165, 217.486, 141.1087, 113.0105, 
    118.703, 126.1676, 90.83533, 74.9175, 85.22266, 86.1847, 108.5499, 
    97.74491, 85.57736, 64.07814, 40.13272, 24.09916, 78.24743, 80.76043, 
    124.5104, 132.6886, 90.25305, 50.69267, 81.38572, 64.80839, 89.60198, 
    115.1036, 102.3747, 89.09599, 91.98434, 106.8285, 90.62163, 137.0851, 
    183.7695, 40.38134, 27.67106, 11.31515, 23.2658, 37.70986, 46.24703, 
    62.2045, 86.09678, 336.5412, 717.0566, 919.0491, 854.2428, 596.1452, 
    380.2888, 384.9098, 468.5178, 498.7417, 522.8006, 451.6152, 351.5222, 
    233.9609, 161.0052, 184.1114, 234.4022, 294.4582, 302.137, 342.4128, 
    411.9693, 392.7577, 351.6703, 590.9839, 653.2507, 725.2677, 801.4582, 
    656.3619, 55.66471, 28.70166, 97.66091, 137.6178, 146.7572, 75.24693, 
    99.51981, 291.1764, 193.6622, 6.543282, 0, 0, 0, 0, 10.53877, 52.14492, 
    0, 0,
  43.77597, 464.1584, 56.89383, 468.3003, 1272.138, 1580.384, 1018.172, 
    560.8243, 492.4376, 414.2195, 387.2528, 175.9947, 96.38813, 88.09875, 
    109.2793, 71.96533, 25.01822, 58.2986, 73.01802, 38.57325, 49.70271, 
    62.90857, 57.06133, 27.90662, 27.32676, 23.32841, 78.08787, 112.5397, 
    118.9064, 113.533, 66.1688, 38.50869, 78.81353, 50.76294, 38.3057, 
    62.43602, 80.58298, 45.74772, 40.23263, 38.5184, 22.24349, 97.94888, 
    42.41491, 12.44253, 28.08678, 14.85801, 30.86785, 37.11079, 35.73439, 
    33.91776, 124.3871, 381.5867, 780.6381, 921.0138, 807.3401, 514.1893, 
    283.6758, 323.1736, 314.6895, 374.642, 395.0815, 392.9985, 310.7736, 
    226.0156, 184.2313, 147.4343, 164.883, 202.6225, 252.7558, 260.424, 
    307.9431, 309.5395, 311.4832, 401.2553, 517.3415, 550.1964, 679.3637, 
    525.896, 1.616105, 2.896513, 88.79086, 59.5556, 70.75466, 69.71838, 
    122.3319, 154.2911, 15.59744, 0, 0, 0, 0, 0, 27.71455, 6.569491, 0, 0,
  0, 439.4178, 195.6855, 907.5368, 1805.264, 1501.639, 712.643, 483.2295, 
    497.7593, 420.5321, 315.0768, 136.8431, 80.70911, 102.5947, 110.8975, 
    56.06786, 0.2648131, 3.387826, 36.63493, 22.48626, 4.213938, 32.13628, 
    34.12004, 9.394886, 55.34244, 71.22887, 124.1325, 164.2337, 141.1722, 
    73.3173, 29.08077, 2.917876, 50.12897, 16.72008, 8.767165, 20.09276, 
    6.12492, 9.995467, 2.303684, 0.02967453, 7.202766, 15.59999, 0, 4.923676, 
    28.76822, 14.64493, 19.81721, 22.2378, 29.72172, 55.51414, 46.22926, 
    135.3196, 311.9851, 389.0701, 426.3514, 394.7778, 346.0056, 381.4013, 
    311.8159, 286.077, 316.2218, 321.0644, 306.4557, 227.0812, 163.6294, 
    111.7403, 127.4932, 171.2171, 128.8476, 186.4454, 234.3389, 277.8444, 
    263.8623, 387.7439, 507.9923, 593.5289, 671.5868, 151.9244, 0, 0, 
    0.1526855, 11.12141, 27.27045, 5.642293, 0, 0, 0, 0, 0, 0, 0, 0, 
    29.69389, 0, 0, 0,
  336.1212, 283.2744, 280.2505, 1349.746, 1791.143, 1240.253, 581.5303, 
    454.5894, 529.9597, 451.9621, 271.3024, 88.98106, 65.69213, 79.26176, 
    83.76402, 15.86282, 0, 0, 0, 0.01159282, 3.559813, 3.361201, 26.5549, 
    78.995, 104.8708, 111.296, 123.7502, 183.7094, 170.4765, 96.75568, 
    18.82452, 36.92904, 173.0009, 147.0736, 0.6561724, 40.09827, 1.400087, 
    18.67419, 0, 4.921213, 17.68606, 0.02064603, 0, 0.5728964, 18.75198, 
    13.3812, 8.656983, 8.488718, 38.44683, 61.09453, 51.83106, 52.62397, 
    58.6014, 59.39347, 165.6035, 290.221, 454.3603, 531.7468, 356.0366, 
    250.5548, 230.6507, 267.4886, 263.0035, 170.9993, 101.3395, 226.0812, 
    405.6003, 438.8228, 243.4076, 140.5213, 194.1314, 222.0123, 325.5292, 
    476.0626, 621.8958, 708.6229, 614.3857, 5.007009, 0, 0, 0.5131387, 
    10.68596, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 30.96639, 0, 0, 0,
  1014.961, 1059.676, 999.4585, 1486.217, 1353.48, 822.1008, 483.4728, 
    423.429, 432.9811, 400.1913, 184.7545, 59.76541, 51.08024, 32.45238, 
    3.397727, 1.339373, 0.5192116, 1.949396, 6.878533, 0.8359628, 0, 
    0.4469217, 32.46057, 94.17204, 138.7826, 139.0123, 142.075, 170.2651, 
    199.8437, 156.3874, 66.95568, 99.59976, 214.9215, 163.2938, 0, 
    0.00557197, 0, 0, 0, 37.75103, 85.04147, 0, 0, 0, 2.593199, 6.704577, 
    0.9132928, 2.0938, 109.5198, 89.66087, 71.78169, 61.52934, 55.7276, 
    50.0367, 66.96713, 204.8958, 385.6734, 415.6871, 273.868, 163.4537, 
    185.3572, 235.6016, 183.325, 121.5506, 331.4378, 656.7086, 973.7778, 
    936.9366, 698.6102, 315.4651, 158.0312, 304.8352, 599.1711, 767.9793, 
    739.1931, 587.2299, 272.567, 0, 0, 0.0005063568, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.3449626, 0.8638448, 0, 0, 0,
  1276.519, 1596.647, 1710.525, 1532.737, 942.0485, 525.4172, 468.8974, 
    340.8898, 335.7376, 367.5742, 202.7082, 87.97628, 47.15509, 23.6611, 
    2.109894, 16.11546, 63.89506, 99.67946, 35.14595, 6.804534, 11.33926, 
    3.489694, 4.426375, 51.48684, 116.296, 132.7959, 119.1194, 141.0041, 
    206.496, 213.7981, 189.8233, 189.694, 225.2005, 137.5171, 0, 0, 0, 0, 0, 
    51.36637, 209.3645, 35.64569, 0, 0, 0, 0.1678525, 0, 0, 2.154153, 
    17.08876, 89.85088, 131.7713, 127.0772, 66.14963, 54.64122, 98.0938, 
    154.5197, 216.6144, 122.0288, 144.2869, 194.6717, 195.0684, 113.4059, 
    305.1859, 773.1769, 944.6837, 944.9396, 1041.262, 1010.897, 714.8572, 
    441.2517, 615.52, 994.8956, 1017.131, 735.3895, 398.553, 39.48136, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16.48005, 0, 0, 0, 0,
  576.1854, 931.6247, 906.6362, 782.9591, 492.1016, 465.3861, 284.8566, 
    247.166, 278.3712, 328.5902, 197.9191, 70.77742, 37.59184, 12.53315, 
    7.181137, 43.26176, 121.2297, 201.0618, 133.2232, 65.32127, 50.51119, 
    18.33489, 0, 0.11232, 20.32129, 27.82987, 23.76683, 29.30825, 141.2721, 
    243.3896, 253.101, 230.2507, 183.3705, 51.35647, 0, 0, 0, 0, 0, 0, 
    70.44017, 221.9524, 66.5798, 0, 0, 0, 0, 0, 0.3017679, 8.757327, 
    127.2703, 222.3685, 176.8489, 129.8425, 56.31729, 30.53881, 53.13721, 
    56.63842, 85.90793, 110.0528, 170.028, 155.7422, 181.1576, 658.582, 
    891.925, 765.0097, 566.7166, 683.1484, 938.3599, 946.0663, 950.6962, 
    1152.784, 1400.864, 1190.112, 699.8245, 303.8513, 1.38781, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 4.373055, 0.3063857, 0, 0, 0, 0,
  645.5978, 651.4741, 348.0461, 338.1821, 333.729, 297.324, 274.5483, 
    329.6071, 320.4292, 242.4523, 142.7768, 33.2918, 19.17206, 13.50416, 
    14.204, 8.873847, 37.03663, 147.5774, 138.1909, 116.1385, 174.9569, 
    163.6211, 73.71962, 29.18241, 51.88186, 92.01063, 38.92251, 26.84706, 
    114.0117, 203.6541, 270.5715, 215.7726, 151.7382, 14.68677, 0, 0, 0, 0, 
    0, 0, 0, 40.54074, 369.3293, 317.3165, 114.3371, 3.862887, 0, 0, 0.11153, 
    0.006048144, 19.55387, 142.5781, 154.5665, 123.9076, 179.1985, 79.16, 
    14.5393, 34.07465, 42.74265, 97.64807, 169.0159, 219.1613, 396.9012, 
    642.2534, 732.5916, 397.1309, 377.0508, 643.4995, 985.1297, 1109.908, 
    1146.201, 1363.316, 1434.265, 1369.427, 928.765, 436.3409, 111.6556, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5.772016, 0.006933623, 0, 0, 0, 0, 0,
  832.0802, 796.4195, 452.5931, 305.7719, 293.3802, 263.662, 251.0075, 
    350.6158, 214.3606, 118.4772, 23.99523, 9.823727, 0.9374197, 9.133391, 
    30.28316, 31.31364, 7.673902, 30.12636, 73.6406, 163.2412, 282.5515, 
    383.3724, 343.9316, 270.9898, 269.3295, 315.7319, 274.4701, 208.2753, 
    218.7913, 263.5744, 306.8953, 271.2532, 182.3894, 67.36945, 0, 0, 0, 0, 
    0, 0, 0, 0, 5.676641, 71.09753, 100.5261, 93.03223, 0, 0, 0, 0.029983, 
    0.2834589, 5.7791, 29.0103, 202.0174, 299.2979, 245.8783, 10.45641, 
    3.441845, 9.227307, 65.13091, 143.5608, 212.5292, 258.0329, 406.613, 
    314.3367, 276.2676, 445.5888, 781.3271, 1096.255, 1218.235, 1079.923, 
    998.8617, 1214.761, 1232.076, 1011.277, 597.6057, 136.1366, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 2.308824, 17.42456, 0, 0, 0, 0, 0, 0,
  522.8505, 646.8199, 434.2559, 254.1983, 198.1381, 141.3106, 157.4017, 
    202.436, 98.83956, 4.720938, 5.80146, 1.222248, 0.002537446, 0, 6.751021, 
    16.09051, 4.110047, 0, 67.87675, 217.9813, 406.6455, 577.1392, 615.5616, 
    464.1506, 415.4912, 491.5859, 515.1653, 499.5445, 526.2872, 472.2782, 
    484.1233, 346.7195, 209.6823, 28.12877, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.04541712, 0.1208085, 35.22072, 93.14128, 169.8435, 
    92.35309, 0, 0, 0.01013316, 4.865694, 16.84927, 23.22182, 27.02969, 
    119.0616, 246.3213, 518.4421, 657.4585, 736.8021, 1052.213, 1052.852, 
    1112.684, 1157.132, 1119.51, 1128.288, 975.9925, 711.0227, 271.4639, 
    11.86194, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10.20065, 51.1852, 0, 0, 0, 0, 0, 0, 0,
  189.5987, 372.6584, 272.8972, 153.0684, 129.0797, 107.2802, 101.2548, 
    98.52764, 13.1368, 0.6186931, -0.0932398, 0.01887309, 0, 0, 0, 0, 
    5.934471, 249.3546, 496.3241, 641.0406, 712.6684, 883.3423, 769.7581, 
    568.9565, 546.6921, 654.5696, 742.6288, 773.7735, 770.8872, 664.8349, 
    517.9086, 240.3035, 48.13427, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 25.80465, 75.88532, 127.7064, 5.597481, 0.01321575, 0.01744381, 
    0, 0, 0, 0.008600875, 0.2463465, 0, 3.196367, 26.82889, 218.4336, 
    438.3653, 500.2625, 445.5697, 536.2654, 907.6587, 1133.265, 1245.885, 
    1148.132, 918.5613, 905.1179, 873.1757, 565.6349, 139.6936, 9.307497, 0, 
    0, 0, 0, 0, 0, 0, 5.973339, 51.01183, 18.53154, 0, 0, 0, 0, 0, 0, 0,
  66.53913, 126.0707, 158.3924, 101.3495, 129.9872, 153.1423, 111.0585, 
    69.88337, 5.909921, 0, 0, 0, 0, 0, 0, 0, 6.110831, 443.8941, 822.0618, 
    1065.257, 1147.54, 1026.579, 615.9289, 217.0476, 161.5421, 240.8548, 
    308.3307, 226.1226, 224.5132, 167.3122, 91.86687, 2.702835, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 1.687579, 0, 0, 0, 0, 2.009178, 150.2296, 
    137.6718, 53.3191, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01111945, 8.059679, 
    76.88058, 223.2468, 192.0626, 54.48991, 351.7439, 523.5924, 854.4131, 
    841.848, 774.7855, 709.6036, 701.8489, 900.449, 776.0449, 283.2952, 
    20.40456, 0, 0, 3.21502, 41.93052, 145.8842, 257.1946, 238.5102, 
    233.1759, 92.08567, 0, 0, 0, 0, 0, 0, 0, 0,
  10.54719, 38.52236, 89.41316, 88.45621, 129.8748, 140.0378, 1.758609, 
    3.622372, 20.79722, 16.84281, 3.764497, 0, 0, 0, 0, 0, 0, 9.974582, 
    203.0671, 552.9215, 723.358, 628.1764, 114.8102, 1.827135, 0, 0, 
    0.02597354, 4.145141, 11.91014, 1.813728, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 2.070437, 19.12915, 65.26246, 40.89855, 0, 1.946335, 0.4316256, 
    4.962647, 138.3129, 0, 0, 0, 0, 0, 0, 0, 0, 0.7391827, 0.9985219, 
    0.398542, 4.360011, 16.71775, 12.17988, 71.93053, 79.30731, 98.12679, 
    133.4162, 234.3277, 244.6326, 294.9109, 406.4966, 458.4559, 607.9581, 
    806.5295, 651.6235, 97.59635, 26.42796, 0, 11.91634, 142.9294, 523.1003, 
    623.8453, 728.3721, 414.541, 179.0205, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0.2375568, 35.22453, 45.78533, 100.8335, 98.73385, 0, 19.24257, 
    69.95895, 49.19936, 14.10529, 0.5963095, 0, 0, 0, 0, 0, 0, 0, 14.52876, 
    100.917, 29.60974, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.002305, 0, 0, 
    0.049075, 0, 0, 0, 0, 10.97873, 31.62269, 20.17602, 8.189528, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 24.33025, 35.88162, 3.392136, 8.202249, 
    9.667623, 4.784458, 29.97687, 95.48793, 70.86581, 107.1511, 47.01993, 
    186.0479, 250.5408, 327.3635, 495.9941, 663.1337, 707.337, 343.3452, 0, 
    0, 12.89661, 177.2778, 526.8167, 650.3031, 730.8545, 475.256, 140.5307, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0.1563355, 32.96153, 93.6973, 8.055909, 7.271522, 46.84789, 107.1797, 
    96.87433, 65.0823, 5.47474, 1.638984, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 46.7029, 45.70561, 2.701415, 
    1.950268, 1.063997, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1.490511, 10.38847, 0.8451264, 0, 0.1427283, 5.747555, 26.19526, 
    79.84738, 54.79946, 32.89713, 97.37908, 252.4611, 375.3538, 398.1776, 
    596.9442, 749.3185, 517.8513, 3.130794, 0, 0, 92.81933, 348.3482, 
    500.1969, 715.4668, 515.3165, 78.95136, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 23.82193, 117.2348, 1.692671, 2.966081, 75.61375, 119.2401, 
    156.9432, 150.2247, 187.7098, 168.4926, 20.22646, 0, 0, 0, 0, 
    0.008525716, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 112.4393, 
    187.7537, 277.7043, 196.2434, 63.29765, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0.6239529, 13.39494, 0, 0, 0, 1.266546, 41.70436, 
    25.22967, 28.20456, 109.732, 279.7055, 394.6047, 507.9118, 776.3243, 
    775.1523, 364.5099, 50.67634, 5.433064, 185.3506, 421.2495, 414.1049, 
    393.2517, 297.5771, 294.7875, 7.586363, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 2.931184, 22.6025, 0, 26.93795, 109.4093, 139.878, 177.1416, 
    88.31774, 86.30247, 174.0245, 163.1162, 240.8645, 75.69065, 3.21588, 
    0.5801046, 6.936382, 0.1045908, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 1.200257, 139.026, 418.142, 149.2554, 1.2402, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.164914, 0.7948571, 0, 0, 0, 
    0.001168255, 16.67364, 19.89136, 43.50631, 130.2915, 266.5667, 415.8081, 
    554.9022, 713.0673, 638.9822, 273.1252, 216.0703, 123.0732, 400.6276, 
    240.1565, 113.1827, 94.77327, 41.31813, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 12.43825, 0.1656403, 16.24762, 3.12718, 2.06611, 
    13.84467, 122.0781, 227.2487, 363.1719, 217.4649, 58.97001, 0.598401, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4.693333, 86.21237, 
    0.054159, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    9.497975e-05, 0, 0, 0, 0, 0, 4.237197, 6.721555, 63.53002, 114.1027, 
    265.6567, 554.0557, 724.3539, 712.1773, 539.7785, 160.6944, 68.24227, 
    103.9293, 73.31152, 28.09826, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0.03340246, 0, 4.537661, 95.45872, 73.8838, 90.62366, 
    59.25259, 54.20035, 152.8858, 94.76863, 8.248804, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1057689, 19.82886, 
    233.0814, 269.9969, 373.4673, 617.0306, 770.7498, 660.8774, 426.0227, 
    199.58, 211.4468, 198.4001, 14.72842, 0, 0, 0, 0, 15.84741, 3.091941, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 68.96684, 105.0802, 102.1657, 102.4648, 46.12123, 
    0.1862036, 4.137225, 14.37615, 0, 0, 0, 5.570907, 19.88484, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1777319, 
    320.2881, 508.4323, 575.6027, 669.407, 672.3879, 490.291, 289.8031, 
    238.265, 313.8378, 200.7386, 9.265935, 0, 0, 0, 0, 0.1091187, 4.402359, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0.1957944, 113.7033, 75.3949, 52.71202, 37.44812, 
    0.2004635, 0, 0, 0.123569, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    13.78675, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5.807943, 138.4678, 
    425.4565, 693.1362, 582.7962, 419.3349, 270.5754, 275.724, 489.4667, 
    545.7513, 206.3423, 1.7709, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 20.8598, 0.006193054, 2.341495, 0.4137827, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.4644903, 19.146, 0.3230906, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 76.46013, 93.74072, 366.0079, 
    496.2035, 424.2791, 175.4117, 154.8367, 347.1221, 670.9517, 666.6006, 
    261.9197, 13.65668, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6.259748, 
    120.2423, 2.125335, 0, 0, 0, 0, 0, 0, 0, 0, 0.5916959, 0, 2.078349, 
    11.29419, 52.72276, 269.5899, 324.7525, 54.04507, 40.68792, 0.01734185, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    27.23831, 326.5949, 448.5767, 470.8265, 265.0998, 97.36693, 175.0721, 
    356.4594, 464.9758, 296.394, 24.18855, 0, 0, 0, 0, 0, 0, 0, 0, 6.498864, 
    0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 434.9876, 
    549.625, 194.8289, 0, 0, 0, 0, 0, 0, 0, 49.79148, 229.9053, 270.3666, 
    218.3152, 435.0714, 763.8671, 711.7297, 577.2573, 432.7135, 282.8728, 
    35.13057, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 9.57939, 23.93509, 458.746, 758.4965, 540.113, 253.5558, 102.6653, 
    138.8913, 305.0443, 234.599, 15.73475, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    26.66078, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7.860931, 
    705.9603, 764.272, 264.1802, 0.009830754, 0, 0, 0, 26.49382, 30.51307, 
    107.7551, 497.813, 1169.735, 1488.845, 1487.634, 1470.97, 1528.288, 
    1292.458, 1079.739, 876.5819, 425.0653, 38.33871, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9.993676, 78.49228, 0, 
    302.9012, 626.1432, 557.4089, 253.4888, 65.42033, 56.02234, 195.751, 
    71.06109, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.04533782, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 39.38756, 
    486.9271, 529.4836, 132.7024, 0, 0, 0, 188.4812, 192.5964, 498.543, 
    708.6475, 1124.227, 1743.003, 2079.127, 2174.609, 2030.333, 2037.837, 
    1968.742, 1794.981, 1306.613, 536.4325, 38.71229, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.2987449, 0.9965169, 0, 
    24.91258, 299.2193, 349.5217, 135.9241, 25.71449, 1.858234, 83.3325, 
    37.25776, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.5446421, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.008149051, 
    79.37028, 181.9968, 190.1527, 16.7675, 0, 13.55061, 980.6506, 768.5872, 
    1105.977, 1530.174, 1995.253, 2289.703, 2406.146, 2417.229, 2295.283, 
    2278.623, 2349.081, 2062.894, 1572.461, 794.2656, 199.4317, 65.12003, 
    90.86436, 1.968355, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 58.45197, 215.2836, 156.8912, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 1.912825, 3.799026, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    10.55764, 11.55569, 0, 0, 140.3663, 1585.396, 1665.679, 1860.954, 
    2327.909, 2685.942, 2719.711, 2651.773, 2599.41, 2509.09, 2444.553, 
    2411.1, 2231.088, 1777.786, 1073.075, 389.2512, 394.257, 742.5377, 
    431.4628, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 6.323763, 161.9636, 163.3663, 42.97362, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.2813061, 5.751188, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 162.3825, 1830.881, 2420.234, 2799.512, 2933.921, 3054.115, 
    3021.108, 2897.282, 2813.163, 2631.317, 2454.22, 2377.28, 2253.893, 
    1763.675, 967.3515, 294.468, 567.5514, 896.8688, 723.8139, 165.1352, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22.55821, 
    205.1908, 176.4454, 100.5338, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5.576109, 1.351869, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 224.3244, 1715.302, 2661.883, 3042.112, 3078.042, 3083.966, 
    3056.699, 2966.114, 2775.983, 2461.252, 2203.078, 2069.804, 2055.312, 
    1617.411, 858.8635, 63.53865, 565.2546, 820.6309, 464.1451, 208.9816, 
    21.89472, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.308722, 
    41.45142, 0, 0, 39.56498, 1.861557, 0.9454954, 8.430882, 0, 0, 0.2580895, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 15.21186, 1.925179, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 69.28409, 1442.782, 2432.051, 3022.305, 3064.017, 2982.046, 2920.952, 
    2867.871, 2768.787, 2520.354, 2211.113, 1641.312, 1364.499, 1291.194, 
    1387.434, 845.2209, 244.3112, 296.0118, 614.2589, 358.0775, 523.442, 
    111.5307, 0.1241507, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6.110101, 52.63713, 243.9889, 184.6683, 0.4007951, 7.643325, 46.26271, 
    0.01746987, 11.53573, 9.214417, 0, 0, 2.880076, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 20.27884, 0.2822629, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 388.4866, 1897.231, 2823.74, 3016.014, 2869.568, 2752.483, 2647.189, 
    2529.865, 2443.268, 2159.798, 1604.969, 955.6561, 423.3286, 422.3328, 
    778.8141, 553.3457, 156.9905, 464.2124, 635.9963, 351.1034, 437.6381, 
    20.91868, 26.49133, 1.27366, 1.299142, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 3.944896, 32.97338, 270.1112, 460.1797, 328.6203, 29.76436, 98.42758, 
    162.2669, 21.47914, 0.01439463, 0.09217066, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.01224168, 16.85926, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 220.2471, 1591.738, 2466.678, 2747.279, 2660.819, 2426.795, 2163.563, 
    1904.25, 1726.834, 1309.499, 717.4695, 72.1908, 0.01969476, 0, 139.6303, 
    56.38565, 0.01733694, 280.8316, 373.5753, 88.71832, 60.37281, 22.64031, 
    35.58979, 1.627476, 11.44019, 3.820878, 2.149208, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.01889744, 6.854713, 95.4062, 415.7192, 609.9531, 237.4828, 87.95111, 
    174.6365, 179.5905, 1.821839, 0.4608677, 1.038414, 1.955436, 0, 0, 0, 0, 
    0.4032466, 0, 0, 0, 0, 0, 23.75265, 6.992056, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 344.95, 1579.479, 2305.747, 2500.39, 2205.512, 1810.193, 1200.209, 
    851.3199, 495.871, 307.6716, 18.7188, 0, 0, 0, 0, 0, 0.007190464, 
    328.6132, 334.6894, 151.1666, 47.72522, 19.96992, 2.669097, 2.000999, 
    5.087904, 39.56742, 29.48166, 1.290598, 0, 0, 0, 0, 0, 0, 0, 0, 7.210662, 
    34.74933, 341.6028, 763.1323, 677.7067, 334.8472, 120.0849, 233.7542, 
    94.9697, 21.47264, 47.76735, 13.35156, 8.629306, 32.41949, 2.232151, 0, 
    0, 0, 1.06906, 0, 0, 0, 0, 12.63473, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    220.6236, 1349.775, 2132.709, 2395.235, 2048.53, 1480.806, 855.7775, 
    314.9611, 477.5641, 130.0667, 3.648897, 0, 0, 0, 0, 0, 0, 10.08162, 
    642.4855, 281.7012, 101.1102, 60.59174, 61.11189, 54.33709, 36.61767, 
    64.51082, 191.8937, 50.27359, 0.1158935, 0.7644691, 0, 0, 0, 0, 0, 0, 0, 
    127.1192, 404.733, 737.6123, 874.3842, 641.8504, 235.5844, 192.8914, 
    214.4153, 206.9348, 198.1494, 125.9625, 26.56938, 2.941694, 5.601278, 0, 
    0, 0, 0, 0, 0, 0, 0, 4.25005, 1.223589, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    123.0767, 1440.606, 2345.219, 2595.379, 2201.878, 1579.878, 765.6243, 
    263.2791, 17.18813, 95.84882, 0, 0, 0, 0, 0, 0, 0, 18.90151, 14.24182, 
    240.224, 244.171, 170.7711, 72.88946, 36.88171, 3.688538, 30.90802, 
    42.64079, 82.76118, 41.20324, 110.692, 64.07503, 0, 0, 0, 0, 0, 0, 
    116.6442, 851.2905, 1040.522, 1011.616, 761.973, 391.5457, 285.8691, 
    222.6031, 231.2289, 132.9321, 127.5657, 79.20253, 79.93398, 60.85431, 
    7.069205, 0, 0, 0, 0, 0, 0, 0.002840273, 31.90177, 12.23519, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    113.4006, 1133.138, 2195.308, 2608.468, 2239.793, 1572.94, 1003.211, 
    518.9925, 189.4889, 0.6126093, 0, 0, 0, 0, 0, 0, 0.1651795, 133.9569, 
    417.8274, 384.9297, 215.625, 141.7358, 90.05803, 79.19399, 29.33371, 
    2.240706, 12.30619, 0.2534847, 0, 94.7438, 162.481, 149.9046, 37.89026, 
    0, 0, 0, 0, 5.356696, 552.9598, 964.9863, 891.923, 640.1644, 439.5914, 
    361.2435, 278.5941, 283.0451, 244.8269, 280.0539, 219.772, 241.4119, 
    332.4167, 319.8716, 147.7597, 7.835948, 0, 0, 0, 0, 0.3774112, 84.49905, 
    37.25802, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 30.39107, 
    914.6385, 1832.73, 2461.096, 2238.884, 1490.557, 718.7988, 432.395, 
    372.0842, 0.9015442, 0, 0, 0, 0, 0, 105.8306, 357.3896, 523.8076, 
    521.7178, 440.9008, 328.9724, 202.1082, 166.6164, 82.55063, 126.2423, 
    70.6189, 12.28226, 42.67114, 60.72597, 91.16128, 142.8304, 148.7395, 
    152.2123, 97.86357, 0, 0.3341298, 0.6432131, 4.719822, 37.05452, 468.78, 
    599.9188, 399.7013, 211.5083, 353.3973, 316.7687, 280.8083, 341.3538, 
    511.3751, 442.6859, 504.624, 253.1497, 250.1017, 213.2764, 67.04365, 
    3.304585, 0, 0, 0.1683532, 53.87643, 48.47186, 10.75609, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 89.8662, 
    469.3024, 1154.713, 1449.781, 1272.478, 681.3491, 128.84, 4.544834, 0, 0, 
    0, 0, 0, 5.419511, 61.07015, 489.1122, 578.3217, 527.3911, 395.0327, 
    218.0269, 167.6713, 137.974, 115.5373, 0.6435879, 88.33016, 45.21404, 
    6.509036, 44.30594, 115.2863, 242.208, 245.5465, 151.2771, 0.4254271, 
    11.1162, 1.786039, 48.14689, 37.55202, 70.14665, 156.7791, 498.9786, 
    523.2408, 473.1295, 354.968, 545.134, 489.5596, 703.8699, 925.6036, 
    986.3214, 886.7418, 869.757, 604.8533, 197.4831, 113.1076, 12.6825, 0, 
    0.02486209, 6.962315, 96.1065, 54.04581, 0.01545697, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.1216824, 0.9288862, 134.0087, 201.5549, 60.90172, 0.3555474, 0, 0, 0, 
    0, 0, 355.5598, 602.0829, 651.0312, 450.9958, 386.381, 256.653, 158.6886, 
    43.34907, 61.85168, 159.5036, 113.3953, 25.31179, 87.31884, 165.2257, 
    4.966446, 0.1061549, 45.43877, 108.6841, 188.0823, 174.495, 113.4314, 
    0.01686891, 145.4191, 132.487, 172.8789, 193.6581, 150.9564, 166.1918, 
    400.6677, 583.3967, 722.2389, 745.6167, 800.6808, 849.4872, 1009.411, 
    1053.753, 947.8483, 415.5219, 584.1187, 491.2827, 259.1023, 215.041, 
    112.3413, 76.86075, 134.8813, 221.4578, 45.61331, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 3.875198, 477.9095, 533.1882, 461.8639, 235.7978, 
    111.7738, 22.34331, 6.797899, 1.574463, 51.39446, 134.1712, 4.203103, 
    6.980784, 108.1984, 118.4102, 3.881124, 11.86376, 72.39351, 102.465, 
    159.5778, 156.6727, 107.9339, 109.4576, 488.6499, 418.6319, 300.2693, 
    237.9754, 185.1014, 104.7926, 403.3925, 659.502, 1010.157, 881.0416, 
    936.1367, 774.4136, 1186.745, 1002.815, 1015.139, 535.5046, 386.2178, 
    179.3871, 69.36623, 267.0681, 111.3501, 67.82533, 6.994944, 1.526611, 
    3.172025, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 5.725166, 102.8057, 111.4602, 125.5778, 65.69091, 
    11.31183, 6.297175, 5.844241, 2.358717, 171.9062, 167.7866, 43.11033, 
    79.99084, 74.58493, 27.5016, 14.16823, 6.523846, 31.63298, 63.06898, 
    67.15324, 85.22324, 67.61577, 224.0022, 476.0859, 396.943, 309.3507, 
    246.142, 132.8316, 335.7784, 784.7097, 1053.235, 1127.867, 967.6097, 
    771.317, 924.9985, 1333.487, 1034.066, 789.8601, 234.963, 249.6979, 
    81.2932, 14.26598, 163.186, 164.9658, 5.164979, 1.026154, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.19746, 170.4447, 463.7712, 416.7452, 239.2617, 
    79.01589, 6.674962, 0, 0, 49.56345, 226.9828, 192.8199, 164.6065, 
    182.8128, 118.2701, 17.30331, 8.986745, 3.3333, 23.55511, 61.35153, 
    53.04255, 132.2586, 229.133, 315.2996, 329.1717, 262.2387, 250.0072, 
    217.4491, 311.0166, 854.7855, 1325.855, 1237.892, 1063.641, 815.3153, 
    855.515, 1043.939, 1759.73, 1143.116, 371.2457, 14.33288, 2.286062, 0, 0, 
    0.1220521, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 13.13908, 199.9922, 369.35, 332.041, 183.8263, 
    84.41653, 28.31347, 5.11356, 0, 3.346521, 94.1303, 145.3444, 260.3771, 
    308.1046, 216.5467, 65.93798, 66.89045, 91.82342, 129.8517, 169.2161, 
    212.0327, 380.3462, 430.9281, 398.8634, 271.8267, 213.1764, 198.3177, 
    260.7658, 507.0705, 1261.594, 1556.329, 1201.677, 977.4053, 903.3651, 
    1023.128, 1437.7, 2083.172, 1221.35, 86.26831, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 1.492808, 28.12763, 241.1122, 312.6933, 227.4316, 
    40.73929, 3.901017, 60.77868, 29.63254, 0, 37.46666, 47.92201, 90.67201, 
    252.6916, 297.8447, 250.6762, 146.2321, 137.6703, 164.451, 210.1363, 
    267.7924, 336.6427, 471.1196, 486.8597, 425.3645, 315.1228, 279.0462, 
    273.7747, 290.0505, 636.9206, 1410.759, 1544.152, 1250.766, 1127.925, 
    1065.812, 1110.734, 1416.591, 1600.496, 408.8422, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 8.41072, 11.77269, 0, 0, 1.62508, 8.022939, 6.219764, 0, 
    20.28673, 0.6057806, 40.99087, 150.5031, 84.34249, 84.26646, 195.8636, 
    227.4629, 190.5297, 136.6387, 154.2375, 176.6017, 216.4878, 304.6136, 
    374.8836, 462.7287, 472.5354, 402.6108, 307.9417, 327.0253, 306.5867, 
    373.0538, 668.3615, 1415.796, 1557.029, 1306.125, 1279.073, 1162.341, 
    1153.206, 1149.406, 1078.977, 41.16324, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 4.901734, 217.5294, 284.0266, 9.755486, 12.21576, 30.38478, 
    126.8581, 295.4576, 261.4576, 148.2994, 19.41799, 0.001383794, 4.122153, 
    25.35506, 13.69719, 14.41783, 64.17224, 71.70509, 82.17438, 88.62575, 
    143.002, 168.497, 227.1901, 295.2106, 377.9786, 424.9349, 434.2556, 
    359.2029, 243.9208, 256.3825, 320.5891, 276.9689, 544.5539, 1255.969, 
    1424.041, 1287.706, 1179.742, 1196.443, 1053.201, 1167.506, 829.4473, 
    18.81178, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.3367717, 55.36858, 332.4312, 482.9248, 279.4982, 0, 4.759403, 138.2639, 
    246.2088, 336.8652, 256.5343, 116.4693, 7.490035, 1.586183, 5.608893, 
    0.125523, 0.02205558, 0, 18.84512, 43.35651, 73.8119, 134.7575, 190.767, 
    245.426, 262.851, 321.6095, 350.954, 368.8531, 361.5361, 275.9557, 
    193.2714, 264.4291, 287.2755, 295.1925, 454.3226, 894.5059, 1154.717, 
    973.0314, 1099.105, 1148.796, 1120.024, 862.0306, 375.9889, 12.88452, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.2140546, 
    0.1701733, 26.3982, 16.54789, 11.51096, 64.69183, 320.2927, 487.4863, 
    486.2169, 178.1183, 52.80968, 111.4205, 188.5571, 226.6747, 194.1454, 
    121.9309, 19.68636, 0, 0, 0, 0, 0, 0, 0.08443239, 12.21449, 77.40128, 
    139.2317, 232.2935, 274.8673, 306.887, 328.7855, 366.2649, 352.3075, 
    297.598, 212.2141, 162.9654, 161.8156, 294.4319, 331.9783, 424.2078, 
    668.4012, 775.5222, 991.9241, 1072.528, 1282.538, 1139.612, 931.2537, 
    216.4193, 62.45685, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3.731169, 
    99.69241, 145.8221, 164.5461, 190.2277, 222.6298, 352.1655, 453.9755, 
    483.7257, 366.7473, 201.0961, 195.8921, 224.278, 247.8174, 199.336, 
    145.5127, 58.51702, 0.01620398, 1.724691, 0, 0, 0, 0, 0, 0, 3.441099, 
    66.59528, 167.6643, 266.4513, 312.1495, 332.5176, 373.2896, 422.7214, 
    417.7817, 331.4211, 227.7531, 191.2091, 276.8271, 346.7453, 491.9813, 
    515.8571, 477.7105, 837.2191, 1215.665, 1373.787, 1364.735, 1284.096, 
    957.2903, 218.0976, 83.97918, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7.299129, 134.0267, 
    294.2319, 344.9782, 270.6827, 318.7709, 384.5544, 494.1917, 494.657, 
    473.3284, 365.3275, 308.8357, 293.0063, 310.0292, 272.0663, 223.5598, 
    135.7657, 49.15474, 0.05388123, 0.2981069, 0, 0, 0, 0, 0, 0, 0.2216611, 
    69.87698, 190.6432, 286.7062, 330.1897, 367.8758, 406.1044, 450.1877, 
    427.9415, 330.3656, 250.8139, 289.5048, 447.8335, 462.0058, 478.6495, 
    494.2013, 530.5643, 958.8607, 1535.851, 1566.941, 1493.999, 1267.836, 
    1004.899, 187.0762, 37.84942, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.2778322, 1.216981, 0.320554, 
    82.15788, 124.0773, 328.814, 414.2038, 370.9027, 408.5572, 474.0244, 
    515.583, 504.9358, 517.7888, 478.3085, 405.8519, 390.0446, 340.6481, 
    284.1749, 193.1102, 63.77376, 0.2711483, 0.001171568, 0, 0, 0, 0, 0, 0, 
    0, 0.01659026, 97.79198, 225.3099, 301.7682, 358.1664, 393.5924, 
    409.4816, 387.7672, 372.0033, 279.7969, 234.8109, 369.993, 486.2102, 
    487.3097, 453.6224, 565.4487, 638.8194, 1025.565, 1495.267, 1465.116, 
    1353.271, 1132.2, 829.127, 232.6918, 86.18745, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.03872748, 20.11839, 53.78059, 
    33.44499, 88.68514, 177.8256, 19.69762, 253.2851, 404.7767, 437.9373, 
    469.3643, 499.6412, 501.7674, 551.6224, 574.769, 536.6869, 488.521, 
    416.7465, 350.7989, 264.6436, 127.1555, 0.415809, 0.4254224, 0, 0, 0, 0, 
    0, 0, 0, 0.6914847, 19.04652, 131.946, 247.1787, 306.9858, 363.0714, 
    397.9942, 400.0674, 409.7594, 398.0919, 355.8009, 291.4016, 333.1392, 
    498.2859, 440.002, 539.7181, 723.6176, 765.5291, 965.6453, 1312.768, 
    1339.947, 1188.61, 996.9376, 753.3426, 184.1582, 17.82256, 30.13374, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.789168, 70.13921, 107.3934, 180.0283, 
    234.5805, 241.1893, 107.9595, 15.09211, 188.5137, 368.2224, 514.8614, 
    566.2856, 554.1669, 566.897, 608.2187, 604.4344, 543.1758, 479.5136, 
    420.2968, 358.7137, 272.7408, 113.1928, 4.518106, 5.010964, 0, 0, 0, 0, 
    0, 0, 0.7098004, 13.29282, 97.01318, 193.7101, 286.6924, 317.051, 
    366.6038, 397.0652, 432.3381, 481.5545, 519.4891, 467.0329, 436.6177, 
    526.4904, 556.9227, 596.2275, 609.3391, 692.4142, 720.394, 862.9467, 
    1120.028, 1117.907, 1092.196, 985.4866, 917.553, 349.6905, 24.9056, 
    102.5677, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18.45255, 45.57545, 90.12004, 208.861, 
    326.2532, 247.4885, 3.031927, 0.8162752, 62.72859, 240.1284, 478.4014, 
    642.7585, 624.4623, 612.9011, 633.5761, 635.511, 540.0829, 464.6622, 
    389.1842, 327.2373, 250.5822, 128.0566, 4.151914, 0.01724564, 0, 0, 0, 
    0.06221788, 16.14303, 56.51927, 60.10637, 63.71621, 129.8515, 214.7995, 
    265.7689, 302.5134, 336.1973, 365.2288, 442.3849, 504.6011, 502.0141, 
    480.3363, 467.8888, 553.1976, 593.0986, 637.1354, 629.6438, 659.4634, 
    735.4026, 1028.44, 1056.044, 946.681, 926.314, 1064.744, 949.1011, 
    392.1784, 18.68724, 70.3578, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18.13205, 81.59405, 283.5952, 
    99.12554, 0, 2.600603, 22.27865, 40.11892, 259.8885, 493.662, 624.6654, 
    578.1021, 631.7147, 627.2502, 560.2089, 436.4544, 359.2498, 263.4945, 
    198.2276, 96.85187, 8.224985, 0.006419148, 10.41262, 28.47488, 33.42284, 
    63.55798, 89.37606, 117.4287, 123.5775, 113.715, 153.6499, 198.5007, 
    238.3534, 277.4305, 321.2411, 352.9605, 414.103, 455.9593, 452.3423, 
    458.7655, 565.2747, 608.5494, 639.5411, 687.265, 764.0191, 736.5245, 
    987.5319, 1266.858, 1113.241, 848.986, 966.5779, 1123.773, 1059.529, 
    375.9788, 5.606318, 11.23915, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 50.03308, 18.7767, 0, 
    1.26797, 38.3414, 37.16248, 6.458248, 236.8902, 463.1305, 562.8348, 
    578.8032, 630.9438, 520.6262, 426.2543, 325.3188, 244.9647, 138.4487, 
    36.07342, 0.5078325, 2.94648, 57.33051, 95.80891, 105.8, 111.6879, 
    121.1859, 142.7138, 152.8308, 160.8624, 182.531, 201.2338, 222.661, 
    264.4805, 303.7233, 333.4624, 371.3336, 438.1491, 455.2211, 496.9004, 
    597.2755, 643.8214, 617.1034, 691.8447, 823.0101, 988.5286, 1358.407, 
    1648.078, 1373.022, 979.8769, 1118.349, 1293.235, 1281.518, 524.8214, 
    12.07863, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18.53168, 7.44618, 
    0.2774768, 0, 35.85915, 285.9109, 179.5872, 150.5524, 421.4404, 514.148, 
    569.3135, 533.7565, 453.5545, 348.8341, 297.6014, 196.2376, 72.14723, 
    1.141348, 3.445107, 14.83014, 68.87897, 118.991, 129.5745, 158.0152, 
    182.8073, 209.6761, 221.1556, 222.757, 222.7252, 225.1968, 215.3978, 
    252.5812, 274.6012, 313.8231, 378.8444, 483.5266, 526.6315, 559.9622, 
    581.9632, 617.732, 638.4788, 691.2427, 829.9338, 1126.817, 1687.072, 
    1798.549, 1466.908, 1100.552, 1091.336, 1508.885, 1401.512, 703.5411, 
    81.51077, 0.2449444, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15.97898, 137.8128, 2.629696, 
    0.1815157, 0, 28.15523, 299.744, 311.1771, 79.97313, 377.6644, 488.9033, 
    461.6871, 486.7418, 409.492, 350.8954, 279.0941, 180.3749, 25.7736, 
    3.397881, 18.72686, 43.95182, 103.1606, 144.6976, 190.1044, 222.457, 
    259.2217, 285.7209, 287.2361, 281.1645, 272.6286, 249.3425, 225.9028, 
    238.7993, 272.0008, 332.6962, 384.1511, 468.3911, 546.1947, 577.4488, 
    627.5869, 635.5259, 700.1279, 776.9152, 929.8552, 1510.917, 1895.887, 
    1799.537, 1355.943, 1119.573, 1392.253, 1618.039, 1311.142, 575.1276, 
    257.3511, 0.8315546, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8.894205, 72.59029, 14.85453, 
    7.508962, 13.51235, 142.9096, 296.0406, 327.9227, 156.2393, 437.1971, 
    388.5025, 385.3842, 401.033, 394.5582, 335.838, 280.1766, 193.5683, 
    96.386, 35.52516, 58.84515, 86.79417, 122.0659, 181.4595, 237.5804, 
    289.2039, 326.9966, 354.348, 356.1935, 336.6149, 307.5397, 253.4356, 
    225.7552, 236.1096, 334.7573, 444.7771, 494.1808, 514.2294, 524.8425, 
    587.1181, 631.0831, 694.0496, 751.4611, 825.4266, 1097.83, 1658.775, 
    2006.745, 1602.702, 1223.444, 1127.629, 1333.478, 1458.12, 871.0525, 
    466.6771, 267.9041, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01038057, 0, 6.643703, 101.4879, 
    82.98901, 51.23274, 85.14922, 210.2779, 283.6747, 309.324, 233.2301, 
    492.1425, 371.6667, 362.65, 444.5501, 397.6977, 330.4786, 280.92, 
    273.9966, 219.3448, 153.7401, 126.073, 117.5657, 150.8828, 219.6838, 
    283.4588, 333.4008, 374.8239, 400.1253, 395.6437, 375.5026, 312.2456, 
    243.2001, 227.2077, 279.3844, 409.5839, 514.515, 561.0614, 561.6627, 
    541.6973, 592.7158, 646.3815, 705.6855, 755.9585, 820.3306, 1077.465, 
    1725.695, 1795.541, 1577.446, 1249.411, 1148.976, 1319.127, 995.0981, 
    382.848, 349.3625, 65.2517, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 49.50258, 104.9451, 82.473, 
    92.12851, 176.1149, 268.6027, 316.0862, 341.2645, 486.9077, 443.9214, 
    441.7123, 453.1961, 411.6028, 339.4975, 305.282, 294.3625, 287.3364, 
    230.1652, 207.584, 207.6316, 229.0633, 299.8941, 320.3898, 366.2971, 
    403.0446, 399.9144, 400.9593, 372.4525, 306.9135, 239.632, 240.6821, 
    343.6025, 474.4823, 553.2586, 592.0007, 575.3657, 602.5383, 624.6992, 
    700.6254, 727.1317, 764.283, 781.6901, 1065.684, 1631.907, 1692.728, 
    1571.499, 1298.507, 1313.886, 1286.554, 934.9397, 106.3758, 289.6695, 
    15.00103, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11.55675, 115.867, 
    22.48811, 65.3556, 149.1486, 286.7424, 407.3988, 236.5376, 274.9689, 
    357.7444, 443.3862, 421.6057, 401.2734, 343.1813, 298.683, 307.432, 
    300.7722, 291.2484, 308.8382, 334.8492, 323.8983, 337.6805, 341.7525, 
    399.8321, 429.9846, 410.5637, 382.6377, 354.2699, 306.8083, 234.6121, 
    282.1734, 378.2628, 513.45, 570.4268, 609.7987, 630.7244, 657.3438, 
    763.2346, 822.8828, 897.2252, 876.2137, 902.7307, 1085.887, 1506.075, 
    1453.561, 1306.629, 1103.886, 1026.492, 1225.022, 985.5616, 402.682, 
    411.0314, 92.16769, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8.036347, 62.52849, 
    3.547037, 32.43497, 104.1824, 329.8143, 462.2404, 251.2797, 109.8259, 
    300.0777, 382.1133, 340.6129, 357.1865, 326.0741, 305.6071, 339.9389, 
    372.1312, 391.5172, 407.5522, 352.1345, 293.8417, 268.1846, 292.7089, 
    444.7627, 466.584, 417.2143, 374.3411, 349.6299, 313.55, 266.888, 
    336.9229, 432.6651, 484.9139, 546.2026, 630.8204, 650.4514, 755.9393, 
    824.0303, 861.4523, 911.7997, 958.1385, 976.4166, 1254.706, 1563.365, 
    1293.88, 1170.993, 864.0294, 700.7004, 757.6398, 917.2304, 682.3601, 
    402.354, 43.28111, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.05915249, 0.08011421, 0, 
    6.02283, 76.62966, 347.7174, 469.9626, 235.3439, 100.1177, 160.2919, 
    227.011, 263.368, 336.6925, 322.0186, 290.6877, 363.0302, 432.0052, 
    448.0348, 357.6713, 268.9411, 179.2584, 179, 233.9073, 359.2671, 
    464.7566, 411.7307, 372.834, 358.2526, 326.1168, 293.7316, 402.5888, 
    470.521, 497.5835, 578.8224, 635.5013, 674.5109, 734.5461, 763.5286, 
    810.0879, 885.3263, 939.2901, 1104.282, 1317.147, 1582.151, 1373.822, 
    1213.066, 873.9077, 635.079, 382.4486, 656.3605, 884.5526, 664.905, 
    217.4573, 32.62277, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.014362, 
    61.41228, 327.5756, 417.7493, 328.8751, 249.4016, 131.7789, 157.5266, 
    287.179, 367.0403, 311.7421, 237.5124, 263.4082, 315.4411, 318.5938, 
    269.0101, 179.5965, 192.4013, 228.7823, 193.9452, 278.2494, 363.2266, 
    430.6738, 408.0237, 404.8087, 350.7692, 302.6519, 419.8691, 508.0556, 
    530.116, 605.4689, 677.9661, 698.0052, 724.3315, 784.8451, 801.787, 
    928.4433, 1166.382, 1351.242, 1463.7, 1691.588, 1541.213, 1399.71, 
    1026.168, 717.6241, 512.4301, 377.8375, 697.6708, 594.645, 397.4904, 
    142.8448, 0.532489, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.2053152, 
    67.53915, 303.6299, 379.2345, 436.3914, 423.1708, 180.6438, 155.2336, 
    276.7622, 326.9408, 266.7624, 175.7495, 176.1388, 195.9187, 226.1668, 
    186.327, 215.0712, 291.8131, 416.8516, 394.0894, 300.8634, 340.7516, 
    360.322, 408.5583, 425.7607, 360.9985, 326.2549, 435.8652, 544.7354, 
    572.8199, 653.0318, 746.2729, 793.1929, 824.189, 828.2086, 914.1102, 
    1028.284, 1346.432, 1671.313, 1678.606, 1814.529, 1881.197, 1709.896, 
    1406.109, 1219.147, 1059.282, 948.7432, 834.345, 919.3475, 724.296, 
    356.6761, 76.5276, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.8787696, 13.35174, 
    137.5124, 287.6332, 345.7241, 417.4199, 379.3897, 131.3522, 106.2649, 
    169.0464, 272.2558, 288.1475, 201.0602, 176.5896, 223.6827, 266.1863, 
    218.2081, 176.9505, 269.0522, 436.2097, 486.094, 402.9827, 347.54, 
    334.3905, 365.894, 393.4282, 347.4721, 379.8949, 443.5723, 566.2279, 
    602.1741, 676.5858, 812.3363, 900.5889, 908.915, 931.9954, 944.5102, 
    1117.414, 1304.28, 1882.296, 1832.433, 1976.871, 2069.233, 2070.061, 
    1899.477, 1551.457, 1340.278, 1386.592, 1314.673, 1244.868, 1230.34, 
    806.1844, 287.225, 40.42369, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2.817714, 35.69061, 
    138.5443, 281.9023, 361.2498, 453.4521, 359.1906, 222.1722, 156.6933, 
    136.975, 236.7071, 325.3279, 228.1469, 196.3775, 242.6227, 329.216, 
    249.9151, 180.1256, 229.7955, 351.343, 390.6742, 362.7199, 313.2054, 
    299.3227, 315.3665, 337.3273, 403.3815, 440.4469, 459.0341, 544.0665, 
    574.6163, 685.2004, 805.9506, 978.1014, 1079.502, 1060.385, 1335.979, 
    1386.026, 1736.179, 2369.993, 2377.097, 2108.683, 2192.729, 2248.685, 
    2160.981, 1428.064, 1097.215, 1308.715, 1435.482, 1437.344, 1562.363, 
    1290.539, 805.3401, 441.8997, 16.92101, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;
}
