netcdf \00010101.atmos_daily.hfls.tile3 {
dimensions:
	time = UNLIMITED ; // (182 currently)
	phalf = 66 ;
	grid_xt = 15 ;
	grid_yt = 10 ;
	scalar_axis = 1 ;
	nv = 2 ;
	pfull = 65 ;
variables:
	double average_DT(time) ;
		average_DT:_FillValue = 1.e+20 ;
		average_DT:missing_value = 1.e+20 ;
		average_DT:units = "days" ;
		average_DT:long_name = "Length of average period" ;
	double average_T1(time) ;
		average_T1:_FillValue = 1.e+20 ;
		average_T1:missing_value = 1.e+20 ;
		average_T1:units = "days since 0001-01-01 00:00:00" ;
		average_T1:long_name = "Start time for average period" ;
	double average_T2(time) ;
		average_T2:_FillValue = 1.e+20 ;
		average_T2:missing_value = 1.e+20 ;
		average_T2:units = "days since 0001-01-01 00:00:00" ;
		average_T2:long_name = "End time for average period" ;
	float bk(phalf) ;
		bk:_FillValue = 1.e+20f ;
		bk:missing_value = 1.e+20f ;
		bk:long_name = "vertical coordinate sigma value" ;
		bk:cell_methods = "time: point" ;
	double grid_xt(grid_xt) ;
		grid_xt:units = "degrees_E" ;
		grid_xt:long_name = "T-cell longitude" ;
		grid_xt:axis = "X" ;
	double grid_yt(grid_yt) ;
		grid_yt:units = "degrees_N" ;
		grid_yt:long_name = "T-cell latitude" ;
		grid_yt:axis = "Y" ;
	float height10m(scalar_axis) ;
		height10m:_FillValue = 1.e+20f ;
		height10m:missing_value = 1.e+20f ;
		height10m:units = "m" ;
		height10m:long_name = "Height" ;
		height10m:cell_methods = "time: point" ;
		height10m:axis = "Z" ;
		height10m:positive = "up" ;
		height10m:standard_name = "height" ;
	float height2m(scalar_axis) ;
		height2m:_FillValue = 1.e+20f ;
		height2m:missing_value = 1.e+20f ;
		height2m:units = "m" ;
		height2m:long_name = "Height" ;
		height2m:cell_methods = "time: point" ;
		height2m:axis = "Z" ;
		height2m:positive = "up" ;
		height2m:standard_name = "height" ;
	float hfls(time, grid_yt, grid_xt) ;
		hfls:_FillValue = 1.e+20f ;
		hfls:missing_value = 1.e+20f ;
		hfls:units = "W m-2" ;
		hfls:long_name = "Surface Upward Latent Heat Flux" ;
		hfls:cell_methods = "time: mean" ;
		hfls:cell_measures = "area: area" ;
		hfls:comment = "Lv*evap" ;
		hfls:time_avg_info = "average_T1,average_T2,average_DT" ;
		hfls:standard_name = "surface_upward_latent_heat_flux" ;
	double nv(nv) ;
		nv:long_name = "vertex number" ;
	double pfull(pfull) ;
		pfull:units = "mb" ;
		pfull:long_name = "ref full pressure level" ;
		pfull:axis = "Z" ;
		pfull:positive = "down" ;
	double phalf(phalf) ;
		phalf:units = "mb" ;
		phalf:long_name = "ref half pressure level" ;
		phalf:axis = "Z" ;
		phalf:positive = "down" ;
	float pk(phalf) ;
		pk:_FillValue = 1.e+20f ;
		pk:missing_value = 1.e+20f ;
		pk:units = "pascal" ;
		pk:long_name = "pressure part of the hybrid coordinate" ;
		pk:cell_methods = "time: point" ;
	double scalar_axis(scalar_axis) ;
		scalar_axis:long_name = "none" ;
	double time(time) ;
		time:units = "days since 0001-01-01 00:00:00" ;
		time:long_name = "time" ;
		time:axis = "T" ;
		time:calendar_type = "NOLEAP" ;
		time:calendar = "noleap" ;
		time:bounds = "time_bnds" ;
	double time_bnds(time, nv) ;
		time_bnds:long_name = "time axis boundaries" ;

// global attributes:
		:title = "cm5_c96_am5f7c1r0_b06_piC_galb_noiceinit_alb" ;
		:associated_files = "area: 00010101.grid_spec.nc" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
		:history = "Wed Apr 30 14:48:00 2025: ncks -d grid_xt,0,14 -d grid_yt,0,9 -d time,0,181 /home/cew/Code/cmip7-sprint/testfiles/input/00010101.atmos_daily.tile3.nc -O /home/cew/Code/cmip7-sprint/testfiles/00010101.atmos_daily.tile3.nc\nFri Apr 25 14:15:06 2025: ncks -x -v sphum,psl 00010101.atmos_daily.tile3.nc -o reduce/00010101.atmos_daily.tile3.nc\nFri Apr 25 13:47:12 2025: ncks -d grid_xt,35,55 -d grid_yt,30,45 00010101.atmos_daily.tile3.nc var_select/00010101.atmos_daily.tile3.nc" ;
		:NCO = "netCDF Operators version 5.1.9 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco, Citation = 10.1016/j.envsoft.2008.03.004)" ;
data:

 average_DT = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 average_T1 = 0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 
    18, 19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 
    36, 37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 
    54, 55, 56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 
    72, 73, 74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 
    90, 91, 92, 93, 94, 95, 96, 97, 98, 99, 100, 101, 102, 103, 104, 105, 
    106, 107, 108, 109, 110, 111, 112, 113, 114, 115, 116, 117, 118, 119, 
    120, 121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 
    134, 135, 136, 137, 138, 139, 140, 141, 142, 143, 144, 145, 146, 147, 
    148, 149, 150, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 
    162, 163, 164, 165, 166, 167, 168, 169, 170, 171, 172, 173, 174, 175, 
    176, 177, 178, 179, 180, 181 ;

 average_T2 = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 
    19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 
    37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 54, 
    55, 56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 72, 
    73, 74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 90, 
    91, 92, 93, 94, 95, 96, 97, 98, 99, 100, 101, 102, 103, 104, 105, 106, 
    107, 108, 109, 110, 111, 112, 113, 114, 115, 116, 117, 118, 119, 120, 
    121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 134, 
    135, 136, 137, 138, 139, 140, 141, 142, 143, 144, 145, 146, 147, 148, 
    149, 150, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 162, 
    163, 164, 165, 166, 167, 168, 169, 170, 171, 172, 173, 174, 175, 176, 
    177, 178, 179, 180, 181, 182 ;

 bk = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.00193294, 0.00749994, 0.01640714, 0.02841953, 
    0.04334756, 0.06103661, 0.0813586, 0.1042054, 0.1294836, 0.1571101, 
    0.1870091, 0.2191095, 0.2533426, 0.2896406, 0.3279357, 0.3681587, 
    0.4102391, 0.454293, 0.5001689, 0.5468886, 0.5935643, 0.6397641, 
    0.6851825, 0.729505, 0.7723162, 0.8125153, 0.8492141, 0.8817441, 
    0.909788, 0.9332725, 0.9524949, 0.9678352, 0.9798011, 0.9889621, 0.99575, 1 ;

 grid_xt = 36, 37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50 ;

 grid_yt = 31, 32, 33, 34, 35, 36, 37, 38, 39, 40 ;

 height10m = 10 ;

 height2m = 2 ;

 hfls =
  29.90368, 49.35181, 49.9096, 95.12691, 71.87212, 35.03489, 47.63442, 
    50.20385, 53.5752, 11.16579, 14.51125, 27.03942, 11.70793, 14.27759, 
    -0.3786513,
  85.97427, 75.98698, 57.91388, 77.04918, 35.42171, 26.09041, 44.20863, 
    40.81323, 50.58518, 40.09371, 21.50808, 49.16239, 49.14007, 5.695109, 
    -0.3838496,
  77.86563, 86.58753, 82.07342, 79.01974, 63.59566, 5.253563, 42.06587, 
    43.8668, 50.82354, 48.50815, 47.83553, 52.98396, 56.59428, 50.79833, 
    23.60787,
  90.28301, 79.84243, 84.45894, 86.84377, 96.03311, 70.30258, 5.590069, 
    37.44505, 66.14964, 48.09973, 42.62407, 47.77813, 53.16575, 54.2935, 
    40.27913,
  108.1024, 96.88148, 87.83829, 87.85508, 89.05102, 96.91717, 82.45899, 
    7.665728, 23.434, 30.05699, 38.93267, 44.75055, 51.67457, 57.85662, 
    60.49834,
  111.5299, 111.7298, 101.9088, 96.64767, 93.89856, 92.98494, 86.36525, 
    85.89212, 63.87637, 54.17691, 35.88317, 47.81981, 51.35664, 57.47815, 
    59.41167,
  142.48, 126.0268, 119.2533, 111.6749, 106.4043, 106.0936, 105.7216, 
    104.1531, 96.93313, 94.34602, 76.10916, 52.9972, 54.02652, 56.78365, 
    56.2613,
  160.5278, 143.6519, 129.296, 121.3241, 115.8553, 113.2635, 111.5116, 
    110.4745, 105.2159, 105.8064, 92.3639, 59.81791, 54.64816, 56.76723, 
    56.20507,
  150.6531, 140.6597, 129.5796, 121.8886, 115.4403, 112.5857, 109.8309, 
    111.2056, 112.5377, 108.7657, 99.57213, 64.77615, 57.7329, 57.47926, 
    52.13752,
  130.8871, 124.7921, 120.3337, 114.0291, 108.5477, 105.3859, 107.403, 
    107.7126, 95.67406, 57.05529, 68.44485, 65.23853, 54.89882, 53.54874, 
    48.85418,
  19.94387, 68.18848, 35.11386, 77.19118, 53.91861, 27.53799, 39.91742, 
    39.15331, 30.5566, 8.709927, 6.694763, 16.43366, 8.347309, 7.020243, 
    -1.035404,
  94.01846, 63.43055, 68.16828, 77.42448, 37.32515, 15.14052, 46.80177, 
    45.37751, 38.44511, 26.12229, 12.31758, 26.77488, 30.09464, 3.41725, 
    -1.226893,
  136.9446, 119.7449, 95.17655, 95.66568, 65.04585, 2.645418, 37.6474, 
    49.59634, 51.96608, 34.23428, 30.95558, 31.09142, 29.64791, 30.73212, 
    12.87078,
  145.8134, 144.2041, 137.166, 121.9089, 106.4885, 69.11348, 2.082128, 
    35.04427, 61.74097, 39.09015, 32.89597, 32.47304, 30.65792, 26.59863, 
    21.80292,
  140.8575, 139.7991, 135.6308, 130.8493, 119.6519, 108.6756, 80.07188, 
    4.914348, 10.67877, 20.84244, 32.31161, 32.82687, 32.6984, 30.39337, 
    29.32289,
  136.3033, 136.7004, 131.5711, 129.3912, 126.5813, 120.7381, 109.4274, 
    104.0917, 68.36091, 65.57024, 27.8831, 33.6718, 33.63538, 33.11654, 
    30.79506,
  134.0072, 133.4505, 128.346, 124.3258, 121.1189, 119.2733, 115.7979, 
    110.9834, 103.5854, 110.1534, 65.93564, 35.3195, 34.24898, 35.51768, 
    34.48705,
  132.0383, 130.3293, 126.3854, 122.4379, 116.0227, 110.2302, 104.9459, 
    103.797, 107.2649, 115.0891, 82.69083, 37.3639, 35.0563, 36.77258, 
    35.45859,
  121.8291, 121.4803, 118.6989, 116.8132, 114.5379, 112.4398, 110.5155, 
    110.9144, 113.3944, 110.972, 87.62427, 38.8427, 35.22116, 36.03963, 
    32.42701,
  104.0649, 105.2761, 106.6556, 105.4754, 104.2499, 106.519, 111.2164, 
    111.2786, 96.00427, 57.59768, 61.20727, 38.20073, 33.92863, 33.76033, 
    30.82523,
  29.49665, 79.39426, 36.22445, 66.26254, 38.2092, 15.41371, 24.21033, 
    24.48758, 14.63505, 2.524331, 4.54463, 10.4499, 3.422899, 3.775796, 
    -1.475031,
  99.55483, 107.1141, 100.3814, 83.37931, 22.29678, 7.595412, 29.30658, 
    26.37353, 16.6594, 17.80875, 8.695395, 17.84048, 24.64693, 0.227561, 
    -1.737749,
  103.4131, 108.9124, 111.5458, 104.6378, 61.59361, 2.802226, 23.29206, 
    25.85521, 24.45564, 25.46906, 22.63697, 21.23371, 20.75711, 31.25564, 
    7.687753,
  107.2414, 108.6677, 114.9735, 118.6814, 115.5807, 58.64091, 2.099117, 
    19.09479, 31.21553, 24.77027, 22.57123, 22.27404, 20.89271, 18.62674, 
    19.85809,
  112.411, 112.5591, 115.7835, 123.7976, 127.4977, 104.6736, 57.6132, 
    4.565296, 4.721332, 12.36031, 22.25357, 24.86841, 23.59048, 22.24597, 
    20.97233,
  117.1093, 118.8862, 118.9836, 123.8579, 130.4616, 120.5527, 96.96727, 
    89.75337, 58.5301, 62.34965, 23.91878, 25.80862, 24.56903, 23.34992, 
    20.58767,
  125.197, 127.1145, 125.566, 126.8255, 129.7521, 124.0255, 112.465, 
    107.3583, 105.8252, 115.1535, 53.1879, 29.93278, 25.48637, 25.08777, 
    24.93339,
  129.218, 132.7282, 132.9009, 133.1095, 130.4518, 125.4616, 119.5993, 
    120.1405, 120.1186, 124.772, 67.88586, 32.96475, 27.17938, 27.13265, 
    25.45874,
  124.2681, 129.776, 132.8704, 134.642, 131.5636, 124.6623, 120.7146, 
    124.0693, 126.605, 123.8061, 79.37349, 35.25262, 30.18461, 28.38721, 
    25.50344,
  112.2394, 118.5169, 125.1055, 128.377, 128.4959, 124.6787, 121.5553, 
    118.413, 105.4979, 67.91891, 61.62674, 35.53001, 34.50707, 30.05908, 
    29.44142,
  30.186, 69.28781, 31.06088, 58.54395, 15.96561, 4.620884, 14.55353, 
    13.90488, 12.6291, 2.516629, 0.08817343, 6.27221, 2.267228, 1.925579, 
    -0.5842738,
  76.43607, 74.09801, 64.90688, 53.85924, 11.82014, 4.326458, 13.74294, 
    17.06936, 17.14952, 13.72735, 3.454065, 11.49145, 17.80231, 0.1519339, 
    -0.6532018,
  73.31511, 61.42937, 62.24793, 60.46941, 32.29095, 1.437121, 10.94933, 
    19.07415, 24.72638, 20.27587, 16.40111, 12.39819, 12.49832, 17.63468, 
    5.994524,
  64.27818, 56.91526, 64.82674, 67.00723, 61.38698, 29.21724, -0.9560582, 
    8.484658, 19.52128, 17.59842, 13.38289, 12.58552, 12.94139, 11.7723, 
    12.58611,
  56.88434, 59.40531, 66.11562, 66.77129, 60.15685, 59.47005, 60.73809, 
    1.913983, 1.959728, 6.339938, 11.84248, 14.41221, 14.31263, 14.03899, 
    13.24203,
  59.13514, 65.76833, 68.94794, 63.59967, 53.0408, 62.47777, 101.1762, 
    104.3756, 59.04048, 63.25182, 21.98762, 16.94074, 14.82189, 13.24846, 
    13.05468,
  66.43985, 72.16913, 71.20568, 58.61789, 47.93162, 69.23689, 102.617, 
    114.6154, 122.7928, 131.7735, 53.16456, 20.55632, 16.28527, 14.81254, 
    16.99631,
  79.22583, 78.72034, 75.36917, 57.70323, 59.79492, 86.53474, 116.2762, 
    126.0243, 133.4176, 134.9903, 52.05973, 22.9968, 16.82232, 18.68106, 
    18.8256,
  86.39959, 84.33742, 76.67826, 65.11486, 76.66173, 101.989, 121.4774, 
    122.6847, 127.7903, 127.3481, 59.16478, 25.83772, 18.96892, 22.60896, 
    17.56969,
  82.10811, 79.4471, 74.3224, 79.92526, 90.79325, 106.555, 119.7112, 
    119.0771, 104.7615, 64.15684, 44.37476, 26.20104, 26.78516, 22.69279, 
    21.8245,
  36.72674, 81.28628, 42.7725, 62.04868, 12.70072, 3.76093, 16.40561, 
    14.87112, 15.64011, 5.036236, 0.4752112, 5.133053, 1.451237, 1.659036, 
    -0.07729162,
  88.24762, 90.31697, 76.54839, 58.91077, 5.428793, 8.784087, 20.42345, 
    17.18258, 14.91925, 14.53654, 3.636008, 9.195682, 13.24052, 1.155654, 
    -0.03052879,
  88.41698, 79.50895, 65.36109, 62.22869, 44.06359, 2.832501, 18.19785, 
    20.30075, 18.67632, 14.73027, 14.26157, 10.05181, 8.753593, 9.843642, 
    4.233417,
  92.827, 76.27119, 64.16093, 74.79767, 95.81362, 61.10793, 0.7413305, 
    12.99763, 15.36454, 12.65689, 10.6776, 8.94291, 7.449193, 6.694005, 
    7.335553,
  95.04328, 78.2803, 68.45449, 77.66142, 92.79767, 103.6608, 88.86219, 
    1.818138, -0.8169997, 2.180555, 8.341966, 9.496581, 7.581588, 6.61267, 
    6.959939,
  97.1233, 83.79354, 73.23766, 77.5854, 85.7849, 96.5926, 115.8155, 103.431, 
    46.08648, 45.8288, 16.7435, 11.03699, 8.031536, 6.566501, 7.002732,
  103.468, 93.03603, 79.83617, 78.98044, 81.47308, 89.50407, 104.6459, 
    106.0877, 107.396, 114.6892, 45.79217, 14.09298, 8.311985, 6.690997, 
    7.770307,
  113.2272, 100.9135, 83.53759, 78.87901, 81.04982, 91.24094, 110.6284, 
    117.9091, 122.1383, 116.7452, 36.88425, 15.36965, 8.722073, 7.851161, 
    7.529326,
  114.955, 104.7511, 86.78647, 78.46326, 79.75532, 96.0891, 117.7008, 
    117.1062, 117.1589, 111.1448, 41.56239, 15.84196, 9.023249, 9.529157, 
    9.556837,
  106.1012, 91.87922, 78.07041, 76.89349, 82.38218, 96.99767, 118.4921, 
    113.6096, 96.60474, 51.79499, 31.48509, 14.90121, 11.94797, 13.33376, 
    13.79647,
  38.42847, 86.24054, 50.74516, 77.28505, 25.98875, 11.07192, 17.71925, 
    16.68664, 14.39678, 3.697607, 0.7760437, 2.277699, 0.2863366, 1.192304, 
    -0.3061956,
  94.83387, 101.8266, 99.5528, 89.31242, 18.1683, 8.21797, 20.72439, 
    15.52581, 10.16745, 8.871483, 2.075456, 6.024156, 8.96297, 0.6530478, 
    -0.07454053,
  98.64342, 100.9419, 102.7324, 100.4351, 63.25273, 1.982138, 16.34619, 
    15.96945, 10.27515, 9.143429, 6.998737, 5.765967, 7.795322, 9.332646, 
    2.92713,
  106.617, 103.0239, 101.8157, 104.8686, 115.3563, 69.49582, 2.71488, 
    7.231191, 8.275229, 6.174344, 4.700841, 4.115173, 4.105628, 6.653508, 
    5.375134,
  113.7324, 106.4996, 100.6247, 98.5798, 109.3904, 115.075, 88.72878, 
    2.340438, -0.6090736, 0.931077, 3.71731, 4.049097, 3.372426, 5.169108, 
    6.129706,
  121.4625, 108.6822, 98.70801, 92.25932, 101.9606, 109.7147, 112.195, 
    94.00412, 35.01019, 30.77778, 9.600596, 4.315543, 3.819422, 6.572888, 
    7.634212,
  132.5433, 113.4959, 98.57487, 89.82738, 96.96941, 102.0061, 100.4616, 
    95.8113, 84.82072, 81.96284, 29.51884, 5.482117, 3.663484, 6.211717, 
    8.228372,
  136.9637, 114.5358, 96.54081, 90.36079, 95.60961, 98.44691, 100.3844, 
    107.9918, 107.6623, 93.50208, 22.51789, 6.29215, 3.26133, 7.204817, 
    8.026834,
  130.8438, 110.3816, 94.72894, 89.33306, 93.2246, 95.40867, 99.18629, 
    103.9554, 103.4363, 88.22191, 23.56927, 6.958236, 4.935464, 7.890628, 
    10.04526,
  111.6337, 91.8197, 84.34911, 82.35535, 86.10698, 88.0366, 98.55688, 
    102.4768, 83.2356, 38.64003, 23.44515, 7.703847, 5.622465, 7.255063, 
    12.02281,
  32.50927, 81.45358, 43.80713, 71.60387, 12.81567, 6.982353, 9.667059, 
    7.020205, 7.605055, 0.5317229, -0.9479934, 1.495114, 0.8275149, 2.068601, 
    -0.3387798,
  91.1184, 97.6827, 103.4084, 94.75546, 16.56893, 6.65987, 11.51831, 
    7.545704, 6.14158, 6.75714, -0.07978026, 6.261873, 8.234672, 0.8442042, 
    -0.3063043,
  100.7904, 100.0999, 109.7211, 109.7658, 67.59688, 2.290895, 8.849565, 
    7.151902, 5.533168, 7.292179, 7.216505, 7.172476, 9.167984, 9.623001, 
    4.323376,
  110.2588, 106.229, 111.7948, 117.355, 115.0207, 66.79968, 3.239507, 
    2.227865, 3.637924, 4.219467, 4.993548, 4.54461, 6.620676, 7.630599, 
    6.571214,
  122.7285, 115.1463, 116.1139, 117.7818, 111.7654, 99.51218, 66.73161, 
    4.002596, 0.6218349, 1.272291, 3.841454, 5.166663, 5.290385, 9.149816, 
    6.353565,
  137.1347, 123.4726, 120.4826, 118.7013, 110.7266, 94.22355, 81.31451, 
    51.53695, 16.9724, 12.23622, 3.594113, 5.170259, 10.22675, 12.17357, 
    9.564744,
  149.1279, 133.3751, 127.4895, 121.1564, 111.2926, 94.67313, 79.86821, 
    58.64264, 45.60876, 39.25768, 13.85659, 5.801545, 10.11314, 12.16992, 
    12.24926,
  151.9458, 138.549, 130.919, 125.2543, 112.8746, 95.80505, 77.1086, 
    65.81042, 64.69772, 54.3854, 9.961553, 4.563283, 9.22791, 12.68642, 
    12.35505,
  137.3895, 135.6548, 132.2379, 127.1491, 113.7518, 94.57756, 73.16664, 
    59.55267, 62.97247, 53.91339, 9.757659, 3.515329, 7.934896, 13.90606, 
    15.25981,
  114.8731, 113.884, 118.5555, 116.9369, 104.844, 86.97745, 64.56825, 
    51.59933, 50.42272, 20.0403, 15.59557, 3.957745, 6.366655, 11.54648, 
    15.59239,
  30.18808, 84.62022, 43.47585, 63.60222, 9.003234, 2.140717, 6.241577, 
    6.751247, 9.361827, 1.787945, 0.5546011, 3.325044, 1.050202, 1.336251, 
    -0.3785072,
  89.2901, 107.056, 112.5555, 97.24577, 9.210705, 1.825709, 6.087929, 
    7.500794, 7.729077, 8.685429, 1.684649, 7.172385, 9.063536, 0.6593789, 
    -0.3660343,
  96.14007, 107.9689, 122.341, 111.2797, 57.71985, 0.8191461, 2.804862, 
    6.527435, 6.606506, 8.496464, 7.978731, 7.953539, 7.795706, 9.637957, 
    3.809421,
  97.4012, 109.3972, 120.3036, 116.0186, 100.9226, 51.7659, 2.197204, 
    1.652244, 5.18921, 5.277846, 5.755652, 5.979486, 6.740044, 6.920969, 
    6.015733,
  93.2859, 109.5849, 119.8859, 115.7827, 96.33742, 75.78777, 47.55151, 
    3.103341, 0.3949554, 0.6734973, 3.511671, 6.431262, 5.271238, 6.232954, 
    7.017113,
  89.23018, 109.4818, 117.9915, 111.6573, 95.82558, 76.7115, 59.08517, 
    33.2608, 14.47476, 13.9872, 3.431054, 6.833865, 6.161099, 7.151192, 
    5.899425,
  98.00774, 110.4625, 115.2062, 107.4661, 95.04036, 76.5915, 62.00294, 
    41.10871, 35.69903, 37.89821, 17.13119, 8.840962, 7.948787, 7.917403, 
    5.938035,
  105.9171, 107.6985, 109.5422, 104.3143, 95.82286, 77.88793, 62.95683, 
    48.22698, 46.18477, 48.10065, 13.29519, 10.88321, 10.55753, 10.07931, 
    7.368233,
  97.09384, 101.3303, 106.2748, 100.9473, 94.26534, 79.95941, 67.11412, 
    53.08924, 47.90296, 44.94852, 10.68196, 10.87008, 12.11396, 12.03743, 
    10.61857,
  88.62538, 88.4072, 91.07698, 90.8297, 86.56057, 75.29155, 68.15191, 
    58.31402, 44.30017, 20.33135, 18.17934, 10.54808, 12.98565, 13.729, 
    14.36697,
  24.57923, 87.54375, 45.5293, 68.36984, 10.51135, 3.388565, 8.643313, 
    7.343522, 8.642472, 1.565436, 0.1354226, 1.037474, 0.1093328, 0.3236986, 
    -0.7445637,
  66.03447, 107.1877, 130.8473, 120.37, 8.502699, 2.100133, 10.46188, 
    8.150336, 6.572431, 6.325274, 1.254235, 3.032681, 4.606669, 0.2559429, 
    -0.7981956,
  61.08755, 99.68035, 135.1019, 132.9292, 64.70701, -0.8013177, 7.425273, 
    8.847104, 7.398215, 5.81604, 5.07602, 3.267292, 3.568213, 5.569273, 
    1.46137,
  65.62801, 97.86332, 129.3069, 131.4884, 125.4186, 64.50034, 0.6746535, 
    2.226521, 4.782799, 4.206266, 3.163759, 2.478707, 2.421834, 3.53519, 
    2.52588,
  67.70213, 97.5533, 125.668, 124.2423, 112.4326, 105.0493, 67.44787, 
    1.951169, -0.355635, 0.6797235, 3.732384, 3.542207, 2.870119, 2.811302, 
    3.617533,
  68.72215, 99.01833, 120.6139, 114.9863, 103.4812, 93.47498, 90.98562, 
    66.36252, 21.0097, 14.88989, 5.896696, 5.54091, 3.250336, 2.695906, 
    3.472968,
  77.41035, 102.5833, 116.5281, 106.8948, 93.52341, 81.57275, 76.43265, 
    64.22813, 47.40879, 37.97075, 17.2997, 6.924463, 3.255536, 2.801549, 
    2.726642,
  76.54099, 101.5757, 110.2919, 100.1256, 87.11421, 74.26595, 66.52436, 
    60.61691, 64.39285, 57.56174, 11.91743, 7.315583, 3.450686, 2.664583, 
    2.325415,
  70.31889, 93.75163, 104.1219, 92.75918, 79.21854, 68.23678, 59.23326, 
    49.88986, 52.16423, 49.24265, 8.475417, 7.523419, 5.309663, 3.84711, 4.059,
  67.93323, 73.58688, 85.36782, 82.24178, 70.97454, 59.83671, 55.28371, 
    46.8718, 38.73386, 14.93961, 19.63724, 12.15921, 7.461158, 7.223077, 
    6.809978,
  26.47719, 85.46861, 31.56744, 40.74089, 7.722154, 2.261551, 5.036795, 
    4.349507, 7.859059, 0.5124635, -1.049118, -0.4210033, -0.5028114, 
    0.356695, -0.7079582,
  105.5777, 117.1837, 116.1522, 92.40034, 6.315258, 1.103365, 5.304066, 
    5.153759, 4.660228, 4.870198, -0.4541016, 1.545104, 4.368216, -0.3715715, 
    -1.419207,
  109.9012, 111.473, 120.6357, 108.7367, 51.29454, 0.3283034, 2.710755, 
    3.947121, 3.45694, 4.184247, 3.185236, 2.239609, 4.351305, 7.880531, 
    1.335079,
  109.5466, 110.2223, 113.0833, 104.9857, 98.38891, 51.20784, 1.804374, 
    1.058605, 1.724231, 1.663301, 1.35853, 0.8497254, 2.154696, 4.192729, 
    2.590097,
  108.4224, 107.4779, 107.7327, 98.52992, 88.61711, 76.47887, 46.60236, 
    2.728671, 0.5688186, 0.6144986, 0.6512331, 1.064924, 1.841826, 3.136277, 
    5.737541,
  106.1909, 104.7672, 102.5325, 91.69552, 85.74497, 73.91805, 61.00898, 
    39.89679, 9.986721, 6.454754, 2.626477, 1.669256, 1.443214, 3.198856, 
    5.099245,
  100.0508, 101.554, 100.0589, 89.2617, 81.37468, 70.13655, 61.33883, 
    47.35518, 30.81644, 20.66212, 8.993962, 2.462138, 1.733932, 3.318035, 
    6.65327,
  89.29751, 94.89266, 96.01482, 86.53867, 79.63798, 70.52106, 61.46402, 
    52.88126, 43.17549, 34.13777, 6.48778, 3.152555, 2.043488, 3.7796, 
    6.266811,
  75.13184, 84.42372, 92.91314, 83.94262, 74.71026, 65.95347, 58.05433, 
    51.62436, 46.49327, 33.88717, 4.542201, 4.52388, 1.71512, 3.46715, 
    5.833891,
  70.85905, 67.70951, 75.36549, 73.44813, 67.69289, 59.36004, 54.16603, 
    49.34906, 37.14367, 9.934594, 18.45495, 6.934974, 2.587228, 2.019352, 
    4.524894,
  18.78163, 52.77678, 14.90022, 14.59516, 5.93289, 0.9605854, 3.03368, 
    2.898131, 5.360455, -0.7691152, -1.395314, -0.5525165, 0.08213606, 
    0.6453346, -0.2734925,
  82.27737, 73.54359, 57.80042, 39.78855, 4.272964, 0.6006019, 2.471731, 
    3.74517, 3.173373, 2.207945, -1.644575, 1.952385, 4.281771, 0.05585356, 
    -1.083858,
  86.27838, 68.86145, 58.49443, 47.59401, 21.96551, 0.4693513, 1.189526, 
    2.880363, 3.071236, 2.178289, 0.5825414, 2.390519, 5.917029, 9.506378, 
    2.369711,
  87.53782, 68.60797, 57.92356, 45.58937, 40.29551, 24.07293, 1.390242, 
    0.5794807, 3.438195, 2.258563, 0.8166333, 1.460459, 3.351725, 5.83935, 
    3.906226,
  87.6755, 73.34155, 63.54002, 51.13981, 38.86657, 36.26987, 22.59074, 
    1.842122, 1.340012, 1.826331, 2.456657, 1.968187, 3.239811, 2.014405, 
    6.575009,
  97.17207, 84.75861, 74.2229, 61.23966, 47.24783, 32.87975, 32.20639, 
    31.69081, 7.027502, 5.677295, 2.993354, 3.910709, 3.601695, 2.348301, 
    5.274329,
  112.6707, 100.8946, 88.19744, 75.48951, 61.24736, 41.68485, 29.67625, 
    32.5138, 29.98355, 20.04575, 7.942853, 9.602835, 11.69892, 5.334942, 
    7.946824,
  118.1627, 111.0942, 99.89064, 86.17458, 70.8885, 55.67154, 41.00448, 
    34.87667, 40.8327, 30.91412, 6.064475, 8.9467, 11.96924, 10.02819, 
    12.53911,
  92.75445, 95.06287, 93.87996, 87.25611, 74.63335, 59.32275, 42.71797, 
    34.45713, 42.58983, 30.40879, 3.159762, 6.107217, 8.336852, 13.0379, 
    12.56552,
  39.55753, 45.69468, 57.62575, 64.87571, 66.90756, 58.24409, 46.98421, 
    38.7984, 34.37933, 18.54759, 14.1199, 6.09305, 5.813642, 10.29587, 
    17.05504,
  13.30149, 32.53336, 8.355282, 7.407232, 4.22814, 1.048014, 0.7153053, 
    0.5866193, 1.625545, -1.428348, -1.940767, -0.9561903, -1.127535, 
    -0.09182524, -1.584681,
  68.3721, 56.88147, 40.11684, 26.03813, 4.508847, 0.5273022, 0.9635403, 
    0.3278145, -0.0009985565, 0.6875437, -2.445827, 2.52393, 6.510187, 
    -1.549051, -2.793425,
  81.39851, 65.60841, 47.99545, 39.95062, 14.0932, 0.810169, 0.7681339, 
    0.7338738, 0.5268404, 0.6401086, 0.1434827, 2.424726, 7.236571, 10.65053, 
    3.623119,
  88.70378, 73.79662, 60.76027, 51.87826, 39.78304, 19.37771, 1.885115, 
    0.5253685, 1.039932, -0.08564169, 0.03022117, 0.8721144, 4.214062, 
    8.791627, 7.751519,
  101.6248, 84.05923, 72.09203, 58.90822, 42.36943, 30.58704, 29.08043, 
    2.308074, 0.9087524, 0.1503799, -0.453934, 0.01041596, 2.467347, 
    4.409618, 10.49641,
  124.374, 100.4672, 82.80069, 65.71591, 50.5032, 35.18113, 39.07077, 
    32.55652, 4.37772, 3.244015, 1.955873, -0.1146376, 0.9613274, 2.619037, 
    8.54131,
  145.0918, 121.5093, 95.17712, 72.43375, 54.97179, 43.27481, 46.91421, 
    47.55139, 21.87001, 12.02665, 0.9822231, 0.4269893, 0.7771398, 1.805971, 
    5.175327,
  84.00933, 95.23468, 92.83062, 82.95136, 67.74385, 53.99934, 52.55643, 
    55.76779, 48.22968, 20.26272, 1.448886, 0.6188775, 0.9310435, 1.857559, 
    5.942267,
  29.90461, 28.22689, 39.70499, 47.87196, 56.61988, 56.90285, 52.57628, 
    50.88248, 49.68959, 25.42119, 0.7054198, 0.6385462, 0.4554259, 2.111306, 
    9.812976,
  47.57483, 30.0147, 18.88925, 16.17144, 22.56445, 34.83792, 45.58129, 
    45.74036, 33.89213, 10.32452, 9.544725, 1.571931, 0.5819535, 1.788452, 
    11.1174,
  13.57814, 34.1977, 12.2607, 9.249291, 0.5059137, 0.7741088, 3.914135, 
    1.709165, 0.8641163, -2.033188, -1.920604, -1.175854, -2.425058, 
    -1.072011, -2.287942,
  74.78226, 60.23242, 41.62208, 24.98189, 1.29598, 0.8391411, 1.800985, 
    5.049444, 0.5213516, 0.4465938, -1.461738, 2.136908, 6.219481, -2.815194, 
    -3.692159,
  104.0417, 75.02303, 54.88061, 47.97498, 9.977523, 0.9378572, 1.874602, 
    0.6005602, 0.1346452, 0.2656295, 0.5669618, 3.213577, 9.15824, 6.46928, 
    1.046759,
  111.0852, 91.2922, 68.40704, 57.97689, 34.92154, 19.50797, 1.576279, 
    0.3586957, 0.9098591, -0.1441196, 0.6145869, 1.436572, 6.872272, 
    9.558455, 3.188888,
  112.609, 96.64046, 80.47746, 64.25097, 49.81643, 27.98478, 25.65077, 
    2.555064, 1.333963, 0.8687795, 1.896384, 0.2914441, 2.005431, 4.037496, 
    5.690548,
  127.1416, 105.1932, 87.03973, 69.5534, 54.22186, 31.27092, 33.49612, 
    20.94199, 5.129068, 1.758508, 1.192667, 0.2278414, 1.043189, 2.727348, 
    5.636965,
  143.252, 115.2759, 92.98357, 75.30956, 59.79359, 40.08524, 36.57541, 
    33.77793, 23.47128, 9.547459, 1.881151, 1.342453, 0.9182288, 1.058129, 
    4.482892,
  129.3354, 114.8389, 97.59138, 82.43187, 69.3362, 52.93929, 42.8776, 
    44.81554, 40.03536, 20.41593, 3.822012, 2.024852, 1.172462, 0.8066443, 
    5.054892,
  83.22093, 87.92197, 84.60986, 74.09715, 66.51075, 57.17056, 45.71261, 
    42.73257, 43.8128, 19.65173, 5.719695, 2.500978, 1.216195, 0.8742379, 
    8.876205,
  49.56099, 50.45634, 54.73209, 51.43567, 46.83803, 39.51837, 35.63923, 
    30.77153, 20.21692, 11.56435, 13.89837, 6.384721, 2.708577, 1.359933, 
    2.586909,
  23.41496, 49.97394, 21.3794, 17.12297, 9.025062, 4.073584, 5.569523, 
    3.969945, 0.1256429, 0.1748729, 0.1838249, -1.81349, -2.532548, 
    -1.070713, -1.295746,
  102.8972, 113.078, 101.1623, 63.43551, 4.357746, 2.141901, 5.054039, 
    5.89582, 1.016136, 0.123897, -0.3247503, 0.1553202, 0.9931154, -2.406762, 
    -2.305177,
  131.1096, 107.578, 105.7801, 91.31606, 32.81245, 0.49412, 1.669903, 
    4.069776, 0.966688, 0.4910338, 0.8994322, 3.041832, 4.777748, 2.005229, 
    -0.1447813,
  124.8587, 100.9399, 92.42648, 84.71326, 68.12788, 25.80164, 1.089392, 
    0.9511096, 0.551167, 0.2553824, 0.4369473, 4.464934, 4.321387, 3.827909, 
    0.8551162,
  120.2555, 98.7739, 83.09498, 68.2732, 53.19942, 38.30709, 23.57843, 
    0.7229719, -0.1056403, 1.294129, 0.910893, 5.231286, 3.469577, 1.549408, 
    1.553757,
  117.8531, 102.2303, 83.61473, 65.45231, 50.02188, 37.28321, 31.27781, 
    13.15704, 4.682369, 2.492971, 1.844992, 5.442476, 2.79801, 0.3859285, 
    1.249109,
  122.7208, 106.3293, 88.25124, 71.63872, 59.36905, 49.06512, 45.49749, 
    34.44044, 10.49614, 7.618894, 4.471473, 3.554519, 2.136803, 0.257809, 
    0.5811884,
  126.7441, 107.3773, 92.54943, 79.67731, 70.74802, 61.4152, 54.72653, 
    48.96899, 36.64364, 10.6842, 5.784152, 3.475363, 1.692901, 0.2138115, 
    1.19219,
  120.0001, 106.3708, 97.67731, 84.4561, 74.64599, 67.32226, 57.91807, 
    50.4833, 42.52057, 8.942161, 3.080378, 1.727621, 2.347973, 0.7866868, 
    1.549434,
  105.3979, 91.47171, 85.90102, 78.07801, 68.15745, 59.60543, 53.51885, 
    43.82676, 19.27892, 4.433223, 15.33205, 12.64189, 6.926015, 3.822307, 
    1.624696,
  22.22833, 41.37538, 26.72543, 18.32915, 7.438858, 1.596839, 5.425286, 
    2.449892, 1.986639, 0.7831967, 0.08850629, 0.001944832, -2.485955, 
    -1.065739, -1.748997,
  91.24485, 115.6091, 113.8874, 65.07887, 4.520698, 0.2312146, 5.564359, 
    4.209386, 3.166172, 2.751459, -0.1489739, 0.9640814, 2.42536, -1.007937, 
    -1.325,
  123.2562, 130.4299, 142.3843, 126.6546, 48.81153, -1.261877, 1.284333, 
    5.18229, 5.850114, 1.7462, 1.701533, 3.880837, 3.872205, 4.79714, 1.124696,
  124.9263, 130.1762, 135.0383, 130.4988, 115.7138, 46.80382, 1.172284, 
    1.626661, 0.8985941, 1.27995, 2.013076, 5.829338, 3.696787, 3.810457, 
    3.563014,
  127.5713, 129.1324, 128.0264, 119.7102, 104.8124, 86.13882, 40.59246, 
    1.370446, 0.6574772, 0.8781065, 2.284708, 4.543116, 2.786208, 0.4796868, 
    3.941795,
  130.1723, 129.5411, 123.8853, 111.4149, 97.59155, 80.6694, 63.58323, 
    25.23462, 6.342264, 3.1422, 1.922023, 4.164571, 3.01382, 0.03829878, 
    3.104929,
  136.105, 130.1023, 117.1698, 101.8401, 87.08183, 71.64167, 60.77864, 
    44.38995, 20.78153, 8.88689, 5.473445, 4.665816, 3.763793, 0.2467589, 
    1.909569,
  134.9875, 121.0809, 106.4883, 91.64308, 79.61833, 65.30515, 56.09495, 
    49.81306, 36.52143, 5.017908, 1.399805, 3.910501, 5.261173, 2.439451, 
    0.2336047,
  118.4609, 109.0607, 99.55521, 82.19293, 69.74351, 62.12638, 55.14629, 
    48.93284, 42.53249, 8.116418, 3.57538, 7.980077, 7.450477, 4.076424, 
    0.8442473,
  96.87086, 82.99832, 76.27638, 68.51903, 61.49507, 56.25101, 53.88441, 
    48.39561, 22.9142, 6.003797, 12.9489, 9.511526, 5.841746, 3.440416, 
    1.272064,
  22.6576, 32.4407, 18.17668, 11.54107, 3.767122, 0.6167119, 2.206626, 
    1.242267, 1.02083, -0.7703428, -1.128839, 0.30199, 0.2912996, 1.08073, 
    -0.7883871,
  104.5952, 102.4739, 90.40776, 36.42833, 2.40574, -0.2851488, 1.943156, 
    1.327826, 1.461751, 1.114768, -1.799542, 0.1077398, 4.438672, -0.2801046, 
    -1.316779,
  134.59, 124.3738, 125.5938, 102.6243, 39.6147, -1.008629, 0.4807245, 
    0.8904589, 2.473561, 2.526087, 2.62651, 2.219491, 3.614229, 5.362515, 
    0.9192011,
  127.8646, 118.3296, 114.8677, 114.6179, 105.9822, 42.28569, 1.23608, 
    1.014671, 0.5810108, 1.670663, 3.58618, 5.066324, 2.401541, 6.277529, 
    2.598217,
  116.82, 110.0764, 105.7363, 104.7175, 101.714, 89.84661, 47.13345, 
    1.814595, 1.092597, 0.9263912, 3.462831, 5.695686, 4.510716, 6.316182, 
    4.13028,
  109.3323, 106.2468, 100.7064, 98.01514, 95.51157, 88.2784, 73.84159, 
    28.1215, 4.637388, 3.252171, 2.072342, 5.487834, 6.244354, 1.758876, 
    4.931785,
  107.6027, 105.5856, 98.34628, 92.20093, 90.53793, 83.53003, 75.43031, 
    58.51278, 32.12598, 7.967865, 4.807187, 4.652191, 7.83581, 2.331764, 
    4.884169,
  102.7907, 98.10677, 93.18297, 87.43872, 86.05378, 81.12525, 72.84167, 
    67.84283, 53.13207, 6.824866, 3.561195, 6.098897, 6.900964, 5.395291, 
    3.982335,
  87.96717, 88.31148, 88.83035, 78.97267, 72.97, 72.61009, 68.49818, 61.1498, 
    53.6131, 16.7996, 0.8701842, -0.4665387, 3.903913, 2.39498, 2.630861,
  65.93203, 63.70838, 64.57483, 61.38929, 58.09587, 56.21888, 56.8648, 
    54.0829, 34.17706, 6.281018, 9.603544, 0.8643194, 0.07140119, 2.834181, 
    1.59824,
  17.08274, 22.79878, 12.19366, 6.518814, 0.9467631, 0.6370949, 2.524407, 
    2.412424, 3.345431, 1.178244, 0.5990047, 1.947864, -3.061199, -0.3629045, 
    -2.075095,
  89.72498, 78.88132, 70.80174, 19.49694, 0.8558829, 0.2982442, 0.5296374, 
    4.013184, 5.226988, 5.396495, 2.585808, 5.731801, 4.715858, -1.312606, 
    -1.986089,
  125.9799, 109.1019, 105.8027, 77.85902, 28.76685, 0.3009539, 0.7404091, 
    1.241367, 3.300524, 3.742934, 6.396356, 8.760115, 9.395368, 7.533149, 
    2.697002,
  126.5396, 111.0333, 101.0616, 95.2252, 86.14955, 32.39393, 1.476258, 
    1.1478, 1.847766, 3.035673, 4.693535, 9.132061, 10.54852, 10.21661, 
    4.947008,
  123.994, 110.3615, 99.37972, 90.56306, 84.56766, 75.50903, 39.64746, 
    1.908824, -0.1341741, 1.216959, 3.030031, 4.887264, 9.314935, 9.321968, 
    8.712398,
  118.4656, 110.6659, 97.24171, 86.96208, 80.12447, 74.22636, 66.38262, 
    29.21091, 4.293637, 1.129684, 0.6290677, 2.606295, 7.735639, 8.159175, 
    10.53386,
  114.1842, 108.3779, 94.47625, 83.08455, 76.17387, 68.49342, 65.19955, 
    53.25021, 27.70503, 4.474119, 0.8748928, 1.706829, 6.735674, 7.688566, 
    9.97698,
  108.1836, 99.39413, 89.15707, 79.99306, 73.23821, 64.03442, 57.10177, 
    52.6415, 38.28222, 7.933767, 0.7634932, 1.308966, 3.388895, 4.429898, 
    9.216691,
  87.18431, 86.3454, 84.96982, 73.35369, 64.98226, 59.65019, 52.29439, 
    44.0552, 39.48341, 15.87989, 2.627708, 1.461246, 0.444689, -0.5053429, 
    6.303177,
  47.43485, 47.05842, 48.2165, 46.88092, 43.49154, 37.90566, 35.46536, 
    32.77933, 20.92215, 7.014334, 13.57057, 4.201021, -0.2979303, -0.3725488, 
    3.212216,
  10.53724, 16.54176, 7.117758, 2.504647, 1.682591, 0.4128057, 0.2766299, 
    0.09710203, 0.6932734, -0.9842138, -0.5500378, 2.870814, 1.543371, 
    0.6008071, -0.3279994,
  74.27631, 63.69739, 51.66106, 10.81565, 0.7135787, -0.0780296, 0.7539436, 
    0.5714356, 1.062332, 0.9171147, 0.0526816, 5.926825, 6.276806, 0.4043359, 
    -0.1970292,
  102.1033, 82.89684, 68.58689, 42.45002, 15.7169, -0.04038233, 0.9750904, 
    1.097207, 0.6391953, 1.610436, 1.511192, 6.331003, 5.515947, 5.363008, 
    1.909152,
  94.2893, 73.99242, 59.22892, 53.97691, 53.13985, 25.88139, -0.5031691, 
    0.4601661, 0.6478425, 2.041674, 0.4924111, 4.852791, 6.516751, 4.714964, 
    4.085649,
  91.00934, 73.39039, 63.3561, 60.73801, 63.66508, 58.23418, 34.45382, 
    -0.2865628, -0.4529567, 0.6246152, 0.4340631, 2.115819, 6.811916, 
    5.050382, 3.940291,
  91.50684, 80.97996, 72.70546, 69.38122, 66.99736, 61.93395, 49.38157, 
    19.98278, 1.467786, 0.8163297, 0.4999828, 1.111216, 6.37607, 5.176373, 
    3.410509,
  102.2583, 93.00263, 81.38353, 73.52991, 67.73954, 55.82565, 44.06916, 
    28.2466, 8.091382, 1.590002, 3.603325, 0.4251748, 8.575987, 7.192189, 
    4.129333,
  117.3091, 98.69096, 84.92051, 74.10898, 63.5275, 47.44484, 32.31718, 
    23.53262, 11.17871, 1.414122, 2.255944, 0.8335972, 5.082013, 8.726713, 
    5.790557,
  116.3438, 98.79052, 86.3037, 64.16962, 46.22614, 35.11141, 26.80191, 
    19.49836, 19.52842, 2.802256, 0.3982889, 1.860684, -0.3052516, 9.17203, 
    7.959656,
  85.03412, 60.63144, 43.46054, 30.9631, 23.43472, 17.54529, 13.05361, 
    11.47727, 5.306835, 1.182497, 6.138447, 4.773204, -0.1487855, 0.1926806, 
    6.418915,
  7.246726, 7.722124, 2.542367, 1.151054, -0.07612758, -0.8464163, 0.5221314, 
    1.700409, 3.198539, 0.3243846, 0.08580402, 0.6634401, -0.1916987, 
    -0.2634647, -0.6662365,
  58.2199, 37.29919, 22.75604, 4.520345, -1.917446, -2.903551, 0.4648795, 
    0.8115535, 2.708542, 2.76171, 0.7949862, 2.166757, 1.796563, -0.5174991, 
    -1.155372,
  79.22413, 50.22612, 38.10333, 37.55997, 9.458339, -4.661607, -0.5554881, 
    0.6033998, 3.045292, 2.915061, 3.225939, 1.227774, 0.9243242, 1.7286, 
    0.5306609,
  77.64022, 52.14898, 45.12033, 57.78852, 63.11992, 21.69567, -4.955317, 
    -0.8598396, 0.1724278, 3.034958, 1.172018, 1.126351, 0.8137801, 1.893374, 
    1.500754,
  76.92761, 59.07192, 56.1985, 64.07368, 69.28941, 57.11776, 18.87615, 
    -0.393273, -0.392643, 0.05242146, 0.9163216, 0.9349968, 0.889462, 
    1.348927, 2.945161,
  80.68804, 72.46483, 65.87189, 63.92653, 64.63512, 53.8386, 32.24916, 
    6.037809, 0.4705498, 1.151992, 2.375057, 2.528286, 0.6164359, 0.7661468, 
    2.62862,
  87.63432, 79.33015, 67.46415, 62.40193, 60.74817, 44.32622, 29.77818, 
    16.20581, 3.666794, 2.050765, 4.515259, 1.164024, 1.153472, 0.6023744, 
    1.416373,
  107.0292, 88.11824, 74.2562, 66.67204, 58.00711, 37.96879, 23.13296, 
    16.79456, 7.003991, 4.458494, 3.97069, 2.632654, 1.545469, 1.077764, 
    1.10984,
  120.0127, 100.9114, 87.51768, 66.10465, 44.65312, 29.81259, 21.70095, 
    12.85546, 20.47687, 7.983472, 5.416316, 4.646871, 3.401493, 3.171158, 
    0.6614599,
  116.0796, 90.63185, 68.54478, 51.21669, 34.01461, 25.30859, 15.53687, 
    18.15434, 10.32999, 2.254669, 7.632349, 6.066761, 6.463171, 3.882585, 
    1.426278,
  11.09611, 10.35876, 4.550984, 3.553478, -0.3129986, -1.001043, -0.3654585, 
    -1.909333, -1.253081, -1.521389, -2.075215, -0.9933099, -1.139876, 
    -0.4398958, -0.5344399,
  61.02659, 48.06143, 38.10545, 7.428717, -3.03936, -3.080598, 0.07463632, 
    -2.917236, -2.01302, -0.3237132, -1.566895, 0.343835, -0.2687302, 
    -0.8874721, -0.7694766,
  102.2306, 80.73547, 72.74444, 59.77872, 11.72549, -6.219584, -0.9898472, 
    -1.439836, -0.8284131, -0.4333771, 0.7292968, -0.4291794, -0.009113139, 
    0.7599922, 0.5420966,
  107.7566, 90.48556, 79.81256, 78.41113, 76.17835, 21.98814, -6.907546, 
    -1.613366, -0.7476686, -1.373742, -1.124215, -0.07554233, -0.02159486, 
    1.448426, 0.8455588,
  100.816, 91.61137, 83.3195, 80.33856, 77.1692, 62.42758, 22.78151, 
    2.472059, 1.319631, -3.535224, -1.603065, -0.6341151, 0.5534724, 1.07504, 
    2.444677,
  97.00207, 90.35598, 83.10506, 77.17623, 70.48801, 61.35701, 46.10346, 
    12.26883, -1.569687, -1.045488, -0.7801447, 0.4420822, 0.5284873, 
    0.7073554, 2.70805,
  117.2422, 102.9123, 87.42103, 76.73817, 69.58231, 60.27348, 53.95155, 
    40.01564, 10.7631, 0.563759, 0.2021647, -0.01071768, 0.4107583, 
    0.2465282, 2.026705,
  134.3343, 114.3648, 98.56543, 85.10333, 75.54594, 65.06734, 53.71107, 
    44.37587, 15.56352, 3.592594, 0.1145135, 0.08604349, 0.8994926, 
    0.6351922, 1.927069,
  125.7478, 115.8997, 107.6107, 85.74478, 72.18227, 64.81384, 54.3349, 
    26.85908, 27.24333, 7.301414, 0.920945, 0.6371266, 0.7114252, 2.835636, 
    1.795042,
  102.4674, 92.4741, 83.31606, 76.30054, 70.70908, 51.52143, 25.69902, 
    25.90574, 13.18707, 3.061278, 10.52678, 3.170315, 0.8643384, 5.493074, 
    1.271303,
  14.58924, 16.78651, 10.6947, 8.427719, 1.065692, 1.286234, 2.688967, 
    0.5406233, -1.103798, -4.557888, -5.559404, -4.7809, -3.58154, 
    -0.3985161, 0.08429023,
  63.89902, 64.33423, 68.15115, 23.23631, -1.381936, 0.4095814, 4.436946, 
    1.387655, -0.4176323, -2.481973, -4.805069, -3.039433, -2.310397, 
    -0.902095, 0.2273798,
  100.4755, 102.544, 105.2819, 89.39794, 22.39526, -3.385552, 6.246519, 
    2.007766, 0.2501453, -1.418857, -1.83044, -2.676917, -1.890622, 
    0.3202477, 3.138744,
  94.44328, 96.11738, 96.97085, 101.8043, 99.63952, 37.9515, -5.252584, 
    1.93853, 2.157538, 0.9811754, -0.5571719, -1.343664, -0.8591319, 
    1.149935, 6.47956,
  88.68691, 87.99039, 90.73826, 96.89995, 99.25885, 91.00958, 47.88388, 
    -3.710571, 5.539172, 0.7220715, 0.985905, -1.424792, -1.023717, 
    0.8506967, 7.915033,
  90.99182, 90.4763, 91.69444, 93.82588, 93.943, 89.95068, 78.79163, 
    39.35892, 2.719269, -1.518754, -2.093357, -1.078406, -0.8990402, 
    1.104421, 7.991939,
  105.8016, 104.9553, 96.90771, 90.13425, 86.89614, 78.24458, 72.35986, 
    58.15146, 31.03196, 4.111075, -0.2803243, -1.075849, -0.4818511, 
    1.675105, 9.507362,
  107.1344, 99.29503, 89.72141, 78.418, 72.18621, 62.51011, 52.66475, 
    48.25158, 28.13189, 3.673615, -1.328251, -1.215957, -0.06426112, 
    4.294222, 8.811193,
  90.27811, 85.33817, 83.36359, 61.23458, 48.87893, 43.47573, 40.93189, 
    28.91154, 27.32003, 5.934484, -0.6122813, -0.8283917, -0.1801715, 
    7.123547, 8.089182,
  76.29438, 59.90445, 50.89516, 42.09608, 36.43325, 25.21506, 18.30215, 
    24.93946, 20.5172, 9.006474, 11.31887, 2.105595, 1.458268, 11.84436, 
    10.06992,
  15.72382, 19.07047, 10.70595, 7.113619, -0.6367933, 1.363595, 3.806137, 
    -0.2206943, -1.613441, -1.564519, -1.055347, -0.4605925, -1.327691, 
    -0.4374749, -1.302706,
  62.23787, 67.84962, 74.99915, 28.27457, -3.28436, 3.188649, 7.877884, 
    0.60919, -0.6572022, -1.339212, 0.8426532, 3.191484, -1.094352, 
    -2.434501, -1.815938,
  125.7949, 124.0461, 126.0558, 106.2739, 18.06061, 4.509028, 12.26436, 
    3.356738, 0.8128174, 1.42373, 4.641937, 1.424961, -1.052207, -0.3982835, 
    2.00405,
  135.1759, 131.3084, 125.604, 121.8303, 114.664, 47.97168, -2.910938, 
    6.12469, 8.305097, 7.596898, 4.87257, 0.9738377, 0.9320605, 2.058074, 
    7.833517,
  138.3601, 134.2627, 126.9165, 121.4669, 116.163, 103.3968, 54.09521, 
    3.516146, 4.112544, 6.704878, 5.296577, 0.3917941, 1.435472, 2.512043, 
    9.978131,
  129.419, 131.443, 128.7714, 119.5501, 110.619, 96.38457, 76.9692, 43.10973, 
    7.056839, 2.640622, 0.4069771, 0.9048219, 2.178325, 3.39434, 8.868921,
  117.5053, 124.1768, 118.0266, 110.1082, 97.46327, 79.39495, 61.92112, 
    39.97672, 19.38669, 6.607297, 1.081368, 0.8099793, 2.017826, 7.226653, 
    11.05634,
  104.5738, 100.1254, 96.15104, 89.78866, 80.24786, 65.37197, 44.86188, 
    30.39183, 17.83506, 2.98122, -0.962851, 4.089853, 3.27943, 11.71073, 
    9.343472,
  91.6655, 87.76267, 86.63747, 67.34834, 58.8918, 52.90306, 36.70835, 
    21.57247, 15.76316, 4.457379, -0.02230215, 4.856136, 6.428777, 15.64835, 
    7.751491,
  68.79224, 56.1526, 48.44509, 41.20295, 38.58993, 29.03275, 16.46228, 
    13.00393, 9.805787, 2.6528, 11.01609, 9.077023, 13.82538, 19.40878, 
    12.06738,
  20.60157, 30.32688, 19.89192, 15.88396, 2.453444, 6.697354, 12.18001, 
    2.74144, 0.6514192, -1.074935, -0.3154721, 0.6796522, -0.1562666, 
    1.455447, -1.414905,
  68.29458, 82.65501, 82.98494, 42.02277, -0.6128617, 14.4743, 22.7748, 
    5.11364, 2.850668, 0.9826097, 0.5877157, 5.08845, 4.513945, -0.6439924, 
    -1.483436,
  123.899, 145.898, 155.5166, 133.6622, 29.59651, 0.4474408, 31.42752, 
    10.40829, 2.882557, 1.965476, 3.908322, 4.813197, 5.317468, 2.042396, 
    2.154827,
  87.04647, 112.8011, 130.3719, 144.513, 150.7506, 67.82391, 1.031154, 
    14.67446, 13.43662, 4.940795, 5.153761, 6.765351, 4.549097, 4.390751, 
    8.450621,
  52.67962, 61.86754, 77.87392, 101.2584, 125.0484, 137.7057, 90.30102, 
    2.356297, 3.353236, 10.72205, 12.78035, 6.095914, 4.626577, 5.371455, 
    10.88862,
  38.24305, 38.59344, 40.7076, 52.74179, 71.71147, 94.86112, 118.6036, 
    94.47249, 16.92625, 7.052399, 6.424479, 5.805183, 5.191628, 9.314658, 
    7.60779,
  41.93066, 37.36334, 26.95583, 26.85499, 32.28986, 45.95699, 62.85778, 
    82.65483, 67.14292, 17.50184, 9.85369, 5.877537, 5.700848, 12.14485, 
    8.841957,
  47.59095, 35.06035, 23.88915, 18.40948, 18.12976, 25.71507, 29.21385, 
    41.80032, 36.72779, 16.42183, 11.18068, 6.265831, 10.91283, 12.15478, 
    4.963975,
  63.56519, 57.4529, 44.70818, 23.2788, 14.65771, 16.59018, 25.2606, 
    26.94181, 23.28276, 19.42702, 12.92336, 10.4985, 13.11523, 11.61774, 
    4.606426,
  65.46201, 56.60966, 41.9995, 26.29555, 15.37045, 6.685363, 7.679442, 
    13.22472, 15.76409, 11.76514, 22.25762, 15.66688, 18.20195, 14.46988, 
    9.143884,
  22.31285, 41.82386, 23.81147, 19.84408, 1.913201, 7.394906, 15.21095, 
    2.941142, 1.371723, -0.745594, -0.5474017, 0.8977721, -0.05770789, 
    0.340385, -0.4151376,
  60.24287, 76.22002, 67.01897, 33.8489, 0.08519208, 17.09135, 24.19915, 
    4.906903, 2.703791, 1.536101, 1.021081, 3.028128, 1.920331, -0.2932227, 
    -0.1344599,
  129.073, 139.5308, 151.3822, 128.5015, 30.57735, -0.766568, 28.06095, 
    9.183539, 4.207488, 2.278802, 4.007248, 2.195721, 1.527375, 1.34636, 
    -0.6190421,
  71.36657, 130.7758, 146.0695, 160.6456, 158.6333, 62.49929, -1.411533, 
    12.44693, 11.30653, 5.460469, 4.152697, 3.486592, 2.78645, 3.450991, 
    3.013888,
  19.32068, 76.99693, 117.6985, 135.3599, 155.0155, 142.1637, 91.00884, 
    -1.471523, 0.3412119, 7.764553, 12.71935, 5.746925, 3.715983, 6.524325, 
    5.59503,
  49.47943, 41.90141, 83.13833, 101.7558, 121.6066, 126.553, 126.9997, 
    90.95529, 19.34705, 7.405837, 7.564253, 9.83874, 5.752183, 5.678336, 
    3.028652,
  86.1485, 58.89543, 58.26816, 74.37655, 93.902, 102.0984, 104.5146, 
    96.96236, 72.1911, 22.33753, 12.01586, 7.443448, 6.58411, 4.833464, 
    2.50026,
  113.4389, 74.77645, 47.49895, 43.21021, 56.47236, 67.45911, 70.78571, 
    75.81577, 64.91847, 16.34413, 12.06474, 10.6332, 7.060524, 1.812683, 
    1.59411,
  134.8289, 116.9446, 89.39108, 52.38294, 33.32264, 28.78196, 35.29733, 
    41.1111, 34.26794, 15.21102, 9.442139, 14.66119, 5.44729, 3.259635, 
    2.266409,
  117.2437, 108.7467, 97.17236, 78.41349, 62.59727, 40.71472, 15.35693, 
    17.45927, 14.42144, 12.34039, 17.30555, 18.46424, 11.18237, 6.489121, 
    8.142972,
  19.89256, 38.32197, 23.92707, 16.20843, 0.1235649, 4.226707, 9.525249, 
    0.9393094, 3.09822, 0.01007217, -0.5800887, 0.8250026, 0.1331111, 
    -0.1268196, -0.2605721,
  55.4377, 66.36122, 55.91887, 24.03334, -1.471316, 11.40703, 10.69614, 
    1.457098, 0.8986131, 1.900687, 0.5258155, 1.554246, 2.064913, 0.0321008, 
    -0.2022071,
  139.9185, 118.7841, 127.4246, 90.10793, 23.28973, -3.109636, 8.88983, 
    2.146485, 0.6237631, 0.620444, 3.061792, 0.2374202, -0.08518, 1.155644, 
    0.09802637,
  138.7178, 138.8376, 148.6567, 161.5416, 138.7313, 47.10777, -3.120254, 
    2.008982, 1.993137, 0.709151, 0.6035123, 0.3502293, -0.0004253625, 
    0.8147698, 2.333973,
  120.8029, 126.7297, 137.3749, 149.0183, 153.7443, 132.3467, 81.57898, 
    -2.065093, -2.273005, 1.589857, 4.034198, 2.718947, 0.9015378, 1.882506, 
    3.78464,
  105.729, 116.7153, 124.7765, 131.653, 140.1079, 134.7871, 129.0983, 
    83.74647, 20.76351, 8.892305, 9.277593, 6.082729, 1.574183, 1.358453, 
    0.7865368,
  99.74789, 108.0068, 111.3518, 115.5965, 120.994, 119.4792, 116.5507, 
    104.6818, 79.20172, 29.50753, 12.8985, 3.873017, 1.844878, 1.403048, 
    0.2956401,
  106.0831, 95.43082, 96.10548, 99.86343, 104.737, 104.9484, 99.24001, 
    99.0429, 79.9278, 18.85373, 6.013254, 2.924318, 1.924449, 0.2722466, 
    -0.5743543,
  109.3908, 92.57372, 89.33399, 81.73631, 83.99887, 86.65121, 87.77892, 
    84.01328, 62.5155, 9.605803, 2.018128, 3.640275, 1.184665, 0.02972057, 
    -0.6723465,
  118.5799, 93.41724, 74.78822, 61.09295, 59.93667, 55.70576, 47.02143, 
    44.05295, 27.64898, 4.355146, 20.8393, 11.43981, 4.431174, 1.808198, 
    2.046512,
  20.99783, 34.96086, 19.54382, 11.34887, 1.211518, 1.701319, 9.63632, 
    3.670358, 6.784611, 1.711643, -0.2112006, 1.409892, 0.05721566, 
    -0.1645085, -0.5037336,
  63.27058, 69.04553, 59.93394, 17.27278, -0.539054, 3.159139, 4.322719, 
    2.373714, 2.456975, 5.384324, 0.2043052, 2.294691, 4.096256, 0.002093374, 
    -0.3678253,
  146.8741, 118.4246, 114.6226, 59.11048, 20.66039, -2.599115, 1.537438, 
    1.069307, 0.9125943, 1.108115, 3.738207, 1.476287, 0.9181105, 2.023468, 
    0.1710481,
  166.4726, 159.787, 154.1886, 140.2215, 109.0107, 36.95096, -1.684811, 
    -0.510194, 0.4456949, 0.3688377, 0.2544344, 0.4800326, 0.341624, 
    0.837231, 0.8030855,
  160.7214, 153.2652, 148.9286, 144.3466, 132.2302, 111.0273, 72.36047, 
    -0.6806368, -1.104578, 0.5506509, 1.100345, 1.599476, 0.3967465, 
    0.9456145, 1.53078,
  161.1817, 148.8614, 141.5025, 134.8767, 129.4132, 121.2184, 105.1389, 
    60.90562, 17.07412, 10.03014, 3.388005, 2.480997, 0.5734553, 0.3286156, 
    0.5311942,
  160.6834, 156.5592, 139.9457, 127.0052, 121.4512, 113.5024, 103.786, 
    86.42385, 63.31908, 23.57274, 6.351859, 0.8659413, 0.6260529, 0.2638762, 
    0.02923573,
  157.9491, 144.1775, 132.8425, 122.1266, 113.5636, 106.471, 93.27217, 
    86.82108, 67.68479, 13.71044, 0.9636956, 0.1246292, 0.4871922, 
    -0.07826704, -0.1344487,
  141.8503, 136.0471, 134.2692, 114.6693, 101.83, 94.73858, 85.71942, 
    78.26839, 59.29343, 3.759375, -0.3686389, 0.5323474, 0.2991954, 
    -0.151412, 0.08454645,
  112.7322, 107.3674, 102.1606, 91.31337, 87.60993, 76.61287, 60.09325, 
    51.21246, 11.30759, 1.20857, 11.84962, 2.734981, 0.7090364, 0.474739, 
    0.6024845,
  22.23557, 31.86886, 16.60464, 12.37874, 4.077756, 1.152878, 5.734324, 
    2.26664, 7.314206, 1.098366, -0.9157621, -0.01312651, -0.2673116, 
    -0.001310782, -0.521365,
  78.35322, 64.58408, 60.62361, 20.76217, 4.31933, 0.05428689, 2.273893, 
    1.229744, 1.269176, 5.978805, -0.6641939, 0.9222888, 4.413029, 
    -0.2352125, -0.5051381,
  146.9324, 109.49, 106.9174, 43.38867, 30.00633, -1.562005, 0.3198791, 
    0.9749001, 0.9638099, 1.392915, 2.60321, 0.7150165, 1.256325, 2.322798, 
    0.3247022,
  182.0668, 167.938, 152.2977, 116.7198, 89.17094, 39.09883, -0.196683, 
    0.2328766, 1.116352, 0.2832803, -0.001485779, -0.3052641, -0.2137082, 
    0.2538901, 0.3330145,
  181.2013, 164.3027, 145.9015, 134.4036, 114.7405, 90.38945, 61.93287, 
    1.18782, -0.2507572, -0.30248, -0.2397035, 0.07863513, -0.2816444, 
    0.028429, 1.020561,
  187.3037, 163.5353, 141.3132, 125.2299, 115.9747, 101.7845, 80.3368, 
    46.59472, 16.14249, 9.915348, 1.265805, 0.8271359, -0.2130556, 
    -0.1396713, 0.5810201,
  192.9508, 173.0439, 142.7937, 122.384, 109.3453, 101.1221, 90.67538, 
    76.4241, 53.09095, 19.24258, 3.534718, 0.314263, -0.1946273, -0.2789749, 
    -0.5259003,
  191.6284, 163.6473, 138.6517, 119.4478, 105.75, 97.9306, 88.52231, 
    84.07422, 50.8004, 8.81254, 1.037233, 0.5060514, 0.06616116, -0.6467129, 
    -0.6022408,
  177.6573, 157.3645, 141.5645, 113.9118, 97.00634, 85.96732, 79.54613, 
    71.48424, 45.66077, 2.469692, 0.9841859, 1.492721, 0.9228254, -0.447767, 
    0.2154918,
  152.5922, 134.033, 115.3111, 95.84639, 85.08085, 71.62435, 56.33461, 
    46.95739, 5.874403, 3.73544, 8.057158, 1.174014, 0.7223753, 0.7775673, 
    -0.1122638,
  15.87134, 18.76693, 8.131706, 8.242081, 3.347142, 0.6719509, 2.564712, 
    1.420087, 7.469917, 2.131357, 0.1379902, 1.462156, 0.6622924, 0.407781, 
    0.01095961,
  61.58652, 40.36055, 36.06594, 13.7854, 3.197062, -1.009471, 0.242777, 
    0.3142565, 0.8181628, 6.600163, 0.4639015, 2.737119, 5.284531, 0.388549, 
    -0.1621939,
  114.4022, 71.91082, 66.90151, 27.19086, 22.72086, -0.8458874, -0.7628998, 
    0.245169, 1.534502, 2.81328, 2.833883, 2.183099, 3.269195, 3.670285, 
    0.5326001,
  144.7977, 125.3666, 107.7047, 70.9413, 54.74907, 26.07757, 0.8888339, 
    -1.084572, 0.9244533, 1.857922, 1.553599, 1.339986, 1.626328, 1.804221, 
    0.5858628,
  150.7523, 132.5568, 112.3114, 97.93046, 79.83254, 58.59063, 36.56096, 
    0.7614123, -1.642516, -0.1647211, 1.161354, 1.977741, 1.037422, 
    0.7029938, 1.329924,
  161.7714, 139.1353, 114.0029, 98.62347, 91.32633, 82.46001, 67.61968, 
    40.37791, 13.98211, 9.887424, 0.6553971, 2.058656, 2.246067, 0.9230723, 
    2.053214,
  177.8549, 153.09, 121.7386, 101.3309, 91.36643, 87.53484, 85.46003, 
    74.94579, 50.33876, 19.64761, 5.294463, 3.060111, 2.522828, 1.587924, 
    0.8527647,
  189.5227, 155.9552, 124.6182, 103.8313, 91.05861, 85.92097, 80.11664, 
    79.29354, 39.04864, 10.95281, 4.532603, 2.362721, 2.75802, 1.687791, 
    2.593197,
  184.7265, 157.3777, 137.3161, 106.1584, 88.28087, 79.49378, 74.92304, 
    66.16909, 35.10575, 3.628879, 3.096787, 4.341189, 2.096451, 1.533079, 
    4.770424,
  164.3042, 139.0993, 116.9511, 94.88786, 80.84007, 68.55215, 52.82988, 
    42.53783, 4.156323, 2.425681, 8.466454, 2.578623, 1.914096, 0.9313082, 
    4.20955,
  6.918462, 11.30589, 4.783022, 8.69015, 4.768448, 1.038756, 2.790328, 
    2.589309, 5.931563, 1.362358, 0.01560024, 0.5925379, 0.2112717, 
    0.7091407, -0.5106096,
  33.27906, 24.22874, 23.6187, 12.52046, 3.160642, -0.2595853, 1.336006, 
    1.877489, 2.086587, 5.29507, 1.073556, 2.557749, 4.674639, 0.211956, 
    -0.3366299,
  66.98876, 44.38277, 48.4646, 23.19744, 20.2512, -0.08458579, 0.0195942, 
    1.80874, 2.512485, 3.583096, 3.728193, 2.05739, 2.469242, 2.492198, 
    0.5137846,
  81.02215, 71.12636, 64.85213, 49.43845, 42.07266, 23.68692, 0.9287721, 
    -0.03818915, 1.402941, 1.427831, 0.9624852, 0.3414597, 0.6625904, 
    1.626881, 1.63386,
  80.31509, 66.34386, 56.23251, 55.61992, 53.63073, 43.01221, 36.50462, 
    1.089334, -0.3449547, 0.0481331, 0.1600429, -0.02580942, 0.07104061, 
    2.055907, 1.797926,
  84.46951, 68.27753, 58.98163, 57.04462, 58.12016, 58.02185, 46.09645, 
    27.17335, 11.92252, 6.886523, 1.102544, 0.9043821, 2.054952, 1.63114, 
    1.199638,
  97.10349, 83.99274, 72.23737, 66.48504, 65.54422, 64.80518, 63.54066, 
    56.14337, 36.10329, 16.47599, 7.805425, 2.817779, 3.149524, 1.727736, 
    0.4304023,
  111.714, 94.03904, 83.57626, 77.36305, 72.64751, 72.5695, 69.74502, 
    70.58344, 31.25874, 12.88601, 7.05876, 6.251244, 3.722001, 2.951324, 
    3.671376,
  118.7129, 105.0685, 101.132, 86.33358, 77.4146, 74.11215, 73.00768, 
    63.03328, 36.00825, 12.99251, 9.210077, 8.12495, 4.353728, 1.092728, 
    3.167009,
  116.1531, 102.1497, 95.80022, 82.74215, 78.20937, 64.57455, 51.88446, 
    43.58713, 16.92286, 8.909548, 14.94246, 4.641979, 3.18861, 1.091094, 
    5.082088,
  6.866405, 12.11227, 7.440466, 7.557224, 4.192243, 1.041064, 2.527581, 
    3.49837, 9.989483, 4.059295, 0.7319483, 1.412251, 0.00743485, 0.5891928, 
    -0.5462293,
  33.39428, 25.84284, 23.35131, 12.64, 3.152363, 0.03681581, 1.838713, 
    2.42672, 2.962511, 9.301719, 1.132095, 4.568504, 8.271872, 0.6829286, 
    -0.6231328,
  74.53683, 49.05962, 54.76242, 26.08775, 20.35403, -0.4757505, 0.609773, 
    2.37357, 3.543193, 4.735531, 5.736291, 3.236716, 5.324316, 6.268993, 
    1.075771,
  86.70895, 83.66671, 84.12639, 61.58627, 51.69527, 24.59933, 0.464794, 
    -0.2430109, 1.850308, 1.817282, 0.9601849, 0.8730577, 2.616858, 4.156607, 
    2.992189,
  80.39858, 77.28609, 79.4409, 82.1995, 72.66193, 55.49557, 42.76293, 
    1.217695, -0.2517184, 0.1942339, 0.9318044, 1.030453, 1.55189, 3.018736, 
    2.421076,
  74.72267, 70.36242, 69.028, 70.83138, 71.21909, 67.92098, 48.08621, 
    24.21361, 12.97038, 12.0619, 1.496627, 2.336644, 3.127031, 1.366861, 
    1.327822,
  70.14317, 70.26904, 65.92292, 64.57822, 63.61613, 65.46491, 59.46345, 
    44.84966, 30.92755, 14.32806, 8.216029, 4.576352, 3.724916, 0.2453773, 
    0.4877162,
  68.01521, 69.17648, 65.38541, 63.42719, 59.53327, 61.70404, 57.48721, 
    58.38144, 26.24035, 11.09135, 7.315159, 5.867043, 3.843086, 1.832813, 
    2.370294,
  72.47325, 72.38429, 73.85424, 65.43279, 59.07335, 57.65696, 55.32922, 
    48.44593, 25.63393, 9.270832, 6.72471, 6.658771, 4.758523, 1.899341, 
    4.302763,
  76.81453, 69.99756, 66.92525, 59.07172, 55.8156, 45.4808, 41.87849, 
    41.00342, 18.69978, 11.42786, 13.04423, 5.782802, 1.541925, 0.8644131, 
    3.986528,
  6.388035, 8.90411, 4.962897, 4.139628, 1.943253, 1.350938, 3.135601, 
    4.140835, 7.17861, 2.240658, 0.709874, 2.173063, 0.8170034, 0.09931247, 
    -0.5647999,
  25.75513, 19.19607, 14.94981, 6.481943, 1.980212, 0.2751198, 2.613648, 
    4.42171, 3.64321, 5.947108, 1.086976, 4.270164, 7.530069, -0.02620844, 
    -1.133828,
  68.41074, 40.94712, 39.49126, 17.41117, 16.62776, -0.0742311, 1.041465, 
    4.233152, 4.297518, 3.995972, 5.500649, 4.027871, 5.123505, 8.494543, 
    1.807762,
  84.04762, 68.12806, 60.70402, 45.54222, 46.05194, 24.82908, -0.3182441, 
    0.3090553, 0.4179733, 0.8659896, 1.156277, 1.057529, 2.291552, 3.354586, 
    5.267365,
  79.82899, 62.36317, 55.444, 60.55046, 70.627, 62.06534, 49.56425, 
    0.7589381, -0.6031016, -0.1922876, 0.5572335, 0.8089683, 1.144537, 
    2.498991, 3.236842,
  82.05742, 60.95105, 50.19255, 53.02166, 69.75645, 74.07005, 55.64823, 
    29.89597, 15.72624, 17.33043, 3.082911, 2.042516, 0.9659197, 0.7868986, 
    1.45302,
  90.76971, 68.03381, 51.27436, 51.53168, 60.48287, 71.09749, 68.1192, 
    48.22852, 29.40718, 16.00048, 9.578324, 3.637832, 1.315687, 0.1304238, 
    0.3802457,
  94.19666, 70.73887, 55.31953, 51.98014, 54.12405, 60.81882, 60.51667, 
    61.67469, 25.23521, 10.39421, 6.610447, 3.282655, 1.285171, 0.1427898, 
    0.3759757,
  88.18517, 76.79643, 67.95038, 55.78798, 50.40701, 50.52664, 51.24622, 
    46.14695, 18.48466, 6.013133, 4.631451, 3.451361, 1.142103, 0.4416799, 
    2.017945,
  68.82475, 65.08752, 58.61722, 49.71735, 44.45569, 35.97164, 37.32862, 
    37.18366, 11.6181, 11.69871, 12.59933, 3.654423, 1.814511, 1.480222, 
    2.239727,
  4.388189, 5.709753, 3.275817, 4.545206, 4.005537, 1.692399, 1.695522, 
    1.977994, 7.584723, 3.321341, 1.320626, 2.62773, 0.5780239, -0.2434583, 
    -0.6588875,
  19.54116, 15.21366, 9.333258, 4.051891, 1.564445, 0.3647751, 2.50382, 
    2.529792, 5.16563, 10.08803, 3.865289, 5.933836, 8.623833, 0.0781113, 
    -0.882863,
  63.86889, 43.11731, 35.07822, 13.29846, 9.447755, 0.3447632, 0.4391579, 
    2.552718, 5.004588, 8.020439, 8.178792, 4.06084, 4.826558, 9.230638, 
    2.609009,
  91.56107, 79.43638, 66.25795, 42.07096, 34.76308, 17.58269, 1.161399, 
    0.8782402, 2.99053, 3.620505, 2.558389, 0.2890934, 1.1295, 3.316309, 
    6.546983,
  96.24668, 84.19604, 75.2868, 65.51451, 57.80898, 46.41997, 43.7305, 
    2.139687, -0.2280078, 0.4420246, 0.60956, 0.1849463, 0.5101025, 2.600175, 
    4.471726,
  101.8371, 87.89344, 80.18446, 69.64695, 62.5693, 57.87349, 47.34915, 
    27.69484, 16.69691, 19.65109, 4.726748, 1.25349, 0.4518113, 0.5157449, 
    0.7601919,
  108.7448, 93.66865, 79.57963, 67.82495, 62.03089, 62.24409, 60.34958, 
    42.26848, 30.03499, 15.57199, 9.226762, 2.728594, 0.8791099, -0.1059055, 
    -0.03699078,
  105.755, 82.97324, 69.71866, 61.26823, 58.04163, 62.13078, 63.22522, 
    65.12022, 27.13642, 7.506483, 3.423671, 2.166056, 0.8241341, -0.2111501, 
    -0.3894435,
  91.98398, 70.78197, 59.30465, 50.15725, 49.13982, 53.82518, 58.84792, 
    48.13334, 10.7264, 2.146027, 0.9437912, 1.831651, 0.7519641, 0.1378007, 
    0.7936348,
  70.52986, 51.20567, 36.87776, 31.63184, 34.71836, 36.86619, 39.20161, 
    29.62205, 4.867118, 6.938465, 13.6, 3.359471, 1.96418, 1.880352, 1.297778,
  4.044114, 6.816444, 2.591328, 3.341135, 2.977991, 1.061741, 1.683389, 
    2.072923, 5.544252, 1.414718, 0.1695678, 2.416718, 1.508582, 0.03083469, 
    -0.2535711,
  20.78418, 17.72585, 9.642958, 3.396045, 1.480908, 0.2798037, 0.3274716, 
    1.322605, 2.812196, 4.997379, 1.637199, 5.17753, 7.512562, 0.1208669, 
    -0.326828,
  80.41451, 58.03146, 42.65614, 14.10658, 8.784615, -0.1013111, 0.2998252, 
    0.1962056, 1.633297, 3.477793, 4.650483, 4.02741, 4.53861, 5.023382, 
    1.809947,
  129.2487, 109.3778, 91.0023, 57.75541, 37.91636, 15.55416, 0.5197056, 
    0.3381503, 2.200316, 1.086949, 0.6325354, 0.5314354, 0.844766, 3.603487, 
    4.797509,
  142.2511, 117.7249, 100.3143, 85.74317, 71.43305, 41.65548, 43.24298, 
    1.176609, -1.221175, 0.3158872, 0.4032465, 0.4754507, 0.4596883, 
    2.188372, 4.132111,
  154.6587, 127.9421, 108.6336, 89.15532, 73.53083, 50.48246, 48.82312, 
    34.62307, 17.03575, 17.83146, 7.612364, 2.495625, 0.617137, 0.4563054, 
    0.8530292,
  168.7473, 146.8099, 117.9049, 91.71568, 74.40262, 52.22624, 48.55627, 
    38.5601, 29.69434, 16.53453, 10.13646, 2.450294, 1.074703, 0.204908, 
    0.3505172,
  174.245, 144.4797, 116.1113, 92.47206, 73.87418, 58.18258, 43.51696, 
    48.29106, 25.47779, 5.600669, 2.412003, 1.579889, 0.6247523, -0.1213053, 
    -0.2287036,
  161.0893, 135.01, 117.8717, 89.03242, 69.99001, 52.90858, 41.89174, 
    30.9488, 3.421309, -0.4220638, 1.124134, 2.172003, 0.5699536, 0.04365128, 
    0.1990537,
  128.4202, 106.845, 87.41223, 65.43203, 52.7134, 31.5861, 18.62258, 
    12.98102, 0.8293166, 4.063568, 14.12666, 5.07519, 1.920794, 2.749535, 
    0.9467462,
  14.55886, 16.60509, 10.59774, 8.299086, 3.463044, 1.173187, 3.684113, 
    2.849663, 4.408836, 0.8552094, 0.439912, 1.152976, 0.3831888, 0.1364698, 
    -0.1279447,
  26.49326, 28.49026, 22.98479, 13.21264, 2.421565, -0.03705001, 1.410222, 
    1.184445, 2.380005, 3.463023, 0.9818017, 3.768773, 4.403581, 0.08725008, 
    -0.1738581,
  78.56872, 81.49058, 61.45955, 31.7697, 13.58117, -1.288976, 0.1987442, 
    0.4304881, 1.365633, 2.810546, 3.299643, 2.245838, 2.784974, 3.399297, 
    1.216147,
  135.2973, 143.6265, 144.2414, 105.165, 70.1602, 22.22945, -0.2664168, 
    0.1321648, 0.4227335, 0.7584792, 0.7588061, 0.5889272, 1.575834, 
    2.631922, 3.176378,
  134.873, 144.8641, 152.7446, 153.5213, 136.9306, 87.12828, 55.70242, 
    0.7168612, -1.026034, -0.02191875, 1.047182, 1.299143, 0.5948645, 
    2.10823, 3.098607,
  137.0857, 146.1478, 153.0368, 149.6087, 140.7331, 119.0614, 87.04352, 
    39.554, 13.56976, 14.00337, 10.31241, 3.716467, 0.5048596, 0.1646888, 
    0.1363548,
  141.2507, 158.7949, 156.6927, 146.0507, 135.9337, 117.5361, 96.63229, 
    50.94432, 28.03129, 13.27633, 10.55942, 2.286835, 0.8982582, -0.03143292, 
    -0.247006,
  134.7119, 148.5623, 154.1508, 146.1526, 131.8513, 115.1963, 88.50205, 
    70.79274, 27.83645, 8.05227, 2.678135, 1.586658, 0.5943199, -0.5030316, 
    -0.5328822,
  120.2707, 139.0359, 157.8953, 145.3652, 126.6838, 102.7665, 81.90085, 
    47.70535, 2.819022, 1.151671, 4.035663, 5.124688, 1.126728, -0.3183497, 
    -0.6377057,
  92.88868, 108.1187, 125.096, 117.2876, 105.6353, 72.67341, 49.33298, 
    17.38741, -1.125652, 0.996522, 12.10302, 9.217152, 6.228098, 3.211774, 
    0.1747036,
  9.359711, 11.05099, 14.00344, 10.5895, 3.771117, 1.77404, 5.003469, 
    2.803015, 4.071799, 0.619143, 0.2035917, 1.676034, 0.3604806, 0.133038, 
    -0.2233906,
  10.08576, 15.52411, 20.85332, 11.63595, 1.791251, 0.366443, 1.063257, 
    0.8512682, 2.032284, 3.295501, 0.9763303, 4.263405, 4.514638, 
    -0.02770502, -0.2838835,
  27.45222, 33.79779, 36.80569, 26.45945, 18.28937, -1.29635, -0.1167192, 
    0.5073723, 1.142544, 3.044527, 3.05782, 3.302544, 4.033011, 3.136504, 
    1.280124,
  54.04808, 63.13784, 96.67687, 94.26723, 63.16162, 27.40109, -0.2738751, 
    -0.2678546, 0.2802677, 1.444661, 0.8855215, 1.124036, 1.943436, 2.809242, 
    2.706087,
  54.14397, 58.71478, 101.7011, 149.0736, 146.1932, 94.85861, 65.01464, 
    0.7948853, -1.268608, -0.003814073, 1.295211, 1.52725, 0.7339991, 
    2.02069, 2.959548,
  59.96632, 59.48887, 91.94228, 137.4881, 156.2213, 147.4291, 104.8511, 
    44.02245, 13.96584, 16.0402, 10.10425, 4.404938, 0.6095792, 0.625601, 
    1.09404,
  68.47215, 67.17393, 87.24362, 126.3329, 141.8921, 142.9786, 130.2811, 
    62.18128, 27.39512, 15.2422, 11.70349, 2.592869, 0.9247746, 0.1183376, 
    0.3746546,
  70.18999, 62.10947, 80.71021, 116.2985, 132.4234, 132.093, 122.0757, 
    105.5466, 43.6262, 4.821988, 2.290868, 1.479908, 0.8221701, -0.3191255, 
    -0.04507909,
  61.83972, 56.03202, 81.89761, 111.8281, 122.4777, 116.9855, 109.4424, 
    86.3607, 11.37132, 0.471317, 0.8673828, 2.235812, 0.7680944, -0.2824779, 
    -0.4952983,
  44.54456, 41.33125, 61.87999, 88.78664, 100.3192, 89.33984, 73.04132, 
    33.68549, 2.164055, 3.817274, 16.62353, 7.678683, 4.073222, 1.24646, 
    -0.0002392718,
  5.404897, 8.487907, 5.315319, 3.563461, 1.646193, 1.098958, 5.541072, 
    3.471275, 4.955183, 1.044714, 0.4324035, 2.138086, 0.780611, 0.283708, 
    -0.2702653,
  2.165627, 5.983566, 5.533259, 5.268647, 1.904035, 0.2359195, 0.9517161, 
    0.904033, 3.216601, 4.088559, 2.021407, 4.880505, 5.170397, 0.03081079, 
    -0.2668653,
  28.74813, 12.01199, 9.783665, 15.8192, 16.8573, -0.8991542, -0.09182227, 
    0.6437547, 2.458055, 3.561493, 4.113936, 3.946652, 3.973447, 3.729563, 
    1.245814,
  57.22603, 34.88296, 35.326, 53.30899, 55.37593, 28.28452, -0.4980192, 
    -0.2021589, 0.7558404, 1.751584, 1.730412, 2.146008, 2.379544, 3.019785, 
    3.068314,
  61.75705, 36.32748, 37.17508, 91.89911, 102.0839, 75.94101, 63.94812, 
    0.8292408, -1.112996, -0.07514083, 1.141065, 2.542381, 2.134119, 
    3.033406, 3.448534,
  61.31998, 42.05828, 34.56693, 79.24259, 124.8896, 121.8721, 94.26723, 
    43.29134, 15.02395, 20.31949, 10.61833, 4.887038, 2.670412, 1.887479, 
    1.664036,
  53.62528, 46.00749, 33.22266, 66.66516, 111.9665, 120.4312, 113.5221, 
    51.59859, 24.31259, 20.89156, 14.1416, 4.166949, 2.818989, 1.22363, 
    1.358363,
  47.03439, 42.46827, 30.6738, 62.27616, 106.1074, 116.4902, 115.2927, 
    97.83349, 38.53641, 8.164229, 4.771861, 2.842199, 1.926087, 0.6547892, 
    0.8034915,
  43.93756, 46.09156, 33.86147, 63.88824, 102.002, 105.5986, 110.8208, 
    91.49403, 15.72137, 1.342314, 1.455084, 2.57056, 1.628764, 0.3454459, 
    0.2870009,
  41.35513, 33.95655, 25.20681, 60.30651, 88.57633, 87.41327, 75.60003, 
    34.6511, 1.738208, 3.908272, 16.47932, 5.951554, 3.472338, 2.074309, 
    0.9644018,
  12.34895, 23.72948, 16.95962, 9.878695, 0.6679932, -1.05396, 2.872085, 
    3.445674, 6.585554, 1.205214, 0.07100741, 2.049047, 0.6086206, 0.2973502, 
    -0.1855525,
  20.05295, 23.57977, 18.97778, 8.325895, -0.8929101, -1.323132, 0.3703938, 
    0.8752767, 3.970492, 4.943547, 1.950812, 4.722537, 4.736569, 0.188696, 
    -0.09056067,
  59.01222, 46.62051, 28.9908, 13.2154, 9.575144, 0.7798293, 0.1197056, 
    0.5853129, 2.342686, 3.842464, 4.182871, 3.663407, 3.381278, 2.997191, 
    1.115695,
  77.25736, 73.01712, 67.31779, 43.44421, 38.577, 28.41826, 1.600067, 
    -0.198049, 0.6989279, 1.589285, 1.73758, 1.994432, 2.084929, 2.555553, 
    2.66598,
  68.50197, 62.60684, 63.49672, 68.01614, 58.40202, 60.09602, 55.62456, 
    1.763298, -1.260073, -0.1724547, 1.051453, 2.424623, 2.254079, 2.611152, 
    2.619644,
  47.61856, 49.89893, 54.11147, 61.52852, 86.07258, 92.47985, 70.46204, 
    34.0975, 15.2597, 24.30936, 11.69364, 5.142875, 3.357468, 1.819349, 
    1.370107,
  33.54693, 38.50911, 45.90456, 53.47615, 80.75874, 95.82201, 77.83356, 
    33.64388, 19.63742, 28.40892, 16.5892, 5.519827, 3.795207, 1.556324, 
    1.043219,
  47.08414, 37.4615, 43.01911, 54.21694, 81.76984, 96.63639, 92.35482, 
    80.64072, 30.20992, 7.724949, 5.027131, 3.886546, 2.997612, 1.176997, 
    0.6731918,
  62.57632, 51.70843, 56.54266, 67.57208, 88.67961, 88.04257, 93.71989, 
    87.59763, 13.80927, 1.830784, 1.726526, 3.143086, 2.285978, 0.9743386, 
    0.314999,
  55.88556, 48.05275, 56.46151, 67.78201, 82.72865, 83.65289, 75.49938, 
    33.98481, 2.896862, 4.038934, 15.02788, 5.033606, 4.224604, 2.806138, 
    1.725357,
  11.38116, 24.2413, 15.36138, 11.34831, 4.402399, 1.915132, 4.670912, 
    -0.1791007, 2.046124, 0.4612974, 0.4832015, 2.467858, 0.6645582, 
    0.2374889, -0.2195697,
  18.89774, 13.70928, 11.51379, 6.917161, 0.4816031, -0.4234578, -0.9065337, 
    -1.571236, 0.4073871, 4.412258, 2.658629, 5.448883, 4.732843, -0.0682177, 
    -0.3144331,
  43.90399, 31.6975, 21.27318, 5.178652, 2.873506, -3.031407, -1.370559, 
    -0.06736714, 0.136452, 3.523693, 5.180663, 3.91813, 3.101057, 1.931496, 
    0.5061494,
  53.45724, 54.36798, 55.24842, 41.37078, 29.14405, 18.07778, 0.2433975, 
    -0.8256311, 0.348949, 1.490141, 1.860195, 0.939934, 1.002515, 1.17886, 
    0.6895242,
  48.56254, 42.59452, 50.04825, 66.57832, 49.18287, 46.43287, 41.32749, 
    -0.07078708, -1.023355, -0.02950838, 0.7139902, 0.9331197, 0.7702572, 
    0.9060776, 0.7420447,
  44.89578, 34.49855, 40.97416, 63.76461, 88.18393, 77.77001, 53.47974, 
    28.28688, 15.70396, 24.32817, 13.61855, 4.163005, 1.936447, 0.5139781, 
    0.3514528,
  42.09401, 31.71765, 39.11277, 64.08595, 86.96937, 86.42196, 69.01888, 
    28.08468, 19.93396, 32.91476, 20.97504, 5.107639, 2.478744, 0.4627276, 
    0.1288947,
  47.49926, 35.60483, 48.46841, 74.52361, 82.31356, 85.63415, 76.26558, 
    60.30485, 22.56143, 6.502588, 3.668226, 3.434296, 1.907518, 0.4140908, 
    0.1137049,
  93.53347, 76.49297, 82.31866, 83.79047, 81.98648, 73.93304, 70.71094, 
    64.18654, 6.811677, 1.257604, 0.5246304, 2.696961, 1.779478, 0.7065251, 
    0.3333307,
  126.4319, 102.3365, 92.29211, 81.84277, 74.89867, 72.86861, 61.74554, 
    34.00574, 3.976048, 3.192465, 12.78266, 4.624208, 3.494203, 2.15305, 
    1.460148,
  13.83617, 25.94479, 19.25668, 16.78261, 7.600307, 6.853483, 11.80828, 
    5.844065, 3.142127, -2.357169, -0.9584278, 1.924985, 0.5590072, 
    0.3432139, -0.6671764,
  20.67979, 10.02046, 10.1259, 6.128447, -1.134687, 0.3003163, 1.557444, 
    -0.5843254, -0.7728994, -0.1459848, 0.1090207, 5.840993, 6.294119, 
    -0.6658747, -0.6942703,
  38.06145, 27.02188, 17.53258, 4.754651, 2.821937, -3.121923, -0.5931786, 
    -1.08818, -1.89172, -1.090536, 1.589399, 2.762485, 3.219573, 4.384929, 
    1.535175,
  43.91561, 38.84271, 34.69165, 19.15962, 14.24852, 14.366, -2.349682, 
    -0.8828033, -0.6170915, -0.8806016, -0.5449321, 0.7699458, 2.292385, 
    2.923526, 2.905548,
  57.08944, 35.02924, 26.62428, 25.58481, 18.04945, 28.24698, 25.68878, 
    1.846705, -1.411829, -0.3384869, -0.02351947, 1.657039, 2.643474, 
    3.316209, 3.050165,
  73.70503, 43.84743, 25.02929, 16.33171, 25.57077, 41.20292, 34.36587, 
    20.12507, 10.9604, 17.85535, 10.21513, 4.181758, 3.402912, 1.695614, 
    0.7198355,
  100.7815, 87.64117, 44.47017, 30.37009, 48.13451, 63.54127, 53.92683, 
    21.61746, 13.77804, 27.35834, 19.08873, 6.432719, 3.403971, 1.154366, 
    0.3013713,
  105.9972, 108.571, 97.47346, 84.28847, 82.19557, 79.1996, 71.38497, 
    54.7188, 15.30219, 4.022578, 5.030489, 4.147271, 2.313595, 0.5010047, 
    0.2007132,
  101.7465, 98.67638, 97.25077, 89.6267, 80.46864, 70.81818, 71.21621, 
    57.75574, 5.631276, 0.5062013, 1.697488, 2.280216, 1.280911, 0.2912831, 
    0.4232097,
  99.90714, 92.38465, 88.55293, 80.25062, 71.60961, 66.25438, 58.67944, 
    30.72969, 3.482317, 2.098287, 9.653114, 2.874056, 2.191787, 0.7981873, 
    1.071755,
  5.183647, 12.72801, 8.686093, 10.1685, 3.876512, 6.888312, 12.94714, 
    4.864653, 1.492113, -1.173732, -0.2964106, 2.256327, 0.2866695, 
    -0.06687397, -0.8869894,
  10.38618, 9.655508, 7.722704, 5.324511, 0.1497669, 5.126477, 5.931157, 
    1.15372, -0.2251447, 0.2862049, 2.173511, 6.889573, 5.426901, -1.171602, 
    -0.8501444,
  34.01496, 21.46774, 13.81747, 8.756476, 3.708832, -1.433366, 2.281929, 
    1.506517, -0.01103867, 0.5946547, 3.762893, 4.186195, 3.61023, 2.919265, 
    0.7757559,
  59.25295, 57.30571, 47.73619, 24.98057, 10.69937, 11.73436, -1.497935, 
    -0.4029495, -0.3808522, -0.005865283, 0.56893, 1.124302, 0.8598834, 
    1.255444, 3.409332,
  67.47971, 63.59373, 57.71818, 38.94672, 20.31402, 22.34825, 24.44481, 
    1.744249, -1.487697, 0.1535186, 1.098534, 1.144915, 0.7355295, 0.9820973, 
    4.21455,
  72.46187, 77.00417, 71.57227, 59.30402, 40.34632, 29.67512, 26.67362, 
    15.71203, 9.735662, 14.79052, 11.2427, 3.990831, 1.73896, 0.2594633, 
    0.7509582,
  69.20894, 90.30524, 87.58894, 81.16476, 76.23361, 63.34146, 45.4051, 
    13.42008, 6.573867, 17.60049, 16.52743, 5.058398, 2.899371, 1.092824, 
    1.744892,
  62.21234, 79.46809, 83.87737, 82.89995, 82.15086, 78.98485, 68.93133, 
    44.04487, 5.798854, 0.8609774, 2.676554, 2.592448, 3.143722, 1.448665, 
    1.256547,
  65.25019, 72.8667, 82.04556, 81.97169, 79.0891, 71.77863, 71.31044, 
    45.6724, 3.593518, -0.1287052, 0.7006037, 2.481032, 3.360813, 2.274962, 
    1.153378,
  67.74423, 65.95383, 71.81374, 74.01299, 69.66163, 63.60931, 54.18094, 
    26.35069, 3.064302, 1.391166, 7.916646, 4.329821, 5.401638, 4.175929, 
    2.736255,
  3.899038, 9.17772, 5.761263, 10.69158, 5.396436, 2.727552, 6.928013, 
    4.602211, 2.988006, -0.466958, 0.7963279, 3.504035, 0.6924875, 0.6660094, 
    -0.7557452,
  6.648255, 4.342385, 3.847083, 8.34293, 2.646766, 2.873374, 3.380169, 
    2.613879, 2.168083, 2.553164, 4.972426, 8.102619, 5.963445, -0.5647514, 
    -0.5868906,
  21.8222, 29.47264, 13.2507, 6.05553, 5.407341, -0.8542578, 1.344201, 
    2.160426, 1.303005, 1.840725, 6.362077, 6.336686, 3.803827, 3.366808, 
    0.938206,
  28.06132, 48.28136, 62.04911, 47.35456, 13.3193, 5.798284, -0.5296165, 
    0.47923, 1.74609, 0.423499, 1.432031, 2.501482, 2.476824, 3.858428, 
    4.148554,
  30.17177, 41.24666, 59.73441, 69.56509, 50.51907, 36.43223, 15.33461, 
    0.9014785, -0.1413856, -0.576661, 1.749107, 3.965732, 3.099115, 4.694294, 
    5.985976,
  39.98779, 40.19173, 58.15473, 67.97734, 70.54916, 63.42082, 37.28935, 
    17.73143, 7.190026, 8.761929, 7.479939, 5.152677, 5.589265, 2.816618, 
    3.101128,
  55.38453, 47.78082, 59.24928, 63.34394, 66.35192, 65.34595, 56.4798, 
    24.27891, 11.88127, 9.442648, 9.255536, 5.569592, 5.259742, 2.562783, 
    2.776191,
  60.92366, 53.31963, 59.89239, 59.1121, 61.85505, 61.14209, 54.43132, 
    35.17119, 7.457906, 0.8870412, 2.513535, 4.53313, 4.983537, 1.494376, 
    1.680545,
  57.949, 61.08184, 66.79913, 58.33969, 57.82745, 50.78621, 46.76939, 
    29.76441, 3.134448, 0.5116138, 0.888831, 3.313326, 2.363811, 2.065266, 
    2.766559,
  55.48414, 62.52527, 59.02903, 51.84928, 48.92208, 43.27856, 29.23684, 
    15.44535, 2.867059, 1.467955, 3.276219, 3.920672, 5.080344, 5.743951, 
    5.568815,
  2.435209, 1.499518, 1.040914, 0.1595782, -0.6345119, -0.1744883, 4.714468, 
    2.097344, -0.5553514, -3.053376, -0.8289124, 0.7122684, -0.2814075, 
    0.1930377, -0.3476243,
  7.351909, 0.7018722, -0.3369588, -1.406151, -3.136816, 0.3074705, 1.527739, 
    0.7096329, -0.3100904, -1.927197, -0.3944449, 3.159023, 2.988323, 
    -1.052958, -0.7505062,
  38.8214, 28.67903, 11.87147, 0.3597491, -3.368663, -5.513414, -0.8082934, 
    0.4221407, 0.01756535, -0.7601136, 0.7804992, 2.291548, 1.213281, 
    1.151809, 0.2293782,
  46.81808, 49.40308, 59.82494, 46.18501, 14.11111, 3.17097, -3.300416, 
    -2.180513, -0.291216, 0.05891332, -0.1590987, 1.193045, 1.355539, 
    1.600671, 2.564805,
  50.18024, 51.86064, 59.28167, 64.73302, 46.61271, 30.5472, 11.04847, 
    -2.364887, -1.482873, -0.0430776, 0.6779694, 1.624109, 0.8505027, 
    1.967148, 3.485492,
  67.96906, 66.32769, 66.3128, 62.36168, 57.80955, 42.6006, 20.14351, 
    6.021194, 2.219466, 7.117272, 3.906554, 1.720248, 1.953739, 1.337427, 
    1.296786,
  81.14077, 78.29267, 70.48584, 59.35223, 49.11701, 43.47285, 41.67857, 
    6.770081, 2.684553, 10.10499, 3.368714, 1.492151, 1.985837, 1.747409, 
    1.830149,
  74.66233, 77.99712, 66.54198, 59.14003, 44.80952, 46.12711, 48.17435, 
    18.71973, 3.146075, 3.153499, 1.324597, 1.025485, 2.157059, 0.9869643, 
    1.029231,
  70.4637, 71.6287, 70.24158, 64.60006, 42.98298, 40.32517, 50.24158, 
    16.34215, 1.929987, 2.138925, 0.9733394, 1.156568, 0.9525593, 1.544628, 
    2.055114,
  50.54245, 43.58863, 50.13107, 55.59089, 37.90025, 37.1836, 35.79466, 
    5.233744, 2.345862, 2.293691, 2.437469, 1.531, 2.962146, 4.640205, 
    5.039995,
  1.75976, 3.15207, 1.780996, 1.254351, -0.3531309, 2.040078, 5.921021, 
    2.892453, 2.817059, -0.08675341, 2.39088, 2.067647, -1.31549, -1.379833, 
    -2.514129,
  6.828779, 2.569663, -0.01877049, -0.2749247, -0.9954996, 4.956987, 
    4.286738, 1.911723, 2.084765, 1.845596, 1.472567, 4.168598, 2.925955, 
    -1.801167, -2.370799,
  22.09287, 26.90104, 16.68692, 4.62763, 0.3800509, -0.481227, 5.099034, 
    4.145948, 4.785136, 1.539754, 2.123123, 7.245882, 6.949527, 7.09549, 
    2.427346,
  36.52017, 40.43914, 41.96263, 40.81761, 14.52163, 2.005637, -1.341529, 
    0.4519238, 3.674053, 4.459483, 3.742679, 4.563221, 7.430385, 7.506978, 
    5.315083,
  46.24939, 30.52752, 36.21714, 50.60452, 49.1669, 44.41604, 7.026293, 
    -2.319753, 1.972545, 1.429634, 3.485823, 3.486864, 4.50065, 6.087221, 
    4.820377,
  43.73701, 26.2527, 33.95047, 49.89194, 55.91448, 57.43909, 37.75434, 
    13.5756, 7.994363, 10.57634, 2.664799, 5.344742, 4.739399, 3.622988, 
    2.468236,
  42.55763, 34.03909, 35.60477, 41.23074, 48.81012, 53.76504, 53.67685, 
    15.30097, 8.972592, 11.696, 4.10859, 2.533807, 4.381945, 1.819244, 
    2.087968,
  41.18981, 38.41803, 37.69562, 37.32046, 45.18844, 49.59167, 45.26008, 
    24.16005, 7.220518, 5.642119, 1.815897, 1.421811, 1.076081, 0.2475117, 
    -0.1472333,
  38.96841, 38.51645, 43.5158, 37.28323, 38.00712, 35.44163, 37.24181, 
    18.58155, 3.342819, 2.119658, 1.351051, 0.67397, 0.7215001, 0.1337224, 
    1.071651,
  27.09497, 19.93931, 26.69957, 26.28618, 27.98245, 26.2296, 21.74064, 
    7.966285, 2.512035, 2.541886, 2.717835, 1.352167, 1.186508, 1.822415, 
    2.276566,
  1.813704, 3.233923, 1.42038, 0.8710449, 0.9309641, 1.522079, 3.369287, 
    -0.3714291, 1.860776, -0.7279969, 0.3405536, 2.48272, -0.5630535, 
    -0.4231899, -0.9576259,
  12.94027, 3.282207, 0.8623229, 0.7945129, -0.2858466, 1.443991, 1.016557, 
    -0.903657, 1.595984, 0.8944393, 1.426157, 3.540465, 4.153048, -1.071944, 
    -0.8471001,
  51.39279, 25.97791, 9.906734, 2.649966, -0.01392651, -2.902716, 3.534369, 
    1.847623, 1.56935, 1.697822, 2.918848, 3.82763, 3.629143, 6.112501, 
    1.769353,
  58.07429, 33.68622, 19.87171, 16.4403, 5.761203, -0.7022638, -2.301128, 
    -1.253146, 1.001728, 1.573573, 2.107579, 4.471217, 3.237418, 3.663099, 
    4.316433,
  56.22093, 23.22289, 16.17121, 21.1525, 23.08997, 13.3852, 4.555724, 
    -2.329021, -1.595542, 0.3280798, 3.322966, 3.84945, 3.262823, 3.145422, 
    7.21811,
  40.84507, 14.47975, 13.82396, 21.88189, 28.8143, 23.5573, 13.53786, 
    5.613025, 3.350636, 1.539751, 3.724298, 3.770087, 1.963499, 2.115255, 
    1.297411,
  40.07626, 25.51195, 17.00105, 12.30455, 29.22553, 26.36129, 27.28509, 
    8.98771, 7.761366, 3.230379, 3.863431, 2.082626, 1.547749, 0.207461, 
    0.07938775,
  38.482, 25.70419, 21.38906, 18.47438, 30.68266, 29.23041, 23.47178, 
    13.91358, 7.671986, 2.767738, 1.346714, 1.806335, 1.637243, 0.5773134, 
    -0.2078891,
  33.09498, 23.80731, 29.43639, 25.79855, 27.27843, 14.7153, 23.428, 
    15.06896, 9.159411, 2.517804, 1.701407, 1.588092, 0.5893769, -0.09988259, 
    0.1385928,
  23.09861, 17.68579, 22.22136, 22.43556, 17.1166, 12.4227, 13.56156, 
    13.12247, 11.40312, 0.9617061, 2.115476, 3.493823, 1.164714, 1.269663, 
    0.7063378,
  6.575338, 6.432883, 5.418181, 4.692688, 1.660913, 0.1987141, 1.532393, 
    0.04169042, 2.956045, 0.6849058, -0.5398725, 1.856838, 0.8340239, 
    -0.441386, -0.8446481,
  16.07882, 8.331029, 6.300362, 3.24943, 0.930096, 2.774775, 3.984691, 
    -2.340515, 0.9000363, 1.61772, -0.03579338, 2.956389, 3.783712, 
    0.07773563, -0.3962367,
  52.99281, 26.65591, 13.87701, 3.79846, 1.563375, 0.3269563, 5.923834, 
    1.454613, -0.3102602, 1.521006, 1.768864, 1.741721, 3.514367, 5.881544, 
    2.999811,
  62.69874, 38.33881, 28.03369, 20.46, 6.055729, 2.429345, -0.4092607, 
    -3.160959, 1.71267, -0.5792942, 1.319132, 2.702005, 1.929079, 3.351481, 
    4.347421,
  60.48857, 30.62448, 22.34435, 20.19608, 15.93394, 15.7582, 3.846551, 
    -0.2937633, 1.235642, -0.6556017, 0.8781714, 1.436438, 1.310595, 
    0.7952416, 1.153039,
  53.34589, 28.20593, 20.6624, 16.92747, 19.54651, 22.50174, 15.35082, 
    4.752454, 2.856608, 2.951216, -1.135097, 0.6584123, 0.617467, 0.1742976, 
    0.2268053,
  49.9691, 30.33211, 22.62495, 17.2753, 24.50376, 26.32432, 27.03874, 
    10.28474, 7.575606, 3.716303, 1.17684, -1.600904, 0.05190624, -0.7273785, 
    -0.7341955,
  48.85194, 35.97629, 29.43616, 25.78283, 29.75191, 28.82881, 20.80861, 
    14.98266, 8.090235, 2.726654, 2.455, -1.458659, -0.3237881, -1.362072, 
    -1.479417,
  51.41874, 42.77354, 35.73101, 24.88937, 19.81708, 20.10754, 16.78421, 
    11.25112, 8.539948, 5.734523, 3.952251, -1.621395, -0.8462371, -1.847281, 
    -1.887854,
  49.38015, 35.07935, 17.52637, 22.75365, 22.56615, 19.73224, 10.14246, 
    3.488858, 9.247434, 2.383208, 3.712861, -0.1987698, -1.064581, -1.870129, 
    -1.166813,
  12.22508, 14.01371, 10.55903, 5.251404, 1.961942, 0.7817435, 1.760427, 
    0.5178299, 3.481184, -1.150722, -1.287246, 0.03928632, -0.5484998, 
    -0.1726217, -0.5957912,
  22.8591, 18.86709, 8.781142, 2.060932, 0.8685549, 1.817579, 2.003814, 
    2.583795, 0.6694894, -0.04367967, -2.227202, 0.3560876, 1.417251, 
    -0.8509544, -1.083931,
  56.15536, 33.5559, 21.87171, 5.928852, 2.422089, -0.2192911, 3.648763, 
    3.257291, 2.126432, -0.1197812, 0.6363172, 1.320962, 1.424607, 1.043934, 
    -0.5362309,
  73.09976, 60.7655, 50.5693, 33.72653, 13.15106, 4.014913, 1.088654, 
    1.484929, 1.56562, -0.4281753, -0.4162622, -0.4136262, 1.540546, 
    1.637417, 0.8682584,
  70.62804, 50.89082, 46.21961, 47.12318, 47.41882, 43.09353, 15.34427, 
    -0.05361024, 3.126911, 0.9477517, 2.840892, 1.602696, -0.2599959, 
    -0.8831921, -0.04135275,
  62.68394, 52.8858, 52.08575, 53.29713, 56.65408, 51.76535, 38.50487, 
    13.44943, 12.30747, 4.600828, 3.165449, 0.143951, -0.7430436, -2.650143, 
    -2.427988,
  64.46273, 63.24615, 60.34185, 51.11412, 52.03843, 49.09736, 43.97701, 
    21.91533, 11.40303, 7.068031, 3.206474, 0.2635052, -0.9757362, -2.471223, 
    -3.879834,
  73.00603, 72.39917, 65.66953, 49.31604, 48.79176, 44.44981, 28.86527, 
    19.41625, 10.63785, 5.86399, 4.034077, -1.551673, -2.871127, -3.733658, 
    -5.410429,
  88.75619, 82.76125, 68.7824, 45.41068, 30.93999, 23.98317, 21.73852, 
    14.20187, 9.373736, 4.282205, 2.621496, 0.001373522, -1.954821, 
    -5.103332, -5.800098,
  81.30153, 61.73955, 45.77644, 23.83769, 16.5107, 10.55713, 13.35587, 
    4.853877, 11.26841, 3.636683, 4.39241, 2.029356, -0.3994178, -2.688092, 
    -3.973614,
  7.850387, 11.39418, 7.551475, 3.677087, -0.2523759, 1.001588, 3.711318, 
    1.513677, 0.3686389, -2.381731, -1.086272, -0.3081718, -3.447302, 
    -2.371452, -3.397798,
  17.96573, 11.11967, 7.434206, 1.170885, -0.1163275, 1.230591, 2.912275, 
    1.821283, 1.013014, -2.29414, -1.237043, 1.198811, -0.7908339, -4.008371, 
    -4.470683,
  41.93896, 24.28555, 19.80186, 5.747272, 2.178439, -1.57813, 4.557709, 
    1.797949, 2.98475, 0.9967035, -1.125303, -0.2281228, 0.4758794, 1.263509, 
    1.400398,
  62.80862, 60.41133, 58.02987, 40.0605, 14.74758, -0.5184395, -3.893912, 
    0.4526912, 4.902908, 4.967141, 2.874815, 3.936849, 4.62953, 4.909822, 
    2.959107,
  72.46993, 57.56159, 53.64738, 53.38183, 52.60046, 44.63266, 16.06561, 
    4.292862, 12.58871, 4.26583, 9.261398, 7.193728, 4.788824, 3.680939, 
    3.898804,
  79.40703, 64.70467, 57.67032, 53.49766, 55.41567, 52.44248, 41.4352, 
    14.55321, 13.82872, 4.393772, 4.877415, 6.192197, 5.312916, 6.176622, 
    5.313393,
  85.20586, 75.07565, 63.12983, 53.10936, 47.90722, 44.51086, 35.27472, 
    17.78139, 8.943485, 4.180688, 7.248631, 7.716616, 7.346115, 7.045784, 
    4.796766,
  78.31598, 72.3533, 61.35637, 47.32912, 40.73555, 34.32608, 16.58623, 
    5.481494, 6.779449, 8.993547, 9.077344, 7.792743, 8.803036, 6.226724, 
    6.893404,
  76.13242, 69.62039, 62.26483, 44.15334, 30.46054, 14.1625, 5.400001, 
    2.342519, 10.14131, 18.0301, 16.22876, 5.938043, 3.734259, 3.13833, 
    4.194368,
  62.9539, 50.96459, 43.68787, 25.42104, 10.20332, 1.009764, -1.208714, 
    1.08524, 12.84785, 5.857971, 25.2241, 13.68259, 5.97333, 3.538811, 
    3.091584,
  9.018078, 10.77715, 11.04554, 7.453901, 1.108978, 2.762038, 7.002882, 
    -0.6503437, -1.536595, -3.019669, -1.575047, 0.2672043, -2.239011, 
    -1.794592, -1.659637,
  16.01173, 14.22042, 9.239686, 4.077148, 0.1600491, 3.734255, 6.592985, 
    -0.3411807, -1.047285, -2.178634, -1.410621, 1.458638, 0.7391939, 
    -1.470661, -1.696468,
  38.19559, 25.00936, 19.6281, 9.585414, 5.089429, 0.593056, 8.044885, 
    3.772893, 0.4452186, -1.372459, -0.3847176, 0.04525021, 1.332554, 
    0.7441847, -1.613763,
  65.522, 60.83107, 59.59883, 43.81694, 22.15567, 7.638948, 1.780224, 
    4.471048, 1.596539, -1.519086, -0.02040853, 0.1594061, 0.3389495, 
    -0.283601, -1.503618,
  80.58009, 63.46978, 59.13079, 57.62725, 54.66072, 45.52105, 21.43842, 
    3.21863, 2.25485, 7.74108, 10.44473, 0.3508781, 0.1155617, 0.6057773, 
    1.741912,
  93.06045, 75.54879, 64.05084, 54.76829, 54.36369, 53.78077, 51.91803, 
    19.56646, 6.483203, 9.267973, 7.886806, 4.487195, 3.643326, 2.014488, 
    0.8005832,
  100.8877, 84.89015, 69.5838, 56.36555, 55.87269, 54.48233, 53.1521, 
    38.5017, 14.98616, 10.22228, 8.225001, 5.512803, 3.412123, 2.139031, 
    0.4484325,
  92.80727, 79.3015, 67.14082, 56.68347, 54.06336, 54.41021, 46.20864, 
    34.42593, 15.0808, 8.200409, 9.315218, 5.654869, 5.737627, 2.600223, 
    1.21774,
  82.32118, 72.36709, 63.74429, 49.27013, 43.56567, 35.58694, 35.3182, 
    25.17199, 13.5621, 16.52664, 19.60349, 9.255196, 3.973143, 1.419564, 
    1.556426,
  61.91172, 48.70434, 42.09173, 31.61938, 23.44073, 21.34387, 23.15768, 
    13.63381, 16.97772, 11.278, 20.98499, 9.986096, 3.764356, 2.033145, 
    0.8272324,
  7.643978, 9.235319, 10.15579, 7.827963, 1.970072, 1.41857, 2.889863, 
    -1.526411, -1.339511, -1.975543, -0.5376485, 1.643853, 0.2351148, 
    -0.4128199, -1.490507,
  10.96478, 9.150533, 8.35072, 4.428903, 0.2530223, 1.844547, 4.181346, 
    -0.9527066, -0.5089256, -0.5451484, 0.5212233, 2.908957, 1.662556, 
    -1.301691, -1.94733,
  43.6748, 25.53168, 14.25606, 6.142734, 1.767628, -2.687583, 4.996476, 
    3.255873, -0.2244196, -0.8003115, 1.232925, 1.437861, 1.547228, 2.7576, 
    0.2869851,
  63.57059, 56.72898, 47.04182, 30.00669, 8.073073, 0.2412503, -1.832915, 
    2.904889, 2.092639, 0.4461304, 0.8298481, 0.5038842, 0.4132968, 
    -0.4811483, 0.1547062,
  65.80724, 47.72176, 38.19818, 29.61188, 22.96041, 13.40199, 5.845812, 
    -0.4594698, 2.019348, 3.454977, 3.365364, -0.4398556, 0.09699421, 
    -0.07197373, 2.092665,
  60.39717, 46.66221, 31.78154, 23.48742, 23.05187, 21.80632, 17.85914, 
    12.8472, 1.897609, -0.3777013, 1.477907, 1.05799, 2.736135, 3.077568, 
    3.471955,
  58.04517, 45.27096, 30.00443, 20.5348, 20.60451, 21.09889, 23.02508, 
    14.44758, -0.9386146, 0.184706, 1.180655, 2.289254, 3.612411, 4.175875, 
    3.650101,
  50.88394, 35.25235, 24.06096, 20.80255, 17.85658, 24.50613, 18.81511, 
    12.82308, 1.956903, 2.434424, 2.15794, 2.362243, 4.532862, 3.73765, 
    3.379681,
  38.24327, 33.11184, 24.81027, 15.46826, 14.33457, 13.03548, 15.89174, 
    8.751036, 8.471144, 13.14837, 19.73645, 5.454602, 2.930194, 2.651608, 
    4.429123,
  26.68371, 16.25958, 13.14424, 9.515829, 8.223699, 11.89366, 8.537031, 
    8.322426, 14.26101, 8.943339, 22.4901, 5.013624, 1.833764, 1.884833, 
    2.46417,
  1.626505, -0.157152, -2.587794, 0.1977393, -2.365137, 0.6808322, 0.4363789, 
    -2.863973, -4.626109, -5.282138, -3.834164, -1.679859, -1.299588, 
    -0.4116406, -0.7168422,
  1.076251, -1.923954, -0.1793424, 0.9558343, -3.036156, -0.07858675, 
    -0.1941225, -2.7723, -4.351609, -4.693684, -2.592196, -0.9884319, 
    -0.5648823, -2.447341, -1.792405,
  16.39749, 2.73616, 0.9160926, 2.822285, -0.9227214, -2.640282, -1.75264, 
    -2.135846, -3.386327, -3.058849, -0.7416697, -1.146829, -0.9414723, 
    -0.04988914, -1.335372,
  27.39722, 13.35059, 10.48034, 2.954791, -0.1037834, -2.043643, -1.175703, 
    -3.315588, -2.735032, -0.9743633, -1.099424, -1.045072, -0.3118467, 
    -0.7934534, -1.089383,
  20.92707, 7.451521, 4.440421, -0.7851969, -3.821951, -3.826364, -2.053238, 
    0.6282496, 0.5919082, 0.3871288, 3.020656, 2.231344, 1.466076, 
    -0.6892903, -0.8279525,
  20.76311, 10.70467, 1.058484, -3.491356, -2.977879, -1.710162, 1.182781, 
    2.355821, 2.656244, 3.048964, 2.505289, 3.349787, 1.885191, 0.8210471, 
    0.4431589,
  18.47518, 9.144469, -0.08488012, -4.226247, -2.746601, 2.834538, 8.149645, 
    7.596794, -0.7854706, -0.382321, -0.6938693, 1.271089, -1.095223, 
    -0.1410411, 0.7036033,
  20.66465, 7.81869, -0.4774307, -2.30922, 0.1645658, 8.649256, 10.12191, 
    10.9256, 4.010998, 2.419244, 3.492096, 0.1299944, 2.375196, 2.091136, 
    0.4706825,
  12.58478, 5.260535, 2.639871, 0.5342295, 3.8884, 3.989344, 9.206285, 
    9.60856, 7.718661, 7.036959, 7.635525, 4.665065, 4.233239, 0.8802065, 
    2.819674,
  5.816957, 1.155093, 2.222514, 0.2008693, 1.214052, 3.420396, 4.750662, 
    3.530115, 6.790024, 3.34013, 12.44898, 9.182978, 2.870599, 1.482044, 
    0.8482374,
  4.903165, 5.998007, 2.363876, 1.31142, -2.964505, -3.071554, -1.406302, 
    -3.188286, -5.689812, -3.990845, -6.924283, -6.275736, -7.003881, 
    -2.95203, -4.030611,
  8.34295, 3.937001, -0.944772, -3.43071, -3.988939, 1.946086, -1.239746, 
    -6.919049, -7.849659, -9.855776, -8.785881, -5.706223, -4.858743, 
    -4.229399, -3.474815,
  54.69243, 26.38986, 10.33014, 0.4711803, 2.71939, 1.541544, 7.298374, 
    -6.981695, -9.06566, -9.048694, -6.840137, -5.548235, 1.161948, 
    0.1550977, -0.2225691,
  79.30001, 64.38274, 49.18232, 25.06607, 6.00966, 6.002729, 4.784188, 
    -1.999281, -4.810891, -4.941515, -1.905724, 2.713062, 1.391408, 
    -0.4060074, -0.4945868,
  89.54347, 60.63388, 44.14243, 32.37734, 22.9546, 15.85623, 6.69173, 
    5.792382, 8.14572, 9.316611, 11.20369, 5.925487, 1.960713, -0.2761218, 
    3.27299,
  94.1323, 65.93013, 41.3963, 26.18207, 20.46601, 14.97147, 9.615466, 
    4.81168, 3.637586, 10.06447, 5.095219, 2.340595, 1.157685, 2.743717, 
    2.648859,
  79.38768, 60.19711, 36.95291, 18.63198, 17.28156, 12.24056, 11.19394, 
    9.02281, 3.532353, -1.071153, -1.086932, 0.1216355, 2.069445, 3.479093, 
    2.129116,
  67.82021, 51.83459, 32.06626, 17.28247, 11.58634, 12.32793, 8.676758, 
    7.292012, 2.030042, -1.771412, -2.314343, 1.769676, 1.274908, 3.115482, 
    2.789776,
  61.09227, 45.57125, 29.80877, 9.221329, 5.424506, 2.000367, 3.412956, 
    1.408714, -1.213799, 1.277075, 5.54247, 2.450085, 2.222856, 2.72857, 
    3.894973,
  40.4322, 24.36454, 14.43414, 2.893696, -1.733174, -1.591292, -1.712387, 
    -3.527731, -1.195574, -2.415206, 4.664673, 1.306085, 3.955405, 2.297874, 
    2.073648,
  6.984534, 11.73732, 7.719885, 4.877561, -0.9635597, 0.1371802, 4.981512, 
    1.675785, 3.214798, 1.287914, 2.105367, 2.052469, -0.793635, -0.3916246, 
    -1.75676,
  17.75848, 12.36057, 1.015459, -1.773596, -2.614132, 6.411448, 10.12586, 
    4.237305, 3.795216, 2.013545, 1.438633, 2.439005, -0.006047727, 
    -1.187926, -2.466514,
  84.88357, 59.7076, 27.93799, 4.791508, 10.7142, 7.497671, 20.89803, 
    12.18564, 6.753211, 3.78937, 0.3964724, -0.4618669, 0.7860574, 1.075681, 
    -0.4312948,
  113.05, 101.3821, 85.42408, 66.6934, 32.58694, 13.76767, 7.967448, 
    21.40243, 6.238531, -3.061912, 0.01065032, 1.358978, 1.62467, 1.198058, 
    -1.137567,
  129.1444, 99.1372, 81.96249, 70.76983, 59.17099, 37.82913, 20.99562, 
    5.420468, 11.88976, 6.883071, 7.891559, 1.822116, 2.115934, 0.4189573, 
    -1.154777,
  133.5298, 103.4775, 80.77534, 65.08003, 54.67845, 39.56319, 29.84733, 
    16.59066, 6.164475, 7.086111, 5.471366, 2.276669, 1.224151, 0.3255824, 
    -1.607568,
  114.7221, 94.48264, 71.42841, 48.08504, 38.77205, 30.50669, 24.4695, 
    14.96484, 7.809525, 3.549786, 2.410255, 1.426457, 0.5204886, -1.132837, 
    -1.390476,
  97.51422, 80.02534, 59.228, 37.19104, 26.02057, 23.20504, 11.61088, 
    6.50558, 3.126206, 0.44941, -0.1026707, 0.2764811, -0.4220562, -1.982721, 
    -0.219417,
  95.81113, 78.58762, 56.51763, 29.53951, 18.73184, 8.28157, 7.706101, 
    4.033734, 1.785909, 1.037547, 1.502794, -0.5257959, -2.314677, -2.608016, 
    -0.2297243,
  66.95355, 48.36655, 34.10338, 13.61543, 6.924318, 4.879791, 3.702683, 
    1.704093, 1.562057, 3.953677, 2.587463, -0.318615, -3.039964, -2.601941, 
    -0.5939938,
  8.433226, 14.76523, 9.931136, 13.84939, 4.595325, 5.056677, 7.54457, 
    1.39725, 2.25457, 0.6846545, 3.832284, 2.816854, 2.043978, 3.68303, 
    2.986075,
  24.44161, 18.62675, 5.091505, 3.243083, -0.5083394, 14.59779, 27.93085, 
    9.404482, 4.3372, 3.525371, 3.986953, 4.879425, 3.903668, 1.29563, 
    2.376209,
  107.2721, 79.11096, 37.98656, 10.92586, 2.102499, 7.763313, 42.86227, 
    16.10644, 5.082078, 3.76889, 3.270571, 3.974495, 4.171533, 4.664287, 
    3.733107,
  132.5238, 128.6175, 114.4006, 96.44434, 43.50419, 6.728018, 6.458217, 
    30.19988, 19.00261, 7.087803, 3.773136, 0.9930974, 3.510649, 4.491348, 
    2.234997,
  139.4191, 118.0734, 105.6508, 92.3395, 83.74704, 52.93619, 28.30206, 
    5.478143, 14.02979, 8.537084, 15.64136, 2.040949, 2.349695, 4.030582, 
    -0.3074164,
  135.8859, 115.8104, 98.78111, 86.68181, 79.96814, 68.80487, 56.00101, 
    31.59575, 8.528331, 9.463281, 8.118515, 1.201321, 0.8904682, 2.844539, 
    2.586166,
  111.5596, 100.524, 82.75582, 67.03834, 64.02609, 59.57596, 54.06664, 
    41.33876, 23.05293, 3.993142, 2.612886, 1.539085, 3.628761, 3.029142, 
    1.975479,
  103.0773, 91.11559, 77.61054, 60.93111, 52.483, 52.75173, 41.73192, 
    36.06158, 22.31095, 5.603849, 2.370614, 0.7347124, 0.5392958, 0.4027804, 
    1.363778,
  98.90613, 91.86177, 80.16806, 54.50221, 38.59829, 28.08579, 29.14231, 
    26.17961, 15.26084, 9.441341, 12.11848, 2.734362, 2.836132, 2.760169, 
    0.2164001,
  85.65278, 80.22507, 72.57728, 48.7252, 29.75609, 18.96057, 10.87392, 
    6.343828, 5.785064, 8.761722, 11.60802, 8.302004, 3.263608, 0.3915396, 
    -1.428494,
  8.598839, 12.60285, 8.82789, 11.8054, -0.9651868, 4.090631, 7.466276, 
    0.3335201, -0.4603038, 0.07416751, 2.354001, 2.625161, 0.5373743, 
    -0.418413, -1.01712,
  29.32501, 13.98756, 5.366831, 0.783029, -2.003118, 11.70432, 23.2676, 
    2.438988, -0.3588927, 0.08873336, 1.647132, 2.810888, 0.4834746, 
    -1.997543, -1.109092,
  91.24198, 78.95042, 48.42895, 14.76437, -0.7778364, -0.8827861, 48.57378, 
    14.71005, 0.9907182, -0.6955885, 2.540988, 2.158676, -0.4018443, 
    -0.137693, 0.507758,
  83.14867, 96.427, 101.1141, 97.14822, 41.56054, 5.385226, 2.954977, 
    36.75001, 15.08702, -0.1767632, -0.7799471, 2.699054, 3.02222, 3.564715, 
    3.805798,
  60.61082, 52.12328, 59.497, 67.70856, 75.59782, 51.81737, 29.24124, 
    6.640471, 11.07547, 9.862411, 17.02239, 7.116921, 3.518059, 1.926052, 
    0.9759572,
  60.95817, 42.01963, 32.60752, 29.2443, 33.56203, 38.56037, 44.5044, 
    38.26422, 2.80108, 4.473489, 6.353438, 8.48274, 6.365528, 4.364683, 
    2.705247,
  81.9411, 66.12932, 54.50425, 46.17118, 47.45642, 46.97384, 50.46146, 
    48.68244, 33.77202, 6.305119, 7.954051, 7.499958, 5.026536, 3.608469, 
    3.010875,
  111.0779, 94.99518, 81.97506, 73.77521, 72.33942, 70.8806, 56.93114, 
    46.06016, 32.08177, 2.213649, 3.860754, 2.472544, 2.746574, 2.035348, 
    1.45874,
  126.5454, 117.5681, 104.887, 87.31127, 76.97518, 63.9777, 52.74137, 
    42.48478, 22.34432, 10.44001, 25.98902, 7.59622, 4.623483, 0.763741, 
    -0.1560046,
  118.8097, 112.3504, 104.8298, 85.87143, 66.84686, 48.52433, 28.16592, 
    12.35269, 13.51187, 9.724479, 18.21206, 8.850883, 2.020109, -0.09405952, 
    -0.4601309,
  10.9514, 17.58259, 16.61627, 17.5868, 1.232492, 4.033365, 9.206289, 
    -1.286613, -2.451065, -2.726454, -1.794955, 0.2845971, -1.449125, 
    -1.339469, -1.850559,
  34.29975, 20.2452, 11.20235, 4.602374, -2.014219, 14.69912, 25.53616, 
    3.694875, -1.895076, -1.703998, 1.30982, 3.324961, -0.2005305, -2.894871, 
    -2.151715,
  56.15651, 50.448, 45.13408, 14.90881, 1.101234, 0.5788496, 43.56945, 
    15.66062, 1.187028, -1.581149, 4.356527, 1.401173, -0.2896102, 
    -0.5815083, -1.215201,
  52.28486, 48.0868, 48.91588, 53.3501, 33.96002, 4.929929, 2.039088, 
    32.76545, 19.79228, 1.851014, 1.338186, 1.794279, -1.658955, -0.9735625, 
    -1.174687,
  54.59466, 41.54119, 36.90854, 37.00881, 37.66311, 36.54256, 26.87868, 
    3.29043, 6.708549, 11.92383, 13.44654, 1.799009, -0.8448159, -1.66616, 
    -1.597265,
  74.56741, 56.91481, 49.56064, 43.00965, 43.2901, 32.9485, 43.11827, 
    36.91218, 5.484413, 0.5770407, 4.935421, 3.607596, 2.978589, 2.917304, 
    3.166155,
  90.80222, 76.6973, 59.31364, 50.23574, 50.90833, 52.14195, 40.76438, 
    36.55199, 25.30531, 8.33453, 4.522566, 6.017321, 3.504299, 1.967942, 
    1.443788,
  96.09171, 88.43172, 73.59711, 60.69981, 55.12657, 53.49904, 46.72903, 
    40.81102, 27.64492, 2.219496, 0.4371805, -0.3080081, -0.9157287, 
    -0.9954056, 0.02645,
  87.93005, 89.29797, 82.89723, 70.26093, 66.24009, 61.88292, 57.78361, 
    51.12474, 30.14552, 20.37409, 41.73618, 4.638021, -0.572404, -1.508417, 
    -1.910929,
  70.74546, 77.08968, 77.84695, 64.21171, 59.19159, 47.59967, 26.08377, 
    12.56047, 14.8853, 10.61998, 24.60779, 7.121814, 3.054089, 1.985719, 
    0.9971849,
  9.324906, 16.69868, 13.96491, 18.25063, 2.554796, 7.021338, 13.65743, 
    4.146435, 0.666465, -0.1922874, 2.558734, 4.268527, 1.931365, 1.03482, 
    0.4309795,
  27.9847, 22.50804, 13.02631, 7.807407, -0.5744366, 19.58294, 29.89682, 
    8.427144, 1.569432, 0.3690257, 6.816765, 10.23121, 4.520355, -1.478583, 
    -0.5634794,
  50.08276, 39.31733, 36.52443, 10.5202, 1.875208, 1.754473, 40.14448, 
    20.86116, 7.937434, 1.966771, 8.588349, 7.148789, 2.999469, 2.745234, 
    0.9317961,
  50.65396, 47.67327, 50.34447, 51.17544, 23.10808, 3.730291, -0.1435679, 
    26.49561, 19.16544, 3.591655, 6.266503, 7.332445, 4.088881, 3.869726, 
    1.895801,
  51.45573, 39.89571, 38.78256, 41.43379, 43.51101, 30.07928, 17.55989, 
    3.952733, 10.6856, 8.255809, 14.0484, 5.624501, 2.744027, 1.535325, 
    1.58158,
  64.03122, 49.73091, 40.56884, 35.82761, 36.48739, 39.37555, 44.66961, 
    28.41446, 3.072989, -0.5219243, 0.5885051, -0.7488438, -1.293101, 
    -0.2444824, 0.5021273,
  80.51273, 67.6141, 53.40797, 48.50321, 48.08891, 46.84576, 48.0011, 
    45.57572, 27.60418, 5.552867, 1.549825, 0.7469596, 0.8511103, -0.2434367, 
    -1.117394,
  103.3358, 91.40045, 78.73042, 75.26903, 75.06483, 74.74384, 64.58522, 
    58.82447, 32.13204, 4.540134, 1.59696, 1.30769, 0.7852826, 0.1789705, 
    -0.3937433,
  119.3757, 111.757, 102.4609, 94.42988, 89.09182, 79.57234, 71.73164, 
    53.74294, 25.49446, 15.4818, 25.44591, 1.990078, 0.3691415, 0.1209832, 
    0.0864189,
  103.3761, 100.6836, 97.04888, 82.71478, 69.85825, 51.04074, 27.31229, 
    17.91287, 17.44399, 9.443393, 14.98931, 0.8871168, 0.7284331, 0.6647623, 
    1.410578,
  9.636248, 18.53181, 17.8991, 18.41269, 2.594181, 2.961803, 12.41312, 
    2.187389, 0.1507019, -0.924073, 1.30465, 4.661441, 0.813588, -0.6463923, 
    -1.070585,
  21.51109, 18.40498, 13.91358, 7.288987, 4.452792, 25.26661, 29.81849, 
    5.436512, -0.6340856, -1.150665, 3.617606, 9.327283, 5.141623, -1.077569, 
    -0.351234,
  49.65343, 37.99233, 34.35171, 10.2187, 4.844835, 3.965756, 37.15806, 
    16.57026, 4.826535, -0.998875, 6.811653, 5.403562, 0.9898329, 2.039024, 
    0.6420643,
  54.57508, 48.39342, 47.95551, 37.6662, 23.13886, 9.837066, 3.559628, 
    22.81029, 11.83185, 1.345773, 3.304636, 2.645577, -0.08900806, 2.066498, 
    2.10437,
  65.90444, 58.81204, 57.28429, 56.86474, 36.14133, 29.69939, 18.81632, 
    3.902354, 7.702297, 7.125417, 14.61763, 7.792048, 1.524594, 0.9575947, 
    0.246574,
  77.91571, 74.75957, 70.1835, 70.80016, 77.02394, 51.37048, 36.07191, 
    23.85742, 3.759778, 1.449831, 2.980891, 2.360238, 1.555035, 0.4058156, 
    -0.7616412,
  81.25413, 82.06901, 73.17374, 73.63916, 83.69462, 92.18371, 84.09587, 
    55.91685, 23.42458, 4.133821, 1.923625, 0.4650187, 0.42904, -0.9166317, 
    -0.480867,
  82.7374, 73.09833, 61.98402, 62.68536, 68.73109, 78.54485, 76.56322, 
    74.28017, 31.29856, 8.672359, 1.719594, 1.053408, 1.064021, -0.2022473, 
    -0.9776288,
  87.29636, 70.22615, 60.01299, 56.52241, 58.66514, 57.60682, 52.40772, 
    36.06271, 18.96962, 14.36251, 16.09633, 2.265358, 0.1053375, 0.06190119, 
    0.07955436,
  92.00948, 70.17563, 60.08638, 44.70596, 38.26158, 29.69507, 17.95294, 
    13.97866, 12.60489, 7.763633, 8.167176, 0.7049639, 0.9859377, 0.5439801, 
    1.330531,
  9.532152, 15.07024, 10.17675, 14.09601, -1.466819, 3.016914, 10.19523, 
    1.000336, 0.7237169, -0.8104279, 1.421367, 3.575162, -0.006445527, 
    -0.5851552, -0.922075,
  32.29867, 22.71077, 7.98823, 4.667947, -1.391326, 16.49268, 20.73861, 
    2.364363, -0.04056245, 0.623805, 4.56824, 9.345811, 4.955382, -0.6983109, 
    -0.6778686,
  57.09753, 52.84748, 34.59722, 3.547364, 2.375182, 2.777515, 27.00433, 
    8.734971, 1.227926, -0.5066484, 11.03157, 8.698533, 1.506434, 1.772234, 
    0.2450126,
  50.75285, 56.55313, 47.77981, 35.20155, 16.08528, 3.439861, 0.9009537, 
    12.76919, 7.25918, 0.6244166, 3.671712, 4.822048, 2.155133, 2.450563, 
    3.334762,
  74.57838, 70.32983, 55.79291, 46.83341, 36.07377, 19.45507, 8.349995, 
    0.4790759, 5.121462, 4.929121, 10.85987, 3.953933, 3.07485, 3.300693, 
    2.635084,
  112.6278, 97.93974, 70.9129, 48.26275, 53.52996, 47.91853, 37.86052, 
    18.16743, 2.805291, 1.741678, 4.164302, 4.869164, 1.177387, 1.182161, 
    1.311607,
  136.8904, 112.3687, 76.60861, 47.47672, 51.96491, 70.8413, 81.6526, 
    66.77481, 25.67349, 8.96559, 5.909829, 1.689631, 1.47276, 0.4335572, 
    1.262715,
  135.598, 102.187, 59.79013, 54.45629, 57.41259, 65.62025, 63.59294, 
    51.82744, 16.50178, 6.667192, 3.505495, 3.144705, 3.014321, 0.5775229, 
    0.9144019,
  146.5731, 123.1042, 97.23866, 74.51564, 61.48671, 47.87324, 42.43169, 
    26.8125, 12.80769, 11.57434, 12.33461, 3.750223, 0.9901108, 0.7279097, 
    0.2506637,
  161.111, 131.0173, 112.7525, 79.2656, 59.40571, 33.23883, 18.69444, 
    11.43204, 7.779245, 6.483746, 6.177783, 1.014662, 0.4925878, 0.2088311, 
    1.002726,
  9.919583, 17.30066, 13.33459, 13.46007, 2.021158, 6.802731, 15.07888, 
    0.1479663, 2.973409, 1.73219, 3.186131, 5.873537, 2.262995, 0.6032555, 
    -0.3786741,
  24.7067, 13.68934, 6.596042, 3.371925, -0.5432887, 19.86605, 23.23781, 
    3.361459, 1.969206, 4.285196, 7.62679, 11.62411, 7.950454, 0.9147947, 
    -0.2572634,
  52.51332, 46.78766, 30.74556, 5.9697, 3.520129, 0.7515644, 25.26168, 
    12.10259, 2.339298, 0.03238342, 14.84769, 11.22279, 4.573127, 4.009881, 
    1.437504,
  56.53345, 62.41013, 69.09586, 56.95918, 26.83195, 6.569636, -0.6496505, 
    9.960818, 6.519596, 2.170712, 2.61076, 2.729575, 2.843359, 3.107018, 
    3.641677,
  68.08393, 73.92796, 75.47882, 69.65369, 61.86928, 37.134, 8.600003, 
    -0.05769422, 2.204556, 1.938686, 4.506897, 0.6559052, 0.2765961, 
    2.994403, 2.678076,
  118.9202, 105.9989, 88.89292, 69.44013, 52.24389, 45.43345, 47.53197, 
    18.27439, 2.168753, 1.065404, 0.4851954, 1.299094, -0.8249782, -1.667298, 
    -1.443798,
  147.0782, 128.5827, 102.7159, 73.27668, 55.07247, 50.03984, 54.90751, 
    50.07997, 13.63427, 5.466974, 1.850582, -0.6116993, -0.7319043, 
    -1.462537, -2.096854,
  173.2031, 148.1383, 122.6028, 99.81889, 92.83425, 90.36578, 79.34074, 
    68.27064, 20.41072, 6.043579, 2.552256, 1.535738, 0.4711268, -0.382011, 
    -1.052914,
  203.5812, 175.6058, 155.0753, 126.31, 103.1597, 79.64197, 50.98777, 
    37.31024, 19.60047, 11.44101, 5.159283, 1.655578, 0.8168426, 0.1090562, 
    -0.3112368,
  179.1599, 152.1294, 130.8291, 75.67622, 47.0814, 28.08339, 22.19984, 
    20.5327, 11.40032, 6.42815, 2.575958, 0.6490391, 0.3062659, 0.2124477, 
    0.2630271,
  3.043342, 8.365808, 5.369421, 9.215887, 1.966169, 5.611006, 11.43017, 
    4.556148, 4.304733, 1.715453, 1.145565, 2.67446, 0.3744179, -0.1641784, 
    -0.3257529,
  17.54303, 7.558211, 5.650983, 4.139949, -0.004418987, 9.244152, 12.23877, 
    4.201063, 3.849452, 4.863791, 4.308456, 7.194433, 3.962681, -0.2330336, 
    -0.4167754,
  50.90778, 38.47618, 17.40399, 3.772252, 3.804351, 1.491036, 10.87245, 
    6.746195, 4.619035, 6.398775, 14.11361, 8.660316, 0.6244587, 1.351249, 
    0.1347473,
  38.13242, 37.74413, 51.46238, 38.57705, 15.71435, 4.829234, -0.3523106, 
    6.344265, 6.979866, 5.856353, 6.800614, 6.469513, 0.93029, 0.8285818, 
    1.844436,
  80.40564, 76.0312, 68.30048, 60.88083, 47.34915, 24.37303, 8.356426, 
    0.222752, 1.713577, 3.350927, 4.852377, 3.40659, 1.425452, 1.403393, 
    1.331456,
  125.7306, 108.1225, 94.80416, 81.04377, 72.10369, 57.38212, 39.74213, 
    19.89432, 7.552169, 6.879227, 4.095043, 2.802652, 2.094643, 1.052696, 
    0.1091699,
  143.397, 131.5803, 113.9259, 100.4089, 93.43165, 81.93346, 61.1445, 
    35.74632, 11.61308, 9.740399, 4.916357, 1.017124, 0.008159536, 0.8099894, 
    0.8727504,
  156.709, 147.9612, 131.81, 121.6289, 112.4514, 105.3272, 79.9861, 62.3393, 
    13.18185, 1.543528, 3.235308, 1.842857, -0.07243426, -0.3327206, 0.1456727,
  150.1356, 142.3047, 135.2259, 118.7727, 84.22401, 60.89654, 50.22097, 
    33.9062, 11.11467, 3.16426, 4.912498, 2.115764, -0.3344897, -0.8898684, 
    -0.7113947,
  125.951, 116.6237, 105.5057, 57.44862, 31.01858, 16.82476, 14.81504, 
    19.35372, 9.990909, 1.6057, 2.145909, 0.4759702, -0.1684238, -0.05160339, 
    1.022957,
  3.703366, 5.328925, 2.409638, 5.203924, 3.516695, 6.945303, 10.52868, 
    2.919256, 1.092333, 3.061877, 2.841709, 5.492331, 3.245187, 2.272308, 
    1.115501,
  20.0192, 13.02908, 2.694352, -0.2348914, 1.077765, 10.69617, 9.990748, 
    4.132512, 1.939239, 4.15437, 6.028474, 14.4713, 12.5657, -0.701148, 
    -0.2512487,
  40.53384, 40.49393, 22.05552, 1.244189, -0.07679018, -0.8206546, 9.389323, 
    6.139486, 4.717746, 4.205225, 13.26749, 8.180907, 4.643218, 6.03524, 
    1.733894,
  50.30874, 33.35743, 41.96211, 43.28929, 11.14722, 3.954144, -0.5897752, 
    3.793497, 3.745774, 2.17082, 2.821061, 4.318365, 2.319355, 3.622356, 
    3.664846,
  119.4392, 95.3829, 65.39652, 33.85017, 43.61244, 25.07795, 9.049622, 
    1.005051, 0.8478833, -0.1652538, 2.64957, 1.710611, 1.073408, 1.686107, 
    1.306363,
  133.7411, 130.9825, 121.6312, 89.47735, 60.07737, 46.35794, 37.62235, 
    15.39829, 6.866483, 6.932343, 4.723991, 4.127508, 2.260173, 0.5512128, 
    0.2708068,
  129.875, 130.7195, 130.8659, 126.2543, 120.4123, 96.29472, 59.5789, 
    35.27776, 12.69217, 13.12875, 7.091452, 1.964399, 1.148754, -0.09505803, 
    0.2529273,
  126.2949, 120.6446, 116.8556, 117.1977, 122.7118, 120.6154, 90.62038, 
    55.10666, 10.41197, 2.326861, 1.847398, 2.208391, 2.110735, 0.3502366, 
    0.2155268,
  122.3575, 119.4451, 121.6735, 113.8707, 76.31185, 61.00161, 50.04784, 
    29.99663, 11.46244, 3.637101, 1.695829, 2.365681, 1.06745, 1.664598, 
    0.6937389,
  117.2753, 103.5383, 97.72542, 52.43141, 24.28182, 13.8316, 12.37644, 
    18.36254, 10.92406, 0.8243782, 0.6450568, 1.536807, 2.16355, 2.038485, 
    2.132248,
  5.404662, 5.548995, 3.48376, 4.579548, 2.449775, 4.55773, 10.63186, 
    6.497167, 8.299306, 2.032952, 0.2111214, 8.194454, 5.147171, 3.70605, 
    1.61638,
  15.37467, 4.978432, 3.500475, 1.197817, 0.8857738, 8.226168, 12.17997, 
    6.550169, 2.867821, 10.00323, 4.864781, 13.55169, 14.97183, 1.108641, 
    0.0625532,
  71.00584, 24.69325, 13.41101, 1.072333, 3.071448, 0.1189457, 9.238224, 
    8.41756, 4.390395, 7.350257, 13.64221, 7.055607, 4.363616, 9.204147, 
    4.212916,
  125.3304, 68.39661, 41.69936, 42.84666, 8.470553, 5.404868, -0.3771086, 
    4.43244, 4.89044, 3.0748, 4.135899, 4.909578, 2.24617, 5.130326, 8.702857,
  138.0486, 124.1039, 61.27312, 43.60243, 55.47449, 19.68179, 12.21521, 
    -1.646871, -1.164386, 0.7872146, 3.490983, 3.789318, 2.544544, 3.844365, 
    6.536257,
  120.3097, 132.8836, 121.6302, 60.59538, 55.89475, 65.39383, 43.72617, 
    19.4368, 11.33265, 12.25248, 10.52455, 8.709432, 4.435757, 0.7043632, 
    0.639948,
  120.4004, 127.0722, 136.3846, 109.3294, 70.86607, 64.02545, 54.99581, 
    45.26957, 18.48922, 18.65232, 13.46588, 6.391707, 1.803993, 0.9900978, 
    1.588242,
  126.3867, 123.0048, 126.7984, 122.0542, 105.6477, 80.1215, 54.47491, 
    32.6825, 9.806539, 3.821202, 1.111728, 5.182357, 2.857636, 0.2141911, 
    1.534527,
  146.8946, 135.0059, 131.907, 118.6689, 68.66545, 48.27018, 32.4186, 
    15.55002, 3.88831, 0.8870779, -0.4581871, 3.042228, 2.160665, 0.6764488, 
    1.609753,
  133.8706, 120.3392, 103.957, 50.53819, 19.19444, 11.57842, 9.344169, 
    13.72622, 4.995981, -1.097878, -0.7836344, 2.981674, 2.463599, 3.92635, 
    4.051002,
  3.061623, 9.935167, 3.182284, 8.601567, 6.007753, 4.955175, 15.09131, 
    8.362559, 9.421849, 2.450495, 0.9297222, 3.726008, -0.7765248, -2.501439, 
    -3.580653,
  32.34975, 8.585974, 5.917196, 4.335653, 1.687588, 5.683316, 8.645703, 
    4.663864, 1.762085, 11.05885, 2.186305, 10.32763, 11.07622, -2.637249, 
    -3.309569,
  115.3409, 58.21879, 17.58278, 4.596961, 3.868526, 0.3529231, 6.256145, 
    4.09295, 1.996274, 7.655152, 10.63347, 2.201042, 1.757927, 8.052748, 
    1.832955,
  133.1365, 114.108, 80.22078, 48.4216, 12.92784, 9.483373, -1.017406, 
    0.1537119, 2.152223, 0.9898846, 0.1820195, -0.05799042, -0.6312618, 
    3.685024, 9.085467,
  136.9311, 115.3339, 93.33306, 71.13115, 56.38411, 24.7161, 17.75023, 
    -1.685235, -1.481161, -1.312224, -1.598098, -0.556206, -0.06713495, 
    3.253809, 7.969224,
  144.8104, 131.5429, 110.8139, 81.15955, 72.75014, 69.00186, 38.98925, 
    20.18613, 14.19769, 16.12295, 5.927698, 2.41379, 1.645448, -0.04448749, 
    -0.1920199,
  152.2795, 151.5925, 127.71, 99.46967, 82.73849, 77.40237, 71.90533, 
    46.79424, 23.50245, 28.55996, 15.57052, 4.829176, 2.825353, 0.851712, 
    -0.7309126,
  161.8659, 159.3571, 138.894, 115.6721, 96.04369, 77.58031, 67.60442, 
    51.06643, 13.2613, 6.335359, 4.27108, 4.83948, 4.602006, 0.9942273, 
    -0.1390413,
  168.4556, 165.7915, 156.2322, 117.0866, 53.92212, 43.05979, 35.72849, 
    21.42727, 8.254116, 3.462464, 3.241389, 5.26355, 2.281567, 0.5472095, 
    1.277106,
  138.9886, 128.0429, 112.0602, 49.29536, 18.8522, 12.57961, 12.70736, 
    22.94083, 9.206445, 2.536146, 4.685773, 3.822316, 3.40547, 0.7706236, 
    2.715749,
  2.988695, 10.68878, 4.812542, 6.796207, 2.280535, 5.098886, 16.68489, 
    8.260121, 10.27993, 4.400008, 5.09793, 7.662319, 2.211668, -0.09167443, 
    -1.926595,
  37.46715, 13.90726, 7.546229, 5.844191, 1.429928, 3.145568, 13.70928, 
    9.739537, 5.340526, 13.55306, 5.888784, 13.04649, 13.52344, 0.4975284, 
    -0.9580925,
  88.60468, 48.38886, 19.96867, 6.03303, 3.545408, -1.249829, 7.379891, 
    6.943944, 6.046851, 11.14251, 9.492773, 6.377231, 6.187712, 8.322006, 
    2.338556,
  112.5458, 95.98917, 86.3651, 61.1755, 15.44929, 15.90929, -0.5142096, 
    2.197108, 4.318505, 2.131122, 2.398215, 2.325512, 2.530718, 8.058232, 
    9.427196,
  128.1574, 105.4604, 97.60448, 98.17224, 70.93217, 36.48241, 33.04419, 
    -1.50028, -1.278496, -1.270542, 0.2614288, 1.802472, 3.602487, 5.525944, 
    9.650279,
  144.7057, 122.4088, 108.2948, 100.9612, 109.0533, 94.14673, 41.19624, 
    22.74452, 15.41737, 15.12023, 5.861205, 4.854538, 4.353373, 2.635706, 
    2.20961,
  158.7811, 140.6536, 119.0758, 104.409, 109.1863, 109.3083, 92.82559, 
    45.05149, 20.67967, 28.96074, 15.5394, 4.929102, 2.452058, 0.2838337, 
    -0.3332829,
  170.078, 147.98, 123.8432, 105.5147, 102.7632, 94.57954, 83.68662, 
    54.83899, 6.588829, 2.68788, 2.909161, 1.33106, 0.01399682, -0.3491144, 
    -0.01370925,
  166.5055, 149.9943, 133.5864, 88.99371, 48.89985, 45.23363, 37.0808, 
    15.12213, 3.046529, -0.5109892, -0.9228903, 0.3754868, 1.293017, 
    0.7489223, 2.526384,
  127.6838, 106.2238, 83.8574, 30.72374, 6.731597, 3.061593, 4.394678, 
    15.48422, 3.902503, -0.09801307, -0.570269, 0.4017186, 2.465174, 
    0.3002842, 3.156206,
  0.7899338, 4.575413, 1.780321, 5.360276, 1.025493, 3.587324, 7.667677, 
    5.006925, 6.74924, 1.292111, 0.7698832, 7.357461, 3.953676, 2.383729, 
    -0.4447821,
  38.23088, 9.719289, 3.309002, 2.5491, 1.13868, 3.488976, 7.348588, 
    2.782895, 0.8213834, 6.603689, 2.220237, 12.19481, 17.03778, 2.558912, 
    -0.6425495,
  108.0762, 64.33129, 26.8918, 11.13461, 15.45371, 0.1665143, 2.096756, 
    -0.08141546, -0.158044, 6.523411, 8.539541, 7.653617, 11.93951, 14.39084, 
    4.4688,
  138.1736, 130.3413, 118.7677, 69.25672, 26.63862, 24.5829, -0.8386088, 
    -2.161829, -0.3704646, 0.2515953, 2.192067, 3.490644, 4.836611, 9.658442, 
    10.59946,
  133.9267, 119.9264, 115.9913, 108.0926, 53.9598, 31.53693, 28.33328, 
    0.2080507, -0.1494615, 0.8308439, 0.8337133, 1.921846, 1.52099, 7.626162, 
    11.28213,
  120.7359, 111.4906, 102.274, 93.83176, 90.09401, 61.95076, 24.65998, 
    19.47858, 13.57546, 19.35438, 5.971211, 4.189891, 2.696282, 2.84146, 
    1.403776,
  106.4425, 102.5116, 91.75366, 81.12626, 83.55528, 80.82541, 65.38277, 
    29.15407, 21.4608, 25.80549, 10.48247, 4.477657, 3.262295, 2.038724, 
    0.2330539,
  100.4746, 98.03016, 87.24811, 77.2887, 77.79671, 70.28101, 62.41821, 
    41.50972, 10.89768, 5.37367, 2.688962, 2.328418, 0.8185675, 0.8990702, 
    -0.103413,
  89.6946, 91.30871, 89.60931, 67.12952, 40.25208, 34.95858, 30.44538, 
    10.47873, 2.356475, 0.3722575, -0.03275099, -0.05601056, -0.07182936, 
    -0.06304086, 1.509454,
  61.32689, 57.39396, 52.57165, 20.24905, 9.354373, 4.387329, 5.3309, 
    6.569396, 1.205815, 0.3604477, 0.08012602, 0.0727319, 0.3872516, 
    0.1607266, 2.395898,
  5.673601, 11.63837, 5.664033, 5.573139, 3.822894, 2.787962, 7.303291, 
    7.701485, 11.80382, 6.082405, 2.69853, 5.997936, 1.970697, -0.1624503, 
    -2.681576,
  38.48741, 17.37552, 10.62248, 7.681941, 3.693772, 0.11239, 2.303665, 
    3.239144, 7.409675, 15.70318, 5.586512, 12.26287, 10.76519, -0.234419, 
    -2.169636,
  77.47474, 45.52302, 20.75062, 9.451737, 11.06845, -1.183607, 1.727966, 
    3.84601, 4.444406, 8.408164, 9.418921, 7.104014, 9.337223, 8.116943, 
    2.604858,
  94.35476, 88.63383, 80.42104, 43.06142, 16.93812, 14.70293, 0.7821622, 
    -0.7375525, -0.03014299, 2.701111, 5.13627, 5.328602, 6.038811, 5.884924, 
    6.46787,
  92.60941, 82.7131, 80.08508, 72.59095, 33.41475, 24.08871, 22.41379, 
    1.334594, -0.0444024, 1.004017, 3.27095, 1.794034, 4.048741, 3.749029, 
    5.200914,
  69.48475, 65.59474, 61.87865, 58.13654, 58.67712, 45.90973, 18.86834, 
    22.47316, 11.31627, 14.42587, 1.461923, 2.964928, 2.088866, 2.022695, 
    0.8196942,
  50.45742, 50.1705, 44.23718, 41.48241, 51.10054, 57.35799, 51.75927, 
    25.53228, 17.36204, 15.39815, 3.836805, 2.624846, 1.30087, 0.6709396, 
    0.4697837,
  48.55468, 49.06136, 43.15909, 40.67619, 48.96564, 49.32332, 43.54312, 
    27.32493, 5.916618, 3.714964, 1.599302, 1.960805, 1.889458, 1.398737, 
    0.3001082,
  55.53613, 59.86457, 56.08726, 42.69505, 24.66681, 20.08923, 18.05309, 
    6.001796, 2.751878, 2.335023, 0.8628984, 0.04528611, 0.9368213, 
    0.6135628, 2.667342,
  44.83483, 39.60159, 32.79221, 9.988139, 4.614219, 2.069551, 2.172424, 
    2.129323, 1.701478, 1.378016, 0.1449208, 0.07738672, 0.4564783, 
    0.3463978, 2.882521,
  3.807262, 10.65962, 6.088942, 9.247755, 8.424295, 4.150636, 6.576757, 
    5.122167, 12.20291, 6.662595, 3.037291, 5.810923, 4.128937, 0.6036286, 
    -1.600672,
  15.91818, 7.365229, 7.17765, 6.170622, 3.915471, 0.2004982, 6.294865, 
    4.912925, 8.752883, 14.45077, 2.677036, 10.91493, 18.72832, -2.355054, 
    -3.429125,
  47.72126, 22.38335, 10.94606, 5.620122, 6.231019, -0.7638651, 4.423758, 
    4.910983, 5.703192, 9.159429, 5.191825, 8.835026, 16.13761, 13.89504, 
    1.649734,
  59.8266, 51.5264, 45.08557, 28.85809, 13.00891, 14.49243, 0.7770862, 
    1.578783, 9.688672, 6.999934, 5.620124, 5.908081, 9.612594, 8.01161, 
    7.551116,
  70.09881, 53.83348, 44.58155, 41.46489, 22.83873, 25.42594, 22.72285, 
    -0.5970554, 4.955249, 7.493343, 4.02878, 1.886892, 4.392962, 4.381302, 
    9.17795,
  87.26139, 71.92995, 58.87762, 45.70492, 38.35206, 38.37043, 20.47924, 
    20.98756, 14.01325, 12.25667, 2.629669, 2.12003, 0.6345705, -0.4071553, 
    0.8689408,
  88.14307, 77.65264, 65.81824, 50.17055, 41.18291, 36.61623, 52.41901, 
    29.28051, 19.69386, 10.65981, 4.290544, 2.090034, -0.2635911, -1.335444, 
    -1.84508,
  74.47139, 61.19081, 49.08209, 40.09215, 42.75396, 41.92321, 41.56329, 
    28.39035, 10.86794, 8.486175, 5.037026, 2.633173, 0.8711451, -0.2336554, 
    -0.8818481,
  66.9439, 50.50374, 44.43298, 36.81223, 23.12269, 18.45275, 16.18618, 
    5.99614, 5.859745, 7.246586, 4.458266, 1.662878, 1.379327, -0.2693075, 
    2.107361,
  53.4633, 37.71749, 33.76222, 6.370066, 2.90202, 1.002344, 1.311635, 
    2.582903, 2.598416, 2.623667, 0.3239742, 0.7589166, 0.5902497, 
    -0.3580109, 1.490278,
  5.970777, 12.04284, 9.969385, 8.883695, 8.090846, 1.760396, 4.24878, 
    1.55993, 4.548876, 1.349956, 1.452004, 2.979613, 0.2985502, -1.268135, 
    -0.113153,
  29.40181, 11.96063, 8.90564, 7.589459, 3.243542, -0.1222754, 3.627908, 
    2.752867, 4.288167, 7.647427, 5.618585, 8.054809, 8.180506, -0.8063442, 
    -0.4872782,
  80.99802, 36.5196, 13.85992, 4.031024, 5.341089, -1.11948, 3.168245, 
    3.679539, 3.535969, 8.298427, 9.973845, 7.579525, 5.886652, 8.909203, 
    6.487288,
  86.5119, 78.79455, 74.15643, 43.35979, 10.4289, 5.082088, -0.3415588, 
    3.29023, 5.778468, 3.742826, 9.726416, 7.090722, 4.539525, 3.537922, 
    12.02358,
  83.78008, 57.22052, 62.35383, 57.60373, 18.07155, 13.50328, 14.2921, 
    0.1776404, 2.19602, 1.455992, 2.105608, 1.961362, 2.338878, 2.538415, 
    9.701479,
  83.56735, 58.39245, 62.93098, 60.12107, 52.81957, 42.1082, 16.01365, 
    12.65804, 7.631045, 5.894701, 1.084252, 0.5687811, -0.1582994, 4.464565, 
    5.143251,
  93.81342, 77.49091, 75.93842, 65.90534, 75.50696, 80.09862, 68.09823, 
    27.04657, 10.45184, 4.573747, 2.349161, -0.3277874, -0.2066951, 3.759228, 
    4.299592,
  102.9003, 88.0678, 83.36039, 85.03275, 102.7213, 97.94154, 80.05118, 
    30.77123, 8.126666, 2.257672, -0.4272868, -1.439368, 2.686309, 3.568018, 
    2.095468,
  105.5293, 95.5341, 105.2243, 94.94392, 58.51999, 48.03277, 34.73695, 
    11.92268, 6.457448, 1.477303, -0.4142101, 0.6201785, 2.082223, 3.032688, 
    4.289776,
  94.96902, 89.17733, 90.43118, 22.2816, 11.32724, 7.387245, 6.709749, 
    11.56002, 4.963806, 0.8278776, -1.019371, -0.2752171, 0.9143337, 
    1.012303, 1.923231,
  10.8473, 18.16075, 16.59517, 10.46447, 3.204747, 4.739457, 8.835649, 
    2.442744, 2.887864, 0.6173652, 1.053265, 3.324991, 1.062063, 0.8838992, 
    -0.7328515,
  21.29783, 15.93943, 16.44745, 8.000452, 2.989288, 6.943119, 8.307812, 
    2.762227, 3.068642, 5.11371, 3.577806, 6.110896, 7.106818, -0.3100891, 
    -1.032779,
  54.82008, 35.23146, 27.30505, 12.47789, 8.971059, 2.482983, 8.068266, 
    3.397163, 1.320232, 5.432103, 3.98285, 1.654284, 4.170973, 7.739233, 
    2.805328,
  55.71623, 71.17043, 87.46861, 64.81257, 15.3501, 8.065226, -0.06081075, 
    0.5850395, 1.381314, 1.256742, 1.282837, 1.424591, 3.295589, 5.167778, 
    5.247733,
  50.95375, 47.22168, 60.9451, 67.82958, 31.9623, 15.90691, 14.30326, 
    1.654236, 0.9137887, -0.02624129, -0.4257951, 0.6080714, 2.593694, 
    4.269022, 5.625473,
  99.0628, 86.59691, 82.52103, 79.42303, 69.30188, 40.58114, 13.96982, 
    19.29168, 10.01495, 8.228806, 0.9657458, 0.9109624, 1.761126, 3.407151, 
    3.826215,
  141.8063, 129.9046, 111.7458, 94.77632, 94.68422, 94.54005, 67.88239, 
    21.79366, 7.441621, 4.155895, 4.35167, 2.19973, 1.990655, 0.6810285, 
    0.2449064,
  173.7704, 164.7486, 145.819, 126.6018, 127.4205, 117.6832, 87.8119, 
    29.09389, 5.507992, 2.444004, 1.671912, 1.497142, 0.271037, 0.08805656, 
    -0.00937655,
  196.6922, 189.5668, 174.1656, 125.065, 81.12553, 62.63584, 37.53814, 
    12.89812, 2.476467, 1.373136, 0.3917704, 1.146111, 0.8633564, 0.8570692, 
    2.186048,
  167.6246, 154.3451, 118.1628, 25.85355, 14.3624, 6.27533, 5.45688, 
    14.38298, 3.3496, 2.276276, 0.3936279, 0.8438295, 1.234116, 0.4296832, 
    1.894847,
  6.717868, 14.90379, 17.14935, 13.941, 1.994292, 4.404149, 7.665853, 
    1.166133, 1.295968, -0.1485356, 0.5828787, 1.494596, 0.2919521, 
    0.8382845, -0.004525182,
  15.7201, 15.94295, 16.23755, 9.69235, 3.009358, 7.261256, 5.398427, 
    1.065801, 0.5411004, 1.451902, 1.002917, 3.737195, 4.133713, -0.1292174, 
    -0.1905923,
  45.57643, 30.42903, 20.37746, 11.90903, 11.49738, -0.395142, 1.686651, 
    0.3560112, 0.1053782, 1.873847, 2.677229, 2.576149, 4.858668, 8.568286, 
    2.793417,
  56.73268, 69.4944, 85.09476, 62.25507, 22.78151, 17.29721, -1.40381, 
    -0.06827955, 0.5209522, -0.05564907, 0.8634862, 0.9394608, 3.965825, 
    5.446682, 3.83549,
  97.27412, 90.56219, 104.0787, 107.5739, 35.63, 18.52357, 18.25853, 
    -0.2944423, 0.1548417, 0.2628221, 0.468281, 0.5465664, 3.446313, 
    4.586314, 4.689394,
  137.5724, 128.2232, 119.4812, 111.1593, 85.62065, 41.68147, 8.847628, 
    10.93466, 4.230277, 4.358967, 0.8688876, 1.248802, 2.677544, 3.275026, 
    4.016756,
  151.036, 145.9497, 125.9809, 104.9364, 99.03716, 82.59054, 39.32248, 
    11.01635, 4.372634, 3.721895, 1.929913, 1.419456, 1.276283, 0.8721017, 
    1.543148,
  153.2684, 145.1635, 124.6664, 104.5877, 99.86815, 85.78118, 58.66644, 
    18.11948, 5.11406, 2.13169, 0.4457825, 0.4439321, 0.1632933, 0.07973691, 
    1.35773,
  160.6536, 150.8909, 131.5316, 97.21337, 70.25398, 51.61681, 25.20997, 
    8.094605, 2.392662, 0.843794, 0.06382936, -0.1905777, -0.2162997, 
    0.2735058, 1.737774,
  133.0045, 119.6874, 81.69778, 15.82498, 6.351663, 5.499237, 2.951801, 
    6.4422, 1.911971, 0.4387189, -0.1613601, -0.2964325, -0.2403323, 
    -0.04749517, 0.777725,
  3.656258, 7.167528, 7.540684, 6.446011, 1.642161, 3.612134, 7.435907, 
    3.122318, 3.38802, 0.02068568, 0.09810527, 0.6005309, -0.09561584, 
    -0.07191042, -0.7605262,
  9.288404, 7.027572, 6.80075, 4.344369, 2.072933, 2.838658, 3.727733, 
    1.913186, 0.2935774, 1.429502, 0.6956308, 1.771896, 1.140498, -0.8472306, 
    -1.066647,
  47.14822, 24.84071, 13.25029, 9.203364, 12.95606, -2.453154, 2.50193, 
    1.348795, -0.2246843, 1.124301, 1.444334, 0.8036211, 2.283727, 4.171575, 
    1.090504,
  62.57385, 73.37763, 72.2149, 44.55949, 21.87885, 18.81751, -1.351005, 
    -0.4842702, 0.3821291, 0.3600661, 0.8547824, 1.645294, 3.36919, 5.996624, 
    3.942664,
  86.64374, 79.28466, 90.00928, 91.0856, 24.9072, 16.67237, 20.10452, 
    -0.3761629, 0.3669469, 0.4834587, 0.9901174, 0.8748327, 4.101905, 
    4.184525, 5.247979,
  109.7096, 98.999, 96.70618, 92.29388, 62.55156, 28.13688, 8.667454, 
    10.54852, 2.642658, 1.400823, 0.7575825, 0.884762, 2.68405, 3.637408, 
    3.587086,
  126.9679, 119.5393, 104.5848, 89.07006, 81.88863, 65.84589, 26.13843, 
    2.886411, 1.456634, 1.286935, 1.188196, 1.136019, 1.351161, 0.9505464, 
    1.936031,
  131.7411, 119.748, 97.63679, 81.40974, 77.37193, 65.70816, 45.67576, 
    13.90806, 2.560983, 1.198634, 0.5230988, 0.3552896, 0.1789786, 0.1609935, 
    1.828872,
  131.3989, 117.7366, 98.90179, 73.7401, 55.97231, 39.2348, 19.11161, 
    4.267552, 1.884445, 0.7582474, 0.1009862, 0.02927023, -0.08787226, 
    0.3520556, 1.618823,
  107.5871, 94.96961, 58.3739, 8.617567, 2.826733, 2.324134, 3.193919, 
    2.216947, 1.066565, 0.2896398, 0.09608596, -0.1108482, -0.2029659, 
    0.02361427, 0.6186045,
  5.19751, 8.486818, 4.814653, 2.940401, 0.5431216, 0.3018713, 2.738617, 
    3.486621, 7.241432, 3.48326, 1.129009, 2.709696, 0.4705891, -0.1446217, 
    -0.8162465,
  10.55801, 3.2642, 2.194049, 1.353446, 0.06791573, 0.2297352, 5.253278, 
    5.046925, 6.136176, 8.078125, 1.104558, 2.632577, 2.401822, -0.3592823, 
    -0.4176695,
  31.97244, 15.17405, 5.653316, 2.2239, 8.328739, -0.7099618, 2.230315, 
    2.619374, 2.159065, 3.93473, 2.380321, 0.4067617, 0.9667298, 1.65126, 
    1.572274,
  53.24646, 59.46415, 55.30265, 28.98717, 15.00034, 20.11322, -0.4503989, 
    -0.6714479, -0.2784406, -0.4618838, 0.1025366, 0.5695838, 1.574734, 
    2.995717, 3.04537,
  78.65922, 70.41429, 75.19558, 70.95703, 14.50677, 17.2427, 21.6966, 
    -0.09512186, -0.1235256, 0.3450509, 0.7004942, 0.6768405, 1.831092, 
    2.6988, 4.456103,
  88.00204, 84.00136, 82.79287, 78.66214, 51.31026, 21.94109, 8.438101, 
    12.66038, 3.2736, 2.812805, 0.544319, 0.4020651, 1.187011, 1.929428, 
    3.70929,
  88.92047, 93.62904, 88.1881, 79.784, 81.28005, 69.34258, 26.11041, 4.43259, 
    1.387761, 0.8789319, 0.4081855, 0.2506776, 0.2754418, 0.2538801, 1.076859,
  83.86174, 90.6964, 82.13145, 74.67203, 79.40794, 74.64634, 51.57473, 
    13.2099, 2.817374, 0.8985233, -0.06597362, -0.2152603, -0.3174117, 
    -0.2154959, 1.574007,
  79.37604, 84.79029, 81.25388, 71.72398, 62.9432, 47.5089, 22.63457, 
    6.021813, 2.542269, 0.7049531, -0.1362174, -0.283403, -0.3833803, 
    0.1072144, 2.447974,
  80.21519, 78.61595, 55.27074, 11.44846, 3.528527, 2.752672, 6.921828, 
    3.80952, 0.993763, -0.04957977, -0.3746369, -0.3040196, -0.02427871, 
    0.0263174, 1.09318,
  5.67055, 9.725774, 7.669638, 5.136595, 2.579179, 0.2979728, 2.457583, 
    2.368788, 4.80913, 1.530809, -0.02524396, 1.072637, 1.319449, 0.3467499, 
    -0.4481342,
  14.39752, 5.83843, 6.260094, 4.475141, 1.979375, -0.1946894, 2.631612, 
    2.859612, 5.27788, 9.096496, 0.2910242, 1.653879, 3.426524, 0.1933549, 
    -0.09262436,
  52.0363, 21.5927, 8.741211, 5.180288, 8.092701, -0.8470914, -0.4659574, 
    0.09124587, 0.576705, 3.267192, 2.531073, 0.4695855, 1.4314, 1.90883, 
    1.502699,
  67.14145, 64.9388, 56.43419, 25.40125, 9.227283, 11.43916, 0.2541684, 
    -1.065523, -0.06995848, 0.5073367, 1.686889, 2.303581, 4.479073, 
    4.604462, 2.459281,
  77.92933, 64.82967, 65.71933, 52.29609, 8.873663, 9.297225, 13.30322, 
    0.7865784, -0.7780553, -0.198835, 0.3903871, 0.9232666, 3.475113, 
    4.263199, 5.319134,
  90.11845, 76.10561, 69.75836, 55.43331, 35.52626, 16.11519, 8.671752, 
    12.90069, 5.985867, 4.021914, 0.3338702, 0.574201, 1.66519, 1.918205, 
    4.327782,
  101.5985, 93.17658, 79.86345, 62.96686, 65.33945, 61.5106, 24.24233, 
    8.836763, 5.064083, 3.005413, 1.417763, 0.7030746, 0.3472625, -0.3294203, 
    0.9399443,
  114.1845, 104.2142, 84.27591, 70.32843, 76.27316, 71.62971, 50.23944, 
    12.41875, 4.566344, 1.605396, 0.3840801, 0.1312973, -0.1670596, 0.108404, 
    2.34409,
  121.1992, 108.3613, 97.4715, 82.50688, 69.10529, 48.73384, 18.7709, 
    6.883577, 3.867786, 0.8506292, -0.1220345, -0.2182516, 0.02834091, 
    0.7004718, 4.196331,
  115.8486, 108.2527, 72.02443, 24.8007, 8.179914, 6.056065, 4.423459, 
    6.072254, 1.984586, 0.01090452, -0.5587403, -0.2808461, -0.001063216, 
    0.204336, 1.826964,
  11.54867, 17.37876, 8.063355, 7.860371, 3.999559, 0.3109089, 0.5689675, 
    0.2822036, 3.052584, 0.9097395, -0.1150491, -0.1321779, 0.1177961, 
    0.7095652, 0.1228292,
  21.1428, 12.34083, 9.747813, 6.026583, 2.644008, -0.6791436, -0.1852928, 
    0.03401369, 1.883022, 4.316, -0.1882009, 0.4122207, 2.102487, 0.1905383, 
    -0.1160363,
  71.3574, 25.35953, 7.462311, 4.770664, 4.795106, 0.1118171, -0.1075549, 
    -0.07416849, 0.646031, 2.158161, 1.5458, 1.259321, 3.272127, 3.578202, 
    1.541879,
  84.11239, 72.84257, 49.10973, 18.35873, 6.259519, 6.961913, 0.8495733, 
    -0.1540351, 0.1256157, 0.3361664, 1.033255, 1.365934, 4.148954, 4.606797, 
    2.681902,
  82.7017, 61.35749, 55.96498, 43.39519, 7.56679, 10.26333, 10.21464, 
    1.259433, -0.0954951, 0.3436172, 0.3889436, 0.3328735, 2.681817, 
    3.837993, 5.1575,
  90.34059, 66.30574, 56.15143, 46.72179, 31.81917, 16.57863, 10.32136, 
    10.37988, 4.12169, 3.327969, 0.5509236, 0.3129369, 0.6347235, 2.240233, 
    4.307891,
  100.3274, 76.20246, 61.37107, 52.08746, 56.41391, 48.37729, 17.26945, 
    8.281069, 4.854741, 2.854274, 1.615025, 0.3979927, -0.2194347, 
    -0.2684039, 0.848268,
  107.6398, 77.49471, 65.5695, 58.96395, 62.00769, 53.18819, 32.05578, 
    7.687101, 3.744697, 2.092644, 0.8045279, 0.2660027, -0.3313507, 
    -0.2421832, 0.8665036,
  105.6097, 85.97968, 84.54659, 68.85693, 54.97475, 35.92559, 11.58811, 
    4.857293, 3.143354, 1.124414, 0.2541626, 0.01306429, 0.02686094, 
    0.8197756, 1.880534,
  100.419, 90.60516, 64.21002, 20.74092, 7.431217, 4.880765, 3.753916, 
    3.956063, 1.449094, 0.2595717, 0.02604047, 0.05242974, 0.1345348, 
    0.4503486, 0.8572792,
  11.83619, 22.99591, 12.36693, 14.84892, 13.10919, 3.693322, 4.173384, 
    4.25271, 8.515423, 1.532866, -0.2435024, 0.07870225, 0.004271477, 
    0.2770025, -0.1017341,
  19.50448, 16.19491, 16.21157, 14.78753, 8.915738, -0.4193445, 0.421266, 
    0.2212876, 2.062337, 3.771689, -0.1256625, 0.1706998, 0.9723972, 
    -0.007753437, -0.3007939,
  67.19077, 22.1488, 14.92296, 14.19353, 11.95963, -0.9090081, -0.5610941, 
    -0.4232486, 0.175795, 1.256115, 0.8851469, 0.667051, 1.818213, 2.209314, 
    0.9972326,
  79.15439, 81.35339, 64.94257, 24.69242, 12.27971, 13.16549, 0.1849137, 
    -0.435004, -0.1639811, 0.6681167, 0.6434435, 0.8942712, 2.51711, 
    2.588857, 1.88757,
  72.07687, 67.84425, 71.39023, 52.29934, 8.027168, 11.02086, 13.63384, 
    1.083637, 0.2285142, 0.5551902, 0.5845169, 0.5672135, 2.099679, 2.765115, 
    3.857199,
  73.97555, 67.15411, 61.75819, 47.82977, 28.65155, 10.30993, 8.473467, 
    9.164921, 2.873649, 1.310981, 0.5352521, 0.2718397, 0.6062523, 1.744136, 
    2.773165,
  78.49584, 70.20548, 61.58579, 48.2364, 49.62294, 44.58906, 15.66588, 
    6.133017, 2.242143, 1.085201, 0.6055212, 0.1849464, 0.08927092, 
    0.4724765, 1.083649,
  78.94669, 62.76155, 56.73933, 43.33948, 48.02684, 54.00951, 34.44335, 
    6.227245, 2.001958, 0.6992696, 0.07335107, -0.0701769, -0.2028826, 
    0.3515594, 1.651679,
  63.07409, 48.41979, 55.33009, 46.68198, 41.67961, 32.44452, 11.10764, 
    3.536266, 1.268302, 0.5148509, -0.01234477, -0.1591747, -0.1405032, 
    0.5044838, 0.9399914,
  65.28851, 65.236, 45.36783, 12.87227, 4.832604, 2.77896, 2.479931, 
    1.783077, 0.4284729, -0.01031226, -0.104773, -0.04862448, -0.01024742, 
    0.2709261, 0.890308,
  10.8392, 23.21521, 12.56945, 17.47039, 25.44368, 8.186007, 6.53209, 
    8.798946, 22.01563, 9.200668, 2.004982, 4.127731, 1.77433, 1.399245, 
    -0.2551858,
  15.50376, 18.90195, 17.34176, 28.74774, 25.67242, 3.863486, 5.702753, 
    6.390363, 12.54282, 17.29476, 3.101218, 4.8781, 7.460557, 0.7814217, 
    -0.4133363,
  53.22631, 22.10369, 20.62799, 27.91838, 26.59956, 2.081108, 2.181812, 
    3.501578, 5.276311, 7.835544, 6.057002, 3.451842, 4.735728, 5.949153, 
    1.719577,
  82.15392, 96.11846, 73.99022, 32.01351, 22.43459, 21.38559, -0.1357147, 
    0.2669183, 0.5456308, 0.6203493, 0.4724799, 0.6771669, 2.428495, 
    3.277301, 1.578358,
  82.02149, 79.20547, 89.00423, 62.72267, 14.10935, 13.43366, 15.40137, 
    0.5202878, -0.2200069, 0.1832183, 0.2684982, 0.7977595, 1.317373, 
    2.021243, 2.239004,
  80.1842, 72.31213, 72.96432, 57.06808, 34.49603, 11.17569, 10.3083, 
    10.25164, 3.117356, 1.318091, 0.7348217, 0.6641459, 0.7924606, 1.249391, 
    1.840172,
  93.46763, 77.99214, 62.35846, 49.86139, 54.42788, 43.26928, 13.13167, 
    4.02714, 1.805032, 1.212473, 0.6631275, 0.2012716, 0.137136, 0.7355942, 
    1.200694,
  106.0354, 105.9277, 79.63313, 52.22376, 45.51665, 45.14109, 21.37033, 
    3.047945, 1.055532, 0.1171535, -0.5078809, -0.5689842, -0.6346155, 
    -0.1452589, 0.6766188,
  78.66259, 90.46304, 61.49598, 41.68807, 39.43059, 24.65677, 5.984545, 
    1.965793, 0.8886191, 1.249473, 0.7979415, 0.3172632, 0.2400873, 1.074226, 
    0.3525315,
  51.87991, 56.40879, 39.53695, 11.04988, 3.61424, 2.947459, 3.757467, 
    3.586523, 2.168127, -0.1207415, 2.588243, 3.743545, 0.856315, 1.740583, 
    1.422594,
  4.861222, 15.72794, 8.713657, 13.87104, 28.10395, 8.412468, 3.401807, 
    5.312284, 12.45551, 5.430481, -0.3722726, 1.841876, 3.440318, 3.334133, 
    0.5342036,
  5.774328, 12.7903, 12.84588, 33.15369, 28.07406, 7.556361, 5.44016, 
    5.456695, 9.284754, 13.81939, 0.9448144, 4.85483, 12.3669, 2.732349, 
    0.1659373,
  37.72918, 19.8348, 19.14215, 36.63178, 30.1344, 3.363928, 5.483388, 5.731, 
    7.249324, 8.090333, 5.738497, 5.021003, 8.674994, 14.26111, 6.517949,
  73.50238, 85.81784, 65.58782, 31.68972, 31.66522, 24.45702, 0.6530718, 
    2.892592, 2.925189, 3.932106, 3.41364, 4.25672, 7.62671, 9.091498, 
    8.308447,
  71.13004, 65.51322, 72.9939, 40.91003, 16.80278, 18.53588, 17.55744, 
    -0.1641239, -1.557237, -0.5303828, 0.4029958, 0.9742602, 4.191885, 
    6.414646, 6.76476,
  74.98309, 53.65291, 46.3551, 30.98924, 17.93388, 8.669602, 9.815477, 
    10.69413, 2.878281, 0.9714341, -0.1267242, -0.4928004, 0.6096256, 
    1.877695, 3.726814,
  86.84468, 63.65748, 42.98892, 28.22618, 31.22551, 21.67572, 4.559857, 
    2.212714, 1.6271, 1.227969, 0.7491938, -0.06552706, -0.2772889, 
    -0.3335385, 0.8545909,
  76.75304, 56.19761, 47.66187, 35.12498, 37.88404, 39.89046, 18.84997, 
    1.343487, 2.461893, 0.6637682, -0.4372057, -0.5894601, -0.6160679, 
    -0.6372433, 0.1305282,
  71.32171, 64.25014, 46.22392, 34.89961, 30.77222, 24.76188, 6.841307, 
    3.661548, 1.81673, 1.136982, 0.8942366, 1.183867, -0.1093379, -0.3874333, 
    -0.6871905,
  76.6328, 69.32568, 44.71354, 14.40037, 6.881322, 5.364603, 3.974302, 
    4.010021, 1.722203, 0.123343, 2.164967, 2.935886, 1.216502, 1.592733, 
    0.1165873,
  -0.4273238, 3.276105, 0.03714529, 7.815932, 22.56041, 8.368209, 2.229458, 
    -0.2223839, 2.402169, 1.407232, 0.5042242, 1.851164, -0.4084104, 
    -0.2439892, -1.987758,
  0.8666633, 2.445336, -0.05024532, 17.47935, 18.34064, 4.691138, 4.701615, 
    3.912, 2.774121, 3.363321, 0.6883966, 0.8212711, 4.624248, -0.2235038, 
    -1.426507,
  21.96124, 8.570964, 0.9271173, 13.6664, 15.92388, 2.285938, 3.932944, 
    5.683958, 6.296341, 5.112996, 0.4483516, 0.6825258, 2.532755, 4.929281, 
    1.41396,
  70.73785, 61.11496, 19.70867, 5.593863, 14.19547, 11.39392, 0.502667, 
    2.616303, 4.110201, 4.609333, 4.581661, 3.259047, 3.052796, 3.512667, 
    2.781576,
  83.0798, 53.03295, 31.71466, 7.657673, 4.27426, 7.55847, 8.891111, 
    0.5593026, -0.6344045, -0.1175535, 1.130353, 2.003499, 4.986237, 
    5.095906, 4.598041,
  88.2558, 53.68273, 19.18872, 9.671991, 7.041349, 5.102061, 5.994498, 
    6.053902, 1.773229, 0.9824852, -0.2370408, -0.1562546, 0.6675343, 
    3.864242, 6.073554,
  82.28978, 46.82551, 28.08831, 19.98647, 21.08026, 17.62513, 5.865068, 
    2.353285, 2.198824, 1.509286, 0.6788749, 0.1268783, -0.05238351, 
    -0.1083458, 2.810174,
  63.82428, 46.81022, 43.69988, 31.15797, 27.85072, 28.36303, 12.84109, 
    3.661087, 2.947954, 2.551395, 1.125887, 0.3208056, -0.05918572, 
    -0.2778388, 0.396659,
  58.48931, 53.84549, 49.07985, 27.82285, 19.38963, 12.41728, 3.331457, 
    1.673977, 2.304894, 2.01459, 0.5831644, 1.657123, 0.6305035, 0.06151982, 
    0.2031639,
  54.33384, 47.43537, 27.93066, 6.326366, 2.756556, 2.605112, 2.145129, 
    1.223187, 1.154724, 0.7802762, 0.6078269, 0.9487783, 1.209023, 0.2221872, 
    0.3256447,
  3.684631, 4.08075, 0.2859094, 0.8814225, 3.670865, 1.482001, 0.06676659, 
    0.4260716, 3.098648, 3.423337, 1.571887, 2.57142, 1.200672, -0.3889331, 
    -1.156935,
  8.090662, 4.995725, 1.237493, 3.172431, 3.413388, 0.1351701, 0.7175878, 
    0.9980589, 4.476013, 5.141616, 2.422787, 4.043149, 4.86408, 1.703099, 
    0.649738,
  28.14509, 11.06774, 4.303152, 4.353348, 3.84983, -0.05945795, 0.4164984, 
    0.8683228, 1.853719, 2.922011, 1.690247, 2.106673, 4.567719, 4.659844, 
    2.916863,
  76.15073, 78.01968, 47.31974, 7.551461, 3.509595, 3.027906, 0.3226441, 
    0.5768516, 0.6866046, 1.00811, 2.055053, 2.561825, 2.849086, 1.399809, 
    1.482209,
  89.46608, 74.28904, 70.88906, 23.9317, 2.239194, 2.048493, 4.06191, 
    0.6275893, 0.140651, 0.2652193, 0.4978381, 1.270947, 3.132858, 3.093828, 
    2.558681,
  98.51198, 82.23742, 60.99824, 31.44277, 7.151089, 2.523163, 3.451585, 
    4.578448, 2.423858, 1.198637, 0.335195, 0.3899222, 1.247271, 2.423773, 
    4.988541,
  100.6584, 92.73135, 74.49662, 43.98015, 33.49788, 15.67307, 5.273983, 
    3.104388, 2.937211, 2.847014, 1.049616, 0.5768713, 0.4482953, 0.66857, 
    2.445466,
  98.1997, 90.89803, 76.41012, 50.41419, 36.13034, 27.51586, 11.66159, 
    3.276643, 2.460793, 2.818633, 1.43196, 0.2702031, -0.01547746, 0.2239985, 
    1.392993,
  90.26559, 85.62133, 72.52638, 42.96567, 24.17389, 8.20799, 3.419057, 
    2.925812, 3.483984, 1.735618, 1.228108, 0.2986873, -0.0743221, 
    0.08416065, 1.16037,
  75.9727, 69.05685, 43.4494, 6.573717, 1.028726, 0.3326435, 3.746036, 
    4.241874, 2.156991, 1.42913, 1.467996, 0.556071, 0.124756, -0.0443415, 
    0.8406942,
  2.351553, 4.009615, 2.252579, 2.773167, 3.418243, 0.7811267, 0.3033568, 
    0.7897016, 4.51555, 3.922743, 1.947094, 2.780937, 2.385322, 0.5208082, 
    -0.2309592,
  7.033609, 4.907873, 3.99912, 5.865242, 5.584814, 0.2020098, 0.3694468, 
    0.5192615, 2.066455, 4.119112, 2.518719, 6.638576, 5.903725, 2.023, 
    0.06259236,
  14.65076, 11.42974, 7.06249, 12.19302, 11.7059, 0.2011797, 0.3500323, 
    0.5695592, 0.926734, 0.9757853, 1.233881, 3.961579, 5.72313, 8.545634, 
    4.072796,
  52.2044, 54.09664, 47.34865, 21.73653, 16.98277, 11.42955, 0.4346025, 
    0.2204999, 0.3791922, 0.5076889, 0.5198283, 1.650355, 3.076025, 3.758928, 
    2.228349,
  62.53919, 51.51494, 62.72518, 45.48926, 14.68581, 10.9688, 10.12974, 
    1.36328, 0.2758661, 0.2082997, 0.3471243, 0.8529164, 2.091373, 2.453037, 
    2.797,
  73.36969, 59.65648, 49.83633, 47.68164, 26.11435, 8.893585, 5.215225, 
    3.406776, 0.9360161, 1.153316, 0.2727052, 0.5604218, 1.179755, 1.867801, 
    2.812186,
  73.85642, 69.85751, 59.67293, 49.28366, 57.87881, 36.09228, 2.929753, 
    0.5257015, 1.314473, 2.111635, 1.029456, 0.4297367, 0.6258087, 0.750742, 
    1.669497,
  65.48328, 65.07365, 59.5294, 50.8446, 61.0148, 52.30626, 7.315322, 
    0.9297743, 2.25244, 1.496498, 0.447577, 0.8896948, 0.2274915, 0.2583407, 
    1.781682,
  52.554, 56.53284, 52.99469, 41.20096, 40.08561, 17.01281, 0.8471344, 
    1.373711, 1.865311, 1.322642, 0.1417222, 0.9669469, -0.006519757, 
    0.08748209, 1.892817,
  45.02328, 42.18379, 29.76134, 8.988804, 4.740166, 2.59306, 0.3842889, 
    2.5689, 0.5976768, 0.08462161, 0.8771222, 0.396146, -0.02472048, 
    -0.06328566, 1.138373,
  2.300995, 2.361568, 2.426171, 2.753386, 3.254011, 1.419723, 0.3907295, 
    1.480547, 6.723227, 2.931984, 2.458729, 4.384097, 3.375063, 2.510935, 
    0.3267907,
  3.477895, 2.291207, 2.419004, 5.856915, 5.035282, 0.738941, 0.3723212, 
    0.6994641, 2.767679, 5.497154, 2.627797, 7.957488, 8.407701, 0.2391775, 
    0.5286603,
  8.39947, 6.221568, 8.420113, 12.41463, 13.57286, 1.054223, 0.8038583, 
    0.3653117, 0.5799308, 0.7570009, 1.852075, 4.971475, 5.331409, 5.89567, 
    1.715951,
  23.42164, 32.53154, 37.64045, 18.74732, 14.3918, 13.952, 1.054239, 
    -0.03430216, 0.07490564, 0.4031581, 1.061761, 2.234338, 2.754371, 
    2.228328, 1.192048,
  29.22384, 32.09546, 52.83768, 34.63951, 11.39, 10.87491, 16.20868, 
    0.3930405, -0.3128931, -0.04455961, 0.04794206, 0.5209416, 1.378732, 
    1.50446, 1.38361,
  33.18467, 39.53269, 48.71627, 40.64257, 21.31288, 9.947336, 10.56124, 
    9.979589, 4.886375, 4.122796, 0.1381256, -0.05657944, 0.50638, 1.328853, 
    1.624983,
  31.35317, 51.01718, 57.55498, 46.51522, 44.36878, 31.41408, 6.657743, 
    1.979375, 3.734653, 4.597652, 1.683388, 0.1253376, 0.443267, 1.001837, 
    1.754642,
  34.6623, 55.59682, 60.47985, 49.39672, 53.44055, 46.13645, 12.62778, 
    2.198033, 3.163447, 2.047927, 0.444139, 0.505592, 0.1049719, 0.451748, 
    2.535789,
  35.42574, 56.28335, 61.58158, 46.97224, 45.6629, 29.00507, 5.040436, 
    2.841676, 2.768405, 0.8075979, 0.3009181, -0.003995119, 0.002969628, 
    0.3315992, 2.392484,
  28.99605, 37.72072, 36.60376, 9.796973, 2.215836, 4.19385, 3.002904, 
    4.589749, 1.887634, 0.1943022, 0.1585017, -0.03325316, -0.004004086, 
    0.03311896, 1.416927,
  4.883693, 4.102324, 2.75677, 3.156696, 1.764416, 0.9792817, 0.6125085, 
    0.4776635, 3.001575, 2.534261, 3.342364, 5.290596, 2.974765, 1.283951, 
    -0.6221771,
  8.595101, 4.666385, 3.254221, 5.106872, 2.499079, 0.4799702, -0.3225281, 
    0.04333827, 2.159887, 4.401349, 3.655995, 8.066654, 10.38057, 0.1424071, 
    -0.6209782,
  16.4099, 3.804045, 5.426168, 9.423949, 8.677708, -0.09701408, 0.3049491, 
    -0.01387185, 1.294527, 2.577166, 5.258713, 6.871713, 8.670003, 8.689172, 
    2.520248,
  37.11533, 34.73862, 30.98181, 19.57974, 10.09529, 7.470888, 0.6704596, 
    -0.09582085, 0.204854, 1.528606, 3.874446, 6.405844, 7.001568, 6.043038, 
    3.018545,
  43.14322, 40.28235, 58.90965, 41.12901, 5.278722, 4.867928, 12.01766, 
    1.32122, 0.4448565, 0.9084683, 2.130006, 4.247341, 4.700891, 4.641981, 
    3.063535,
  57.99453, 58.21171, 59.69763, 44.87881, 11.50875, 4.056562, 5.896285, 
    11.05785, 9.159115, 8.26519, 2.153447, 1.914432, 2.184474, 2.585407, 
    1.674746,
  77.95793, 83.74498, 78.25047, 47.58453, 29.50572, 22.99711, 9.364751, 
    8.816206, 7.301561, 7.467116, 4.714387, 2.329598, 0.4463904, 0.8447622, 
    1.690895,
  96.53639, 92.40634, 79.69035, 48.04139, 43.52765, 48.53591, 17.44327, 
    8.275489, 5.465236, 3.684618, 2.09626, 1.249537, -0.2039489, 0.5911705, 
    2.086097,
  101.4362, 96.08561, 76.37713, 50.45122, 52.06279, 35.97363, 12.98441, 
    6.783604, 3.196595, 1.024756, 0.5562966, 0.151096, -0.2694436, 0.5284119, 
    1.919554,
  92.11091, 81.27283, 60.18583, 14.59058, 2.935287, 7.479004, 8.520308, 
    5.169296, 1.781313, 0.2967876, 0.1051744, 0.09877828, -0.08473895, 
    -0.007272923, 1.223932,
  4.668708, 6.849855, 6.42121, 4.674072, 1.564188, -0.4880522, 1.817666, 
    2.882821, 4.445787, 1.952995, 1.410568, 2.08726, 1.137238, 1.258354, 
    -1.472813,
  5.830475, 5.749892, 6.120476, 4.86586, 1.267497, 1.021889, 2.18447, 
    2.672678, 4.02611, 2.684999, 1.278315, 4.809789, 7.477136, -0.2392289, 
    -0.9640595,
  12.61083, 7.921938, 7.337439, 7.754283, 11.44298, 2.194594, 2.004274, 
    2.018594, 1.302177, 0.416637, 1.478555, 3.886358, 6.639899, 8.897132, 
    3.867942,
  45.0276, 45.25999, 36.8357, 20.71714, 19.51031, 14.38188, 1.345029, 
    0.5466756, -0.3194268, 0.2642373, 1.390062, 3.589552, 6.200471, 7.13942, 
    5.556482,
  66.96138, 59.03704, 72.73389, 46.94592, 19.1413, 15.72889, 15.72932, 
    1.909995, 0.05380915, 0.4565151, 1.845281, 3.449103, 6.069872, 7.640751, 
    8.031403,
  92.7716, 84.33831, 75.89066, 59.0121, 31.71758, 13.84073, 13.14981, 
    10.5321, 5.652829, 5.240585, 2.508447, 3.575984, 4.628502, 6.024165, 
    7.255136,
  108.2574, 102.4792, 90.29147, 67.28561, 60.00935, 43.19684, 12.60972, 
    9.185802, 6.617886, 6.565799, 5.173086, 4.316753, 3.711812, 4.717747, 
    6.422554,
  113.3079, 105.3056, 94.24276, 79.52562, 79.60015, 68.40063, 16.88849, 
    8.494495, 6.281794, 4.512864, 3.977029, 3.2905, 1.600385, 3.010233, 
    4.502589,
  101.4707, 101.2459, 94.47416, 80.59113, 76.22179, 46.33571, 13.42437, 
    8.170601, 4.79352, 2.746018, 1.702099, 1.517549, 0.1362019, 1.77257, 
    2.112885,
  77.76922, 77.12516, 65.1589, 26.04194, 6.098595, 9.766381, 8.691834, 
    6.603673, 3.535313, 1.08321, 0.1616936, 0.5088454, -0.08313687, 
    -0.08930721, 1.293219,
  3.100008, 4.099173, 6.133759, 9.541554, 11.57551, 3.299335, 2.485725, 
    4.432418, 5.736284, 3.638894, 3.029941, 5.889144, 3.796546, 3.29522, 
    0.6332447,
  3.844487, 3.429998, 3.371543, 13.66193, 10.21906, 2.997845, -0.01868136, 
    0.5383117, 0.9276854, 1.661077, 0.5970407, 4.462331, 6.04478, 1.800521, 
    -0.12504,
  18.28401, 3.608126, 3.580051, 11.68506, 14.95634, 0.971024, 0.6138013, 
    0.6070004, 0.6556183, 0.3046237, 2.065961, 4.49679, 6.315914, 8.341487, 
    4.436844,
  55.13063, 65.32529, 52.32653, 20.45237, 23.38254, 17.97648, -0.3967291, 
    0.05149603, 1.182914, 0.5454715, 1.085775, 3.531743, 6.041306, 8.475038, 
    6.699168,
  65.88514, 68.60415, 83.06216, 43.74836, 17.27627, 24.22329, 20.22432, 
    0.6013698, -0.9046689, 0.2042826, 1.848462, 1.869702, 5.392762, 8.379976, 
    8.711992,
  72.3456, 73.88579, 77.43362, 59.28424, 28.77593, 20.93573, 23.71957, 
    18.85182, 8.196144, 3.396592, 0.7246168, 1.143585, 3.290339, 5.237389, 
    5.163613,
  71.78493, 80.18375, 86.14674, 77.00641, 73.81576, 45.456, 18.44542, 
    14.23652, 8.536168, 4.510201, 2.040801, 1.824845, 2.559567, 3.656407, 
    5.05996,
  69.10917, 74.71553, 80.36491, 85.32169, 95.73299, 73.33387, 15.44874, 
    10.08299, 7.975521, 4.980104, 2.257447, 2.261472, 1.797465, 3.897358, 
    5.665244,
  66.03913, 69.08877, 68.91737, 68.62911, 70.60031, 35.88372, 10.60319, 
    8.452637, 7.003137, 4.869344, 2.687916, 3.006421, 2.758023, 4.521598, 
    4.214575,
  59.67851, 55.26898, 42.98279, 16.29581, 4.988076, 5.49485, 6.567346, 
    7.42759, 5.244138, 1.516068, 0.5355871, 1.759651, 2.141913, 2.268962, 
    2.770617,
  3.786617, 0.8278634, 0.7791872, 0.9905252, 3.362811, 1.338477, 0.3684489, 
    0.471951, 1.658003, 0.2158145, 1.808434, 2.153279, 1.414801, 0.9828026, 
    1.637991,
  5.184176, 0.4311159, 1.231067, 2.838351, 4.474618, 0.7996763, 1.079712, 
    0.1315162, 0.7755572, 1.087053, 0.5803766, 3.663506, 3.790093, 0.1825817, 
    1.220953,
  9.171069, 1.749374, 2.905763, 4.618219, 8.355799, -0.2220231, 1.362524, 
    2.495358, 1.674017, 1.714796, 2.648196, 5.009607, 4.799857, 3.159851, 
    4.934968,
  28.12668, 38.21116, 38.48243, 8.401937, 15.37255, 10.99036, -0.4236094, 
    1.446497, 2.675229, 2.81153, 5.121954, 6.299585, 6.207986, 5.184294, 
    6.591967,
  29.68461, 30.5533, 50.15492, 29.95018, 10.91608, 15.40176, 13.51394, 
    -0.4063004, -0.4143673, 1.774595, 4.856896, 5.330851, 6.795208, 5.870798, 
    8.145043,
  31.01435, 25.59237, 35.26314, 37.00967, 21.02713, 14.27472, 15.00632, 
    8.829243, 3.436631, 3.264296, 0.9343172, 3.404771, 5.817935, 6.173594, 
    6.362609,
  28.70747, 24.5754, 29.88685, 40.75003, 50.58478, 29.75536, 10.84933, 
    6.25296, 3.084437, 2.133439, 1.010957, 1.56967, 3.181698, 3.250814, 
    4.603945,
  28.22808, 20.76215, 21.60999, 38.2442, 57.41748, 43.34024, 7.951873, 
    4.681819, 3.239569, 1.142235, 0.1608018, 0.595297, 1.031427, 1.630651, 
    2.585516,
  24.29605, 18.38501, 15.90413, 24.03548, 42.64967, 17.14012, 5.46073, 
    3.30488, 2.804355, 1.236741, -0.1602671, -0.01561482, 0.2735596, 
    1.143487, 1.990149,
  15.26146, 9.212502, 5.018726, 3.109477, 7.247283, 2.925599, 2.814787, 
    3.641155, 2.274778, -0.02461991, -0.5624911, -0.4997331, -0.1748355, 
    -0.1148544, 1.005016,
  -0.6028699, 1.517733, 7.588304, 5.87142, 2.129146, 0.9563702, 0.3062836, 
    0.4904389, 2.333215, 1.108399, 2.381243, 3.288762, 2.498851, 2.230231, 
    0.06299105,
  -1.633554, 3.61223, 9.695563, 6.872405, 2.585436, 0.8588639, 0.2582201, 
    -0.1892339, 0.5751101, 1.710769, 1.402354, 3.244408, 5.698324, 0.3604001, 
    -0.3354633,
  -5.067599, 6.494913, 12.54507, 8.85272, 7.89408, 0.5430618, -0.05197317, 
    -0.775255, -0.09861023, 0.4866236, 1.725611, 3.204885, 3.079217, 4.05607, 
    2.925479,
  0.2354597, 25.60706, 41.09566, 15.04557, 11.56073, 8.328782, 0.5339527, 
    -0.3435651, 0.3658124, 0.8942069, 2.10204, 2.900415, 3.808108, 3.998188, 
    6.072144,
  10.87835, 26.81026, 61.75676, 38.87823, 14.54752, 13.37702, 10.27526, 
    -0.04838913, -0.5429714, 0.141965, 0.8197838, 2.219501, 6.228166, 
    7.604512, 9.522365,
  27.37496, 32.56651, 51.29385, 59.10408, 31.22532, 17.42676, 15.9252, 
    8.637461, 1.942776, 2.421789, -0.4220669, 1.989762, 6.720506, 7.898459, 
    9.875306,
  40.61568, 49.72939, 64.57462, 78.43969, 76.80183, 39.7756, 15.07228, 
    5.673485, 2.109687, 1.838778, -0.004289802, 0.9692703, 2.682272, 
    4.077904, 6.794394,
  54.3243, 62.11516, 70.81566, 91.73597, 96.19634, 61.8841, 12.95025, 
    6.172598, 2.469671, 0.6730853, -0.2067067, 0.0808302, 0.3139282, 
    2.205702, 3.876223,
  61.07602, 67.85934, 74.40559, 92.56882, 90.46246, 35.54125, 10.48653, 
    5.437595, 2.387531, 0.1851862, -0.6221381, -0.5429806, -0.4323131, 
    0.7340401, 3.911272,
  57.4537, 58.22273, 57.0379, 45.99911, 20.0841, 9.128695, 5.91441, 5.456153, 
    1.472142, -0.9368068, -1.497058, -1.383981, -0.6783106, 0.1359821, 
    2.997884,
  7.318686, 10.84064, 6.729604, 5.433356, 5.80046, 3.105603, 1.86235, 
    0.072451, 0.6814735, 1.068785, 2.127643, 3.146497, 1.831392, 1.042432, 
    -0.3510335,
  18.1126, 10.11779, 8.081397, 6.218411, 4.937365, 2.155654, 2.136831, 
    -0.4588808, 0.0185537, 0.1728484, 0.7100097, 2.375489, 3.881108, 
    -0.3877048, -0.7312545,
  64.48603, 16.19795, 10.12402, 10.46791, 9.678364, 0.2211054, 0.4764669, 
    -0.1013228, 0.8620815, 0.1454703, 1.038417, 2.287936, 2.375898, 3.954909, 
    1.932591,
  93.79971, 83.24054, 54.83145, 18.02868, 22.30338, 15.98337, -0.0486377, 
    1.502033, 3.638739, 3.675715, 2.940939, 2.746523, 3.206758, 4.52855, 
    3.150389,
  106.0666, 91.95938, 94.41954, 42.57404, 23.60519, 23.54159, 20.41924, 
    -0.7922622, -0.6994917, 2.887318, 4.340294, 4.982509, 6.37614, 7.749938, 
    9.141271,
  115.828, 100.4216, 88.0771, 56.97961, 32.03094, 23.11051, 22.86636, 
    17.5422, 5.99636, 4.603033, 1.922287, 3.856361, 5.139132, 5.94202, 
    8.060028,
  118.88, 113.1295, 100.4654, 75.4794, 74.52648, 33.86583, 19.03415, 
    12.30143, 7.055051, 4.925736, 3.489358, 3.458104, 4.065313, 4.14416, 
    5.842474,
  122.9565, 116.7438, 106.7367, 94.69292, 99.78172, 54.39201, 16.28388, 
    10.58971, 6.386002, 3.379349, 2.402856, 3.509658, 2.634903, 4.090534, 
    4.960438,
  122.568, 119.7371, 114.6406, 102.5154, 89.97865, 33.33917, 13.96584, 
    8.226449, 6.879876, 6.010885, 2.381555, 2.111883, 3.20966, 4.418206, 
    8.385304,
  117.5825, 113.7722, 102.4789, 55.98895, 21.13209, 12.99303, 6.482527, 
    13.99813, 7.651762, 2.25122, 0.9960874, 1.873787, 2.331853, 3.847841, 
    9.104542,
  4.824709, 7.36099, 10.97393, 10.15679, 1.943771, 1.522736, 0.2311996, 
    0.5992182, 0.5546879, 0.09974568, 0.5680224, 1.426171, 1.729578, 
    1.943739, -0.1633599,
  5.767891, 2.044913, 9.106802, 10.18109, 5.229106, 0.9267544, 1.111531, 
    0.339122, 1.044386, 0.4706256, 0.6310326, 1.97287, 4.237631, 0.9372703, 
    -0.01042539,
  35.19564, 6.163779, 6.621233, 17.05257, 15.35847, 0.1039428, 1.426925, 
    1.547173, 2.107789, 1.497252, 2.012168, 1.956168, 2.414199, 4.803495, 
    2.814204,
  66.6483, 65.5153, 45.71462, 22.25013, 27.92909, 18.39972, 0.8234559, 
    1.891659, 2.946154, 1.995354, 4.080049, 3.492318, 2.680469, 4.24701, 
    3.700963,
  81.49687, 75.99548, 79.7112, 34.34558, 24.68509, 24.79478, 20.86877, 
    0.06591882, 0.3148839, 0.869074, 2.434841, 3.937008, 3.945552, 4.077097, 
    5.046245,
  91.9594, 84.89751, 76.25156, 50.50771, 34.74559, 23.33096, 19.48069, 
    11.09611, 4.907143, 1.503306, 0.7292252, 1.179138, 5.109678, 4.153013, 
    4.187423,
  99.46354, 101.3562, 94.25571, 76.53255, 79.43056, 32.03046, 17.75087, 
    8.227773, 6.509311, 5.017823, 1.107644, 1.162715, 0.9593285, 2.175733, 
    3.289807,
  105.6655, 109.2395, 108.6018, 103.0275, 106.7792, 48.14185, 16.12048, 
    6.45777, 4.02384, 6.04216, 3.744202, 1.045004, 0.7574002, 1.467597, 
    1.573552,
  107.5763, 113.3946, 117.3164, 112.7635, 79.12921, 28.47614, 17.83411, 
    8.119097, 7.792799, 9.897443, 5.312364, 2.048369, 0.8791103, 1.654514, 
    2.20784,
  102.2295, 106.6313, 95.88714, 41.98183, 15.0934, 15.34169, 12.47494, 
    26.59154, 17.86773, 6.380649, 1.609595, 2.004822, 1.487556, 2.149907, 
    3.25196,
  5.285139, 3.748814, 4.532318, 5.670751, 1.951017, 1.567717, 0.9676319, 
    1.942033, 1.736056, 0.5214776, 1.034697, 1.493221, 0.5350586, 0.8531367, 
    -0.07032847,
  3.874789, 1.433203, 7.987153, 9.625844, 4.591314, 1.996761, 0.9818811, 
    0.806678, 0.9000989, 1.67931, 1.389567, 2.066661, 2.353095, -0.346195, 
    -0.3980517,
  23.67856, 3.11483, 3.092916, 12.88925, 13.72591, 1.472495, 1.136783, 
    0.782811, 1.031044, 0.6069379, 1.105001, 1.425665, 1.550608, 3.219422, 
    1.553978,
  60.72243, 52.48366, 35.67108, 12.34489, 21.27707, 11.33092, 0.4966468, 
    1.433536, 2.455431, 2.05977, 2.28374, 2.009116, 2.139485, 4.279339, 
    2.59477,
  81.73034, 74.71846, 74.13635, 28.47614, 19.03768, 20.13288, 13.91847, 
    0.05407612, 0.15927, 2.811097, 2.334413, 2.023052, 2.065185, 4.141603, 
    5.171132,
  97.16325, 88.22865, 77.59306, 45.52495, 31.71294, 22.08353, 16.25514, 
    5.504369, 3.679429, 2.93278, 1.042741, 2.377719, 1.638199, 3.896314, 
    6.079379,
  106.9651, 105.9587, 100.0325, 76.57029, 79.0815, 28.05847, 15.78863, 
    6.787226, 6.179605, 4.536752, 1.482008, 1.909627, 1.272145, 2.031934, 
    5.441141,
  113.7856, 114.5183, 112.5392, 107.7332, 103.8542, 36.42612, 16.13631, 
    8.977583, 7.422339, 5.15835, 3.166581, 1.516614, 2.199187, 2.147871, 
    4.257576,
  113.491, 115.8434, 116.8499, 104.2326, 55.63613, 18.63796, 13.937, 
    12.13492, 12.72903, 11.72709, 3.98648, 1.05267, 1.265082, 2.042032, 
    4.113522,
  103.6393, 102.1735, 80.69353, 28.0724, 10.85872, 11.35567, 11.11989, 
    37.05957, 25.48475, 10.38622, 1.54705, 1.041537, 1.19467, 1.949237, 
    2.82735,
  7.528659, 6.394569, 4.231641, 3.536368, 4.196097, 2.061661, 0.9271627, 
    1.0963, 1.600368, 1.960997, 3.58461, 4.664391, 3.01344, 2.846281, 
    0.4142387,
  7.993546, 3.666073, 4.593429, 4.009929, 3.723494, 1.097299, 0.591141, 
    1.209564, 1.371129, 2.217343, 3.748157, 6.196518, 6.563229, 2.144306, 
    0.167623,
  29.98208, 4.065713, 5.905755, 6.937643, 7.304817, 0.837226, 0.8524007, 
    0.9684073, 0.9398182, 0.571797, 1.720054, 2.86982, 3.215818, 3.794856, 
    1.58367,
  56.16795, 47.80771, 29.25559, 8.83627, 17.85647, 8.510339, 0.3268602, 
    1.34399, 1.264472, 2.031605, 2.137275, 2.569014, 2.943532, 3.652306, 
    2.143026,
  69.84217, 63.45285, 62.67034, 18.3849, 12.9831, 13.86917, 8.647532, 
    0.2810959, 0.1868224, 3.371208, 4.076894, 2.588528, 1.982133, 2.301776, 
    3.350608,
  68.85592, 63.88346, 55.77436, 31.57676, 22.3257, 14.38694, 10.97648, 
    6.086995, 3.374323, 1.854836, 0.7273425, 1.529891, 1.4074, 2.367737, 
    2.930608,
  65.2249, 67.88283, 66.16308, 51.42847, 56.32231, 17.32176, 9.317806, 
    6.18602, 5.212429, 2.859483, 0.8890572, 0.951853, 1.217256, 1.678709, 
    3.695765,
  63.20224, 68.47717, 71.18243, 71.16914, 67.00467, 19.17788, 8.466969, 
    5.748768, 4.655041, 3.196281, 1.465516, 0.9458634, 1.172117, 1.42414, 
    3.645888,
  56.90355, 62.30481, 68.29637, 60.77003, 28.74366, 9.709247, 6.660195, 
    6.322032, 7.76182, 6.782423, 2.428527, 0.6934484, 0.7310641, 1.998205, 
    3.383957,
  53.20149, 54.14106, 47.03406, 17.78683, 6.719689, 6.276511, 6.546012, 
    29.55685, 18.97895, 5.082357, 0.6260036, 0.4148763, 0.4207712, 1.81785, 
    2.755612,
  4.850502, 3.715029, 3.484643, 3.544889, 2.215552, 1.942088, 0.9461548, 
    0.7573617, 0.8786879, 0.4369748, 1.966389, 3.350972, 1.90194, 1.686576, 
    0.7870319,
  4.418643, 2.230198, 2.574523, 2.493595, 1.313597, 0.8688964, 0.5062152, 
    0.7215922, 1.169587, 0.9094969, 0.8174405, 2.346475, 3.431905, 1.553638, 
    0.589952,
  19.17283, 2.467386, 2.21903, 4.696699, 4.107194, -0.3587637, 0.8172749, 
    0.379269, 0.5776908, 0.3294183, 1.081334, 2.806901, 3.660981, 3.595542, 
    2.56513,
  48.5038, 41.94487, 22.30172, 3.726253, 9.04313, 4.919139, -0.6156572, 
    2.194817, 1.642743, 2.166386, 2.698266, 2.499055, 1.961941, 1.940864, 
    1.495513,
  68.53171, 64.14784, 63.00041, 11.59189, 9.036364, 7.442227, 6.424255, 
    -3.036725, -0.6791197, 3.707416, 8.093385, 5.591036, 3.11158, 3.352319, 
    3.765277,
  93.50875, 76.48975, 53.05798, 22.17395, 18.95177, 12.30842, 10.55849, 
    5.068061, 2.744432, 2.57493, 3.15262, 5.967537, 4.107214, 3.610545, 
    3.426885,
  103.3982, 83.55264, 65.51006, 45.33494, 55.7642, 19.60227, 9.303172, 
    7.491072, 4.532809, 4.384219, 3.814455, 4.630567, 5.097586, 3.406405, 
    3.417827,
  96.2045, 78.97001, 75.01481, 71.02224, 69.97356, 22.80568, 9.395497, 
    7.174377, 5.494128, 4.570037, 3.893882, 3.307354, 3.462529, 3.60433, 
    3.027348,
  81.61256, 79.76242, 84.40027, 69.63884, 32.68226, 13.52172, 10.93357, 
    10.91395, 9.858034, 7.531061, 4.426867, 2.670925, 2.95838, 3.463207, 
    1.479509,
  67.24663, 68.06326, 57.68629, 23.46097, 14.07249, 11.6113, 11.69521, 
    34.65848, 23.66191, 4.731172, 3.336362, 3.559617, 0.9704375, 2.307102, 
    0.9573624,
  0.9883307, 1.080438, 2.087926, 1.615033, 0.9280567, 1.632521, 1.492245, 
    1.016651, 0.9453088, 0.2364622, 0.8729611, 1.32013, 0.4410416, 0.6848392, 
    0.1128265,
  1.147584, -0.4424507, 0.08025589, -0.9951419, -3.003913, 0.1115374, 
    1.604519, 3.298189, 2.180052, 2.305278, 3.106663, 3.923657, 2.331158, 
    -0.3035396, -0.1532522,
  26.84565, 3.562199, 2.241441, 1.216942, -2.826556, -0.5721899, 2.126301, 
    2.373783, 3.18741, 2.602002, 2.426391, 3.298259, 2.470993, 2.180933, 
    1.154505,
  82.90778, 70.49482, 31.53517, 4.000267, -1.025565, -1.420977, -0.4311159, 
    3.820894, 4.620136, 4.683168, 5.768, 3.864054, 3.646432, 4.883905, 3.25469,
  98.5244, 68.93769, 48.5838, 4.014882, 3.235893, 4.230677, 4.589463, 
    -1.161544, 0.9521347, 7.511703, 11.84921, 7.181654, 5.390148, 4.681074, 
    5.515906,
  97.33441, 58.8721, 20.67627, 9.07215, 12.44233, 6.264477, 5.698705, 
    1.713189, -0.1906358, -0.5806182, 2.695682, 7.127763, 6.511882, 6.715789, 
    6.102044,
  89.65833, 54.90863, 33.67859, 33.15928, 46.21794, 11.00114, 3.586214, 
    2.934413, 2.826959, 2.597646, 1.84384, 3.082066, 5.12649, 5.17448, 
    5.056757,
  73.41934, 57.16958, 54.84872, 60.17173, 55.21128, 15.4347, 5.661821, 
    4.381782, 3.741886, 1.890396, 2.127206, 2.873435, 4.616548, 4.212647, 
    3.812542,
  72.06872, 70.02728, 70.35423, 56.86324, 24.97804, 10.44588, 7.571742, 
    9.896577, 11.67283, 16.28549, 8.163043, 3.960906, 4.352692, 4.895405, 
    2.413567,
  70.60476, 66.49147, 50.85108, 18.93768, 10.39917, 9.610326, 10.46256, 
    30.51844, 26.10915, 8.601774, 8.991468, 4.343666, 1.400139, 3.755486, 
    2.476792,
  0.9731301, 0.3718249, 0.5944481, -0.0008970905, 4.73108, -0.2146392, 
    4.833642, 1.365021, 1.886499, -0.6463867, 1.896559, 2.260355, 0.7840748, 
    0.9176442, 0.5169712,
  2.345938, 0.05703383, 0.7144285, 1.329552, -2.375367, -2.578068, 3.094835, 
    2.896504, 3.344388, 3.103351, 5.807034, 7.961399, 6.286482, 2.575931, 
    1.85043,
  50.01178, 9.521712, 6.234345, 4.426964, 0.9193082, 3.002578, 4.479799, 
    5.79635, 3.722157, 3.069706, 2.914883, 5.19529, 5.042544, 4.66607, 
    2.114428,
  90.86244, 87.73253, 53.80875, 5.580637, 1.935054, 6.171917, 2.952215, 
    4.04834, 5.808293, 5.749458, 6.154044, 4.3865, 4.195712, 4.608287, 
    5.199652,
  98.54713, 66.85395, 40.33101, 9.81486, 11.81558, 7.988523, 5.842246, 
    0.9098969, 2.323466, 6.765242, 11.78488, 6.516198, 4.345763, 4.244966, 
    5.628799,
  79.59863, 36.91941, 15.63009, 28.59671, 16.84852, 4.927894, 3.219029, 
    2.435232, 0.8780584, -0.3604071, 2.516979, 5.950199, 5.048316, 4.812806, 
    5.061022,
  50.60142, 25.48916, 47.49709, 30.928, 41.10728, 7.211793, 2.554702, 
    1.62325, 0.5524995, 0.3890103, 0.7336062, 1.855902, 2.628482, 2.395838, 
    1.984065,
  36.35589, 58.81057, 44.98701, 48.31343, 48.42033, 10.02787, 4.772476, 
    2.968031, 2.192621, 1.375933, 1.122221, 2.104425, 2.541085, 1.585461, 
    1.806059,
  70.59795, 63.74699, 58.08544, 46.96217, 19.11234, 9.159964, 6.928482, 
    8.698941, 11.05844, 13.19687, 4.38787, 1.555785, 3.204401, 3.071176, 
    0.3806412,
  82.49471, 67.52493, 46.25892, 15.56119, 8.745009, 9.295753, 7.887672, 
    23.33418, 22.44018, 6.956616, 7.362689, 1.682884, 0.2022299, 2.53904, 
    -0.007378838,
  5.937538, 6.305572, 4.322502, 1.37244, 0.4938816, 2.232822, 6.728917, 
    3.513563, 2.310299, -0.1696083, 0.5774165, 0.8316671, 0.7628711, 
    2.716136, 3.166397,
  10.15029, 6.882953, 3.916265, 2.202524, -0.3775803, 2.123917, 1.172223, 
    0.1699456, 0.1096677, 0.4884017, 0.2179096, 0.5167186, 0.5133069, 
    0.9974283, 2.193728,
  32.30763, 8.938284, 4.997713, 3.744852, 2.790122, 2.523584, 0.8112922, 
    0.4831456, 0.7020801, 0.6576236, 0.6626107, 0.6423431, 1.031002, 
    0.7739263, 1.23676,
  61.75907, 62.84497, 57.62858, 16.16411, 4.974273, 3.053246, -1.258246, 
    1.622446, 2.007194, 1.833875, 2.215497, 1.755143, 1.460495, 1.364617, 
    0.2636522,
  75.89421, 64.36103, 63.16822, 13.20879, 3.478745, 3.635364, 1.148712, 
    -0.5745736, 0.1228955, 4.144567, 8.117682, 3.797458, 1.883925, 2.058336, 
    2.464998,
  86.72151, 65.62926, 41.11961, 14.62837, 6.465036, 0.06917249, 0.6121171, 
    -0.4347376, -0.7761884, -0.4424909, 1.169821, 3.514153, 3.192312, 
    3.01385, 2.162414,
  86.30855, 67.12823, 44.52944, 22.28353, 22.30773, 1.601747, 0.6238034, 
    1.403731, 1.563106, 1.124226, 1.707807, 2.929781, 3.860103, 3.299892, 
    2.565926,
  73.81803, 57.89239, 47.14967, 33.546, 27.23651, 4.136489, 2.854042, 
    2.883674, 3.079797, 2.047841, 1.743688, 3.00709, 2.941306, 2.300826, 
    2.7495,
  41.11039, 50.84583, 51.38219, 32.77885, 11.30726, 4.892712, 4.407865, 
    6.478714, 10.13997, 9.852685, 2.731486, 2.267623, 2.943807, 2.964318, 
    1.881067,
  43.9267, 43.85178, 33.46407, 13.50219, 6.12682, 4.515655, 5.150437, 
    17.63333, 20.0165, 5.965184, 3.730931, 0.5237694, 0.5839024, 2.784193, 
    1.476701,
  4.716744, 5.15873, 5.023942, 3.104895, 0.8585042, 1.295869, 1.875245, 
    0.1399084, 0.7526517, -0.8215626, 1.085841, 1.784386, -0.1293641, 
    -0.3273894, -1.772853,
  7.652506, 4.632188, 4.495714, 2.033956, 0.1771537, 2.586056, 2.002676, 
    0.438918, 0.3748494, 0.1798149, 0.239587, 1.287245, 0.4279779, -1.470806, 
    -1.374268,
  24.22955, 7.904748, 3.989346, 4.262218, 4.585125, -0.4632673, 2.7005, 
    2.266011, 0.3769006, 1.114024, 1.930316, 2.288854, 1.470774, 0.7912278, 
    0.9378165,
  46.94034, 50.07157, 49.91345, 22.43657, 7.497532, 9.0791, -0.6240214, 
    2.261029, 1.873767, 1.978017, 2.959969, 2.696462, 1.85055, 1.157654, 
    1.458593,
  62.23387, 50.99144, 59.05331, 28.79849, 6.445056, 9.406315, 6.402256, 
    -1.937499, -0.1424298, 2.633765, 6.570449, 3.040801, 1.246931, 1.897202, 
    2.38096,
  73.37996, 54.73251, 45.51503, 26.72418, 12.63119, 4.181505, 5.687135, 
    4.26251, 4.134654, 0.6237935, 0.7576794, 1.810121, 1.116924, 1.523118, 
    1.754822,
  75.60751, 63.11632, 50.83038, 31.43295, 32.04863, 3.669123, 1.02432, 
    2.205846, 1.615041, 1.394648, 0.8756307, 0.6465906, 2.20112, 2.300049, 
    1.341564,
  69.10398, 58.81414, 48.24575, 38.92723, 38.5776, 3.467721, 1.056533, 
    1.180803, 1.374444, 1.430549, 1.287225, 2.959297, 2.857121, 1.89502, 
    2.679203,
  53.11034, 50.70695, 49.35711, 33.62244, 7.25505, 3.367058, 3.898704, 
    4.408228, 5.396223, 4.584219, 2.288461, 2.147559, 2.836077, 2.42025, 
    2.14142,
  44.85237, 25.95175, 12.12912, 4.15855, 3.569469, 5.166556, 6.632286, 
    12.37117, 13.51073, 3.3563, 2.059081, 1.16374, 0.6117242, 2.053012, 
    2.510128,
  6.97179, 8.473328, 8.260953, 5.159526, 1.460864, 0.6100988, 0.8795227, 
    1.771169, 2.005049, 1.585453, 2.990865, 6.755682, 4.187778, 4.967916, 
    3.692251,
  8.316617, 6.118778, 5.469402, 2.414379, 0.6564699, 1.927669, -0.005417849, 
    0.3062019, 1.475075, 3.128104, 4.676201, 7.802202, 6.978359, 2.775382, 
    1.695737,
  22.8042, 3.610071, 3.28747, 4.549757, 4.110651, 1.535806, 1.409869, 
    0.4414407, 1.460404, 1.504868, 2.043373, 1.789398, 2.789864, 3.577061, 
    1.901496,
  35.06679, 34.22791, 28.98119, 11.14366, 7.434839, 6.978791, 0.7153062, 
    2.297671, 2.45806, 1.975387, 1.675732, 0.898307, 1.349121, 0.9254077, 
    1.78077,
  41.42165, 36.4784, 31.88983, 16.23014, 5.469238, 7.300159, 7.673354, 
    -1.930296, 0.2869052, 1.649423, 4.871013, 2.460362, 0.5047768, 0.4857584, 
    0.951097,
  45.69893, 37.05814, 27.4302, 20.39886, 11.64172, 4.725463, 4.656454, 
    2.833184, 0.4889927, -0.317599, -0.2745006, 0.2992582, -0.2118175, 
    0.2882505, 0.002054538,
  57.77436, 46.85925, 40.49239, 30.85232, 32.06718, 8.104975, 2.837595, 
    1.354684, 0.1502484, 0.3110676, 0.1542378, -0.3374955, 0.0561825, 
    0.1999422, 0.5067286,
  78.8204, 68.29929, 58.79893, 52.65309, 53.32987, 10.42849, 4.308452, 
    3.116583, 0.6559739, 0.01720612, -0.4419246, 0.4286579, 1.429446, 
    1.589608, 1.515105,
  98.53683, 89.17432, 79.13008, 58.35683, 22.4869, 10.74093, 8.84655, 
    8.79024, 7.067042, 5.513819, 1.862811, 1.502138, 2.039402, 1.027941, 
    0.6656837,
  110.308, 91.95644, 61.11036, 19.84615, 12.55558, 11.50317, 9.01223, 
    18.86876, 11.08036, 1.67197, 0.4682118, 0.1905358, 0.3666477, 0.6135273, 
    0.6356544,
  4.160027, 4.586697, 9.274728, 6.514206, 2.463774, 2.553691, 7.729863, 
    8.158063, 8.617881, 6.990738, 5.269188, 7.040046, 3.040633, 2.628419, 
    2.057083,
  5.9206, 7.300184, 7.599895, 1.958245, 0.1929478, 4.213069, 3.194656, 
    0.5248065, 5.277707, 6.823534, 8.679059, 8.500693, 7.858272, 1.363165, 
    0.6219943,
  34.10173, 12.72907, 8.381871, 6.48763, 4.394839, 2.839454, 4.089733, 
    3.230683, 0.9589726, 2.077628, 2.419225, 0.2166737, 0.780066, 0.7741818, 
    1.293822,
  67.16784, 68.35654, 60.66537, 25.75596, 9.567767, 4.60991, 0.568832, 
    2.690186, 1.635064, 1.279318, 0.1596563, 1.001941, 1.102104, 2.173998, 
    2.032252,
  87.58175, 78.82859, 84.49123, 35.95831, 13.20619, 10.95598, 6.161593, 
    0.5783809, 0.919099, 1.735943, 3.440017, 2.176421, 1.561654, 1.761667, 
    2.764574,
  105.3115, 91.21653, 80.16167, 43.32114, 20.22636, 12.52642, 9.941882, 
    6.54377, 4.744534, 3.474154, 1.999701, 2.883343, 3.101236, 3.236555, 
    2.882727,
  117.1913, 109.4801, 96.55862, 59.02219, 48.62256, 13.11574, 10.5133, 
    10.27842, 9.769902, 8.219139, 6.374357, 5.451779, 5.492411, 4.931026, 
    5.349729,
  120.2549, 114.2906, 102.5718, 93.68229, 77.98672, 14.50444, 11.30259, 
    9.434158, 9.124426, 6.689562, 5.285571, 6.235288, 6.103418, 6.042924, 
    5.719238,
  115.2013, 108.8004, 98.85052, 71.91947, 24.57799, 10.55879, 8.438096, 
    8.537345, 6.769842, 3.087331, 0.5262995, 0.9149148, 1.40213, 1.214355, 
    1.253802,
  95.14699, 86.03129, 53.80653, 12.32921, 6.228151, 5.001123, 4.649474, 
    13.61299, 6.894752, 0.6524461, -0.01138695, -0.3360703, -0.239038, 
    0.02891872, 0.3933912,
  1.087937, 0.5502371, 2.494855, 2.709439, 2.88655, 7.075269, 10.79565, 
    6.303271, 4.697691, 7.727278, 7.229247, 8.51133, 5.3558, 4.655726, 
    4.367366,
  1.186525, 0.7194525, 0.1631539, 0.4477427, 0.7069143, 8.748765, 9.388798, 
    4.212044, 1.042505, 1.353114, 4.371141, 6.715565, 5.072834, 2.170435, 
    1.075122,
  38.68798, 6.668305, 0.7481418, 0.4266492, 0.9455038, 3.376653, 9.760843, 
    5.682912, 3.906456, 3.023446, 3.736398, 4.975507, 2.466371, 1.833511, 
    0.4495694,
  77.21099, 70.94633, 52.10038, 13.55392, 2.98498, 4.146758, 0.8062451, 
    5.267113, 8.747134, 6.261388, 5.449243, 4.593559, 3.762469, 2.788573, 
    1.105057,
  93.76833, 73.91801, 67.0296, 18.49985, 6.222656, 8.15122, 7.78415, 
    0.3124375, 2.524092, 6.572063, 9.203359, 6.60309, 4.984631, 4.334185, 
    3.385242,
  93.72858, 74.17405, 53.06562, 21.11496, 9.845778, 6.875267, 7.535035, 
    6.788743, 5.722797, 5.614832, 4.187018, 6.670662, 6.715157, 7.412227, 
    6.69558,
  88.13131, 76.49547, 56.48246, 24.27653, 30.01388, 6.949121, 5.279763, 
    6.847844, 6.216441, 5.898899, 4.434446, 4.433773, 5.739051, 6.188897, 
    7.376545,
  74.07816, 58.66056, 42.25734, 66.39984, 57.41656, 6.07821, 4.263055, 
    4.46616, 3.709394, 2.858965, 2.047588, 2.513915, 2.471574, 3.620574, 
    5.566427,
  67.51485, 65.70714, 84.43806, 81.95083, 20.57637, 4.356122, 2.942687, 
    3.10084, 3.847634, 3.172922, 1.464911, 1.603256, 1.19395, 1.342769, 
    3.461938,
  82.10021, 78.16814, 65.34999, 21.83143, 5.399924, 3.125486, 3.221883, 
    9.057036, 6.59949, 1.109305, 0.6091262, 0.334787, 0.008506588, 0.3605321, 
    1.632255,
  1.322678, 2.123792, 4.164842, 1.45896, 0.1275659, 1.275448, 3.170033, 
    0.2886815, 0.3526458, -0.5833734, -0.02441043, 1.19933, 0.6495506, 
    2.139575, 4.482076,
  2.004382, 1.065488, 0.82715, 1.055127, 0.1638094, 3.297366, 2.101003, 
    1.19283, 1.016736, -0.8883684, -0.2899148, 2.267725, 1.556001, 1.672394, 
    2.486608,
  20.76229, 6.926438, 1.915214, 0.9570093, -0.9160673, -0.5248804, 2.632175, 
    2.391387, 0.7001362, 0.7465469, 2.368631, 2.968931, 2.688945, 1.759952, 
    1.281275,
  52.56932, 46.48169, 35.14451, 10.84596, 0.008860965, 1.114074, 1.039699, 
    1.745105, 4.272821, 4.754217, 4.791212, 3.457026, 2.749883, 1.821966, 
    0.2042372,
  57.83919, 50.79058, 55.99577, 19.45569, 3.152509, 5.920071, 5.189651, 
    1.926142, 2.1653, 3.2871, 5.228909, 3.670093, 3.08927, 2.001475, 1.291043,
  61.54322, 58.44996, 56.14491, 29.19585, 14.9017, 10.02247, 9.925682, 
    7.393608, 3.434526, 2.151645, 2.227674, 3.555789, 3.3797, 3.006686, 
    2.56038,
  113.4034, 115.3435, 112.5219, 55.87261, 40.82108, 16.86116, 9.284957, 
    5.330311, 2.749285, 2.105038, 2.292758, 2.582649, 2.464363, 2.92193, 
    3.576437,
  156.6646, 149.8633, 134.1249, 116.2657, 61.83635, 11.46171, 6.065669, 
    3.593014, 2.851645, 2.393826, 1.940459, 2.080788, 1.718402, 2.610148, 
    4.372986,
  163.4815, 149.9184, 129.3388, 80.72134, 20.38715, 6.987159, 4.35626, 
    3.694618, 3.95719, 2.878648, 1.718822, 1.66307, 1.781418, 2.466476, 
    4.158681,
  125.4008, 112.473, 69.33456, 14.86604, 5.665285, 3.968363, 3.669911, 
    11.19304, 7.143874, 1.125681, 1.848114, 1.51351, 0.8254482, 1.380596, 
    2.654655,
  5.184154, 10.4012, 10.77939, 9.504035, 7.414597, 2.779443, 2.981009, 
    2.123757, 4.128672, 3.467206, 5.337275, 10.59754, 4.972414, 3.905413, 
    1.762937,
  7.894533, 8.907721, 10.39915, 13.3287, 14.8465, 6.441638, 3.543865, 
    2.539921, 3.764867, 6.645877, 4.420756, 7.599854, 6.510765, 2.572308, 
    1.181229,
  37.23787, 15.28241, 11.211, 11.98707, 13.49964, 3.548388, 5.228603, 
    3.852262, 2.266169, 4.876801, 5.858673, 3.640619, 3.482469, 4.444963, 
    2.321303,
  57.7307, 65.20927, 61.71103, 23.10632, 9.518402, 10.15612, 4.798563, 
    7.395302, 6.540289, 5.315745, 3.676048, 1.688911, 1.328981, 0.9034364, 
    -0.45923,
  68.54419, 64.70197, 74.61343, 29.72099, 6.875449, 9.50428, 15.07704, 
    3.985679, 2.78906, 2.125562, 3.616982, 2.045898, 0.8453902, 0.618242, 
    0.06585244,
  89.91651, 84.39545, 78.36874, 33.69728, 16.89509, 8.43806, 5.777116, 
    8.467237, 3.862755, 1.954482, 1.080285, 1.574874, 1.091559, 0.857919, 
    0.5204855,
  87.26546, 85.96262, 74.09392, 28.8024, 18.84216, 9.258579, 6.515335, 
    3.654363, 1.977989, 1.90059, 1.248518, 1.052168, 1.68168, 1.940245, 
    1.727611,
  71.01513, 66.08773, 56.71876, 44.078, 20.69141, 4.428043, 2.994734, 
    2.452662, 2.055293, 1.857108, 1.264445, 1.397522, 2.086542, 3.055534, 
    3.587206,
  75.5746, 69.63298, 63.84282, 42.48516, 8.238497, 3.532988, 2.650404, 
    2.459729, 2.599751, 3.948255, 3.874433, 1.754641, 1.297025, 2.39574, 
    2.31244,
  79.90501, 73.75326, 51.54237, 7.170615, 2.753691, 2.272519, 1.244608, 
    3.555784, 3.171737, 1.601562, 5.797743, 1.697822, 0.2161006, 1.504457, 
    1.338078,
  5.851404, 13.20418, 16.44506, 15.28454, 14.6142, 3.842422, 4.016097, 
    5.644266, 6.84875, 6.248717, 7.576801, 12.18638, 8.225635, 2.43858, 
    3.033328,
  9.915243, 13.24953, 14.95967, 30.32431, 22.57847, 4.938068, 1.045076, 
    2.117066, 4.871033, 7.795453, 6.738258, 9.12789, 6.512569, 2.008884, 
    1.710109,
  53.41221, 28.18104, 23.4825, 33.03344, 23.83605, 3.751148, 1.007419, 
    1.261094, 5.000661, 8.00227, 7.346055, 4.552041, 4.584992, 8.037123, 
    7.970729,
  71.89898, 88.29851, 91.24792, 39.72113, 28.10325, 16.43694, 2.760245, 
    1.764783, 2.888948, 3.06766, 4.569711, 1.738808, 2.891261, 3.211987, 
    7.824443,
  70.21291, 72.31601, 89.29205, 32.82484, 23.36751, 24.63191, 17.59468, 
    3.179342, -0.2781606, 0.7787404, 2.686516, 0.860285, 1.071338, 1.739503, 
    4.169616,
  65.64422, 57.68931, 52.61151, 18.61243, 18.2989, 20.36704, 20.97094, 
    14.21741, 5.968769, 2.898597, 1.31937, 0.880502, 1.426054, 0.9842529, 
    1.865098,
  76.19357, 59.34848, 40.23378, 11.54833, 13.58963, 14.43704, 13.95962, 
    12.59019, 8.639886, 6.38184, 2.492861, 1.307615, 0.6327702, 1.427597, 
    1.457496,
  92.66783, 80.41936, 60.19171, 32.58891, 17.2213, 5.543457, 5.75283, 
    7.59988, 6.143927, 5.305562, 3.598323, 2.052817, 1.00524, 1.800457, 
    2.500075,
  101.7919, 96.35878, 82.41, 46.24577, 13.48097, 6.551675, 3.274623, 
    3.040076, 4.224718, 3.941929, 3.068573, 2.313309, 2.020118, 2.091336, 
    2.545387,
  43.8055, 32.34571, 21.28072, 10.35725, 6.668612, 8.396729, 3.748792, 
    1.919505, 1.570578, 0.6406033, 3.366325, 2.187899, 1.864318, 2.50037, 
    2.031224,
  1.531133, 1.078259, 2.166166, 5.020624, 24.80695, 10.7894, 1.730217, 2.646, 
    3.578845, 8.81739, 12.06463, 11.94094, 9.388659, 5.345649, 3.855946,
  4.27143, 1.388392, 0.7295358, 10.44947, 16.83053, 6.329895, 2.575503, 
    3.221339, 2.417585, 9.235346, 11.00083, 12.76283, 6.618962, 3.8243, 
    1.709981,
  26.33061, 7.19471, 3.86634, 10.91765, 10.74065, 4.377716, 2.980933, 
    2.326699, 4.81414, 6.522428, 8.287464, 6.203538, 6.112091, 6.437729, 
    5.59505,
  43.12186, 38.46487, 39.32754, 10.57838, 12.69277, 7.998024, 4.695981, 
    5.230376, 3.96837, 4.190134, 3.597017, 1.417874, 3.909355, 6.143681, 
    5.734393,
  59.8429, 37.107, 36.77884, 5.175008, 9.876561, 12.51432, 3.893995, 
    4.322541, 2.673418, 0.5866979, 1.57855, -0.3351623, 2.769705, 3.489688, 
    6.016744,
  78.05318, 51.55544, 26.15628, 2.517675, 7.235917, 10.72631, 4.998803, 
    2.171864, 1.87915, -0.5414635, -0.8197181, 2.417581, 3.076067, 2.113792, 
    4.155154,
  94.60332, 74.64199, 43.17618, 7.033528, 3.389569, 8.188538, 6.419537, 
    1.097793, -0.4420864, -0.1226995, -1.412983, 2.751209, 3.276476, 
    4.453021, 5.794816,
  111.61, 94.80289, 64.3786, 27.8003, 5.338083, 4.460488, 4.417305, 1.829085, 
    -2.195684, -1.939556, -1.044423, 3.510343, 3.380529, 5.304296, 7.525681,
  127.5346, 107.7408, 79.80571, 30.31748, 7.05999, 8.330577, 2.790274, 
    2.4511, 0.5983832, -2.34073, -0.169365, 3.622088, 3.47604, 5.041762, 
    6.43079,
  129.3702, 115.8463, 69.93726, 18.05674, 3.920355, 6.157795, 4.409606, 
    1.657547, 1.06208, -1.023567, -0.6063229, 3.086423, 2.970793, 5.792549, 
    8.417458,
  5.392992, 7.10312, 3.074578, 6.214971, 2.285697, 0.7410472, 1.285361, 
    2.60697, 4.831236, 8.151539, 3.879118, 4.88413, 3.487341, 2.410195, 
    -0.5805813,
  16.40239, 14.25385, 9.361386, 3.60464, 2.660492, 1.492021, 0.7564152, 
    2.965994, 6.046965, 1.662202, 5.078314, 6.192488, 10.1504, 8.287816, 
    -1.121171,
  75.39969, 38.81816, 16.89114, 9.479999, 1.251772, 0.05498458, 0.7237055, 
    0.7998354, 3.286242, 3.496372, 7.28543, 8.154481, 8.127668, 7.254055, 
    5.121826,
  109.8681, 109.6727, 86.02099, 22.42844, 2.689581, 0.5020962, 1.36329, 
    0.7382814, 3.995782, 4.450266, 4.393402, 5.498856, 8.504573, 10.00264, 
    11.47569,
  128.6496, 123.0953, 105.4701, 20.2325, 5.288925, 1.298015, 3.098219, 
    2.579057, 1.46534, 0.6694022, 4.930083, 8.026071, 10.80359, 11.30696, 
    10.86942,
  142.7725, 139.6605, 103.2128, 24.29509, 11.86294, 2.435861, 1.693551, 
    2.382753, 1.892304, 4.232513, -0.2543254, 9.596797, 8.925919, 5.861864, 
    5.736435,
  157.9521, 160.6952, 126.0356, 42.38845, 19.77561, 2.359786, 4.907101, 
    0.7287047, 0.6247162, 6.913689, 3.392831, 5.928944, 5.185967, 6.135111, 
    6.657076,
  169.3437, 174.4378, 143.0173, 100.4274, 33.80375, 1.967181, 1.524508, 
    2.982308, 1.696904, 5.742179, 3.20001, 4.504247, 4.467327, 7.426926, 
    6.019959,
  171.3329, 178.3788, 156.0607, 103.286, 23.03964, 2.740684, 0.8060032, 
    1.635835, 3.783175, 3.993806, 3.11034, 5.055525, 5.987531, 6.888416, 
    5.986832,
  133.298, 124.805, 84.78484, 29.07913, 12.26606, 3.796831, 1.616182, 
    4.667257, 3.680499, 2.796976, 4.250107, 4.159015, 7.561662, 5.71216, 
    7.567675,
  1.544467, 2.087695, 1.32849, 1.990486, 11.02511, 6.896401, 4.661807, 
    8.029529, 12.41466, 10.12422, 9.766298, 7.847055, 9.061702, 11.53012, 
    6.224305,
  7.253767, 3.106004, 1.629433, 3.310472, 11.33531, 4.397444, 3.294017, 
    7.283557, 7.588115, 8.85457, 8.42948, 12.55433, 18.22574, 8.529901, 
    6.996657,
  73.92358, 34.90188, 9.547541, 3.981495, 3.716835, 4.643897, 2.063211, 
    3.504686, -0.1008381, 0.592003, 9.494267, 14.68769, 15.74755, 18.84682, 
    13.68632,
  97.96046, 92.98058, 76.07868, 14.85817, 2.838658, 3.0083, 3.339872, 
    0.4116389, 1.597472, 3.046897, 5.888569, 12.80221, 14.54755, 16.01468, 
    19.0575,
  109.6934, 94.53535, 81.31237, 11.15026, 1.824545, 1.924889, 3.845844, 
    -0.06600938, 1.267144, -0.1293221, 6.003521, 11.82702, 13.16989, 14.8366, 
    16.44559,
  117.7986, 101.7622, 69.66949, 15.64401, 8.895355, 2.968563, 3.800458, 
    6.664581, 3.526735, 8.460585, 2.337968, 12.6455, 12.127, 11.62063, 10.1331,
  119.2155, 112.9171, 87.46294, 35.36578, 13.49704, 2.915179, 2.969805, 
    2.592125, 3.43943, 5.837554, 10.77615, 13.05644, 11.37345, 7.166646, 
    5.22565,
  116.6421, 112.8864, 97.47898, 71.5264, 28.89347, 3.374111, 0.8891766, 
    3.347916, 1.117153, 9.091572, 8.846946, 7.513453, 6.523007, 4.105535, 
    3.021631,
  114.4991, 114.5759, 107.3089, 61.78621, 16.22955, 4.262167, 0.2021916, 
    -0.1026734, 9.336631, 7.213042, 4.49162, 5.055476, 3.388853, 2.729587, 
    3.655685,
  82.12142, 75.05859, 47.63642, 18.78416, 7.271586, 1.327584, 0.2344884, 
    1.018197, 8.299723, 6.774635, 4.337028, 2.243717, 2.545465, 1.809838, 
    4.428433,
  1.07215, 2.990634, 1.643653, 7.7667, 8.169886, 6.258756, 3.197139, 
    9.110783, 9.626805, 6.879174, 6.76707, 11.39769, 8.728559, 8.742643, 
    4.955742,
  4.110196, 1.247227, 1.961161, 8.804523, 9.093617, 2.198006, 2.013281, 
    9.116291, 5.915938, 10.05828, 5.349485, 16.21955, 22.26495, 9.341016, 
    5.438158,
  36.02866, 18.79485, 12.02032, 14.75469, 6.502272, 5.919912, 0.9768114, 
    7.935176, 6.313883, 8.667553, 9.72227, 14.64304, 21.83322, 26.66927, 
    17.70331,
  45.14111, 49.39048, 55.53159, 23.70643, 12.93986, 6.588696, 2.840415, 
    3.640269, 6.120068, 6.319683, 5.342984, 6.809323, 10.93035, 15.52055, 
    23.76548,
  47.79293, 46.02852, 48.23108, 15.38804, 13.18086, 13.74103, 8.534646, 
    1.856274, 1.773016, 3.120964, 4.861354, 3.730255, 6.069005, 7.737846, 
    14.33922,
  50.56912, 45.96446, 36.19939, 16.73396, 15.80511, 15.12319, 16.65932, 
    14.95581, 8.730628, 11.68512, 4.08628, 3.679972, 2.718155, 2.787049, 
    6.132087,
  49.64563, 52.65963, 44.10058, 23.52427, 14.17659, 11.95562, 8.036961, 
    7.536204, 9.145402, 7.958412, 4.912844, 3.292777, 2.619113, 1.997356, 
    2.741044,
  48.1285, 52.27493, 51.41608, 39.34318, 21.06142, 8.852675, 4.766313, 
    4.077987, 3.093341, 3.345087, 2.499325, 2.119914, 1.821534, 1.52589, 
    1.657996,
  47.48716, 50.92958, 52.9671, 30.95028, 15.0258, 7.29037, 3.143961, 
    2.106585, 1.534937, 1.016678, 0.8408984, 1.342133, 1.25219, 1.09655, 
    2.609094,
  33.85039, 29.9387, 20.98465, 11.25379, 10.6791, 8.723095, 2.780656, 
    1.73596, 0.6826808, 0.255316, 0.9457123, 1.00047, 0.9248466, 0.7307764, 
    3.887084,
  5.430496, 2.656425, 2.934492, 2.695522, 3.112795, 2.109907, 1.685515, 
    1.715166, 2.946063, 4.160662, 4.238678, 10.7377, 8.029756, 7.926235, 
    4.019492,
  3.208178, 3.268411, 2.484337, 3.205456, 7.636982, 2.74253, 2.698115, 
    2.278799, 2.954989, 5.987885, 4.638035, 7.836297, 13.70111, 7.139671, 
    4.706598,
  4.990718, 4.701018, 3.815387, 6.47988, 5.666598, 3.025068, 5.159425, 
    3.706108, 3.554162, 3.260877, 3.712324, 6.990311, 12.40148, 13.75058, 
    10.27984,
  7.863513, 18.18764, 25.5132, 9.857221, 7.511977, 6.22355, 3.293742, 
    3.660969, 4.378118, 3.701264, 2.775709, 3.053614, 5.902493, 8.524112, 
    11.24262,
  13.30505, 18.37437, 31.0695, 8.039486, 10.20428, 11.68548, 12.25267, 
    2.740296, 1.357745, 3.55765, 4.567912, 2.160627, 2.568948, 3.682211, 
    9.063853,
  22.20489, 24.66743, 27.89694, 12.48334, 19.25469, 17.38879, 18.50911, 
    18.88975, 11.50199, 9.19774, 4.670687, 3.467453, 1.32446, 1.967883, 
    4.040304,
  31.58784, 39.56049, 46.98375, 37.04245, 26.27177, 15.67152, 15.39475, 
    13.25814, 10.20726, 9.1445, 4.841232, 3.749395, 1.388519, 0.9392329, 
    2.819039,
  46.5642, 55.68031, 61.67252, 64.57757, 47.12326, 13.92815, 11.61231, 
    11.82545, 7.803073, 5.54513, 4.493846, 3.639294, 1.547931, 0.4637979, 
    1.151181,
  58.32315, 67.52096, 76.63924, 42.01188, 23.76044, 13.07598, 9.76196, 
    10.96766, 7.270822, 3.862808, 3.336233, 4.453131, 1.988994, 0.6188375, 
    1.721694,
  48.21098, 49.0313, 39.4785, 18.44148, 15.84967, 11.45533, 9.458151, 
    12.76051, 9.34308, 2.334214, 5.389732, 5.117229, 1.328113, 0.7526156, 
    2.008554,
  4.862671, 8.197927, 8.58928, 8.632913, 12.08425, 14.31383, 14.57296, 
    12.23147, 9.503485, 5.573126, 10.31037, 8.531377, 4.575723, 5.82917, 
    5.33141,
  11.38033, 10.68192, 9.115034, 11.9404, 16.68057, 12.49888, 15.31023, 
    15.16156, 7.696202, 6.596527, 7.246071, 8.8599, 10.04253, 5.111023, 
    5.021148,
  41.60959, 40.50496, 29.06922, 17.08721, 9.410078, 10.21932, 19.55936, 
    17.0442, 7.745421, 3.63822, 6.611332, 8.17079, 10.99574, 13.88164, 
    10.50342,
  58.53876, 72.51099, 89.79483, 36.72615, 12.03507, 10.16941, 5.069192, 
    18.241, 17.22429, 4.563772, 4.84123, 7.222148, 8.264648, 11.50543, 
    15.26337,
  67.08158, 69.72504, 88.20722, 27.65404, 20.45389, 16.30889, 10.45448, 
    2.649469, 11.67313, 11.11186, 3.917963, 4.208713, 7.509652, 11.57795, 
    15.65003,
  70.6562, 75.0041, 74.28895, 28.76848, 35.98701, 32.62075, 20.47143, 
    16.14425, 12.99373, 9.667359, 3.2873, 3.781112, 7.363853, 7.988725, 
    10.21926,
  68.70419, 82.03535, 85.90082, 65.95271, 39.69341, 20.98352, 22.25481, 
    17.77547, 11.06721, 6.039762, 4.676897, 4.187486, 5.133415, 4.950686, 
    4.3149,
  59.83649, 79.86295, 84.36034, 83.53894, 51.52629, 13.90021, 13.1248, 
    15.09265, 14.37841, 12.19771, 2.138852, 5.362439, 4.3734, 1.87194, 
    2.764188,
  48.5408, 67.2935, 73.29723, 35.15401, 18.22858, 9.227415, 9.812243, 
    11.63841, 15.65965, 12.82213, 7.385444, 5.095074, 2.496601, 0.9676537, 
    0.9942026,
  29.4277, 35.61985, 26.37409, 11.10352, 9.293483, 6.310747, 6.168753, 
    19.26593, 19.78505, 9.46373, 4.966846, 3.329596, 1.149862, 0.9561023, 
    1.940352,
  2.185654, 3.295396, 3.503964, 3.447723, 8.101805, 4.47787, 3.723436, 
    3.954555, 7.305046, 7.497001, 6.922509, 6.250088, 3.586005, 2.328387, 
    5.321836,
  2.535334, 4.690339, 2.062159, 4.701542, 9.383555, 3.859227, 5.933184, 
    7.64292, 9.889399, 9.015483, 2.448064, 6.291701, 3.657611, 2.823868, 
    0.7772301,
  16.21359, 15.59737, 10.4349, 4.798595, 2.941506, 2.35494, 11.35046, 
    9.898454, 10.92611, 8.492952, 7.42719, 5.097867, 6.785001, 9.631906, 
    3.802249,
  16.79363, 23.31626, 26.81675, 7.907197, 3.12273, 1.463861, 1.91976, 
    11.26478, 15.83474, 9.535234, 7.461492, 9.086025, 10.63216, 7.373973, 
    8.455014,
  16.04245, 13.17811, 17.91264, 2.595324, 2.914947, 3.576977, 3.357837, 
    -0.3103769, 6.462055, 10.98003, 7.07399, 4.837254, 8.406094, 9.962164, 
    11.3741,
  13.94076, 6.475413, 3.167701, 1.127657, 6.835409, 6.701187, 4.128849, 
    4.526775, 5.044464, 5.089999, 2.231476, 2.95228, 3.548718, 5.330081, 
    8.890325,
  11.70381, 6.611411, 3.073562, 1.799109, 4.011123, 3.124867, 3.117274, 
    3.200021, 3.287116, 3.974345, 4.042793, 4.008316, 3.17822, 3.697816, 
    5.091951,
  15.43057, 8.739462, 2.030895, 0.4710679, 4.360097, 2.315045, 1.774252, 
    2.601051, 2.788431, 3.340801, 3.454815, 2.963329, 2.495057, 1.896265, 
    2.028047,
  23.19872, 16.53645, 5.410735, 0.1140938, 3.086895, 2.917728, 2.303107, 
    3.000983, 3.760577, 3.600348, 2.684103, 2.853504, 1.971998, 1.785691, 
    1.902284,
  15.21884, 6.000307, 0.3392942, 0.3713567, 1.592116, 1.747717, 2.476525, 
    5.436633, 6.106544, 2.042729, 2.198955, 2.966434, 1.117558, 1.100083, 
    3.008123,
  4.507793, 6.86301, 5.147821, 2.755777, 2.012081, 2.085034, 2.11511, 
    1.05248, 1.35888, 0.5587899, 6.969561, 9.258104, 6.281995, 4.162966, 
    1.451036,
  6.183812, 9.754218, 4.660101, 1.411546, 1.346591, 1.002577, 0.7455794, 
    0.4631866, 0.7071003, 1.759782, 4.82418, 10.00292, 11.3067, 6.558167, 
    1.329319,
  9.002967, 9.986646, 7.057298, 3.002881, 1.117365, 3.979897, 1.080436, 
    1.18328, 0.373367, 1.495904, 3.998015, 6.983577, 10.54894, 15.09812, 
    12.20202,
  21.52468, 22.09698, 20.94165, 5.747143, 2.593776, 1.423217, 3.549464, 
    0.8651205, 1.338251, 1.622158, 1.708515, 4.704922, 8.80357, 12.14365, 
    12.63282,
  34.2441, 25.74604, 28.86388, 7.169082, 4.877475, 3.767886, 2.364406, 
    3.569916, 4.280862, 5.741333, 4.442442, 4.020899, 6.24017, 10.1717, 
    14.48308,
  46.60497, 35.63313, 24.53602, 9.387211, 10.76296, 6.795468, 4.529414, 
    3.77472, 3.826755, 3.277727, 1.628566, 1.571759, 2.386353, 7.233619, 
    11.85766,
  56.17752, 50.00061, 35.81004, 23.36695, 16.18975, 8.607845, 6.211532, 
    8.005191, 6.855396, 5.419368, 2.831987, 0.3003073, 2.171335, 5.573012, 
    8.835835,
  62.77597, 56.59643, 42.14393, 30.86049, 20.77591, 11.84206, 8.121896, 
    10.44164, 8.439621, 8.648725, 5.109609, 1.987559, 4.647085, 6.757268, 
    5.511618,
  61.25751, 55.19579, 44.65454, 20.03787, 13.46713, 10.47675, 9.943113, 
    10.45841, 11.98672, 11.83254, 6.711522, 6.034197, 6.319945, 5.124641, 
    2.979795,
  38.60883, 28.02277, 20.69193, 15.30311, 12.83812, 11.47574, 10.09606, 
    13.26868, 14.06204, 8.659932, 6.74556, 4.889194, 3.87467, 1.431709, 
    0.9504742,
  2.881394, 8.736198, 13.43569, 12.6596, 12.33491, 13.23385, 10.20724, 
    4.236462, 6.183592, 5.874156, 7.115574, 6.72578, 6.245918, 7.923496, 
    6.274902,
  0.8198931, 6.426811, 9.886168, 10.39687, 10.20473, 12.32701, 9.75843, 
    5.682397, 5.044305, 5.479272, 5.069458, 7.0643, 8.350929, 6.646269, 
    6.182791,
  -2.507138, 4.088897, 8.592834, 7.73794, 10.32536, 10.64919, 13.75608, 
    9.057183, 9.695284, 9.566417, 10.27078, 7.361718, 6.189159, 10.23969, 
    9.087637,
  -2.75457, 4.646664, 11.53543, 6.039237, 5.519374, 7.121274, 8.064709, 
    8.061245, 10.79648, 15.2914, 13.39247, 9.33596, 6.662205, 5.99086, 
    7.513615,
  -2.929192, -2.343942, 6.967244, 0.9934083, 4.533331, 6.634311, 5.525456, 
    3.982596, 9.795732, 16.60034, 16.47005, 12.16336, 8.337921, 7.250272, 
    8.35574,
  -2.674703, -4.619043, -1.920466, 0.5999869, 9.052237, 6.794258, 5.051827, 
    5.625656, 4.655973, 7.187147, 7.980967, 12.13842, 7.5142, 3.750374, 
    1.771577,
  -3.061074, -1.633921, -2.18662, 0.2911763, 5.815282, 5.542179, 4.532947, 
    5.206798, 4.623103, 6.654486, 11.03862, 10.55909, 10.10905, 4.123791, 
    4.929831,
  0.5909364, 1.360021, -2.063891, -0.9612098, 4.517266, 4.073059, 4.429997, 
    4.882267, 2.24817, 2.862254, 8.471854, 8.299404, 7.926065, 6.675158, 
    6.77227,
  2.667364, 3.077454, 0.6873364, -0.1018106, 2.107971, 3.532266, 4.412507, 
    4.522281, 4.14853, 2.698275, 2.340304, 3.827747, 4.251781, 2.496605, 
    3.103616,
  -3.747858, -3.367479, 0.351918, 5.691972, 5.256416, 4.494318, 4.856214, 
    6.826885, 7.932067, 3.406953, 1.241649, 1.352838, 0.9961576, 1.379219, 
    2.007988,
  -3.062284, 3.353079, 5.820369, 2.249537, 1.7512, 1.697058, 1.234061, 
    1.640337, 5.629883, 11.45099, 9.014266, 10.28798, 9.379801, 3.767337, 
    5.794563,
  -6.996556, 5.169112, 6.317901, 3.405718, 2.094221, 2.586413, 2.136274, 
    1.240597, 1.489426, 2.05731, 8.004048, 9.890061, 9.742509, 5.322901, 
    3.077203,
  -12.67662, 4.059248, 7.69, 6.23035, 2.564513, 4.095087, 1.526637, 1.506197, 
    1.656975, 1.688932, 6.641018, 10.26173, 9.034347, 8.164462, 4.693578,
  -7.615162, 9.710073, 18.90732, 9.88353, 3.875032, 2.061631, 3.018545, 
    2.55638, 3.490787, 5.451431, 6.933038, 5.974592, 7.394292, 7.607588, 
    5.950253,
  0.843915, 6.092087, 22.52425, 11.74532, 7.263287, 2.854669, 2.32328, 
    1.297651, 2.068781, 7.229664, 5.792607, 5.448836, 7.770357, 8.760791, 
    9.24736,
  10.2957, 7.489223, 17.5736, 15.85173, 13.22528, 6.197799, 2.980661, 
    2.775271, 2.047493, 1.933439, 3.072391, 4.21726, 6.752596, 6.585618, 
    7.795026,
  18.32187, 18.67555, 25.89332, 23.99622, 19.82565, 9.215453, 5.70759, 
    3.467103, 2.282207, 2.575821, 3.456251, 3.742357, 5.346025, 6.509552, 
    3.404184,
  25.07792, 27.68949, 31.06569, 26.19583, 23.35193, 11.23616, 7.515803, 
    6.586007, 4.008044, 3.600106, 4.156508, 4.69917, 4.614934, 4.569488, 
    4.157092,
  28.01575, 30.21822, 30.84817, 16.01024, 13.31253, 12.51225, 10.8592, 
    9.520554, 5.801706, 5.421232, 5.152856, 5.044979, 5.223949, 4.642862, 
    4.350308,
  10.54393, 13.52696, 15.72836, 13.51063, 13.98276, 14.80164, 12.34835, 
    11.75001, 10.47546, 5.174981, 6.349761, 7.258062, 4.472754, 4.705554, 
    3.795896,
  2.841259, 7.988783, 12.61235, 11.91574, 11.43779, 11.23471, 3.954237, 
    3.355638, 3.496151, 6.277546, 5.296018, 7.638427, 9.433766, 8.090599, 
    6.492411,
  -0.5011747, 4.787261, 7.07553, 13.34137, 14.58493, 11.48901, 5.382614, 
    2.185736, 2.93866, 3.967714, 7.305147, 9.568355, 8.786737, 6.231173, 
    5.591025,
  1.001657, 4.31248, 14.44714, 13.79311, 16.56147, 15.02635, 10.31158, 
    5.327566, 5.566949, 5.718362, 6.022138, 8.426184, 11.97222, 5.643385, 
    5.481119,
  14.25533, 17.56484, 28.98732, 18.2644, 15.42615, 14.90514, 11.49095, 
    6.39663, 7.996686, 9.378657, 6.857357, 7.421883, 7.754342, 11.8116, 
    12.07361,
  28.28499, 20.11082, 32.27657, 16.94417, 17.78864, 14.6152, 11.56737, 
    8.980584, 11.17022, 13.62265, 10.90449, 7.712538, 6.344635, 7.432448, 
    10.42294,
  44.15793, 30.13121, 30.89543, 26.356, 38.55605, 13.18669, 11.89317, 
    10.36036, 8.170752, 9.547725, 7.279684, 6.589468, 6.535543, 7.441706, 
    6.811846,
  51.08417, 47.21262, 42.67922, 49.30761, 43.31556, 15.62627, 11.1335, 
    8.743901, 8.399725, 7.662001, 7.593393, 9.251077, 7.019889, 6.717224, 
    5.740667,
  59.90534, 59.65398, 54.9374, 51.68674, 35.17572, 14.02525, 9.565447, 
    8.586807, 7.819817, 7.586133, 8.178695, 9.454895, 9.716278, 7.132096, 
    7.328769,
  63.36945, 62.48767, 56.38887, 27.99783, 13.44679, 14.58315, 10.22829, 
    7.818739, 5.936183, 9.027888, 7.385133, 6.929204, 8.446905, 8.763441, 
    7.906971,
  46.8642, 32.94846, 29.3222, 19.26842, 14.41926, 11.5478, 7.701475, 
    14.13682, 13.04054, 5.166982, 3.431246, 4.492945, 5.804305, 7.169309, 
    8.65891,
  7.561979, 10.5785, 13.28607, 11.64753, 10.46158, 11.52289, 9.134056, 
    9.952115, 12.59728, 11.25796, 8.60621, 9.65609, 6.906155, 6.555454, 
    9.266559,
  31.70922, 21.2114, 12.70707, 10.33565, 10.85297, 7.402137, 7.850227, 
    10.77799, 13.5136, 13.84005, 10.01937, 12.13943, 9.417019, 5.420595, 
    9.180529,
  58.03568, 63.27522, 59.16276, 17.20509, 9.74855, 7.767203, 9.950963, 
    7.718219, 9.766683, 10.85283, 10.86824, 12.03679, 10.71041, 12.27326, 
    9.200017,
  70.13158, 76.88829, 79.14274, 20.68784, 7.598713, 6.37426, 3.715374, 
    8.096236, 11.76392, 12.3782, 10.11965, 11.81794, 13.01873, 11.67558, 
    10.76891,
  78.27828, 73.89172, 75.84969, 19.36727, 11.62658, 5.957719, 4.26986, 
    0.6353078, 6.614648, 15.44417, 13.1053, 8.859039, 9.612075, 11.34647, 
    12.31619,
  91.64589, 79.86754, 70.33263, 35.29053, 36.37516, 5.975729, 3.241467, 
    2.433869, 1.491402, 0.9844564, 2.1818, 4.131538, 6.811574, 10.20574, 
    11.19817,
  102.5043, 95.06926, 80.0368, 61.58727, 38.79556, 8.160635, 3.733692, 
    2.576974, 2.051522, 1.160601, 1.800364, 3.122813, 5.982359, 6.933913, 
    11.39157,
  114.1472, 106.0601, 90.61613, 58.39238, 34.54935, 10.16875, 5.524529, 
    4.379939, 3.899431, 2.427327, 2.323598, 2.971032, 4.24797, 5.293612, 
    9.727464,
  118.0147, 108.3176, 83.57051, 24.74678, 13.55949, 13.12133, 7.615272, 
    7.49595, 7.194677, 7.253037, 3.059306, 2.738317, 3.197109, 4.341107, 
    9.875411,
  88.63766, 59.51375, 43.83028, 15.87599, 10.78613, 13.62701, 10.02984, 
    18.07822, 16.19599, 4.789424, 1.72684, 1.453826, 1.82144, 2.932528, 
    6.300864,
  5.499453, 8.726829, 11.54674, 6.127238, 3.928906, 4.506772, 5.66159, 
    1.990898, 2.296442, 4.441831, 3.684679, 3.467187, 8.881363, 9.685594, 
    7.818371,
  33.29337, 21.55747, 13.07979, 4.755254, 3.246158, 5.414366, 4.099549, 
    2.256679, 2.337595, 3.713462, 2.648931, 3.046508, 4.39339, 5.006205, 
    4.254564,
  73.52367, 69.5163, 52.02278, 8.174847, 4.396859, 5.46748, 6.473722, 
    3.562288, 3.978452, 2.499206, 2.927315, 3.366009, 4.760866, 7.460059, 
    7.616699,
  99.685, 93.60006, 78.23587, 15.73284, 4.317244, 4.150824, 4.9333, 6.062065, 
    5.400423, 4.005831, 3.150311, 3.066239, 4.414666, 5.036112, 7.827782,
  115.029, 96.04568, 80.35657, 11.24857, 5.606457, 4.875593, 3.792017, 
    2.112912, 3.996059, 6.946276, 5.684484, 2.411227, 2.601687, 3.46628, 
    5.5599,
  134.9387, 110.9101, 81.49118, 30.22821, 20.05102, 3.630234, 2.809151, 
    2.608998, 0.4755908, 0.05084966, 0.5149128, 1.406747, 1.875683, 2.69133, 
    4.520948,
  150.5311, 136.2547, 104.032, 59.00658, 27.34947, 3.947368, 2.35365, 
    3.066171, 2.422667, 0.7885829, 1.147089, 1.609577, 2.526404, 2.292016, 
    4.158794,
  163.8034, 155.2028, 126.0463, 64.17219, 28.94842, 7.735057, 5.647287, 
    4.924236, 4.472781, 2.783131, 0.9578558, 1.727751, 2.483281, 1.986893, 
    5.185342,
  164.5967, 158.1429, 111.8428, 34.26023, 15.99206, 9.695072, 7.936027, 
    7.678981, 5.782933, 3.809203, 0.7145897, 1.470772, 1.424672, 2.141333, 
    5.50455,
  119.8574, 81.21732, 62.75498, 29.99428, 15.64822, 11.81383, 8.434342, 
    10.96685, 8.972972, 3.335684, 0.4152024, 1.459174, 0.8876746, 1.762581, 
    4.070777,
  8.60025, 9.002213, 13.26919, 7.844097, 4.755306, 7.166138, 5.566926, 
    6.057733, 6.661591, 6.452715, 3.238002, 1.720872, 4.053388, 4.844605, 
    5.891252,
  67.86707, 38.19833, 16.56716, 9.71252, 6.589056, 6.004233, 4.706165, 
    5.328254, 7.033742, 8.069564, 2.326668, 1.741121, 4.040216, 3.863026, 
    3.176942,
  117.2004, 109.6122, 88.79044, 15.40432, 6.766704, 4.388942, 7.168262, 
    7.70879, 6.758944, 3.870188, 2.985892, 2.676258, 4.945501, 4.484684, 
    1.873682,
  142.3132, 133.6788, 114.1426, 22.56004, 10.41792, 8.70954, 7.255595, 
    8.33451, 5.597026, 4.702219, 3.294883, 2.684442, 4.450986, 3.708818, 
    1.872725,
  155.6479, 134.3035, 112.0644, 17.49621, 9.571495, 7.979961, 14.27761, 
    4.984465, 1.866744, 5.489538, 5.14563, 2.257222, 3.052085, 2.665544, 
    2.399437,
  172.1685, 147.0112, 114.355, 42.49898, 20.09212, 4.370454, 8.686808, 
    16.76372, 7.561567, 4.420062, 3.286273, 2.313531, 1.665398, 2.446575, 
    3.266085,
  181.7325, 171.2238, 138.2692, 69.76372, 26.83731, 4.804699, 5.898106, 
    8.533187, 5.9883, 4.65952, 6.295118, 4.062171, 1.996971, 2.205065, 
    3.264904,
  185.7123, 184.4846, 153.0569, 73.63882, 29.76643, 9.905721, 8.914259, 
    6.536284, 3.115416, 5.380068, 4.569646, 4.113071, 2.161377, 1.420222, 
    3.414776,
  168.1904, 170.7769, 108.3673, 40.01251, 21.79222, 11.69569, 8.725744, 
    4.077286, 1.606377, 2.88329, 2.466753, 2.807827, 1.429603, 1.310026, 
    3.721398,
  95.47284, 72.94338, 51.47762, 29.4625, 15.85362, 11.35995, 7.02543, 
    8.756062, 4.134668, 2.445299, 2.084527, 2.182917, 0.914324, 1.33028, 
    3.925075,
  7.328326, 6.121211, 6.258678, 4.14569, 8.44083, 7.36287, 6.388352, 
    4.957801, 5.8873, 10.02741, 10.7013, 11.65089, 6.978548, 5.871327, 
    2.195255,
  64.51016, 35.17912, 11.72988, 6.508191, 11.84584, 8.846544, 5.81873, 
    5.918783, 6.920636, 10.40532, 9.508422, 8.168675, 8.36772, 2.48082, 
    3.718155,
  92.19244, 85.49278, 74.31934, 13.71828, 13.1618, 8.381676, 5.594738, 
    5.640454, 6.5861, 7.1848, 5.800246, 6.677136, 5.944429, 4.83776, 4.323193,
  99.15993, 95.38464, 98.67122, 26.07488, 16.42313, 19.56247, 7.670455, 
    5.49078, 5.886168, 5.574191, 2.383614, 2.71489, 4.90526, 4.436031, 
    5.691648,
  96.84238, 84.1896, 87.08839, 19.29139, 17.05101, 18.92898, 22.55672, 
    4.145845, 1.698282, 6.00892, 3.743587, 0.2683751, 2.016763, 5.477644, 
    5.67562,
  104.3193, 83.16039, 77.58901, 40.57868, 28.05355, 13.09999, 12.46807, 
    14.36148, 5.294984, 3.660906, 1.280656, 1.364026, 3.379137, 6.695633, 
    5.605469,
  114.1502, 101.2488, 85.30779, 50.98479, 28.01057, 9.940554, 6.856648, 
    5.597165, 4.950172, 2.779768, 1.812234, 1.918743, 5.220222, 7.787095, 
    6.66967,
  117.3997, 112.5516, 86.30108, 47.51235, 26.19162, 10.90839, 5.942521, 
    4.129916, 2.712693, 1.784938, 1.690211, 1.968385, 3.622254, 5.19559, 
    9.082059,
  111.0101, 109.837, 59.70457, 26.80517, 15.31613, 11.09599, 5.852375, 
    3.46231, 2.644133, 3.167474, 1.901918, 2.408542, 2.48878, 3.193586, 
    6.821055,
  66.73417, 49.95588, 31.04224, 19.43809, 11.3269, 10.06573, 6.898151, 
    9.338926, 5.978864, 2.332226, 1.531443, 2.036895, 2.016988, 5.651986, 
    6.952555,
  3.849754, 3.053372, 3.368417, 4.43496, 12.77251, 9.358564, 9.222911, 
    7.890825, 7.486408, 9.266343, 9.691402, 8.267819, 8.458175, 18.87391, 
    18.59392,
  20.76486, 13.82237, 7.019867, 8.434639, 12.82601, 8.635664, 12.22927, 
    9.466063, 11.65254, 15.71316, 10.07443, 10.92097, 19.16342, 11.36895, 
    8.91898,
  42.65711, 50.04939, 52.33981, 13.53567, 9.586612, 4.667419, 12.68806, 
    10.74374, 9.145519, 10.9456, 10.65289, 10.94341, 11.10764, 13.95003, 
    10.32329,
  61.00829, 67.3985, 77.85639, 20.30095, 14.20687, 14.12382, 9.452978, 
    14.46397, 10.40348, 8.085188, 6.527815, 6.964655, 8.749253, 8.321346, 
    6.213634,
  76.78813, 68.89873, 70.39104, 15.27809, 15.06819, 16.9043, 16.25434, 
    5.120355, 3.247671, 8.482716, 6.101467, 2.536915, 3.287513, 5.05205, 
    4.917218,
  97.41567, 79.33905, 72.19421, 33.57134, 24.05188, 11.90638, 11.05343, 
    11.82318, 4.403016, 5.136017, 3.808249, 3.614318, 3.306119, 1.941941, 
    2.607238,
  107.6972, 100.8022, 87.21191, 48.68129, 24.21466, 11.52771, 6.003272, 
    5.977537, 5.228048, 3.320371, 3.331703, 3.901328, 4.801236, 1.231315, 
    4.099072,
  107.0322, 108.9426, 87.50924, 47.18524, 23.46497, 11.29878, 2.702665, 
    5.169593, 4.905815, 3.886457, 4.371002, 3.66636, 3.914898, 6.221284, 
    8.866199,
  98.62885, 100.9306, 54.26655, 26.34493, 14.96682, 7.465344, 4.245193, 
    1.408821, 5.934634, 6.291594, 5.967872, 6.099745, 6.711753, 6.920098, 
    10.19396,
  57.42607, 43.86367, 25.98228, 16.53937, 15.30319, 16.23314, 11.49034, 
    14.93497, 3.802915, 2.946954, 4.160329, 6.494595, 5.915293, 7.522305, 
    7.94818,
  3.566761, 3.87427, 6.728243, 5.884182, 11.05245, 6.228174, 4.078508, 
    4.754014, 10.99527, 14.93788, 15.14072, 9.84854, 9.935251, 8.126615, 
    5.342975,
  28.03857, 11.65374, 7.796602, 10.0162, 13.47486, 5.52739, 4.115419, 
    4.810824, 8.38905, 17.09109, 13.58242, 10.86041, 15.56294, 9.154056, 
    6.338931,
  58.5332, 55.39669, 42.85614, 13.6325, 7.230445, 3.736089, 5.74914, 
    4.312372, 5.545632, 7.618773, 11.12658, 12.63801, 11.15867, 16.77543, 
    12.71747,
  66.18395, 67.20757, 63.98086, 16.53939, 8.699865, 10.124, 4.891482, 
    4.73035, 5.824681, 5.090775, 10.11007, 14.25765, 10.18703, 16.50342, 
    13.99039,
  67.53646, 62.51812, 60.76432, 12.10354, 14.55731, 16.21155, 15.30424, 
    7.061203, 6.036041, 8.266672, 11.65677, 10.26785, 11.80804, 10.85785, 
    13.93024,
  69.55882, 63.89245, 57.57579, 31.86823, 25.61656, 17.44722, 15.2696, 
    16.04265, 9.419142, 7.125101, 7.474017, 8.31655, 9.063935, 8.446479, 
    12.84437,
  70.65202, 72.66086, 62.84706, 37.26368, 21.43703, 16.65172, 14.8164, 
    16.35596, 9.769937, 7.572482, 6.423601, 8.021536, 8.709203, 10.51668, 
    11.52664,
  74.16582, 74.19184, 52.44307, 26.60149, 17.67955, 13.44885, 12.60528, 
    17.53622, 11.57605, 9.172241, 6.974484, 7.661826, 8.279538, 10.03051, 
    10.73678,
  68.01365, 56.15356, 25.49244, 12.46337, 9.510063, 9.442392, 11.46624, 
    15.99475, 13.86963, 8.913006, 6.230647, 7.286419, 8.215082, 8.639404, 
    9.499717,
  32.20455, 15.61025, 8.682547, 5.573016, 4.497946, 9.186203, 11.05717, 
    23.65603, 15.7443, 7.12312, 5.087882, 5.407416, 7.064843, 8.747198, 
    8.840172,
  9.970611, 15.97986, 17.51085, 4.385594, 0.9970059, 4.325548, 3.107603, 
    2.032347, 5.267882, 9.965943, 13.97323, 8.908046, 9.19235, 6.557547, 
    7.066316,
  29.11652, 13.36007, 4.3255, 1.665688, 6.041646, 5.357241, 3.498793, 
    4.282879, 6.795442, 10.35239, 13.49434, 8.33042, 9.176368, 4.135893, 
    4.697537,
  37.30932, 23.22827, 12.4392, 1.585815, 2.135628, 4.641763, 5.221207, 
    7.08053, 8.442834, 9.808507, 11.78244, 10.43777, 4.370228, 8.813113, 
    6.874298,
  29.56773, 24.87879, 23.40627, 5.986911, 6.689305, 4.49867, 4.198097, 
    5.364468, 9.201216, 11.71253, 13.96566, 11.31124, 7.269896, 8.264771, 
    5.405505,
  22.67543, 15.00978, 22.58265, 7.902592, 7.89247, 2.474913, 5.510178, 
    2.717117, 6.745743, 10.27929, 14.13393, 12.68571, 9.546244, 5.622525, 
    6.044777,
  30.09735, 18.16458, 17.38119, 11.59653, 9.681346, 3.625762, 2.920346, 
    5.105989, 4.690075, 7.534822, 8.52477, 10.72006, 9.39475, 6.524132, 
    9.207852,
  35.67212, 27.95454, 20.84762, 11.45211, 8.737482, 6.922668, 2.856996, 
    5.575809, 7.813278, 9.525449, 11.11857, 10.30254, 9.661806, 10.24084, 
    9.97448,
  34.08242, 27.4998, 17.38562, 12.96506, 11.44707, 4.363573, 4.713223, 
    8.24171, 9.95227, 8.083672, 10.6563, 9.57123, 10.01743, 10.12555, 10.50456,
  26.2407, 21.23063, 10.38297, 10.04777, 6.707352, 3.454801, 7.498309, 
    8.925797, 13.01645, 10.27294, 10.10005, 9.627208, 9.024674, 7.508452, 
    8.535956,
  7.12417, 7.123618, 8.301513, 4.376601, 3.423824, 3.579875, 8.930795, 
    19.89916, 15.14746, 7.845837, 7.957963, 8.344316, 11.17095, 6.485116, 
    9.805947,
  4.890178, 8.36952, 12.25101, 4.404466, 4.805227, 6.757946, 3.615366, 
    4.885802, 4.071138, 4.657548, 4.659622, 8.102696, 6.025641, 3.018242, 
    4.286691,
  6.10418, 5.779694, 4.876995, 5.828803, 10.09137, 10.53902, 6.186901, 
    5.312587, 5.227722, 1.810453, 6.090585, 9.928888, 7.540864, 4.354355, 
    1.728018,
  8.058874, 12.18339, 16.50448, 7.853742, 10.86388, 12.63111, 7.486751, 
    7.017419, 1.773554, 1.341855, 7.576833, 10.17557, 9.298622, 12.2966, 
    6.234345,
  11.47497, 22.45592, 30.65296, 11.52489, 7.917209, 8.839954, 7.727059, 
    6.405945, 3.160053, 2.72777, 3.93838, 10.39328, 15.20809, 12.90866, 
    5.018439,
  16.35203, 20.68826, 31.11222, 10.96729, 8.962104, 6.490561, 7.811536, 
    2.143283, 1.190117, 4.329862, 13.3513, 11.6089, 16.27911, 9.995098, 
    8.596031,
  19.4981, 24.52841, 27.02635, 14.26941, 12.28788, 8.073498, 10.1888, 9.255, 
    6.516285, 3.382238, 11.08532, 5.065669, 12.74009, 9.552246, 5.617711,
  17.44376, 24.77666, 21.69642, 14.75412, 11.12673, 8.804317, 10.05119, 
    12.51957, 8.832857, 10.50788, 12.29448, 4.123833, 12.41881, 8.346192, 
    6.887335,
  13.66321, 22.36371, 15.51296, 10.27464, 9.232313, 5.676457, 11.11839, 
    13.55585, 11.28449, 11.85298, 11.72149, 4.245555, 8.233635, 7.572932, 
    7.787826,
  14.42036, 15.9506, 6.721179, 6.200553, 6.503844, 5.70474, 11.16311, 
    15.98806, 11.84591, 13.14684, 10.79438, 4.944166, 9.273602, 9.808477, 
    10.86709,
  3.276735, 1.300131, 4.04726, 4.088091, 6.14043, 5.985323, 11.47903, 
    26.80778, 17.93631, 9.876597, 8.484647, 9.605101, 13.4257, 14.77127, 
    5.850417,
  3.263049, 4.62766, 8.557801, 5.322009, 4.136843, 6.231505, 6.069133, 
    10.79311, 10.12722, 10.99804, 9.190219, 11.06909, 11.58208, 9.46937, 
    9.9856,
  10.7122, 6.94889, 6.631312, 4.659211, 4.93432, 5.118151, 4.079061, 
    3.729159, 8.09825, 9.252338, 9.260014, 11.63809, 10.74586, 8.566541, 
    10.70943,
  13.89577, 18.67985, 14.79441, 3.616826, 3.971192, 6.275032, 4.463066, 
    5.598712, 6.700251, 3.622124, 3.580835, 11.57271, 13.76377, 15.4212, 
    14.49975,
  11.65898, 15.28403, 17.03556, 4.571686, 6.506822, 8.073175, 6.038073, 
    4.706618, 7.430376, 7.902549, 8.769999, 11.77095, 14.37641, 16.36399, 
    13.08145,
  7.422705, 6.425015, 17.53628, 2.67354, 7.512209, 7.086072, 8.964714, 
    4.770696, 8.204809, 13.09609, 16.12298, 12.07735, 15.61726, 13.99909, 
    17.24846,
  4.267732, 4.141009, 13.62621, 6.382339, 8.841192, 5.329917, 7.329643, 
    9.655697, 7.466586, 8.459816, 10.4587, 9.630569, 15.48537, 15.95939, 
    17.73623,
  4.495773, 12.96701, 22.84259, 7.106149, 8.272775, 4.578414, 6.147465, 
    9.207762, 7.960179, 10.39544, 10.69793, 10.3051, 15.37848, 16.88128, 
    17.05769,
  7.116405, 19.92949, 28.24549, 9.618274, 8.002812, 5.688048, 6.476102, 
    9.385939, 8.694263, 13.11047, 11.88796, 16.73848, 18.7516, 17.94102, 
    13.8805,
  9.697922, 19.73104, 16.93647, 10.94364, 7.46316, 3.962421, 6.586277, 
    11.74572, 12.28942, 13.4284, 15.47745, 19.90262, 18.50677, 19.85263, 
    21.14141,
  1.341851, 6.854074, 10.13166, 11.05689, 6.71936, 5.485516, 6.659157, 
    20.04692, 17.23549, 12.56781, 12.94208, 16.06218, 20.23822, 19.05944, 
    24.94065,
  2.428061, 4.767389, 10.6884, 7.906828, 6.333433, 9.117081, 3.95745, 
    5.036367, 8.614313, 13.40126, 12.27934, 10.37899, 12.2328, 9.225894, 
    9.569738,
  3.034466, 5.313538, 10.20881, 9.030788, 15.48862, 10.68589, 5.767509, 
    1.793309, 1.38562, 3.815394, 8.264238, 11.54216, 11.43268, 11.39549, 
    10.41501,
  7.19802, 11.41099, 18.34055, 11.09625, 11.83496, 11.17417, 3.551114, 
    7.140288, 3.010844, 8.282678, 10.48815, 12.37123, 11.08025, 10.22067, 
    9.801101,
  7.515399, 16.82648, 27.56869, 13.50066, 9.374884, 8.506158, 5.108508, 
    6.464664, 9.559613, 11.43905, 12.64779, 12.54269, 11.74279, 12.11889, 
    15.72336,
  10.70897, 17.14866, 24.86811, 11.44863, 7.294089, 8.236723, 8.61191, 
    6.096262, 7.111052, 18.036, 19.72378, 9.27916, 9.596687, 8.932878, 
    11.07216,
  10.72721, 22.80102, 21.84391, 14.35432, 11.15508, 6.775081, 3.147584, 
    6.424003, 0.3839175, 3.3041, 7.908071, 12.64959, 13.06633, 8.092402, 
    9.405892,
  12.40565, 31.64401, 27.88708, 15.43688, 9.030682, 6.668097, 1.675905, 
    3.049578, 1.546535, 3.5642, 7.118373, 13.35764, 15.94882, 12.60602, 
    8.478079,
  16.99381, 39.33361, 29.44738, 15.49414, 6.824984, 5.639039, 0.9580542, 
    1.648452, 3.185537, 5.076983, 8.267848, 16.27735, 19.99493, 20.6433, 
    15.90463,
  16.31865, 38.12187, 18.61556, 7.728917, 8.345243, 2.666736, 0.6795259, 
    3.690876, 6.122715, 11.1991, 11.568, 12.88359, 20.67296, 21.19988, 
    29.27293,
  1.389845, 14.78848, 16.08811, 6.963767, 7.603142, 7.506783, 1.032212, 
    18.33889, 16.7644, 7.825875, 4.03207, 8.795056, 18.89489, 19.47961, 
    30.18831,
  3.102998, 4.357877, 12.7644, 2.107681, 1.859948, 3.242443, 1.459903, 
    1.226448, 1.420359, 6.588012, 5.943287, 1.519664, 10.12604, 12.94362, 
    11.00387,
  11.74495, 6.067078, 5.093845, 1.203454, 4.058632, 3.415967, 0.8944877, 
    1.19951, 1.259244, 1.497597, 0.5027329, 4.343766, 2.018905, 8.339373, 
    8.11013,
  20.09376, 22.0161, 18.33811, 3.022542, 2.493734, 3.009749, 1.724377, 
    1.316962, 0.9138656, 1.778133, 1.077303, 4.196865, 9.828581, 10.6759, 
    8.706294,
  16.73915, 21.23059, 22.33049, 9.91891, 2.853702, 1.993553, 1.981688, 
    3.271491, 3.797257, 4.654199, 3.55047, 8.383936, 11.04272, 13.99707, 
    10.62233,
  16.61185, 11.06449, 16.27404, 10.19516, 5.269343, 4.818093, 6.619477, 
    2.653608, 2.061328, 12.56912, 9.858357, 8.17476, 11.47461, 12.21679, 
    10.58492,
  13.4547, 8.536606, 8.668521, 10.30678, 11.96041, 9.126333, 7.777462, 
    4.99474, 2.3651, 3.441282, 5.186492, 8.457027, 15.39989, 12.07217, 
    11.39566,
  6.234204, 5.246871, 8.085712, 6.463365, 7.473558, 7.029294, 6.547052, 
    7.601271, 8.096537, 5.699979, 6.822537, 8.309536, 11.10545, 16.3121, 
    17.76647,
  5.763628, 6.172034, 6.663489, 5.686531, 7.903007, 7.871511, 8.995727, 
    8.099094, 6.505847, 6.726331, 7.77212, 6.68263, 9.05361, 21.17251, 
    26.46635,
  7.533319, 5.893977, 0.05037434, 1.250563, 3.722174, 5.708616, 7.461498, 
    7.255921, 6.767971, 9.023995, 7.535404, 8.391029, 11.13181, 18.99672, 
    37.7818,
  3.675863, -0.2037102, -1.195224, 1.214914, 2.370047, 5.148553, 5.35533, 
    10.53659, 12.72378, 8.372473, 4.431711, 6.134954, 5.296117, 15.70193, 
    29.29008,
  3.698663, 6.993743, 11.22246, 5.059876, 6.039533, 5.256106, 3.707842, 
    2.519738, 2.197643, 2.641068, 3.920362, 1.488369, 3.674355, 7.518199, 
    6.079666,
  4.928657, 4.673802, 4.462546, 4.170086, 5.288352, 6.272125, 1.57329, 
    5.051361, 3.770569, 0.5615773, 3.224133, 1.653801, 1.12792, 6.381642, 
    5.657463,
  4.168359, 3.374981, 6.108449, 5.047543, 6.721209, 9.914344, 8.024018, 
    6.000731, 4.738085, 2.966486, 2.792916, 2.185208, 3.241462, 7.88799, 
    7.455299,
  2.015721, 1.51993, 3.812742, 4.260083, 6.889945, 7.066133, 5.277748, 
    7.029979, 3.378168, 3.554039, 2.20457, 1.923734, 5.151281, 7.698529, 
    8.494789,
  1.814235, -0.2683868, 2.052361, 2.605045, 4.040477, 4.655022, 4.05384, 
    4.51477, 3.61763, 6.908442, 7.712345, 7.275168, 7.059041, 5.996127, 
    6.396163,
  3.236475, 0.7731532, -0.7810687, 1.438325, 3.636889, 4.261291, 3.504158, 
    3.166973, 5.435647, 7.116991, 6.517343, 6.249733, 7.280231, 5.491056, 
    5.008281,
  4.970069, 3.156476, 0.7418267, 1.336848, 4.044131, 5.131059, 3.386864, 
    3.655378, 4.486467, 4.921389, 4.197061, 3.642584, 4.948885, 5.263684, 
    7.513462,
  3.742634, 3.345432, 2.2659, 1.076696, 4.447221, 4.326276, 4.693994, 
    7.26801, 5.567674, 5.480121, 3.610262, 5.463867, 7.001881, 10.88335, 
    13.49804,
  2.666843, 3.705126, -0.7410621, 2.211224, 4.008677, 4.509508, 7.502392, 
    8.910254, 8.633676, 11.76557, 7.418527, 12.5914, 13.40681, 15.31748, 
    20.49517,
  -0.7159987, -0.900821, 0.1479765, 4.663583, 6.833539, 8.665475, 6.637954, 
    13.67203, 23.58749, 18.34795, 13.72489, 12.54233, 10.7812, 12.32434, 
    15.58037,
  0.1656243, 2.319293, 4.6616, 1.436163, 4.413756, 5.193686, 3.875297, 
    3.08334, 3.790123, 6.220513, 11.80471, 7.808686, 4.174501, 4.850694, 
    5.425972,
  -0.4810048, 0.2339258, -0.02573851, 2.509351, 6.494301, 6.170464, 3.517258, 
    5.724344, 7.29845, 8.398755, 10.49284, 7.870717, 5.806197, 3.527175, 
    3.013306,
  0.09525087, 0.3990347, 1.858006, 2.22869, 6.503281, 8.070031, 7.072868, 
    4.689245, 3.853079, 8.676162, 8.168503, 7.399605, 6.051108, 4.345552, 
    2.510798,
  3.396074, 7.430838, 13.4986, 6.545696, 5.845045, 5.822472, 11.16948, 
    3.665502, 3.3828, 7.581913, 5.995976, 5.7439, 4.811232, 5.000166, 3.107364,
  10.17889, 12.47121, 23.20735, 10.1699, 7.651584, 8.696817, 8.330287, 
    11.31826, 10.79297, 7.29486, 6.683514, 6.315381, 7.486825, 8.274854, 
    8.976293,
  16.10909, 22.72724, 25.21763, 18.95819, 10.98941, 8.652195, 9.420591, 
    10.30316, 9.119826, 7.338478, 6.434547, 4.645281, 4.534564, 4.585266, 
    9.946978,
  20.19512, 32.14788, 35.74609, 28.61042, 12.35305, 8.066519, 7.349457, 
    9.284249, 8.533371, 5.791759, 3.048462, 2.371394, 4.780166, 5.814444, 
    7.43925,
  27.16446, 40.23287, 42.4046, 25.55957, 14.24874, 7.569474, 3.72982, 
    4.817757, 9.813375, 11.83221, 10.62672, 11.34424, 13.22398, 18.93765, 
    21.57236,
  32.93812, 44.02299, 30.73703, 14.96282, 11.03172, 5.874668, 5.194036, 
    11.69511, 16.318, 24.25999, 13.91115, 11.207, 14.61318, 18.87906, 23.68738,
  27.59323, 26.8289, 20.92009, 9.799467, 6.554521, 4.963527, 9.056844, 
    19.48471, 34.27755, 23.0826, 13.31792, 10.44015, 11.54986, 16.24663, 
    20.19979,
  8.268119, 11.67398, 18.74247, 12.7673, 12.9837, 17.57036, 10.88553, 
    12.05954, 13.36845, 18.68342, 15.56008, 10.2344, 8.75268, 9.570903, 
    7.913126,
  26.15542, 24.93779, 12.69706, 12.46959, 20.62157, 15.4435, 9.594753, 
    10.6057, 11.12382, 14.0141, 13.59103, 13.55854, 9.372939, 8.184203, 
    11.64852,
  37.36398, 43.51627, 42.88236, 12.18546, 11.57405, 10.77279, 9.059589, 
    6.976532, 10.91507, 7.467656, 6.236696, 11.50407, 11.88964, 9.252571, 
    9.870075,
  39.7684, 46.66708, 53.53392, 21.16324, 12.2002, 6.876094, 6.595149, 6.5914, 
    8.886246, 12.30085, 5.577707, 5.414877, 5.393193, 11.92928, 11.99424,
  39.80787, 38.48735, 45.46465, 20.0787, 12.90341, 13.6537, 8.95077, 
    4.666912, 9.642086, 14.0267, 8.75152, 5.201325, 2.424131, 2.616125, 
    4.107554,
  38.45251, 35.44275, 31.99342, 24.01562, 17.19767, 6.201495, 11.3804, 
    13.1754, 12.40476, 8.992059, 3.43156, 4.952149, 6.949904, 1.707857, 
    1.664704,
  34.54494, 33.33323, 29.78918, 23.67758, 14.4497, 3.394742, 8.771663, 
    12.66904, 9.694573, 10.88727, 6.231199, 5.818328, 11.128, 7.076066, 
    2.797444,
  30.90437, 29.24553, 25.74581, 16.72448, 15.54472, 3.523092, 8.052455, 
    12.39412, 9.710041, 9.292461, 8.251925, 9.968689, 10.55197, 11.12713, 
    11.81029,
  25.08175, 21.168, 12.85898, 4.783157, 13.03908, 3.411011, 8.908837, 
    15.63343, 17.34891, 25.21638, 13.48447, 14.0674, 7.947894, 8.845376, 
    10.8716,
  10.07691, 5.60551, 8.211735, 5.117954, 9.635515, 5.058187, 6.865208, 
    18.52609, 29.62942, 19.77876, 14.60102, 12.70707, 4.821976, 6.654059, 
    7.499269,
  7.543873, 10.51484, 14.20067, 7.171754, 6.699269, 8.377863, 4.206725, 
    2.394727, 2.795386, 6.337041, 9.179949, 4.039693, 3.841182, 11.18928, 
    10.74164,
  11.73453, 12.52928, 10.37848, 8.139856, 7.306808, 5.350225, 3.813114, 
    4.150894, 4.011644, 3.325429, 3.954359, 0.7292451, 1.090856, 7.928382, 
    11.31894,
  14.78505, 17.74044, 14.30644, 6.697569, 3.440502, 5.833285, 4.681493, 
    5.217937, 6.499227, 4.936364, 4.616441, 3.304236, 2.452352, 3.897513, 
    6.944229,
  13.709, 15.87573, 13.12525, 3.603558, 2.919828, 3.348198, 3.718325, 
    5.692192, 7.882963, 6.16053, 6.965611, 3.71078, 3.016286, 5.401289, 
    2.860288,
  14.66679, 6.053901, 5.749027, -0.05362627, 1.248169, 4.315604, 6.11221, 
    5.330626, 6.118578, 11.84135, 6.776822, 3.11616, 3.564464, 6.132977, 
    3.392307,
  13.03205, 5.668536, -3.658348, -4.098618, 0.9486298, 2.407065, 4.780694, 
    6.226083, 8.185602, 9.498763, 8.484384, 2.307686, 2.589551, 2.807807, 
    5.887866,
  9.460395, 2.07667, -4.722362, -5.377267, -0.4242864, 1.420611, 4.49164, 
    4.560507, 7.180746, 5.702461, 7.745849, 3.331405, 2.250814, 5.359306, 
    6.682524,
  8.01103, 4.0963, -3.91676, -4.208228, -0.4284883, 2.553318, 2.252498, 
    4.625714, 7.778192, 7.171224, 8.339314, 3.29683, 2.012242, 7.983048, 
    9.616318,
  4.524299, 1.639648, -3.750426, -2.004682, 0.4665222, 2.483672, 3.958586, 
    7.521948, 10.57378, 12.42112, 2.698123, 2.674531, 2.093055, 4.164421, 
    13.8059,
  1.427397, -3.107951, -3.241139, 0.5419702, 4.125966, 3.75535, 6.157871, 
    13.05962, 17.3628, 7.08253, 3.706746, 3.277603, 2.664988, 2.965195, 
    12.00215,
  1.244221, 4.470081, 8.300922, 5.190804, 7.324387, 9.419172, 8.741382, 
    9.548864, 7.038557, 5.859206, 6.970069, 6.755681, 7.615614, 7.493334, 
    7.415357,
  -1.313506, -0.1845954, 1.592807, 4.184769, 5.12642, 6.040272, 6.514388, 
    8.883796, 5.558699, 4.43585, 4.098222, 6.121568, 6.930393, 8.837068, 
    7.264675,
  -1.803123, -0.9045669, 1.381377, 1.927863, 4.163505, 10.22108, 10.10711, 
    5.654576, 3.963351, 2.724377, 3.858508, 5.621318, 6.710712, 9.49201, 
    7.064321,
  -0.05637009, 4.524695, 8.331161, 4.668943, 6.262191, 7.389825, 11.22047, 
    6.893852, 8.558782, 11.76393, 7.156417, 7.449942, 7.672348, 9.447997, 
    6.828112,
  5.047029, 7.419824, 15.96922, 9.360303, 9.561107, 9.319517, 6.684943, 
    13.33366, 11.69252, 12.66022, 8.891078, 9.412317, 10.12041, 8.160169, 
    8.319633,
  10.86459, 17.83925, 18.65407, 18.27371, 16.60394, 14.45272, 13.31799, 
    11.30295, 10.76948, 13.07184, 8.713123, 8.759282, 7.298552, 5.90432, 
    4.475357,
  15.82459, 28.2417, 28.98735, 22.13422, 16.42811, 17.25995, 11.79275, 
    13.30018, 12.18856, 3.132445, 5.752433, 5.926584, 5.324461, 6.023223, 
    4.867625,
  22.68285, 37.18311, 33.57843, 19.27213, 15.53847, 14.67737, 15.12586, 
    15.19487, 9.304438, 3.199432, 1.985801, 2.436435, 4.060706, 5.906721, 
    8.795792,
  31.68187, 40.97467, 28.45724, 18.03641, 14.65133, 14.4525, 16.87537, 
    16.79188, 12.8919, 8.601127, 2.196365, 1.462218, 1.900501, 3.878307, 
    13.03079,
  33.15828, 30.58878, 28.26091, 17.14489, 12.48145, 10.31359, 10.59077, 
    16.92417, 17.40353, 5.857203, 1.601991, 1.371948, 2.267248, 4.277776, 
    10.2835,
  10.36752, 21.75031, 25.73421, 17.20876, 17.48476, 16.22233, 11.38585, 
    13.13427, 14.80223, 19.1037, 14.03898, 7.493299, 8.440176, 11.28384, 
    9.476693,
  30.07917, 32.63542, 22.80719, 23.10202, 18.97793, 15.52418, 9.128589, 
    11.60377, 15.10942, 20.87526, 18.15072, 8.791713, 5.885915, 7.293345, 
    5.905128,
  42.03172, 56.66647, 54.79564, 23.52861, 13.06026, 11.92237, 7.930973, 
    8.5783, 14.15322, 18.13033, 19.50916, 11.76527, 3.475718, 7.496347, 
    8.154464,
  48.37279, 62.29063, 72.91969, 29.35015, 11.40493, 9.118362, 5.748271, 
    8.050293, 11.45825, 16.9885, 16.28882, 10.15163, 5.952173, 7.129281, 
    9.657153,
  59.05313, 60.36237, 71.4994, 32.49512, 21.02246, 19.35811, 14.60057, 
    5.638838, 10.52401, 15.62673, 16.61417, 13.46664, 10.60736, 9.966841, 
    13.35141,
  63.83967, 67.36143, 63.88878, 45.61504, 26.36804, 17.22353, 18.31539, 
    16.27094, 12.06798, 6.424187, 6.273992, 9.291859, 11.27382, 10.8861, 
    9.443326,
  67.51764, 74.16679, 69.61843, 41.79775, 18.72739, 17.61614, 14.37636, 
    15.9981, 14.30499, 4.512282, 4.625561, 9.185205, 8.955407, 8.993142, 
    8.254757,
  76.13284, 80.37405, 65.20152, 28.17505, 16.42254, 16.44341, 14.66336, 
    13.38991, 14.28893, 4.634561, 2.759951, 4.873106, 8.139421, 8.476818, 
    13.41592,
  79.91587, 77.21473, 43.22423, 18.31657, 15.24963, 14.53213, 15.08874, 
    16.84451, 15.46071, 12.83811, 3.652556, 2.330044, 3.317807, 3.902057, 
    6.937844,
  69.69057, 51.12549, 31.45366, 17.96336, 14.73926, 12.05872, 14.28434, 
    21.96461, 20.41109, 5.576531, 1.311583, 0.6749693, 3.141037, 3.085479, 
    3.707304,
  7.788261, 12.54239, 16.29298, 12.37994, 13.37633, 8.263979, 4.486209, 
    0.5305662, 2.58313, 13.93897, 17.18447, 16.00582, 17.26668, 19.62749, 
    20.2491,
  36.01708, 25.0232, 13.11654, 15.124, 10.72167, 7.831036, 4.713512, 
    4.261922, 2.708591, 3.142119, 15.56493, 16.76794, 14.96099, 16.40793, 
    15.73848,
  56.91779, 54.91385, 42.45166, 14.26261, 8.575786, 8.147855, 7.611736, 
    8.081338, 6.868736, 7.911653, 15.29162, 17.59083, 15.07671, 11.18607, 
    14.81212,
  67.33114, 66.99439, 65.41519, 21.25418, 8.463194, 7.102389, 7.405868, 
    8.381824, 11.09642, 13.05888, 15.98343, 19.38771, 11.22813, 6.655738, 
    11.99982,
  78.08723, 64.76997, 71.46594, 29.46219, 14.41237, 8.252255, 7.524677, 
    4.0428, 6.997653, 14.96054, 13.72963, 17.13467, 12.55678, 7.158261, 
    8.70034,
  83.4107, 77.31784, 65.58454, 42.91259, 16.0757, 12.15718, 8.771298, 
    5.27845, 4.362533, 6.372791, 7.599556, 11.6662, 15.23296, 11.9879, 
    10.58494,
  83.98241, 84.18285, 73.89082, 38.57868, 15.36672, 14.57227, 8.363623, 
    7.878942, 4.032967, 3.841871, 6.733795, 9.450808, 12.76837, 15.61678, 
    14.27713,
  86.18893, 86.77129, 66.18061, 27.22847, 17.00579, 15.47513, 8.880021, 
    7.805938, 5.676408, 7.026134, 4.924709, 7.126463, 11.73489, 14.9915, 
    18.31984,
  77.02799, 78.5263, 39.79071, 19.74931, 13.04404, 11.04362, 12.43337, 
    15.65325, 12.01128, 11.07171, 12.68935, 10.76204, 9.801614, 14.97896, 
    19.22178,
  54.63742, 42.42622, 26.01818, 18.25164, 14.51734, 13.5083, 10.59087, 
    24.26449, 21.04493, 8.34916, 6.017454, 9.395905, 13.40465, 14.04948, 
    18.35579,
  5.497958, 10.63298, 13.82455, 16.51604, 12.90255, 11.80268, 2.36095, 
    2.277098, 2.138938, 10.44565, 10.33544, 7.026186, 14.18582, 16.45301, 
    5.868669,
  10.71849, 17.43632, 11.9308, 16.23636, 16.41888, 12.29827, 3.037429, 
    3.22322, 3.430655, 2.752931, 5.497829, 15.05231, 13.43055, 16.11197, 
    9.76103,
  22.41759, 37.58424, 35.7631, 13.12041, 10.33181, 11.72251, 4.499533, 
    6.61417, 7.742911, 3.926147, 2.705962, 15.22593, 14.85149, 13.13087, 
    14.87948,
  34.0408, 47.35454, 51.02075, 22.81458, 9.652601, 5.027293, 5.781477, 
    9.741521, 13.92972, 13.79483, 6.712567, 12.88325, 12.73281, 8.176485, 
    11.64019,
  47.12363, 48.00031, 52.5615, 25.76431, 14.79293, 10.45373, 3.724363, 
    3.962574, 6.650102, 16.91203, 14.44213, 11.83243, 13.28423, 10.92467, 
    11.56099,
  53.12973, 55.53384, 48.42036, 32.89751, 20.94374, 16.80771, 8.463005, 
    7.216911, 6.816639, 7.978067, 9.006588, 10.95632, 10.873, 8.043322, 
    8.784369,
  54.55634, 61.28771, 51.69132, 28.44593, 18.32267, 17.67397, 14.18941, 
    15.01316, 10.18778, 8.288295, 11.28289, 11.89467, 10.6828, 10.60747, 
    11.61609,
  57.32635, 64.93594, 45.03381, 18.859, 16.27518, 16.75013, 14.37232, 
    16.08939, 15.1443, 10.64509, 12.33777, 13.38376, 10.95795, 11.80349, 
    14.7345,
  56.4032, 62.90526, 30.1568, 14.65042, 13.00666, 15.48983, 16.30471, 
    23.55122, 20.99109, 20.38221, 16.42139, 14.34084, 12.96846, 8.285271, 
    14.86078,
  46.6337, 39.83, 17.94389, 15.77668, 14.15324, 15.26583, 18.20901, 34.83502, 
    32.35036, 19.39153, 13.72505, 14.23088, 14.92675, 10.97943, 7.511686,
  7.723525, 12.89664, 17.17033, 4.528055, 7.528371, 5.674405, 5.455461, 
    5.31775, 3.553384, 9.766903, 12.82416, 12.36608, 12.15658, 14.22201, 
    11.6998,
  30.84887, 33.69226, 12.21353, 4.679984, 8.104187, 5.859103, 7.765375, 
    7.345448, 4.841114, 0.09290411, 7.439428, 13.63951, 6.703254, 11.26171, 
    9.067771,
  70.85416, 76.17008, 43.22066, 10.80556, 8.686883, 5.884037, 9.981493, 
    12.62571, 12.71708, 6.017685, 0.611897, 11.28273, 7.125917, 11.50421, 
    10.85069,
  82.12918, 77.50759, 61.08959, 22.19265, 14.80148, 4.954791, 9.995506, 
    18.53751, 22.11407, 16.35036, 2.141635, 10.9724, 8.646955, 4.122733, 
    12.11562,
  85.11153, 66.66723, 57.60413, 25.27261, 16.59992, 15.47751, 10.95483, 
    8.555141, 14.91551, 20.46667, 9.455559, 9.620892, 7.833592, 4.523813, 
    9.525325,
  78.74191, 65.92197, 51.36137, 31.90904, 20.56328, 16.42865, 15.18082, 
    11.59523, 9.825571, 9.503582, 7.685043, 11.46527, 9.598631, 9.939899, 
    5.458674,
  70.1334, 65.2062, 52.82906, 26.65571, 18.6771, 17.30482, 15.67264, 
    12.43676, 10.83189, 10.2872, 8.466265, 12.35121, 9.816046, 12.13595, 
    3.590798,
  68.08203, 64.40808, 42.90957, 19.70082, 18.41584, 19.60584, 16.56686, 
    11.14411, 10.70178, 12.22532, 11.24105, 7.326735, 11.21783, 11.56732, 
    10.7167,
  62.66553, 60.48977, 25.83979, 13.57955, 16.9887, 13.03612, 13.33406, 
    20.06588, 18.18107, 20.41701, 12.56583, 8.852895, 4.777715, 6.885974, 
    14.54075,
  52.07021, 40.38333, 14.16873, 12.77323, 14.83105, 7.116243, 12.74642, 
    38.95681, 34.23039, 15.04469, 7.978414, 6.551807, 7.439723, 6.425334, 
    9.298005,
  11.35785, 17.93757, 16.75392, 3.589066, 3.279122, 4.821199, 3.538975, 
    3.398077, 5.227629, 13.14487, 15.37409, 13.1763, 10.78499, 13.91124, 
    17.28684,
  39.93188, 23.90604, 10.35822, 5.181627, 6.911847, 6.170638, 5.357174, 
    8.079648, 7.226909, -0.2031514, 13.47705, 12.0284, 10.31809, 12.31236, 
    16.7494,
  66.87605, 60.62223, 37.50784, 11.07022, 8.753541, 7.014472, 9.745265, 
    10.7747, 9.713295, 6.983955, 5.455486, 11.07452, 10.37136, 10.78256, 
    12.75255,
  63.23594, 62.197, 59.59195, 17.32729, 10.67617, 8.56212, 7.493298, 
    13.58891, 17.57162, 13.37139, 8.413488, 12.78106, 13.2591, 9.4663, 
    8.030831,
  59.28547, 53.8509, 61.5587, 23.90729, 16.07461, 11.61527, 5.848393, 
    8.176632, 16.85364, 19.41058, 9.543209, 14.50158, 12.96873, 11.97238, 
    8.440109,
  50.04458, 49.82516, 52.86028, 33.60735, 18.29867, 12.28313, 5.431341, 
    6.799468, 9.465259, 10.58261, 8.789017, 13.97831, 14.30961, 14.23154, 
    11.22473,
  46.43584, 42.42823, 45.2118, 24.56499, 16.84744, 13.92831, 10.8602, 
    6.379042, 8.344514, 11.31656, 8.001163, 10.01378, 14.01595, 15.85071, 
    13.01869,
  48.01973, 38.51752, 26.46797, 12.71989, 13.71717, 15.65554, 14.86861, 
    8.280451, 7.686664, 10.83334, 9.798966, 8.255592, 10.20977, 17.39069, 
    17.45062,
  48.0521, 39.10248, 14.32099, 8.298391, 7.458748, 11.04567, 16.42772, 
    24.64387, 23.64751, 23.58349, 12.23726, 8.161564, 9.572968, 14.65996, 
    16.15636,
  42.28028, 27.13686, 10.96229, 9.885885, 4.44673, 7.261267, 13.46045, 
    37.08798, 36.02269, 20.10816, 5.568185, 5.290951, 9.539105, 11.17949, 
    13.50675,
  6.877773, 9.037984, 9.104986, 7.109881, 5.704978, 6.094941, 3.25515, 
    9.411878, 11.94612, 13.64448, 16.42357, 10.98765, 10.34775, 11.42545, 
    12.44482,
  13.14207, 8.028597, 9.863694, 13.09799, 12.37592, 7.171238, 3.202533, 
    12.42135, 13.31201, 10.44944, 11.98978, 8.869003, 9.314709, 15.50725, 
    17.07323,
  30.80671, 32.14265, 25.34835, 18.28952, 12.34094, 10.14124, 4.86982, 
    5.71305, 10.02265, 10.50925, 10.67626, 8.402069, 7.492185, 12.41626, 
    15.85843,
  36.15508, 34.08738, 39.98062, 18.81739, 12.13618, 6.230558, 8.854513, 
    8.919893, 14.5953, 13.8439, 10.22269, 9.29283, 10.34161, 10.36787, 
    11.73156,
  46.07389, 30.57623, 39.37285, 23.54445, 15.00002, 13.82146, 12.66904, 
    11.38496, 16.11139, 19.59479, 10.46683, 9.945402, 10.55811, 10.2803, 
    11.31176,
  57.44955, 34.30546, 31.95851, 24.24259, 15.58712, 14.15919, 14.79177, 
    12.65418, 12.4473, 8.837792, 8.112703, 8.700965, 11.32683, 9.630307, 
    10.86571,
  65.69898, 40.15903, 26.43834, 11.46893, 14.18733, 13.99947, 15.89493, 
    17.62473, 15.77666, 11.8176, 10.25569, 10.30039, 11.04058, 10.86047, 
    8.496489,
  73.38629, 46.17716, 18.57071, 4.205355, 13.4908, 12.89226, 16.48267, 
    18.79839, 19.05816, 15.53961, 13.08444, 11.23819, 11.55291, 12.87622, 
    8.456088,
  67.27866, 40.19442, 13.19443, 3.579009, 5.335648, 12.28688, 16.15636, 
    25.9921, 29.07544, 27.04084, 16.81115, 12.65586, 11.56562, 12.19334, 
    11.37902,
  49.91341, 18.26696, 7.585292, 4.710471, 6.341158, 10.14496, 9.891314, 
    37.44408, 37.28421, 21.88426, 14.4512, 11.87831, 10.68866, 10.9725, 
    11.58968,
  6.715446, 12.32842, 15.40867, 13.5513, 11.59027, 11.82118, 10.94069, 
    12.2537, 12.28413, 17.73377, 16.90086, 15.43751, 17.44181, 12.21171, 
    17.78164,
  17.70734, 10.93483, 15.17389, 16.35677, 15.65972, 15.57414, 10.76095, 
    6.667201, 3.705227, 13.39162, 16.44334, 12.08938, 13.7738, 13.42055, 
    15.81255,
  35.43459, 25.01751, 21.38885, 18.77332, 15.44243, 15.40972, 7.542663, 
    5.690144, 8.874345, 14.487, 14.39789, 14.15691, 12.36062, 11.84439, 
    11.17253,
  48.96354, 32.76634, 36.03181, 20.20765, 14.65326, 12.49079, 14.93885, 
    6.875226, 9.13181, 16.90089, 16.40772, 14.27134, 14.52286, 10.31567, 
    10.18725,
  59.98302, 36.29417, 35.81968, 22.06321, 14.08583, 16.25264, 15.05528, 
    11.55524, 14.58602, 22.22334, 19.07607, 15.88473, 14.19593, 8.40904, 
    8.042676,
  62.94639, 41.53881, 31.816, 21.91334, 12.04593, 14.38371, 16.40047, 
    14.97195, 12.50569, 14.32856, 16.41163, 14.70934, 11.76592, 8.495184, 
    8.116351,
  58.74076, 42.3931, 28.86825, 12.40123, 12.77734, 14.38322, 18.00116, 
    18.13213, 17.18326, 17.54985, 17.13127, 14.40718, 12.7266, 11.28407, 
    5.468468,
  54.3919, 42.33194, 19.76437, 9.572264, 12.12735, 11.40301, 17.64375, 
    19.55089, 17.48983, 19.41254, 16.01506, 16.23544, 12.23507, 7.434124, 
    5.984286,
  45.92741, 32.06921, 7.809226, 9.44243, 10.58931, 9.54985, 13.95936, 
    25.2734, 29.087, 29.45703, 21.58056, 16.37145, 13.38892, 5.385533, 
    6.756722,
  32.37474, 14.16473, 7.048883, 9.296768, 9.717568, 4.097017, 10.80062, 
    34.12718, 36.08545, 20.31762, 17.90829, 13.71879, 11.6866, 3.71448, 
    8.768255,
  8.032938, 13.40899, 17.46134, 14.55382, 13.8927, 12.60248, 14.06647, 
    11.57778, 6.212943, 16.84036, 20.15572, 18.08376, 18.59307, 17.50483, 
    20.34146,
  14.15094, 15.83059, 16.80738, 15.31092, 17.03792, 14.64316, 12.82467, 
    3.282656, 2.676466, 10.93109, 16.07293, 13.44213, 10.77262, 11.60975, 
    20.65064,
  29.04327, 33.709, 24.82872, 18.05468, 10.74806, 17.03085, 8.667212, 
    6.448468, 3.290141, 13.33934, 12.1704, 15.54228, 12.62144, 12.23847, 
    13.95635,
  37.4792, 42.73972, 34.58543, 19.54142, 11.91254, 12.80322, 14.46933, 
    8.775954, 5.992656, 7.6039, 12.89282, 14.39744, 14.33007, 15.11819, 
    15.15899,
  50.61591, 42.19562, 31.38528, 17.47073, 9.34383, 8.746971, 9.051016, 
    9.576797, 11.56098, 16.10034, 16.2179, 13.13513, 15.83627, 11.39718, 
    7.911573,
  57.47873, 50.81962, 24.05222, 12.77381, 8.277163, 7.34896, 10.71494, 
    10.21269, 11.75575, 13.64055, 14.86159, 13.71863, 14.44407, 6.721284, 
    7.668416,
  61.46396, 56.14077, 30.6185, 12.49082, 11.37968, 8.764655, 9.78797, 
    11.54253, 12.21446, 11.31664, 8.989518, 11.02408, 16.12036, 8.084015, 
    9.628716,
  67.51611, 64.33193, 28.68892, 12.97747, 12.03119, 9.368281, 7.895267, 
    10.13105, 11.55603, 11.355, 11.10521, 13.39695, 16.42082, 13.65259, 
    14.91258,
  72.66519, 61.98514, 18.9039, 12.65535, 15.56976, 13.16374, 8.6936, 
    10.42161, 13.59324, 17.77401, 11.82845, 12.96494, 13.08655, 12.36268, 
    13.97696,
  61.59923, 36.33981, 19.61254, 21.14592, 17.80334, 12.85232, 10.34087, 
    14.54907, 16.15623, 13.56748, 13.05512, 15.82899, 7.782891, 13.37257, 
    16.93018,
  6.988168, 14.58731, 21.36469, 15.87329, 16.55819, 18.98514, 6.48487, 
    5.748143, 10.17361, 16.85793, 20.13411, 17.75896, 17.18468, 16.31911, 
    18.27447,
  13.14603, 14.73461, 19.53094, 18.19739, 22.31904, 21.99365, 8.283031, 
    5.871309, 3.533367, 5.052707, 7.642642, 10.68006, 9.154794, 14.33224, 
    17.89424,
  32.20904, 33.30395, 22.87098, 15.086, 14.7598, 13.67892, 13.41511, 
    8.261147, 5.752046, 3.779579, 4.820117, 6.423785, 8.890957, 12.05176, 
    13.87286,
  43.2401, 41.81089, 36.675, 18.37753, 10.34746, 11.7197, 12.03605, 13.41238, 
    8.015157, 6.624731, 9.026718, 7.559973, 9.274303, 14.49922, 13.0188,
  59.85962, 46.15721, 50.43934, 27.95314, 14.75616, 12.56081, 11.66955, 
    8.400148, 7.338661, 6.740156, 6.414222, 8.708827, 10.33078, 13.62807, 
    10.64329,
  70.78371, 66.94212, 58.70377, 28.18425, 14.54559, 14.30024, 13.28745, 
    12.534, 11.27554, 8.380885, 6.996848, 10.10637, 12.05523, 10.53325, 
    12.13315,
  80.68179, 82.66698, 67.88811, 15.67459, 11.52004, 8.546787, 8.493925, 
    7.819068, 7.813515, 4.67627, 12.11533, 11.08967, 10.03197, 9.201376, 
    13.22907,
  90.65591, 89.14076, 50.79412, 14.08298, 11.98691, 10.73949, 6.574195, 
    10.51063, 11.50758, 3.085277, 9.857298, 7.959059, 10.18751, 17.09851, 
    23.21509,
  91.80629, 82.54716, 35.17587, 14.06592, 14.89615, 13.17996, 10.21679, 
    13.03515, 12.18792, 4.601978, 7.524978, 5.916307, 8.924169, 22.22228, 
    21.27428,
  76.30461, 60.19405, 29.62939, 21.20521, 17.41319, 12.77367, 8.705235, 
    13.34109, 21.14364, 17.75307, 6.946431, 12.79927, 14.67774, 22.60614, 
    22.09202,
  5.758521, 4.144353, 15.40836, 7.154235, 8.318884, 10.00456, 6.684937, 
    8.629564, 8.519511, 13.71324, 17.23175, 16.61023, 15.32006, 16.20073, 
    17.88052,
  17.97244, 6.165878, 10.25692, 8.78434, 15.91778, 16.85887, 11.03248, 
    8.31284, 9.212755, 11.96214, 14.97437, 12.41554, 11.1913, 14.96146, 
    15.82956,
  27.89193, 25.78156, 15.33184, 5.338192, 9.385045, 17.36632, 13.61965, 
    7.306216, 11.88844, 12.18046, 10.44772, 11.70048, 6.824229, 14.85359, 
    14.33676,
  39.82492, 36.1503, 28.85627, 10.21252, 6.616817, 13.24106, 15.91691, 
    10.94572, 4.839775, 12.42847, 9.137789, 11.4031, 10.59546, 15.14121, 
    11.95374,
  52.76485, 37.26874, 32.64409, 11.17803, 6.369572, 8.626211, 11.58239, 
    10.01306, 9.633202, 8.413174, 14.12192, 10.60822, 9.783205, 17.21995, 
    5.587873,
  61.12614, 50.61601, 27.63655, 16.08952, 12.1036, 9.042233, 9.617579, 
    8.030116, 8.922023, 4.935393, 11.73426, 13.60527, 10.4189, 7.651951, 
    5.035066,
  70.51151, 59.91182, 35.5963, 15.06801, 11.05229, 8.103308, 6.864552, 
    9.055945, 8.437325, 3.462355, 6.688447, 13.19036, 13.73597, 7.310639, 
    10.22237,
  79.30586, 69.73057, 32.66395, 13.81376, 16.25866, 9.875713, 10.17919, 
    12.12691, 8.070483, 14.09785, 9.442122, 8.119615, 14.42429, 10.8417, 
    18.06678,
  83.64369, 68.21067, 22.79014, 13.05622, 10.89057, 6.844739, 9.962316, 
    12.59793, 13.95575, 19.05423, 7.614426, 10.33541, 13.91198, 13.62971, 
    20.87919,
  70.19955, 48.85879, 18.75615, 14.90191, 9.480453, 7.694837, 9.683227, 
    18.28109, 23.41896, 17.13432, 10.26805, 13.40421, 10.24373, 15.69835, 
    17.24927,
  3.41916, 6.399547, 18.82784, 15.36017, 14.27095, 10.07725, 8.130836, 
    6.48456, 7.512996, 17.87113, 17.43375, 12.82426, 16.01165, 11.66127, 
    19.28174,
  5.51868, 5.364141, 8.640143, 10.97676, 20.33237, 17.72381, 6.507685, 
    8.911247, 7.405794, 12.67116, 13.49379, 9.097746, 8.511516, 12.47788, 
    16.3798,
  10.5684, 8.535389, 5.734289, 9.134773, 12.80533, 18.47189, 8.1623, 
    8.924248, 8.796438, 11.067, 8.351424, 7.109838, 8.812653, 8.957376, 
    15.21499,
  24.53983, 19.74155, 15.78221, 3.312295, 3.153027, 9.728602, 15.019, 
    11.14214, 7.279611, 11.29912, 8.347478, 5.233195, 11.348, 6.71005, 
    13.55889,
  43.03109, 27.51895, 21.33971, 4.99752, 4.897422, 4.526624, 6.639979, 
    9.573494, 8.768583, 7.433813, 12.49356, 6.500053, 7.392779, 10.59538, 
    4.798046,
  56.19929, 37.51949, 16.37327, 10.72934, 7.332155, 3.402068, 5.102149, 
    8.082973, 10.55772, 9.216221, 17.21273, 11.5663, 14.17847, 5.702229, 
    8.225226,
  62.46968, 44.52326, 22.8886, 6.648243, 10.00295, 1.573771, 3.914957, 
    6.099509, 10.11058, 8.476004, 15.01202, 11.41865, 12.74573, 5.297674, 
    10.84335,
  70.60891, 55.17264, 22.48785, 7.664191, 10.72282, 4.231557, 3.434581, 
    9.633255, 7.798875, 12.0011, 15.59923, 12.59197, 7.172909, 8.505163, 
    13.81146,
  77.33337, 59.60653, 16.78634, 12.37951, 7.364282, 9.732648, 11.63833, 
    15.45365, 13.27501, 14.49084, 7.570954, 8.280279, 4.959667, 17.00337, 
    12.59407,
  64.3293, 41.51203, 11.46606, 15.39434, 11.10596, 11.36327, 14.73824, 
    23.50173, 14.48728, 16.6015, 7.786547, 12.56713, 5.096466, 12.38565, 
    10.60094,
  3.470348, 1.598784, 4.286116, 2.00978, 4.953644, 5.755564, 4.761757, 
    6.976323, 4.407186, 15.94563, 12.42478, 8.111403, 12.87918, 15.64314, 
    24.05506,
  1.931205, 1.620348, 1.138003, 2.754, 8.181417, 7.480316, 5.592053, 
    7.792187, 5.140991, 11.22696, 17.23702, 5.645305, 6.772675, 14.96106, 
    20.00131,
  6.918729, 6.226316, 3.567798, 6.211318, 8.167244, 10.20765, 6.94675, 
    8.520072, 6.10383, 8.497935, 7.714614, 7.207084, 6.707394, 6.506366, 
    16.57839,
  32.41836, 29.76659, 24.94728, 8.978434, 5.023924, 6.507331, 7.904821, 
    11.04634, 5.869526, 8.261843, 9.68153, 8.361945, 4.680731, 4.542126, 
    11.71207,
  50.73875, 37.22104, 28.47091, 7.916408, 5.340957, 4.057829, 6.047693, 
    9.448908, 10.40038, 8.844907, 11.149, 13.91133, 6.269876, 3.461936, 
    4.675937,
  65.80371, 47.85772, 26.43733, 8.402964, 8.092356, 5.977933, 6.912254, 
    7.496046, 11.67754, 7.759419, 17.37096, 16.59704, 10.5872, 2.700231, 
    4.812826,
  70.47691, 45.01426, 24.39629, 9.575099, 8.485152, 6.672758, 9.777321, 
    4.701339, 8.570476, 6.121338, 19.71607, 16.78115, 15.09296, 7.233111, 
    12.84766,
  73.842, 50.8105, 18.43439, 4.838503, 7.411382, 6.732572, 5.453052, 
    6.679747, 7.18866, 4.50483, 14.86724, 17.95739, 7.101927, 9.65196, 
    18.54373,
  77.81596, 56.04181, 9.562604, 7.403165, 6.917504, 5.547619, 5.945759, 
    9.780274, 12.12716, 6.198795, 19.65711, 16.99339, 5.172892, 14.00076, 
    20.04161,
  66.02103, 42.57501, 13.39648, 13.25265, 6.786126, 7.434832, 9.834175, 
    17.59281, 14.81393, 12.62055, 22.31433, 18.86478, 6.055626, 17.35842, 
    16.52699,
  4.440773, 0.935373, 1.836842, 5.136169, 4.805624, 12.32139, 12.42274, 
    11.13585, 10.00546, 14.8221, 15.35668, 10.60103, 17.1867, 18.0545, 
    24.94994,
  1.335128, 0.4035858, 1.225007, 1.461839, 14.43114, 21.05404, 15.1633, 
    10.74721, 7.030887, 4.979886, 17.15174, 8.44484, 8.978731, 18.4598, 
    17.50628,
  5.732718, 5.54884, 3.289299, 2.031373, 12.7457, 21.05577, 11.96608, 
    3.418024, 8.012986, 3.716095, 11.89727, 10.11971, 8.672002, 7.580273, 
    11.71469,
  29.66675, 32.18366, 26.26745, 12.37096, 6.644321, 12.12986, 20.47025, 
    7.247484, 4.814388, 3.125429, 1.89548, 2.071212, 7.695697, 5.756413, 
    12.17127,
  52.99577, 40.11333, 32.91888, 9.231688, 11.56434, 11.46352, 9.987489, 
    11.40099, 5.459105, 8.754288, 4.195682, 4.817511, 7.159888, 6.330563, 
    7.506321,
  59.96083, 43.57471, 22.52403, 6.040102, 9.66155, 6.105524, 6.197764, 
    5.165223, 9.979511, 9.40985, 11.1813, 5.463935, 6.741442, 9.117826, 
    15.16746,
  58.01385, 40.16736, 21.15391, 5.669014, 7.738391, 8.493499, 6.197567, 
    5.401595, 8.03669, 6.363265, 8.122191, 7.36571, 9.031854, 13.11964, 
    16.15543,
  53.65418, 42.31271, 18.71255, 3.544302, 9.441879, 5.055749, 8.689484, 
    11.50783, 8.766451, 5.689193, 11.74093, 13.06111, 14.80841, 17.97929, 
    18.60157,
  56.9262, 40.20219, 11.14954, 13.12771, 11.85514, 8.119285, 11.90206, 
    14.77882, 11.65609, 6.389435, 12.8622, 14.37332, 15.31828, 17.69933, 
    16.24724,
  49.78788, 29.56965, 7.989432, 10.98966, 8.315238, 9.673043, 14.62434, 
    21.16737, 14.78967, 14.89439, 14.99697, 15.1513, 15.85429, 14.2468, 
    14.5211,
  1.052689, 0.7501506, 2.304278, 6.520503, 9.03481, 10.45967, 9.76571, 
    11.68762, 13.10699, 22.29563, 21.91487, 19.61813, 21.82584, 21.25393, 
    23.95694,
  5.347018, 2.48928, 1.567117, 8.379306, 11.05763, 12.55954, 11.41524, 
    11.97271, 11.9905, 16.91637, 18.32184, 17.37962, 15.50281, 24.7383, 
    24.90141,
  11.82696, 9.254821, 3.571768, 3.671124, 8.77551, 25.10318, 10.18189, 
    8.902757, 11.50325, 8.047616, 11.18657, 13.59886, 9.461036, 8.53809, 
    16.05809,
  19.97728, 23.08619, 20.62702, 3.566925, 1.721893, 7.676376, 22.00702, 
    6.438002, 12.17006, 13.12591, 11.26496, 6.91775, 2.312179, 4.580326, 
    12.12995,
  34.00259, 28.56869, 24.14772, 7.25853, 2.584663, 16.26124, 15.26428, 
    17.72865, 10.89865, 10.07385, 4.452502, 2.635291, 3.263027, 6.193014, 
    13.91254,
  40.67054, 35.08469, 26.02567, 9.967152, 11.24074, 13.09078, 12.05595, 
    8.71802, 9.849376, 5.435528, 5.86449, 3.433906, 8.025795, 10.10168, 
    14.84558,
  43.42514, 36.2203, 33.22927, 10.11053, 10.36821, 9.834541, 8.866509, 
    1.948306, 8.311742, 11.90319, 11.15211, 11.1599, 10.04215, 13.69344, 
    14.88597,
  44.08069, 47.11649, 25.80785, 7.070641, 7.454569, 3.390037, 3.663836, 
    4.851125, 3.612683, 9.46818, 8.89183, 10.30584, 13.2621, 16.57192, 
    18.10151,
  50.11969, 42.54392, 12.30128, 13.18132, 10.55694, 9.530314, 8.521116, 
    7.470567, 6.007597, 10.76812, 11.48088, 11.41694, 15.06773, 16.67263, 
    17.39165,
  43.7768, 30.97469, 11.94502, 14.8698, 11.80369, 10.0062, 8.449228, 
    7.469568, 11.11986, 14.74647, 17.2108, 14.0577, 16.36047, 15.42101, 
    16.7048,
  2.144505, 6.080233, 11.77136, 10.63235, 10.84712, 8.777886, 5.925197, 
    6.006824, 6.056172, 14.97975, 17.06913, 10.86444, 15.12529, 19.03837, 
    26.41262,
  4.324714, 3.248855, 4.269198, 11.75312, 14.89522, 16.16823, 7.092555, 
    6.821553, 6.993706, 10.46843, 15.31244, 10.75604, 9.87288, 22.95229, 
    23.72966,
  14.44616, 15.47274, 12.28631, 4.3065, 11.48192, 16.73623, 8.197906, 
    8.827467, 6.828997, 6.53932, 4.903303, 7.693083, 6.531944, 9.864511, 
    17.83292,
  27.76869, 29.33716, 22.60102, 7.551906, 4.186845, 14.31643, 20.86104, 
    9.005829, 4.254632, 14.79586, 13.02174, 7.047089, 6.689968, 8.532854, 
    12.9825,
  43.70464, 27.53937, 23.58735, 11.00887, 2.926831, 10.04625, 11.55812, 
    11.93144, 11.33844, 12.61861, 12.73752, 8.089684, 8.910219, 6.922346, 
    8.107888,
  44.6056, 36.81124, 28.27929, 10.91459, 5.142582, 10.31083, 10.61095, 
    6.773502, 9.353306, 8.319029, 6.476787, 6.17582, 5.690903, 9.746386, 
    13.07007,
  50.15731, 45.59332, 26.10708, 11.27542, 10.68097, 10.55702, 8.129569, 
    7.231575, 9.371279, 7.022415, 9.401423, 9.522603, 9.287497, 10.68174, 
    15.37757,
  57.92001, 49.67648, 18.65388, 8.40789, 12.57255, 8.703609, 6.032892, 
    5.045874, 1.99284, 8.495312, 7.718342, 8.015544, 11.53883, 13.41586, 
    14.53105,
  51.43838, 44.08336, 12.96223, 14.38689, 13.09901, 6.788805, 2.507638, 
    2.512784, 9.483463, 11.1537, 7.875422, 7.440582, 10.07455, 13.05326, 
    14.95724,
  38.07165, 32.0876, 15.74259, 13.26029, 7.405261, 5.007724, 4.403766, 
    6.736693, 11.77304, 14.58883, 8.139724, 12.23351, 13.05124, 13.96414, 
    14.79467,
  -6.264443, -26.91908, -15.76665, -14.22732, -9.858509, -8.358551, 
    -5.107698, -4.201129, -2.115158, 5.386226, 12.57308, 12.59485, 20.80372, 
    15.4069, 24.27922,
  -18.38193, -18.65717, -13.39192, -10.53487, -14.00443, -3.708397, 
    -3.870043, -0.6874745, 1.677173, 4.733657, 14.41184, 10.46583, 6.928644, 
    21.46854, 20.85795,
  -11.42867, -12.64906, -15.055, -11.10361, -3.624645, 4.983511, 2.076541, 
    2.070671, 5.002807, 6.448273, 7.043623, 6.686728, 4.527479, 2.530141, 
    10.42522,
  -3.110432, -7.104531, -4.042145, 0.365202, 1.057706, 6.749112, 11.30297, 
    4.323905, 5.341418, 5.156525, 4.829545, 3.334956, 14.51175, 14.17705, 
    7.060547,
  8.241092, 6.544611, 16.37358, 11.58074, 5.05667, 8.749697, 15.82717, 
    18.77068, 12.63701, 9.120246, 6.616762, 12.17869, 15.13031, 13.18904, 
    11.14101,
  60.11948, 60.38732, 47.54123, 20.83272, 14.67541, 10.84366, 7.214947, 
    7.644832, 10.11096, 4.429972, 6.977515, 1.881778, 14.95483, 13.03328, 
    9.512226,
  94.09591, 95.78027, 50.21995, 14.34904, 9.104912, 5.580969, 3.991683, 
    5.047433, 14.06457, 16.1166, 12.34384, 7.208489, 8.774491, 10.36505, 
    8.386978,
  102.5459, 95.9594, 30.68114, 8.209728, 7.019981, 17.36933, 11.21885, 
    16.42733, 13.11646, 13.97365, 5.993882, 4.680654, 5.620656, 11.02952, 
    11.60903,
  83.43255, 67.17517, 14.00094, 12.93116, 18.39815, 13.02088, 12.63881, 
    17.56543, 17.72518, 16.12977, 6.029284, 10.73522, 11.40555, 13.88137, 
    11.8197,
  55.26129, 37.79902, 18.34386, 15.96182, 16.33379, 19.56311, 18.5231, 
    17.8549, 15.714, 17.65476, 10.78538, 13.64742, 12.78928, 10.38169, 
    12.59964,
  11.70683, 18.3653, 22.05735, 21.35564, 17.823, 11.51751, 4.735464, 
    1.644286, 0.6695574, 1.7284, 0.05061525, -0.4486395, -1.308524, 
    0.7032454, 1.888583,
  18.97146, 27.81887, 29.98421, 19.7122, 13.44842, 7.678746, 0.9938695, 
    -0.2975031, -0.7553866, -0.8598412, -1.186297, -1.802809, -1.537413, 
    5.004765, 4.362836,
  43.34818, 48.19139, 28.62408, 9.719898, 6.125013, 10.12792, 1.395843, 
    3.173033, 2.980876, 2.706105, 1.875983, 2.172699, 2.459804, 4.02887, 
    8.577732,
  63.40197, 50.46941, 31.787, 13.47458, 2.789614, 4.253912, 15.40375, 
    10.02647, 11.71651, 9.065326, 9.387792, 7.628645, 6.484832, 6.159632, 
    10.56827,
  64.80869, 44.49906, 43.2963, 20.05289, 11.14091, 10.49652, 19.38328, 
    15.83837, 10.018, 13.70175, 10.7021, 9.349363, 9.265002, 11.87735, 
    16.37517,
  60.02435, 63.00847, 55.74553, 24.50939, 17.19982, 14.48721, 11.64689, 
    15.61131, 15.34928, 13.88967, 13.69555, 12.09923, 14.02626, 15.73234, 
    17.01669,
  59.84966, 68.89664, 51.08505, 20.02444, 14.9987, 12.00825, 9.590569, 
    8.552321, 9.06249, 14.59465, 15.66996, 16.18767, 16.59928, 16.53682, 
    16.47891,
  63.06342, 71.44791, 35.47479, 21.75402, 18.09976, 13.70917, 8.010562, 
    6.203384, 5.150041, 8.54986, 8.944345, 12.02746, 13.36598, 15.92315, 
    15.14301,
  63.22895, 56.7981, 25.15486, 24.76536, 23.66552, 23.07464, 14.9363, 
    13.58038, 10.05381, 5.923649, 6.326432, 6.706583, 10.55296, 11.04525, 
    16.36906,
  52.81639, 37.13614, 22.14342, 21.82749, 19.80278, 19.42467, 20.10823, 
    11.49558, 12.55115, 11.77539, 10.3223, 10.45848, 13.3746, 13.66767, 
    11.12703,
  8.61282, 13.19019, 20.99467, 16.19617, 20.3016, 15.36298, 14.3207, 
    13.00137, 14.2318, 19.47133, 20.27602, 16.66297, 21.82516, 18.87853, 
    19.57307,
  8.931422, 15.11815, 20.62332, 15.87441, 19.08537, 23.65466, 16.63254, 
    13.53898, 15.80025, 15.24474, 19.83048, 18.36449, 11.24722, 17.9357, 
    14.3031,
  19.25789, 27.46902, 30.80114, 15.90826, 13.28791, 29.64966, 20.60552, 
    9.186102, 14.88309, 14.16381, 16.24588, 17.43419, 16.31824, 8.04283, 
    7.489881,
  33.37011, 39.16499, 42.05682, 23.48958, 5.646733, 14.72783, 23.27662, 
    13.37562, 12.19009, 16.19726, 16.47249, 17.39671, 15.90833, 5.475546, 
    2.692462,
  60.91443, 50.03797, 50.10135, 13.38111, 3.266021, 3.95399, 18.40044, 
    12.40837, 15.43968, 22.1876, 22.15912, 15.78539, 14.36921, 3.224076, 
    1.365597,
  77.59283, 62.79076, 42.37325, 6.189962, 2.23694, 3.470289, 14.16137, 
    13.99688, 16.2916, 15.16584, 17.86453, 19.82048, 11.02004, 4.586681, 
    3.112336,
  70.79397, 61.76108, 35.25137, 10.60156, 3.9342, 4.566758, 3.913487, 
    10.88775, 9.471572, 5.648141, 7.957106, 15.45097, 7.279519, 5.201444, 
    6.92552,
  60.00951, 51.22642, 21.07968, 13.89341, 13.54323, 13.45732, 5.23887, 
    2.781708, 7.240596, 2.539653, 11.83644, 11.86721, 5.666739, 7.145016, 
    10.83524,
  48.17029, 33.7452, 13.10373, 14.78285, 16.53254, 17.34003, 7.411523, 
    3.329941, 2.412639, 2.471824, 7.20998, 10.91452, 5.743856, 6.59342, 
    13.47913,
  39.17635, 22.23773, 13.06163, 17.83344, 17.48438, 12.3527, 11.97118, 
    5.203453, 4.915187, 8.222867, 9.967899, 8.556453, 7.747008, 7.040644, 
    14.66173,
  20.03617, 28.47845, 22.9596, 19.43888, 12.35705, 7.552725, 7.951385, 
    8.204475, 10.36616, 22.38078, 27.66355, 19.66032, 24.73537, 27.36381, 
    31.12869,
  36.33786, 32.88894, 24.07356, 17.29417, 11.96215, 10.47375, 6.214447, 
    4.58973, 6.385615, 14.19298, 24.66607, 12.97644, 8.538712, 20.45544, 
    24.3003,
  53.00218, 53.16099, 39.07163, 16.74723, 12.08408, 18.64069, 7.005366, 
    5.478376, 8.785187, 8.421756, 7.851758, 10.3525, 13.16957, 16.82614, 
    18.87516,
  70.74493, 70.52991, 58.09069, 30.03556, 12.2431, 20.63652, 16.11272, 
    10.27007, 10.24782, 6.869072, 4.841591, 6.570316, 14.98638, 19.75104, 
    11.69125,
  81.48768, 75.42994, 75.38001, 30.59463, 15.67185, 14.75722, 25.4605, 
    20.36999, 15.87502, 9.386223, 4.801088, 7.147267, 16.55444, 12.89338, 
    3.84858,
  67.9754, 74.98195, 64.1483, 28.48201, 17.92754, 16.86305, 16.5106, 
    19.93697, 17.25578, 17.30004, 13.91673, 10.50238, 14.71941, 4.784759, 
    0.9057176,
  54.70329, 68.24432, 50.05915, 19.93969, 22.77242, 23.77393, 15.28859, 
    13.2588, 15.61072, 14.75333, 4.612092, 13.49261, 12.33383, 3.117588, 
    1.396059,
  45.45616, 55.45109, 30.67289, 20.75136, 19.70855, 17.69798, 10.56267, 
    3.61329, 11.69045, 3.661052, 5.698514, 13.33938, 7.72693, 4.184271, 
    3.755773,
  40.57389, 36.65299, 16.23867, 15.14881, 13.25589, 10.88988, 11.23814, 
    2.641629, 2.408215, 4.397508, 11.70621, 7.958366, 4.879762, 5.678761, 
    8.886791,
  32.68651, 22.5894, 17.56008, 12.96997, 11.41831, 2.084443, 1.97507, 
    2.42297, 3.481315, 11.63773, 8.83126, 8.441237, 7.505974, 12.64687, 
    17.22169,
  12.3696, 11.43908, 16.33296, 27.32851, 29.44186, 26.45038, 18.19617, 
    14.5107, 11.6636, 12.78257, 12.2052, 14.1265, 17.96175, 20.27814, 37.82316,
  6.6684, 8.054525, 15.83793, 25.06632, 33.00315, 32.24537, 18.96839, 
    14.11455, 12.90941, 11.63466, 15.8978, 12.28305, 15.34391, 23.97062, 
    27.87721,
  4.965343, 11.8887, 27.70721, 22.52083, 22.62855, 29.97397, 21.65795, 
    13.96914, 11.10402, 9.861292, 10.0142, 10.54698, 10.48139, 8.413127, 
    16.50465,
  6.393619, 13.01903, 33.59111, 30.12408, 19.66498, 21.61675, 26.6084, 
    21.21212, 14.59842, 9.730254, 10.81234, 9.766061, 6.658182, 5.31481, 
    17.05374,
  6.100163, 11.4166, 31.31106, 19.88482, 17.46712, 23.29917, 25.78482, 
    16.13692, 12.89693, 12.20192, 8.947715, 8.696534, 8.267585, 5.919476, 
    2.787603,
  9.317011, 14.01189, 22.48755, 18.73844, 18.6737, 19.22013, 17.70699, 
    19.72077, 16.17925, 14.77545, 12.40693, 9.768432, 8.042312, 2.154536, 
    0.6904411,
  20.35775, 20.86621, 17.46413, 15.11347, 17.96159, 17.43948, 16.81113, 
    17.61609, 19.20505, 14.48639, 10.64581, 11.40744, 6.702174, 1.546048, 
    1.205845,
  33.50116, 27.61531, 10.99356, 13.38119, 14.7474, 14.79862, 15.79077, 
    16.2347, 16.48611, 11.5688, 12.98801, 11.10876, 6.545703, 2.791526, 
    2.983909,
  45.79203, 27.04623, 6.097048, 9.613022, 13.90335, 14.38704, 13.8635, 
    4.090816, 11.15982, 15.4584, 11.72145, 9.545033, 6.839579, 5.133961, 
    5.931625,
  37.89606, 19.62281, 11.10623, 7.032169, 10.89777, 11.18698, 5.749728, 
    3.454597, 15.48616, 17.56014, 10.52631, 10.93269, 10.71568, 10.4501, 
    13.09787,
  11.53955, 4.584304, 4.004596, 6.578456, 10.80242, 8.202847, 5.775881, 
    6.588036, 19.79609, 25.82554, 21.78052, 20.73399, 26.07714, 25.55074, 
    31.75487,
  2.56271, 1.916862, 3.355546, 11.77007, 16.01582, 10.97761, 5.641521, 
    6.829933, 15.49628, 14.55171, 15.7789, 10.77978, 7.997125, 21.44116, 
    24.06103,
  4.893883, 7.992308, 15.02233, 12.03758, 10.56381, 17.79942, 9.184389, 
    7.480519, 13.57949, 12.81813, 10.62761, 7.043021, 7.40087, 8.3178, 
    11.75899,
  5.914086, 9.519802, 20.79112, 21.24557, 5.641688, 12.31047, 23.06036, 
    12.16288, 13.7459, 15.1533, 12.0651, 6.243584, 5.965768, 7.41121, 9.280957,
  13.50502, 6.534273, 12.67628, 12.8139, 8.969102, 8.822799, 17.46134, 
    14.95861, 14.30583, 19.43762, 13.20758, 5.973072, 6.169975, 7.93812, 
    9.929553,
  27.25586, 10.96496, 3.45327, 7.58877, 13.01471, 14.15108, 12.51193, 
    15.73993, 17.46627, 18.12475, 14.70452, 8.165968, 6.391984, 8.470404, 
    11.57528,
  34.92734, 27.95017, 10.65139, 6.149621, 5.730191, 7.988264, 8.714106, 
    13.12014, 14.2493, 18.06724, 11.9866, 9.625648, 7.901898, 11.50998, 
    12.4963,
  41.62952, 33.36133, 11.67766, 10.24133, 6.294, 5.970921, 6.498485, 
    10.67491, 19.09879, 16.62603, 11.88993, 11.10848, 11.00591, 11.5806, 
    11.11769,
  50.97833, 39.90852, 10.63669, 7.109428, 8.186041, 6.260462, 11.02906, 
    4.084928, 16.882, 17.67501, 10.76051, 12.14578, 11.99203, 11.33028, 
    10.74888,
  38.0696, 31.41508, 15.99712, 8.613798, 4.974508, 8.807147, 12.19332, 
    6.282895, 18.51908, 20.70601, 13.57399, 11.98083, 11.72364, 11.57351, 
    10.61001,
  7.832784, 15.51733, 20.36206, 15.81406, 11.82652, 13.03029, 3.353928, 
    3.476107, 9.31391, 25.0873, 24.85071, 19.58102, 23.80264, 23.02835, 
    24.99666,
  18.63339, 24.91558, 25.88132, 15.16949, 21.17362, 14.92909, 3.293533, 
    5.060398, 4.38993, 21.21821, 20.02078, 14.6996, 16.61095, 22.44303, 
    23.11859,
  32.46791, 37.34135, 33.59319, 13.05697, 14.40037, 16.22461, 6.586367, 
    12.30525, 5.353866, 16.71501, 14.67529, 13.88341, 13.20163, 12.08605, 
    18.23815,
  48.22322, 47.82127, 37.6501, 18.5605, 4.24967, 9.665717, 17.65432, 
    12.36127, 8.119591, 18.18344, 15.31989, 11.97963, 11.03445, 10.65961, 
    13.55728,
  59.10706, 44.28194, 32.73224, 10.14074, 3.267872, 9.099473, 15.18804, 
    20.18185, 14.28772, 19.80173, 12.791, 11.30857, 10.91973, 8.573812, 
    8.353578,
  61.69434, 38.69693, 22.01244, 8.525206, 7.001395, 9.737794, 7.471753, 
    13.61797, 12.09812, 16.54107, 15.31004, 11.38784, 10.17301, 5.7992, 
    4.280759,
  70.92319, 55.34903, 30.35342, 11.14319, 9.207504, 13.70141, 15.1849, 
    17.76607, 9.497787, 14.41115, 11.77877, 10.13908, 8.086697, 4.005731, 
    2.899902,
  77.15557, 62.08293, 25.91095, 16.24067, 19.4165, 17.3907, 15.85449, 
    9.582596, 14.80202, 13.79603, 14.59609, 10.30972, 6.186405, 4.677367, 
    4.301747,
  74.45507, 50.45792, 19.07707, 16.43457, 18.4827, 18.74096, 11.53669, 
    12.19673, 15.20178, 15.90902, 14.19071, 8.074122, 4.971472, 6.439032, 
    3.90723,
  58.00768, 37.44032, 20.68603, 18.49792, 18.08877, 12.81313, 13.0739, 
    16.53733, 17.7355, 18.28947, 16.0418, 8.177767, 4.728948, 5.468945, 
    4.602667,
  20.67292, 26.56934, 23.47156, 7.825364, 9.216705, 11.70887, 6.522962, 
    6.608855, 11.71482, 25.25801, 23.74709, 20.79641, 16.18163, 15.19668, 
    16.94449,
  37.87484, 29.20663, 20.33151, 9.75684, 19.78157, 21.49301, 11.19969, 
    15.26942, 10.14338, 19.44829, 23.08555, 12.90732, 9.230033, 18.12941, 
    17.62198,
  44.79375, 35.39701, 29.74194, 17.28862, 18.40137, 23.56784, 21.528, 
    15.69101, 12.26848, 15.52848, 16.692, 11.41351, 10.13598, 6.100878, 
    9.381322,
  50.43176, 35.28436, 29.80159, 25.44327, 16.85144, 20.45393, 18.07369, 
    14.47473, 12.17739, 17.38238, 14.10551, 12.19654, 7.631859, 6.890477, 
    9.226314,
  51.28371, 32.61539, 30.50114, 17.97676, 15.38342, 17.7725, 18.80578, 
    12.11542, 10.13604, 22.32904, 13.51435, 11.2659, 8.259786, 9.657365, 
    8.75991,
  54.15301, 37.31388, 30.04454, 18.48675, 18.57289, 17.55347, 15.82106, 
    11.66006, 12.9175, 15.62854, 18.17707, 10.88723, 8.956675, 9.8673, 
    9.064577,
  58.7838, 45.51759, 28.29448, 17.20693, 19.59076, 18.28929, 17.01397, 
    15.92901, 12.30023, 13.85371, 14.23008, 12.43202, 9.744147, 10.75056, 
    7.833069,
  65.92616, 49.49175, 22.30115, 19.82412, 20.136, 18.26906, 18.30077, 
    17.79747, 13.94866, 13.12813, 14.78594, 11.93674, 10.24946, 9.705562, 
    6.696263,
  65.51857, 40.58012, 15.52067, 19.59216, 18.99566, 18.72129, 18.05757, 
    19.56, 16.56663, 16.17914, 12.83287, 11.98842, 10.56473, 7.074993, 
    3.998869,
  52.58772, 28.8831, 19.05426, 20.81444, 19.4239, 19.23461, 22.09691, 
    23.84362, 18.58982, 18.17477, 14.23201, 11.86255, 9.178358, 6.593968, 
    3.302645,
  13.30849, 21.23796, 24.67132, 15.3088, 18.35317, 19.88028, 15.53869, 
    14.23194, 14.17015, 19.9379, 21.18303, 19.68615, 25.08701, 24.61969, 
    23.32995,
  25.82377, 26.11526, 24.64007, 20.30181, 27.11903, 27.02014, 16.5522, 
    13.41188, 14.98052, 15.70827, 19.66776, 15.35845, 11.26658, 17.49016, 
    21.91789,
  33.23355, 31.54807, 31.22598, 24.42302, 20.28308, 23.47053, 22.38128, 
    14.69296, 10.37217, 11.12518, 13.53461, 9.407236, 8.566299, 7.120051, 
    10.81052,
  36.86235, 31.09943, 32.91282, 26.91268, 15.52146, 21.70727, 20.20762, 
    17.44453, 12.05737, 13.51574, 10.47309, 8.924372, 8.737784, 7.275603, 
    5.98844,
  35.9502, 29.2996, 35.50156, 21.71711, 18.94692, 16.87445, 18.99889, 
    11.15111, 9.965952, 17.23323, 10.87008, 7.404287, 7.618285, 6.613521, 
    3.796123,
  34.68417, 32.40396, 34.8422, 19.57869, 20.65826, 19.53238, 13.73627, 
    9.605035, 9.175706, 11.32212, 12.3243, 5.563505, 9.083276, 9.363367, 
    5.918387,
  34.07454, 36.35489, 30.04441, 16.78554, 21.34293, 22.45398, 15.47357, 
    10.09307, 9.242736, 7.870856, 7.475092, 4.55808, 6.775396, 11.27333, 
    9.387296,
  35.93103, 41.21257, 23.27297, 20.68091, 22.67832, 22.55381, 15.69433, 
    10.23979, 9.947652, 7.719276, 5.569939, 3.437488, 5.100147, 6.968444, 
    8.893247,
  38.32018, 35.99499, 17.95364, 20.43704, 22.16354, 22.1634, 16.62886, 
    10.7896, 8.216588, 5.688432, 3.743183, 3.451274, 4.23865, 4.790259, 
    6.495662,
  32.68859, 27.81971, 18.2824, 22.40644, 21.84753, 22.9868, 15.19622, 
    11.73853, 7.382404, 7.080549, 5.292193, 3.97531, 4.079859, 4.254381, 
    4.468119,
  12.65716, 19.09266, 20.42741, 18.08443, 17.49421, 23.57756, 14.20006, 
    15.07064, 13.9286, 18.381, 17.49862, 12.85396, 16.64833, 14.47728, 10.4122,
  21.38442, 14.22497, 19.57705, 20.17506, 28.21524, 30.47487, 15.38035, 
    14.08881, 10.45937, 15.36286, 17.39279, 13.39614, 11.76848, 16.8594, 
    12.75409,
  23.42347, 19.51081, 25.46827, 21.6217, 21.57245, 22.7147, 21.81214, 
    13.91344, 9.990849, 12.11442, 14.51061, 14.39674, 13.48238, 12.35741, 
    11.27421,
  23.96582, 27.09156, 32.99677, 26.34299, 16.50054, 16.36147, 16.93416, 
    19.34787, 13.18003, 11.21695, 12.42649, 13.68014, 12.3999, 11.70058, 
    9.590538,
  25.53042, 30.97597, 36.75995, 19.32753, 16.04509, 12.38972, 11.19022, 
    15.20962, 12.97391, 18.75768, 12.54016, 11.37887, 9.487269, 9.299488, 
    8.538425,
  29.48817, 36.75145, 29.6939, 16.32043, 18.08001, 12.13124, 9.284995, 
    8.157001, 12.18583, 11.75763, 11.66641, 11.1839, 8.900006, 8.312118, 
    9.749546,
  34.7758, 42.00829, 22.87277, 15.81701, 16.90415, 13.03114, 10.56665, 
    9.834696, 8.142509, 8.789031, 9.513555, 9.465465, 8.859795, 11.95677, 
    12.30939,
  39.1841, 42.68778, 18.21285, 16.27877, 14.29444, 12.23458, 9.763014, 
    8.693445, 6.974805, 7.533439, 8.496694, 7.560774, 6.406343, 9.254333, 
    8.491739,
  42.62754, 33.8363, 11.78592, 17.74451, 13.31945, 10.67335, 8.193717, 
    6.917278, 4.746682, 4.174281, 5.987788, 5.212744, 3.411124, 2.03503, 
    4.665701,
  35.34274, 21.28841, 12.82498, 12.73258, 9.706232, 9.897425, 7.9382, 
    5.57759, 5.027272, 6.562498, 6.732523, 4.949568, 4.570282, 3.297996, 
    4.968776,
  11.45366, 16.12818, 14.75826, 16.1904, 14.7556, 17.37564, 12.17195, 
    11.26358, 9.68688, 17.66843, 18.08853, 13.98657, 19.48891, 19.3997, 
    11.21605,
  20.99311, 13.71218, 15.04628, 10.45013, 17.66277, 16.71913, 10.87524, 
    10.31149, 7.954154, 9.381289, 15.92948, 13.24141, 12.05661, 19.75101, 
    14.34794,
  24.23281, 17.50524, 18.37535, 10.00453, 12.92319, 13.07283, 10.22563, 
    7.903003, 6.985473, 4.412628, 6.144569, 10.358, 14.00849, 11.37719, 
    14.97447,
  20.95485, 24.17999, 22.44075, 11.66926, 8.830606, 9.311252, 16.02546, 
    9.210466, 6.478034, 3.977426, 4.594916, 8.794719, 14.02353, 11.45328, 
    12.56751,
  21.18426, 20.98461, 24.36827, 10.13003, 9.071306, 6.336375, 7.501396, 
    16.09417, 8.870616, 5.534025, 3.455068, 5.809086, 11.5406, 11.23295, 
    9.376825,
  22.28147, 21.45984, 18.72859, 9.86979, 10.25688, 9.547702, 8.954923, 
    8.030606, 9.873892, 6.030709, 4.646739, 3.701274, 10.25914, 12.31763, 
    10.52681,
  23.69108, 25.22548, 16.37276, 10.5962, 10.04527, 9.059516, 9.092169, 
    7.391588, 6.600261, 5.06871, 3.252232, 2.692637, 9.81918, 12.52461, 
    11.3858,
  29.38786, 30.31938, 17.2303, 9.926304, 8.241608, 7.111389, 6.332052, 
    6.183444, 6.816782, 6.196041, 2.522084, 3.221595, 6.683255, 11.66881, 
    13.16361,
  30.90928, 22.9507, 13.73618, 10.10708, 8.513638, 7.491898, 4.591991, 
    3.204163, 4.091784, 3.576189, 2.249206, 1.76595, 7.914572, 12.22017, 
    16.71458,
  23.78051, 14.21439, 12.61454, 10.78679, 10.54564, 9.223216, 5.897304, 
    1.81244, 3.141726, 8.139982, 5.73622, 2.78832, 7.180003, 11.98434, 16.8078,
  12.59793, 16.16844, 16.95613, 10.37744, 9.640266, 12.65704, 9.316386, 
    7.648838, 6.018374, 9.917238, 11.74652, 11.52074, 21.05432, 12.74947, 
    12.03827,
  15.26968, 13.57114, 12.39008, 6.410087, 13.5642, 14.03222, 8.920505, 
    7.153737, 6.530887, 6.066822, 4.759065, 5.921249, 15.96259, 22.59629, 
    17.09501,
  17.16685, 16.93486, 17.228, 8.496033, 10.65351, 13.49787, 6.730052, 
    4.243608, 4.7362, 6.129112, 1.393678, 6.958644, 15.37743, 13.06019, 
    10.92783,
  18.59482, 24.24876, 22.19997, 9.311351, 6.807811, 7.972583, 9.773348, 
    4.527816, 3.60752, 4.649704, 2.253338, 6.364528, 13.20576, 10.67047, 
    6.796807,
  21.32894, 23.10221, 24.59882, 7.378776, 6.806607, 4.438812, 3.845809, 
    8.023428, 12.22868, 3.933055, 5.405038, 6.670119, 13.31397, 9.23491, 
    3.77979,
  24.11618, 25.44602, 18.16949, 6.039575, 6.07342, 4.34751, 2.055287, 
    3.773426, 7.676521, 6.883921, 7.023417, 6.204734, 10.28231, 7.74362, 
    3.757477,
  27.43529, 31.00689, 13.84078, 6.950288, 6.481699, 4.622325, 3.287326, 
    0.8166238, 3.86471, 6.400523, 4.453972, 6.201047, 9.759119, 8.785497, 
    3.788746,
  33.69465, 35.52215, 8.722841, 7.374172, 7.418831, 6.322882, 8.04504, 
    10.12555, 6.60309, 5.731563, 5.19681, 7.041472, 7.71761, 7.067934, 
    4.493373,
  37.76385, 26.87361, 5.932891, 8.455732, 7.83878, 5.963837, 6.089672, 
    5.945134, 4.643686, 2.931392, 4.923823, 7.317121, 6.949379, 5.574504, 
    5.618864,
  30.17533, 17.09498, 5.863369, 7.637957, 7.495755, 6.270376, 4.814365, 
    2.220619, 2.637145, 6.539342, 7.469469, 9.126403, 6.593007, 6.286835, 
    6.899699,
  8.567593, 8.54374, 11.60991, 8.809821, 6.463219, 4.694684, 3.118199, 
    4.554829, 4.938961, 13.16981, 20.76913, 17.68925, 11.21518, 6.963334, 
    18.65711,
  9.073732, 6.858302, 7.323031, 7.452482, 11.34568, 4.649961, 1.624207, 
    2.348645, 4.920642, 8.321856, 14.84152, 15.43055, 6.318294, 19.4824, 
    16.77904,
  17.23026, 12.32372, 11.82439, 9.421904, 5.940925, 12.0605, 0.9701228, 
    1.952663, 5.671446, 7.056015, 8.492096, 12.62367, 6.932196, 6.931204, 
    7.654322,
  21.03031, 17.18739, 15.47495, 9.122602, 2.462201, 1.334932, 9.274655, 
    6.079445, 6.518226, 8.740311, 10.29388, 12.41125, 10.70413, 7.750091, 
    5.19054,
  28.0431, 20.94212, 18.54416, 5.084989, 2.044286, 0.5183562, 2.76561, 
    16.14866, 11.95251, 12.49708, 10.71152, 10.09588, 4.802048, 4.573822, 
    3.3424,
  36.17215, 27.50083, 13.52403, 4.101087, 4.797705, 2.90161, 3.52921, 
    6.683604, 11.57076, 16.27847, 11.72391, 8.664233, 6.396163, 3.219908, 
    3.064304,
  43.53293, 35.93544, 12.05655, 5.407646, 9.240858, 12.76199, 8.693397, 
    7.724588, 12.74688, 11.68139, 9.741421, 7.975317, 6.907883, 4.416088, 
    4.241112,
  52.62262, 39.28727, 6.079081, 2.578453, 4.460957, 6.926306, 9.585596, 
    9.893123, 9.467938, 9.347692, 8.702761, 7.664449, 7.112482, 4.400968, 
    4.323438,
  53.3215, 25.04185, 1.701516, 2.553516, 4.256514, 5.598606, 5.230043, 
    5.810997, 7.383848, 8.333507, 8.098393, 7.48136, 7.368634, 6.481071, 
    4.161956,
  41.98786, 14.8224, 1.798173, 2.500151, 4.154589, 5.880167, 6.549618, 
    4.3556, 7.930732, 13.4674, 12.55373, 8.42775, 7.963671, 7.071848, 5.182355,
  8.43847, 7.665533, 19.88071, 9.763407, 10.03752, 14.71269, 10.40222, 
    5.305618, 3.518566, 3.665474, 10.76032, 13.36056, 13.35131, 11.49664, 
    22.79476,
  8.117264, 12.77052, 11.61935, 9.89972, 16.01373, 10.88831, 5.95015, 
    5.641889, 2.807858, 3.583671, 7.206583, 10.35769, 2.890402, 22.80975, 
    22.85273,
  25.01507, 24.54656, 19.42073, 10.72633, 12.14735, 14.23838, 1.60958, 
    1.069041, 2.324171, 6.153235, 7.152952, 8.237816, 2.862723, 5.197846, 
    12.03398,
  36.9651, 32.49099, 21.64933, 11.55575, 8.089209, 5.092065, 7.131207, 
    4.928314, 2.744088, 3.617429, 7.554918, 8.423433, 6.413783, 8.309758, 
    5.517326,
  49.56208, 34.19906, 20.4476, 7.032544, 5.251742, 2.332401, 1.401342, 
    16.55868, 14.35192, 5.109431, 8.35854, 7.839812, 6.082312, 3.829111, 
    1.024641,
  55.02913, 36.55446, 17.24504, 6.333887, 3.169244, 1.533851, 1.521407, 
    2.353135, 6.679894, 5.632481, 5.220919, 3.739607, 1.686807, 0.9042706, 
    0.1304474,
  56.03024, 40.75604, 15.68888, 8.435202, 7.486131, 6.761258, 5.075723, 
    5.890526, 3.451956, 2.805005, 7.477798, 6.840862, 1.95156, 0.324746, 
    0.1799474,
  56.14755, 38.93675, 7.823962, 5.055108, 6.762186, 6.302385, 5.413774, 
    4.075044, 3.129173, 4.802251, 3.689919, 2.447497, 0.5464733, 0.262604, 
    0.4411125,
  53.36199, 26.4929, 5.292786, 6.850948, 7.485744, 6.0667, 4.003783, 
    2.604974, 2.843986, 3.304838, 2.694281, 1.298547, 0.7589821, 0.3146514, 
    -0.4831513,
  42.62313, 22.25065, 6.053689, 6.281606, 9.234455, 8.198108, 5.054195, 
    3.270765, 3.753474, 4.240134, 3.295431, 2.387506, 1.245857, 1.191107, 
    0.4111509,
  0.27092, -6.511103, 12.57977, 3.142401, 7.620152, 11.35999, 9.535837, 
    8.258607, 7.638741, 17.2842, 20.19435, 20.10801, 11.55763, 22.70936, 
    27.23103,
  -6.559516, -3.844723, 0.9507602, 6.41038, 16.30573, 19.68503, 17.22047, 
    15.19635, 9.673306, 3.559365, 4.944147, 7.176188, 5.409062, 30.75132, 
    26.75849,
  3.789136, 9.56834, 11.5234, 10.89032, 17.99051, 23.17799, 16.17131, 
    13.9669, 9.551299, 9.324139, 7.544462, 5.833868, 9.058233, 10.26601, 
    14.2354,
  17.11131, 22.32162, 21.01638, 16.87139, 15.81982, 21.6705, 20.27513, 
    13.19993, 7.213296, 9.078578, 4.28314, 6.457832, 12.3142, 14.01498, 
    6.161561,
  38.06559, 30.03217, 26.80264, 16.93306, 15.14508, 15.64734, 14.16045, 
    21.88955, 11.85648, 8.061538, 12.20512, 13.64844, 13.25573, 9.246065, 
    2.079079,
  57.27669, 42.0735, 24.36302, 13.3057, 12.13509, 11.90827, 10.20605, 
    4.799886, 4.04516, 3.102105, 8.799254, 12.26587, 9.616983, 2.949789, 
    0.4056179,
  62.46306, 48.39338, 21.13881, 6.9421, 8.755397, 7.789361, 4.512269, 
    2.639557, 1.381663, 5.187835, 10.08951, 12.85209, 4.131297, 0.5724345, 
    0.2625961,
  50.91619, 38.01831, 6.057644, 6.655156, 5.888712, 6.328432, 6.99123, 
    4.113466, 11.07001, 8.820556, 12.46994, 5.824893, 0.6865296, 0.2165973, 
    -0.4525371,
  35.79502, 19.91251, 6.470825, 5.133379, 6.386581, 4.140378, 3.729975, 
    4.309793, 10.8088, 11.54966, 9.473263, 0.9354373, 0.3009413, 0.03633662, 
    -1.588324,
  25.22402, 13.55481, 5.664901, 7.885609, 6.487161, 4.715539, 7.400829, 
    6.608604, 6.513666, 6.266469, 1.130152, 0.3888564, 0.5788435, 0.2078911, 
    -1.290158,
  2.176733, -11.94272, -2.064931, -12.85594, -5.631726, -0.6703945, 3.36689, 
    7.764378, 7.405427, 21.56738, 32.53291, 21.48896, 18.76091, 17.52499, 
    19.58994,
  -11.76149, -19.53, -15.8799, -6.59666, -0.319781, 10.76974, 14.79476, 
    11.09446, 10.61356, 13.95864, 19.41393, 12.08405, 12.42151, 20.49573, 
    23.16228,
  -8.026366, -8.574936, -3.970496, -2.069314, 6.063198, 28.08202, 21.73236, 
    23.87115, 23.37977, 20.32949, 15.37259, 9.916632, 12.43165, 13.97595, 
    13.72614,
  -4.191896, -1.005988, 6.073674, 8.771507, 10.04778, 24.47206, 31.13068, 
    19.9914, 15.77109, 13.78772, 2.038789, 12.82538, 15.43475, 12.48019, 
    5.185595,
  4.15344, 5.329939, 12.05852, 10.34981, 15.48382, 19.07309, 21.47959, 
    25.93233, 14.82098, 4.654637, 4.924001, 15.09024, 9.293985, 3.350936, 
    0.4738207,
  14.22799, 16.50046, 11.43952, 10.15372, 16.98698, 14.14508, 11.67806, 
    10.38635, 6.599316, 3.963387, 13.6973, 9.349893, 2.988021, 0.3156215, 
    -0.06770415,
  29.50883, 32.5881, 13.77268, 12.02836, 15.33421, 15.8526, 11.82961, 
    11.98067, 7.254375, 9.445777, 12.0851, 3.813476, 0.4536389, -0.1702673, 
    -0.5165606,
  49.28839, 46.41393, 14.78599, 11.66315, 14.96009, 15.3588, 11.31803, 
    5.373975, 10.06064, 9.497027, 9.828887, 1.727405, 0.04080589, -0.4771863, 
    -1.148224,
  57.22205, 42.11052, 16.47914, 11.9228, 14.40946, 13.52595, 11.00788, 
    3.171258, 6.686672, 3.765622, 4.927526, 0.5580705, 0.04558711, 
    -0.3610503, -1.627018,
  46.07793, 34.28185, 19.59406, 13.2283, 13.46993, 13.88681, 12.32219, 
    3.953157, 3.2871, 8.18723, 2.476811, 0.1647802, 0.03880776, -0.1975633, 
    -1.219713,
  -4.147393, -16.43505, -8.412409, -22.57549, -20.28947, -20.83917, 
    -13.64951, -5.669203, -1.935385, 4.423413, 18.93797, 17.0504, 17.90084, 
    17.84129, 11.14418,
  -6.728379, -11.63503, -17.20167, -15.73976, -27.43173, -5.931147, 
    -3.980245, 0.3760605, 1.611362, 6.130231, 16.07107, 16.62704, 9.753775, 
    14.98515, 10.60901,
  -3.810333, -6.579579, -10.28077, -24.11864, -8.458549, 1.507776, 2.756049, 
    4.939929, 9.044388, 11.78728, 15.89195, 11.27222, 5.847999, 6.995395, 
    12.29089,
  -2.612548, -3.545375, -4.686307, -6.395066, -3.17565, 3.680776, 21.97365, 
    14.40767, 11.9733, 14.57472, 5.233856, 7.527257, 9.961079, 11.23799, 
    9.86907,
  -0.450873, -1.960051, -1.965988, -1.905984, 1.490436, 8.43507, 13.87844, 
    22.77344, 13.56278, 9.822192, 13.54012, 11.4395, 8.462229, 4.129997, 
    3.154752,
  1.40567, 1.87845, -1.675985, 0.6708002, 6.346532, 12.48333, 10.65854, 
    13.01593, 14.55803, 9.284698, 8.571388, 5.191796, 3.236097, 0.7122454, 
    0.168148,
  5.922332, 11.13159, 3.842421, 8.187355, 14.27789, 11.87077, 10.78079, 
    9.683919, 13.40759, 4.488038, 2.851832, 0.7511089, 0.009642864, 
    -0.04174066, 0.1857365,
  15.60959, 25.8763, 11.78597, 12.10393, 11.79495, 9.581464, 10.65352, 
    8.785681, 4.647746, 1.632388, 0.2516644, 0.02740831, -0.1512069, 
    -0.1471377, -0.1193526,
  33.96501, 34.75739, 16.51312, 14.10535, 14.2007, 12.41427, 7.451115, 
    5.228532, 3.13677, 0.7795125, 0.01119609, -0.08235431, -0.1590146, 
    -0.2159959, -0.6341516,
  39.84189, 40.30688, 28.80433, 13.10294, 11.09651, 8.883783, 3.653308, 
    4.147968, 3.442711, 1.072461, 0.5396932, 0.2718238, 0.03567366, 
    -0.1975774, -0.9022255,
  3.287091, -0.881871, 27.51654, -2.183754, -3.959461, -4.702731, -2.920518, 
    -3.616134, -8.624144, -9.706544, 7.091648, 8.903819, 9.983317, 3.681126, 
    0.577556,
  -13.81182, -4.384143, -5.04021, -2.563686, -3.14909, -3.952543, -1.672399, 
    -3.870835, -5.318893, -6.208678, 1.221637, 5.337231, 7.378316, 8.961232, 
    12.50447,
  -5.90799, -2.441995, -2.460402, -5.380542, -3.758126, -3.802741, -3.048175, 
    -2.185001, -3.525801, -4.839705, 1.316428, 6.466814, 7.080966, 3.94649, 
    12.57194,
  -1.243535, -2.196008, -2.334274, -2.454709, -3.257234, -3.248444, 
    -0.1002093, -1.241514, -2.487925, -0.2205251, 1.162407, 6.480269, 
    10.18091, 11.35482, 11.31944,
  3.40031, -1.290029, -1.912532, -2.69984, -3.134463, -4.013269, -3.584856, 
    3.769518, 6.325662, 3.296987, 3.480759, 5.219017, 9.113793, 12.00906, 
    11.28361,
  9.241507, 2.085858, -3.336339, -3.144201, -2.049419, -2.337677, -1.283809, 
    0.8323193, 4.39463, 4.805566, 6.125978, 7.371345, 11.6118, 11.06558, 
    7.069271,
  19.89216, 14.33745, 1.753858, 0.4094881, 1.201629, 1.897059, 3.730765, 
    4.741585, 4.223503, 6.698957, 10.0749, 8.997593, 6.110569, 2.920519, 
    3.21504,
  37.50039, 32.27234, 9.147055, 3.879104, 6.862293, 10.44909, 9.355798, 
    9.595165, 11.82243, 7.657557, 5.381583, 2.009965, 1.72818, 0.7947215, 
    0.8476912,
  50.80897, 37.15, 12.64318, 10.17547, 11.09916, 10.60829, 6.028713, 
    2.810813, 2.109066, 1.695677, -0.3852556, -0.08907128, 0.2018689, 
    0.1852647, 0.2244263,
  42.36637, 31.95621, 16.81948, 8.841791, 5.345426, 3.162478, -0.04323757, 
    -1.640614, -0.3480567, 0.3283378, 0.5309427, 0.7568015, 1.968741, 
    3.753271, 1.90594,
  1.618134, -1.517236, 12.90997, -2.480444, -4.166011, 2.074095, -5.584915, 
    -7.204406, -7.341968, -4.908231, 2.212737, 1.152159, -2.175275, 
    -7.254247, -7.004055,
  -3.4014, -1.047895, -0.5992566, -1.637504, -2.692073, -3.202607, -3.239207, 
    -5.743041, -6.805853, -5.357291, -0.6643443, -0.1504623, -3.279357, 
    -5.785015, -5.231091,
  -0.900268, 0.2019615, -0.9166107, -3.050785, -1.867096, 3.625702, 
    -2.231955, -3.990796, -5.200041, -4.115524, -0.2654918, -0.5696293, 
    -3.236187, -5.513299, -3.307013,
  1.461131, 0.8013729, -0.3709798, -1.38018, -2.712719, -2.423266, 1.744738, 
    -3.40626, -2.7525, -1.335583, 0.1915875, 0.8611104, -2.562902, -2.391075, 
    0.02924897,
  3.501828, 2.151463, 2.171224, 0.2129844, -1.212618, -3.228298, -3.460879, 
    1.146727, 4.053803, -1.177502, -0.3773208, -0.4197448, 1.194105, 
    0.7467458, 1.526878,
  5.512121, 4.387985, 1.682631, -0.4211909, -0.1271574, -1.196981, -2.35782, 
    -2.286447, -1.73646, -2.727347, -2.126389, 0.3950771, 2.099711, 2.584181, 
    3.126847,
  9.057566, 9.423124, 1.998252, -0.24812, -0.1746752, -0.2175261, -0.7720022, 
    -1.208753, -2.250012, -2.773932, -2.464443, 0.4393823, 2.233094, 
    2.445789, 3.892203,
  20.03704, 20.09097, 3.242338, 1.351097, 2.324919, 1.190645, 0.1569107, 
    -0.1916415, -0.1668031, -0.1539022, 0.5984135, 2.292394, 2.673942, 
    3.229424, 3.912124,
  31.84216, 18.44663, 2.727938, 3.663011, 5.152979, 5.169881, 5.079674, 
    3.87425, 4.15778, 4.960778, 3.778647, 4.002702, 3.438644, 2.961719, 
    2.943242,
  24.80987, 13.02645, 4.876582, 3.379474, 4.157284, 4.22691, 3.494306, 
    2.320263, 4.12432, 5.032837, 4.904339, 3.50572, 2.828811, 1.462783, 
    1.140365,
  2.568382, -2.596121, 8.570573, -5.118668, -4.721945, 0.6607445, -4.977848, 
    -4.663084, -8.345125, -1.705098, 0.9574661, -0.7383643, -6.538862, 
    -6.436327, -5.187077,
  -2.902987, -2.935104, -1.957354, -2.889476, -2.114466, -4.273256, 
    -4.901767, -3.316114, -4.807358, -1.078782, 0.07309422, -1.199392, 
    -5.147185, -7.051937, -5.69028,
  1.996934, 1.559474, -2.799943, -4.307089, -2.517916, 0.5357499, -3.586151, 
    -2.782742, -2.713039, -1.328678, -0.1220631, -0.997658, -3.10932, 
    -5.611347, -5.405341,
  14.25713, 9.599308, 1.71308, -1.954603, -3.804884, -3.965322, -0.4372431, 
    -1.119108, 0.1713382, -0.681069, 0.1047586, -0.8081093, -1.433064, 
    -4.52937, -3.968328,
  28.94054, 13.15469, 7.095647, -0.2457267, -0.6125674, -4.601802, -6.801643, 
    4.550839, 6.383392, -0.01305341, -0.1312148, -0.9366425, -1.22694, 
    -4.208678, -7.865159,
  38.1482, 18.91143, 4.587734, -0.448559, 0.5188038, -1.295475, -5.596124, 
    -3.946429, -1.569041, -0.9812122, -0.763137, -1.18053, -1.075576, 
    -4.057195, -5.118319,
  49.42927, 32.6926, 4.256866, -0.4377215, -0.1494677, -1.223195, -4.104236, 
    -2.516088, -1.823276, -2.613024, -1.697653, -2.070595, -1.338282, 
    -4.276621, -3.37804,
  62.1712, 44.80917, 5.470869, -0.187463, -0.2733428, -2.341252, -3.282762, 
    -2.42122, -1.503193, -2.516959, -1.532793, -1.220779, -1.51572, -3.41594, 
    -2.365286,
  65.83267, 42.83955, 6.482137, 1.375661, -0.3469162, -1.993552, -1.379088, 
    -1.732409, -2.350254, -1.473097, -0.09053844, 0.4488867, -0.6901276, 
    -1.429336, -0.3757206,
  53.48554, 45.80099, 18.06269, 4.552822, 1.247448, -0.3894298, -1.437979, 
    -2.167591, -0.7926521, 1.0949, 1.706068, 1.662898, 0.4684212, -0.3854696, 
    0.1347782,
  4.370932, -0.2933652, 15.5562, -1.687296, 1.555266, 8.639315, -0.620842, 
    -0.2518605, 0.3433947, -0.489108, 0.741977, -0.3047384, -2.731645, 
    -3.476835, -5.390506,
  0.5272417, 0.210528, 1.153733, -1.019843, 1.896788, 0.6059975, -0.3812947, 
    0.7386543, -0.1611501, -0.1405117, -0.1138449, -0.9939874, -3.176179, 
    -4.712854, -5.935759,
  9.996258, 11.28969, 3.945705, -2.339272, 0.4261184, 10.60312, 0.3518514, 
    -0.2829768, -0.6964426, -0.2461863, -0.02652877, -0.7551466, -3.123709, 
    -5.315659, -10.53403,
  16.17906, 10.87252, 2.680624, -1.08809, -2.214868, -0.516091, 7.380663, 
    -0.2553811, -0.7116102, -0.07407353, -0.2741981, -0.9006311, -3.036454, 
    -5.203269, -5.640512,
  20.93183, 7.236433, 2.780237, -2.737993, -1.865126, -2.094421, -1.671003, 
    5.687954, 0.665873, -0.1076209, -0.1618982, -0.9482761, -3.373237, 
    -5.821029, -10.65476,
  21.53263, 8.054493, -1.399553, -3.865861, -1.40637, -0.1199916, -1.198132, 
    -1.902223, -1.476877, -0.5008059, -0.2910959, -1.299072, -3.834513, 
    -5.113991, -4.951426,
  25.12779, 11.91291, -1.499601, -1.647411, -0.110359, 0.570036, -0.2249326, 
    -1.199457, -1.773692, -0.9520845, -0.6332188, -2.059633, -3.713712, 
    -4.51399, -3.364656,
  28.01296, 17.51425, 0.5690218, 0.3050317, 0.7706268, 0.8185801, -0.4677839, 
    -2.468702, -1.879398, -0.3395211, -0.6064557, -1.926551, -3.214951, 
    -3.538361, -2.385666,
  31.30964, 12.94045, -0.4800107, 0.9254051, 1.604352, 0.3346806, 0.1028297, 
    -1.364894, -0.9897463, -0.2549985, -0.5015321, -1.315123, -2.610837, 
    -2.467548, -1.351764,
  21.75926, 7.274612, 0.5833266, 0.6735986, 0.3994799, -0.3661033, -1.151212, 
    -1.617765, -0.7001847, 0.6856741, 1.029491, -0.5390769, -2.586189, 
    -2.567561, -1.143576,
  4.961019, -3.741922, 12.15192, -5.577336, -0.06927869, 10.2788, -2.494992, 
    -0.8770299, 3.133606, 6.66333, 14.64061, 9.800074, 2.721885, -0.9378346, 
    -5.696407,
  -1.388751, -1.752248, -2.675271, -3.609149, 0.2859588, 4.498477, -2.857816, 
    -0.8653633, 1.52646, 2.614123, 7.56446, 3.470303, 0.9466785, 2.277756, 
    -0.5204603,
  0.06245596, 0.8188241, -0.1726032, -1.99117, -0.1175397, 7.581586, 
    0.3096229, 0.3469546, 0.6365851, -0.008953806, 0.03940203, 0.7013723, 
    0.6766622, -0.2329917, -1.014353,
  6.785868, 5.597761, 0.6490819, -2.670347, -4.531491, -0.986557, 10.99856, 
    0.7463551, -0.4358957, -0.2834357, -0.2190783, -0.2648683, -0.446121, 
    -0.6802471, -1.434088,
  12.90467, 0.271493, -2.719458, -7.430377, -5.629338, -4.899491, -3.081442, 
    18.11914, 11.70194, 0.8121837, -0.1773949, -0.3862971, -0.5559577, 
    -0.9414378, -3.094242,
  6.098626, -2.163714, -7.101274, -8.2833, -3.734939, -2.398386, -2.59791, 
    -0.07981317, 2.189752, 0.3245837, 0.07819828, 0.5158659, 0.7062638, 
    -0.627423, -2.547356,
  5.265429, 2.555361, -2.890774, -3.141018, -0.7165102, 0.0165503, 
    -0.4281736, -0.4056712, 0.5321437, 1.515287, 1.861769, 1.533441, 
    0.03066877, -1.371265, -2.219371,
  11.04347, 16.88262, 0.08062627, -0.4689171, 0.4057806, 0.288435, 
    -0.02625695, 0.5484281, 1.161216, 1.438485, 1.327363, -0.1327724, 
    -0.8722254, -1.675361, -1.784606,
  19.71962, 8.440375, -0.1637067, 0.3618952, 0.6211592, 0.6524211, 0.9764083, 
    1.593054, 1.256098, 0.8284692, -0.08311597, -0.5290591, -0.7124225, 
    -0.1771235, 1.849451,
  11.64792, 5.99645, 0.7120039, 1.153446, 1.169413, 1.113409, 0.6578507, 
    0.970546, 0.3637429, -0.01730341, -0.4277106, 0.6841739, -0.2640811, 
    0.8092532, 3.407258,
  -6.510394, -15.31701, 1.961054, -13.0244, -6.378893, 1.214491, -7.847484, 
    -4.901417, -3.003342, 5.241614, 6.315066, 9.135105, -1.720091, 18.85284, 
    21.34775,
  -18.02115, -15.48446, -13.34642, -11.04692, -7.602328, 0.4856575, 
    -4.489831, -2.095825, -2.846231, 0.1213824, 0.3022175, -0.2988414, 
    1.849848, 12.51901, 13.87056,
  -7.46283, -8.11691, -6.669977, -7.854461, -10.67729, -6.875374, -2.499522, 
    -1.220233, -1.596684, -1.3816, 0.506507, 0.236023, 5.134251, 7.003892, 
    6.946075,
  4.480688, 0.9771051, -1.540044, -3.043377, -5.79477, -3.46904, 2.251105, 
    -0.06112325, -0.3379204, 0.08192348, 0.2369982, 0.2001999, 4.135747, 
    5.913376, 0.8909553,
  8.170977, 1.957807, -0.1829218, -3.552298, -3.224415, -3.591611, -2.301879, 
    11.20892, 9.153218, 0.4872573, 0.1716891, 0.1476424, 2.041971, 4.075759, 
    -0.9368622,
  3.883029, -0.6500434, -2.662431, -4.463251, -3.053229, -2.155818, 
    -3.162465, -2.057711, 0.8227919, 0.2456718, 0.1047777, 2.66573, 4.755736, 
    3.40956, 0.3994907,
  3.926039, 0.04416157, -4.160913, -4.806431, -2.670872, -0.3599988, 
    -0.4415034, -1.028124, -1.052249, -0.6456597, 0.7216188, 1.982564, 
    3.586776, 2.472512, 3.344979,
  5.359735, 3.328457, -4.001319, -3.48671, -1.295168, 0.1255034, 0.508114, 
    -0.1113415, -0.6757913, -0.1140023, 1.011501, 2.836309, 2.500785, 
    2.036186, 5.503997,
  8.942272, 0.482573, -4.118088, -2.009914, -0.9761952, -0.175398, 0.569286, 
    0.8816673, 0.4711385, 0.4948948, 2.528375, 3.749323, 1.597677, 1.274678, 
    9.258679,
  6.728158, 1.394776, -2.484859, -0.6612574, -0.1254686, 0.3334582, 
    0.4261035, 0.1094898, 1.148506, 1.611909, 3.614851, 4.7851, 0.6104379, 
    2.59492, 14.57372,
  0.7196451, -7.975822, 1.788806, -13.52189, -12.06292, -1.540429, -22.77229, 
    -20.27337, -24.04303, 16.21311, 27.46848, 35.91137, 18.73455, 26.42367, 
    28.38704,
  -2.808883, -6.730259, -9.289168, -16.8807, -3.391762, 3.390886, -15.21173, 
    -16.48242, -19.36222, -11.22038, 33.80491, 9.679727, 9.573145, 12.47537, 
    4.370908,
  2.39621, -2.761476, -7.002375, -15.27559, -18.6696, -8.115306, -9.732765, 
    -6.531509, -6.99083, 0.006729853, 4.095418, 6.661496, 8.220447, 3.899725, 
    1.242082,
  11.97808, 1.591869, -5.064059, -9.731519, -13.97282, -11.43167, -3.447256, 
    -2.808286, -0.09184116, 2.112268, 3.035111, 5.410489, 7.55987, 4.760764, 
    1.916755,
  20.35929, 1.680554, -2.522014, -9.650543, -10.15965, -10.2313, -9.224944, 
    1.483384, 8.324732, 1.424763, 2.403156, 4.311026, 7.475469, 4.958546, 
    3.091241,
  18.63408, 6.053243, -1.194522, -7.935789, -7.643531, -6.912182, -6.297842, 
    -3.692837, 1.55383, 1.424369, 5.593338, 7.16558, 7.856499, 6.732728, 
    4.248428,
  17.77586, 11.9261, -1.252705, -5.975002, -7.085229, -6.109332, -5.124907, 
    -1.572039, 0.4850074, 2.50162, 4.578179, 8.634604, 10.86388, 14.15976, 
    13.3607,
  9.408153, 11.9932, -1.577832, -3.974321, -4.550255, -4.256197, -4.034045, 
    -0.6024281, 0.4266132, 3.204192, 3.454881, 6.07896, 11.80489, 13.37578, 
    15.84409,
  5.484, 3.335207, -1.387841, -1.830346, -2.467685, -2.953318, -2.483973, 
    0.3707921, 2.12701, 3.073712, 3.285091, 10.10884, 12.1788, 13.36993, 
    15.38445,
  3.715487, 1.451608, -1.004882, -1.105026, -1.464176, -1.623545, -2.123924, 
    -0.5715244, 1.963288, 2.942073, 4.585232, 11.75314, 11.76991, 14.79094, 
    24.38748,
  8.913525, -4.832813, 7.379843, -7.861134, -6.450587, 5.39198, -8.418597, 
    -17.21495, -20.97104, -9.750216, 16.8848, 26.63933, 22.99306, 29.21691, 
    36.22585,
  4.433646, -3.537243, -4.559417, -8.405585, 1.188743, 3.248339, -8.11386, 
    -9.711308, -13.01089, -8.97878, 30.93805, 8.774287, 7.2017, 5.060055, 
    -2.822627,
  8.268579, 4.825289, -2.927293, -6.185205, -2.951226, -0.09429117, 
    -2.603833, -1.289596, -0.8430613, 1.75815, 8.418125, 6.46937, 3.816463, 
    1.27514, -0.5825682,
  10.62424, 9.361568, -0.564144, -1.647886, -4.880064, 0.5290795, 16.51892, 
    10.81944, 8.585541, 8.155952, 7.854924, 6.322414, 6.034249, 3.29258, 
    4.157983,
  9.342201, 5.206222, 0.7219942, -2.889077, -3.503483, -2.12873, 1.307153, 
    17.98591, 18.0468, 10.66394, 8.708093, 11.50746, 13.58808, 9.910909, 
    10.89845,
  7.802233, 4.798426, 0.3174669, -3.437843, -3.530456, -1.083366, 0.131695, 
    2.492949, 11.90897, 11.87201, 12.27939, 15.73624, 17.07198, 19.5732, 
    16.31425,
  9.932139, 7.244789, -0.1146751, -3.85762, -5.230115, -1.940581, 1.429135, 
    5.997375, 7.809036, 8.115857, 12.20801, 16.91963, 20.32936, 14.99215, 
    18.37665,
  13.48166, 8.334335, 0.6415507, -3.28511, -5.784317, -2.139428, 3.663082, 
    8.294794, 11.62337, 14.74791, 13.92714, 20.23915, 19.16507, 18.83818, 
    17.89914,
  7.398991, 2.388106, -0.9869002, -1.224225, -3.458616, -1.617141, 5.654819, 
    9.226244, 15.89609, 15.6636, 18.69997, 19.45505, 17.56504, 16.98893, 
    17.09458,
  1.955861, 1.421483, -0.5255864, -0.9233766, -2.11635, -0.6794155, 6.324466, 
    9.360941, 12.85096, 22.66145, 21.26464, 17.99607, 18.66988, 18.3579, 
    22.52423,
  1.823607, -7.424862, -0.5306619, -6.066421, -0.5010303, 6.832705, 
    -4.547318, -7.856984, -9.682257, 28.35961, 46.64796, 28.80054, 33.81112, 
    32.31298, 37.7214,
  -10.52345, -7.700259, -6.541845, -5.997666, 9.180605, 8.197957, -3.380248, 
    -4.969745, -6.704763, 2.871866, 34.66692, 7.026197, 4.22334, 1.490578, 
    24.86356,
  -8.573708, -3.408177, -4.62172, -6.580183, 1.438239, 2.733453, 2.345028, 
    0.1894218, -0.7344291, -0.6137437, 4.401941, 1.693473, 0.9741892, 
    3.318598, 7.211857,
  -2.789741, -0.1277146, -2.459475, -3.248973, -8.749462, -0.4514731, 
    12.1228, 3.943524, 2.371354, 1.178627, 1.719349, 5.246585, 6.156436, 
    8.758434, 11.66353,
  3.006144, -1.29037, -1.455726, -5.262969, -5.157847, -4.398675, 1.343606, 
    18.52932, 15.69339, 3.422828, 6.073114, 13.5303, 17.62062, 14.75958, 
    12.11916,
  10.74896, 1.516598, -2.619925, -5.864933, -3.948495, -1.815875, -0.4663392, 
    2.949514, 6.68213, 8.296587, 14.04507, 17.93691, 16.65638, 14.72441, 
    10.93813,
  18.88148, 11.34503, -2.939336, -6.129443, -5.736492, -2.664325, 1.07237, 
    6.437846, 8.173758, 13.42679, 16.53749, 16.63471, 12.99604, 10.62657, 
    10.67417,
  28.83554, 17.98674, 0.3963219, -4.058008, -4.695744, -1.562267, 6.762086, 
    8.354485, 12.48024, 19.83974, 21.76213, 16.23775, 13.99885, 11.14631, 
    8.991014,
  28.6098, 10.82287, -0.6754897, -1.58873, -2.538727, 0.9826137, 8.302863, 
    11.47318, 20.01523, 21.6957, 17.86072, 16.72904, 13.05962, 10.00964, 
    5.610795,
  10.91281, 7.539503, 0.3002036, 0.4381634, 0.5533805, 2.938266, 9.908482, 
    13.93829, 18.36466, 25.2371, 22.59456, 16.34921, 12.99226, 8.942054, 
    6.165766,
  0.7848945, -3.969067, 14.22741, -3.792446, -2.123493, 3.669206, -2.904385, 
    -2.620071, -2.836656, 14.80673, 22.91328, 20.06245, 25.65721, 25.55735, 
    38.41447,
  -0.06865742, 0.9734083, 2.214914, -1.154622, 15.30181, 15.40137, -2.966721, 
    -3.103048, -3.871713, -2.18565, 12.75625, 1.263929, 5.124371, 8.320986, 
    21.35743,
  7.763336, 7.728192, 5.26395, 1.170235, 9.881612, 4.311645, 2.328798, 
    -2.572324, -4.050494, -5.585428, -4.353901, -3.165191, 1.064748, 
    8.503724, 10.89388,
  12.23656, 9.172229, 5.54982, 4.196282, -1.213095, 3.422523, 5.798754, 
    1.745097, -2.295562, -2.691494, -4.339436, -0.7063295, 7.112795, 
    10.22341, 10.5215,
  13.4437, 8.952654, 8.825218, 2.953887, -0.9274853, -0.2582878, -0.6440387, 
    10.34611, 7.735928, -0.3244685, -0.3217371, 3.201384, 10.45978, 12.31378, 
    9.99943,
  21.8742, 15.22506, 7.161778, 0.4756709, -1.029266, 1.740473, -0.7809207, 
    -0.8335601, 3.344539, 1.035892, 2.862604, 8.211963, 12.15566, 13.72397, 
    6.381405,
  20.87677, 15.34555, 0.145182, -4.401241, -4.091627, -2.695747, 2.026048, 
    1.629185, 0.2587465, -0.09453507, 4.581776, 10.61447, 13.73082, 13.51032, 
    8.799782,
  26.34293, 19.61622, 0.2769983, -4.807573, -2.098816, -0.7529991, 3.270832, 
    1.324707, 1.422388, 4.459772, 11.1174, 14.27191, 17.6881, 14.06471, 
    7.875827,
  31.15336, 17.28388, -1.128138, 2.786368, 1.728991, 1.89824, 3.587909, 
    4.004873, 6.889225, 10.89959, 15.30687, 16.91752, 18.88024, 11.35239, 
    7.71986,
  17.32312, 10.85014, 5.331714, 4.0477, 3.220314, 2.584853, 2.285998, 
    6.068783, 12.29908, 21.19501, 23.4604, 21.53663, 10.65138, 4.472248, 
    3.273166,
  -8.33881, -26.73639, -7.368721, -17.25685, -9.783465, -3.308181, -6.853177, 
    -3.936876, -4.026717, 0.3659101, 3.289272, 0.3261576, 7.543603, 14.4277, 
    25.26306,
  -6.806745, -9.613958, -6.615369, -7.330701, 1.619755, 5.556858, 0.1866812, 
    -1.575225, -2.280411, -0.2513773, 8.268064, -2.512388, -5.256567, 
    2.164334, 20.80977,
  8.64445, 9.656073, 6.954939, 0.9523409, 14.06634, 10.94572, 7.997824, 
    4.587051, 0.2383371, 0.5554094, 5.314187, -0.6472102, -5.103109, 
    -4.246277, 7.286836,
  28.18335, 28.10563, 18.50261, 14.97068, 5.126372, 14.95205, 11.76986, 
    7.916452, 1.2917, 3.681133, 1.647254, 0.1138393, -2.321034, -3.10411, 
    -1.496851,
  30.29918, 19.09172, 13.66768, 7.418185, 2.963469, 4.164293, 9.972059, 
    19.05574, 17.18122, 11.05422, 5.389474, 2.885062, -0.3420689, 
    -0.04159615, 1.632408,
  16.99599, 10.32342, 4.663301, 1.310465, -0.2762043, 1.697331, 3.338262, 
    5.826775, 10.81302, 9.584039, 9.209884, 4.706831, 1.599326, 2.045308, 
    4.340075,
  14.72655, 10.35101, 0.7494168, -1.298427, -1.334536, -1.574034, 3.192336, 
    3.72525, 2.378798, 2.898558, 4.039817, 3.588994, 1.456439, 3.973973, 
    6.022289,
  15.30067, 17.55772, 0.7894796, -2.622365, -1.313092, -1.064893, 2.962818, 
    1.638352, 1.141721, 3.043295, 4.053462, 2.112511, 1.761644, 4.880716, 
    8.602533,
  29.34163, 8.492267, -1.835323, -0.6670473, 2.76162, -0.1499191, 2.660597, 
    3.105668, 3.722282, 4.642664, 4.159206, 2.222528, 3.404658, 7.478527, 
    11.55794,
  22.12076, 6.258693, -0.8654261, 3.618958, 4.111524, 1.738101, 2.601567, 
    3.140573, 3.77144, 5.254741, 3.464926, 2.9617, 7.056148, 9.90075, 14.37307,
  9.238822, -1.977131, 33.46371, -12.92393, -0.8452339, 15.64939, -13.9908, 
    -14.97009, -11.31151, 11.91844, 11.72806, -0.6240765, -3.833571, 
    -8.83894, -7.04667,
  6.539925, 4.817078, 5.291521, -0.2668762, 20.3019, 18.09372, -7.642107, 
    -9.77089, -10.78351, -7.152123, 15.13324, -4.373903, -9.255125, 
    -4.006677, -4.840841,
  13.89649, 15.36682, 11.90282, 3.50977, 12.00502, 3.631448, 1.885945, 
    -2.660469, -4.068412, -5.997673, 2.140496, -1.349802, -7.028554, 
    -6.012941, -5.322127,
  31.19027, 36.21841, 26.85789, 21.69637, 3.735967, 11.69305, 15.8055, 
    5.653892, 2.699015, 2.73543, 1.604863, 1.522021, -1.748002, -4.065564, 
    -8.17404,
  30.88286, 26.63219, 32.46252, 20.15965, 7.247006, 4.640059, 8.490844, 
    23.69977, 23.04271, 11.44888, 7.720527, 7.825537, 3.31733, -2.00496, 
    -4.81187,
  24.72655, 24.26026, 17.61006, 8.327372, 3.749499, 5.131712, 4.794313, 
    5.097372, 14.43544, 10.17342, 12.13079, 10.23781, 5.62372, -0.3780084, 
    -2.105638,
  25.06071, 25.52196, 6.527069, 2.516051, 2.239561, 1.206952, 3.804794, 
    5.973567, 5.024543, 7.014791, 8.177003, 7.507563, 3.713946, 0.5982996, 
    -1.412515,
  24.12355, 19.31301, 3.476383, 0.9271459, 1.979526, 0.5643875, 3.189697, 
    5.093317, 3.416073, 6.683426, 7.160124, 4.991545, 1.558648, -0.1091269, 
    -0.792808,
  24.96962, 8.480358, 1.095487, 1.212712, 2.570132, 1.37865, 1.843094, 
    1.792259, 1.929499, 2.708786, 3.345494, 3.150211, 1.799049, 2.617472, 
    5.518963,
  17.32657, 7.041561, 2.161425, 2.891604, 2.389544, 2.976708, 4.420714, 
    6.605948, 4.795909, 4.523962, 4.444817, 3.351276, 3.433466, 5.395309, 
    12.67421,
  8.176683, 4.39013, 24.44608, 3.649145, 9.109997, 23.75352, 5.936916, 
    5.431261, 6.643263, 47.60961, 64.00889, 43.54144, 41.92301, 54.65121, 
    68.27501,
  9.239959, 8.74648, 10.11596, 5.701909, 26.27587, 38.90144, 7.449889, 
    6.725286, 4.137291, 13.5461, 43.39012, 24.61184, 8.170327, 25.87747, 
    51.59131,
  11.08691, 14.3196, 13.2223, 9.062407, 24.04435, 24.67077, 19.60567, 
    5.634683, 4.068923, 3.133593, 7.022612, 4.897765, -1.590685, 0.7008803, 
    10.77965,
  7.385082, 11.06819, 8.646822, 15.90706, 7.163321, 25.90882, 27.5735, 
    9.732686, 10.01906, 7.607781, 3.009487, -2.095328, -2.109119, -1.44371, 
    -0.810066,
  5.352914, 3.905856, 10.14491, 10.99335, 5.014756, 5.325069, 14.37302, 
    20.48741, 20.69181, 25.94593, 0.9143617, -2.511562, -1.809568, -1.842431, 
    -4.16129,
  5.724074, 2.362977, 6.90307, 3.847674, 0.937763, 2.018652, 3.757603, 
    10.0189, 19.77493, 8.69044, 0.09365802, -2.098971, -2.250294, -4.620791, 
    -7.34976,
  8.251154, 5.822141, 1.678624, 0.6925921, 0.8616877, 0.663379, 1.742486, 
    6.980169, 7.22506, 1.045989, -1.044374, -0.9718026, -0.8049871, 
    -1.957145, -2.314036,
  8.969744, 9.617889, 2.958584, 0.3556725, 0.4008829, 0.4375352, 0.8221993, 
    3.376147, 2.672026, 2.176263, 0.3598864, -0.03429336, 1.076823, 1.413269, 
    2.143791,
  13.96972, 7.198673, 0.9808953, 0.7446783, 0.8219213, 0.05076753, 1.132325, 
    2.390825, 2.103014, 1.843581, 0.8458765, 0.7351642, 2.33972, 4.013792, 
    6.778584,
  13.45646, 7.547286, 1.443544, 1.865457, 2.58852, 2.262874, 2.055548, 
    1.926793, 4.46871, 2.576873, 1.833029, 1.732889, 2.93581, 6.044458, 
    9.873237,
  4.506999, -10.22814, 8.067893, -15.98898, -4.356371, 6.498027, -20.7647, 
    -16.6489, -11.91706, 14.51108, 39.19768, 28.58261, 30.40942, 36.1525, 
    40.45944,
  3.950778, -1.754772, -6.828906, -9.795281, 2.997719, 8.147234, -4.437273, 
    -7.836836, -7.2558, -2.590218, 31.45256, 15.48053, 6.947873, 25.48116, 
    31.66662,
  27.09618, 16.16483, 8.138242, -1.299516, 1.109827, 5.832611, 1.856849, 
    -0.6438173, -0.4476835, -1.426932, 3.673469, 1.357575, 1.879599, 5.35536, 
    16.11265,
  48.70646, 41.21472, 21.07233, 13.37549, 0.5159354, 8.865669, 14.33796, 
    4.187973, 3.463931, 2.285736, 1.179491, 0.503481, 4.201794, 2.254535, 
    4.432119,
  46.65388, 38.27852, 33.64263, 15.64253, 1.279682, 0.1819286, 10.45427, 
    21.21609, 16.51129, 12.40848, 0.436837, 1.518301, 4.691846, 0.6819993, 
    -0.6461402,
  42.67638, 35.75754, 24.11729, 9.936125, 3.324455, 2.435499, 2.591563, 
    6.678504, 13.65107, 2.64626, 1.50353, 1.289132, 3.95758, -0.2118194, 
    -0.0372581,
  39.21024, 35.15302, 13.06336, 5.142559, 4.495366, 3.246495, 2.497615, 
    3.756133, 1.955531, 0.7134006, 1.263049, 0.3553453, 0.8198212, 0.5087093, 
    2.1718,
  35.23779, 29.88943, 9.119534, 4.796242, 5.318569, 6.209036, 5.376902, 
    5.53428, 1.971709, 1.797473, 0.1412912, 1.130476, 0.6166385, 0.9243749, 
    2.118587,
  27.49733, 12.24176, 2.699387, 1.237874, 2.217479, 3.428419, 5.67979, 
    4.684037, 1.818129, 1.362694, 2.765263, 2.894587, 1.455687, 1.318004, 
    2.465881,
  14.18764, 6.343552, 1.54003, 0.8972808, 2.361634, 2.854987, 5.049872, 
    4.298646, 1.129951, 3.944123, 2.896188, 2.275786, 3.717991, 2.561419, 
    7.692593,
  8.783351, 1.126383, 23.01756, -1.937707, 1.775887, 19.35512, -16.20685, 
    -27.37823, -25.9231, 34.60514, 34.45422, 8.397607, 36.4497, 19.314, 
    23.42551,
  7.771636, 1.04784, -0.2747752, -2.083687, 19.26577, 23.31323, -5.776835, 
    -14.02988, -19.94863, -12.80137, 12.3482, -16.20202, -13.56606, 12.47261, 
    19.43627,
  20.65558, 13.81419, 2.3646, -1.813711, 8.062943, -7.389494, 4.030321, 
    -3.779794, -11.49664, -23.53679, -22.56152, -18.06847, -16.26453, 
    -4.884269, 9.375942,
  40.72685, 28.93652, 9.179901, 2.350774, -3.917563, 4.352758, -4.956683, 
    -2.558573, -2.972108, -7.650071, -11.63551, -9.892001, -6.422813, 
    -2.534236, 2.864623,
  47.7527, 35.34045, 20.7017, 4.370521, -1.762146, -6.23547, -8.841539, 
    -10.87386, -4.834126, 4.667333, -5.208932, -5.794597, -1.624799, 
    -2.075354, -2.877484,
  53.49956, 37.75536, 26.16868, 4.352927, -2.246194, -2.640651, -7.497859, 
    -11.30659, -1.633203, -4.593372, -2.170239, 0.3766364, 1.522682, 
    0.5809437, 1.541065,
  53.97865, 43.54718, 20.50882, 4.484638, 0.3834527, -1.512302, -2.594483, 
    -4.540064, -5.703581, -3.473988, -1.233123, 1.456524, 2.438689, 2.892722, 
    4.568296,
  46.09804, 41.54121, 21.10943, 6.824957, 4.014452, 0.9298733, -1.665851, 
    -1.330899, -0.3133865, 1.545753, 2.803083, 4.778214, 2.929793, 4.237814, 
    4.728462,
  28.83927, 24.12976, 14.74424, 7.134625, 4.56677, 0.9901208, 1.099582, 
    2.276677, 3.520186, 5.597912, 6.815044, 6.678042, 5.453163, 4.580159, 
    3.750945,
  10.30487, 10.90309, 12.81136, 9.480818, 10.27766, 6.7303, 4.113461, 
    4.08599, 6.768725, 10.22543, 10.97741, 9.166041, 7.741628, 5.715598, 
    5.558072,
  10.52706, 2.78742, 18.97212, -4.223643, -5.380854, 17.00726, -12.74882, 
    -19.61555, -18.60858, 43.26891, 42.82094, 21.05235, 32.08455, 22.11112, 
    28.02687,
  12.80201, 9.069369, 8.587251, -2.064568, 11.56094, 29.68324, -3.115581, 
    -6.792934, -8.531089, -2.33428, 23.08773, -17.63704, -18.41823, 19.38135, 
    19.3291,
  25.15624, 24.52324, 15.54976, 6.429242, 18.95042, -0.7031863, 2.099121, 
    -2.067811, -4.792751, -7.86342, -10.24642, -12.43825, -20.9724, 
    -21.75792, 4.59729,
  35.33384, 33.39656, 21.61065, 15.80776, 7.909419, 12.84857, 0.4394726, 
    -0.7197385, -3.179365, -2.126742, -5.53533, -9.155457, -9.762171, 
    -14.34985, -8.394619,
  29.31226, 29.4223, 26.77158, 12.55313, 5.077404, 4.618428, 5.009659, 
    1.025894, -2.15787, 7.827966, -1.437406, -5.000208, -7.457767, -12.14753, 
    -19.65412,
  23.01346, 22.85874, 22.4522, 7.543766, 4.824805, 3.819819, 3.130197, 
    2.440917, 6.160995, -1.053297, 1.450272, -3.108169, -4.296419, -7.330915, 
    -12.1799,
  23.33409, 20.96055, 14.28001, 3.243609, 5.476511, 4.435947, 2.740995, 
    2.799923, -0.03112328, -2.535302, -3.601331, -3.414121, -3.824174, 
    -4.765811, -7.510549,
  28.73964, 18.50184, 14.25554, 4.093978, 5.992056, 4.921709, 1.897567, 
    2.736612, 0.5687385, -1.080007, -2.278389, -3.424779, -4.216028, 
    -4.162303, -4.982609,
  21.01072, 12.20263, 11.06686, 3.953772, 4.415639, 3.538579, 5.104635, 
    3.650499, 1.090185, -0.4151069, -1.687569, -2.836921, -3.354527, 
    -3.699563, -3.996943,
  9.195654, 8.592856, 9.753042, 6.241288, 7.470234, 6.23734, 6.351833, 
    4.16122, 2.035437, 0.8293924, -0.5853801, -1.547162, -2.484562, -3.03952, 
    -1.405348,
  9.283569, -3.410382, 5.615557, -23.464, -21.67934, -3.122368, -34.43726, 
    -35.27478, -41.5448, 43.06903, 49.29275, 24.70841, 45.43052, 33.4975, 
    56.06009,
  17.22889, 5.883337, -3.667138, -20.82168, 8.323461, 10.87991, -19.19934, 
    -22.59401, -24.50782, -7.405065, 21.79525, -10.71526, -10.63696, 
    26.31244, 27.89314,
  30.59347, 31.56714, 16.15322, -4.68488, -0.6044971, -13.58458, -4.158158, 
    -14.16053, -23.97878, -21.81699, -15.63609, -10.55757, -12.30042, 
    -8.815045, 8.108763,
  45.94678, 42.88017, 29.51938, 18.23229, -3.893125, 2.882535, -7.892148, 
    -6.703981, -11.10495, -9.52961, -11.68421, -6.687077, -4.465934, 
    -3.365241, -6.540054,
  37.05422, 34.66357, 33.69257, 23.39899, 5.250989, -3.590583, -3.652255, 
    -11.59809, -0.1682653, 5.976543, -4.405666, -4.979277, -3.15614, 
    -2.588243, -10.09259,
  25.54669, 20.98624, 25.94023, 17.49182, 9.50454, 3.424869, 0.6869732, 
    1.029232, 6.89183, 3.416284, 8.653063, -1.583371, -2.19488, -1.622304, 
    -3.698783,
  21.57989, 8.574471, 8.679533, 10.20708, 13.5749, 11.7569, 6.29473, 
    5.949222, 4.871881, 2.677306, 2.553352, 0.02258587, -0.6158526, 
    -1.000627, -1.511764,
  22.92344, 5.135534, 2.257733, 7.150038, 10.27864, 10.80469, 7.731019, 
    8.088209, 7.866637, 5.67842, 4.86866, 1.736959, 0.3791873, -0.0527039, 
    -0.6186883,
  23.04024, 7.549012, 1.496955, 2.093375, 7.095438, 9.22483, 9.348203, 
    11.99685, 11.93049, 9.053237, 5.710979, 2.184231, 2.226788, 1.432367, 
    -0.1648342,
  8.95603, 1.92344, 0.2441549, 3.142718, 6.988429, 8.424383, 9.81767, 
    11.55296, 12.96915, 12.5936, 10.40464, 7.082684, 5.002551, 2.743082, 
    2.725956,
  2.410712, -1.942522, 34.81259, -1.026032, 4.479422, 8.826697, -25.92081, 
    -45.13406, -45.81044, 56.50392, 65.20866, 26.17739, 58.23304, 49.07625, 
    88.76222,
  1.012921, -3.085735, -2.081845, -1.831633, 49.20998, 14.17959, -14.89217, 
    -33.58331, -44.38448, -15.13541, 31.40061, -21.07058, -32.1925, 46.53978, 
    66.72239,
  17.87432, 5.234182, -1.080926, -3.288618, 17.43454, -12.34384, -3.049399, 
    -17.00998, -36.7803, -41.60369, -33.01459, -37.75272, -39.97875, 
    -25.42138, 12.82028,
  42.01719, 30.13895, 3.615799, -1.955472, -7.306231, 3.914696, -20.13835, 
    -4.906138, -13.41107, -18.59382, -30.23593, -33.26091, -25.67199, 
    -17.05147, -3.5565,
  57.28447, 39.15798, 21.80513, 2.129856, -2.835824, -14.59327, -14.67744, 
    -37.20589, -16.06759, 6.725023, -16.3041, -24.49639, -21.44041, 
    -14.42536, -17.04887,
  42.9108, 44.45652, 31.52642, 7.272937, -2.395375, -5.53306, -22.36517, 
    -24.69203, -8.065418, -7.273682, -1.704108, -18.32451, -16.8744, 
    -12.01433, -8.097999,
  44.73549, 48.08462, 23.39513, 11.76415, 1.937233, -1.918497, -6.015941, 
    -11.1264, -15.15309, -14.55598, -15.39582, -13.69446, -12.71925, 
    -11.42002, -8.506005,
  47.59138, 41.08615, 22.90215, 16.27361, 11.82917, 1.719893, -2.415322, 
    -6.070196, -9.575216, -9.562228, -9.917851, -8.155359, -7.878132, 
    -7.339599, -8.602995,
  39.75224, 17.15945, 10.61546, 10.40156, 11.87544, 7.054586, 0.3559759, 
    0.02567648, -1.740079, -2.486393, -3.184426, -2.594942, -2.509681, 
    -2.529807, -4.602253,
  17.2882, 6.963691, 4.373751, 6.11458, 13.06264, 10.11943, 5.796793, 
    4.038726, 2.831785, 3.058843, 2.845948, 2.245825, 1.537632, 1.087546, 
    2.153493,
  3.163681, -0.1148655, 16.6295, 1.171271, 7.523092, 28.04642, -0.6350574, 
    -6.44892, -1.986472, 61.31538, 67.60756, 28.82223, 71.03835, 60.8048, 
    117.3155,
  0.4266997, -1.239901, -0.7607331, 0.03691828, 45.90921, 44.75702, 
    -1.886162, -5.39238, -5.337804, 0.06183699, 35.64378, -23.01021, 
    -24.13087, 74.26709, 99.9277,
  11.38618, 6.223752, 0.07030962, -0.3423976, 25.90446, -2.157321, 6.360395, 
    -3.516978, -4.483541, -27.4613, -43.82153, -30.78769, -35.24909, 
    -16.18486, 25.83948,
  35.51102, 22.57857, 1.222785, 0.1991669, -1.926375, 21.04213, -2.757545, 
    3.64329, -5.087921, -15.85838, -37.54645, -35.80604, -30.18942, 
    -18.39124, -1.523378,
  47.31236, 27.80067, 12.70558, 0.3353549, -3.449059, -5.18259, 2.70359, 
    -8.581849, -7.744313, 8.406247, -21.22906, -26.85977, -26.70205, 
    -18.2919, -11.28847,
  32.04221, 35.67815, 18.69378, 2.596593, -1.679235, -4.249856, -9.39783, 
    -9.045596, 2.213144, -2.193112, -0.5193694, -24.27601, -21.40582, 
    -17.11897, -8.174153,
  47.4451, 46.19199, 13.86836, 2.355797, -0.5490658, -2.472077, -7.45305, 
    -8.834955, -11.89811, -12.45212, -17.61066, -22.10048, -19.10714, 
    -17.152, -10.82546,
  54.53809, 48.273, 17.82028, 7.294885, 3.240343, -0.1966553, -5.993449, 
    -9.500063, -12.88028, -13.2091, -12.92623, -17.27656, -17.22673, 
    -16.83039, -12.44643,
  39.80802, 30.93507, 14.84368, 9.561326, 4.210364, -0.5315881, -2.31308, 
    -5.476195, -9.662354, -10.68531, -10.56624, -12.48429, -15.01889, 
    -14.73772, -11.78287,
  19.04305, 20.01595, 10.29216, 12.6389, 12.96039, 3.330249, -1.163898, 
    -3.864909, -5.749431, -8.424107, -9.353343, -10.97929, -11.48853, 
    -11.4431, -10.56309,
  3.540786, 2.598935, 20.33898, 4.58819, 9.477996, 22.32166, -0.2980984, 
    -1.740566, -0.6259034, 44.81991, 71.325, 35.96699, 73.62505, 61.02653, 
    89.08531,
  -2.196887, 0.5748385, 6.423485, 6.067542, 27.71469, 32.77969, -0.2430129, 
    -2.374896, -3.34435, 6.964757, 54.98528, 3.930795, 2.536107, 71.66277, 
    83.79198,
  2.173014, 6.676159, 7.49361, 3.836789, 18.02339, 2.747216, 8.55291, 
    -4.103326, -3.547363, -7.251332, -10.31044, -0.1210544, -8.277349, 
    -7.599751, 29.61217,
  12.94779, 16.46464, 9.489152, 7.212506, 1.552138, 25.67267, 2.630281, 
    7.645096, -3.275418, -8.030193, -17.39736, -13.72806, -9.516129, 
    -10.58768, 7.164935,
  16.03372, 18.81012, 12.37054, 3.755628, -0.4116108, 0.3860964, 7.930712, 
    3.334033, -2.888928, 9.125685, -9.398604, -12.60598, -7.704383, 
    -9.378465, -12.77787,
  13.11731, 24.13904, 13.20375, 1.512056, -0.7079181, -0.6129923, -1.397547, 
    0.09489345, 6.022583, -2.712105, 7.291915, -11.49469, -7.417047, 
    -7.003356, -9.408215,
  19.98664, 34.66796, 9.789346, 0.663168, -0.0707467, -0.4841461, -0.8618392, 
    -1.736901, -5.254347, -14.89423, -13.26754, -10.3067, -8.892595, 
    -7.82117, -8.769135,
  26.58099, 38.34003, 13.43721, 2.702815, 0.6052585, 0.1962099, -0.645403, 
    -1.080709, -4.268177, -11.40062, -10.67041, -11.62847, -10.324, 
    -7.253909, -5.166348,
  21.11982, 27.81017, 12.85135, 4.696507, 0.4065037, -0.07641088, -0.1499249, 
    0.3359508, -2.341281, -6.727863, -7.326422, -10.14646, -9.608006, 
    -8.69521, -4.022734,
  13.95255, 20.6263, 13.53811, 11.23819, 4.998913, -0.1916883, 0.07556101, 
    -0.006485153, -1.726797, -4.27911, -5.636862, -8.301988, -7.717674, 
    -8.02482, -6.884194,
  8.505408, 1.166176, 16.31195, 3.944232, 9.397185, 20.27451, 6.197559, 
    7.199944, 4.202302, 63.24072, 58.96786, 27.24309, 35.79866, 46.43909, 
    101.4929,
  0.3098592, 0.1414336, 0.7613322, 3.546805, 30.74776, 31.30085, 6.439806, 
    5.847007, 1.075507, 15.122, 64.08773, 11.33199, -0.9736633, 45.02871, 
    93.32632,
  0.7079218, 0.3743495, 0.6271619, 3.503035, 22.84511, 19.48786, 14.54798, 
    4.167799, 0.7227295, -0.03574219, 19.52776, 12.37372, -3.98758, 
    -15.22787, 32.63584,
  2.256089, 0.5555296, 0.616933, 6.51719, 7.430949, 31.6597, 17.16877, 
    20.982, 1.510894, -2.899461, -2.079111, -0.3726342, -8.49329, -19.04408, 
    3.120905,
  1.144431, -0.7262238, 5.233365, 10.71468, 9.034482, 11.84904, 26.50241, 
    19.15721, 11.74655, 14.44099, -1.459586, -0.7497969, -6.451662, 
    -19.39128, -23.50856,
  2.549067, 1.955222, 8.933493, 8.542169, 8.64341, 9.599121, 6.412053, 
    15.22744, 19.93791, 14.46657, 9.833583, -0.3961217, -4.544941, -16.20538, 
    -20.33986,
  9.765165, 10.16125, 1.985384, 0.988703, 2.90216, 5.056383, 5.066834, 
    4.703452, 6.190238, 3.241025, 0.8515327, -0.1425847, -4.647602, 
    -13.85817, -17.24264,
  22.03675, 11.8261, 1.423945, -0.6912557, 1.301231, 4.363756, 2.021703, 
    1.714607, 6.796333, 4.380194, 1.7318, -0.3977358, -5.504348, -13.01643, 
    -13.88054,
  21.81513, 4.899354, 0.9547924, 1.943287, 0.359844, 3.254478, 3.635701, 
    4.16113, 6.328898, 4.138492, 1.742875, -0.9455946, -5.746451, -13.07666, 
    -11.81589,
  14.30136, 4.022938, 3.644439, 5.65098, 3.611544, 2.926721, 4.551373, 
    6.517334, 7.575497, 3.993905, 2.940333, -1.151662, -4.724422, -10.92478, 
    -12.09309,
  10.88333, 6.89333, 30.96664, 9.157907, 13.89038, 27.03804, 13.10994, 
    7.15241, 0.6930008, 20.6331, 30.57813, 28.976, 48.32071, 40.42844, 
    78.79162,
  2.301409, 2.080948, 3.263663, 5.422714, 33.87572, 38.09546, 7.688189, 
    10.0197, 1.285419, 4.929044, 33.32828, 9.196508, -1.386133, 43.92007, 
    70.78606,
  1.062887, 2.906348, 2.647925, 1.032501, 22.82162, 18.83229, 14.94208, 
    6.694458, 4.247019, 1.431376, 34.41257, 26.55839, 2.73777, -7.371563, 
    24.29827,
  1.730494, 2.4648, 2.507087, 2.413806, 0.9766299, 20.728, 17.03017, 
    19.64763, 6.472195, 5.219203, 4.886965, 4.176173, -3.976362, -8.193698, 
    7.090415,
  1.860116, 0.6143277, 2.028711, 2.264664, 2.236318, 3.907608, 17.50616, 
    17.85267, 16.97728, 22.0835, 5.834577, -0.5829059, -3.685256, -6.774089, 
    -10.03998,
  3.841636, -0.5401679, -2.494952, -3.160645, -1.005944, 2.722351, 4.574387, 
    11.08345, 19.22344, 23.03929, 25.51372, 2.938745, -2.210304, -6.128382, 
    -9.183692,
  14.11183, 1.813288, -4.664318, -5.208842, -4.192281, -3.129141, -0.1475298, 
    2.142887, 4.990086, 7.66396, 9.485415, 6.09054, -0.9041244, -4.713547, 
    -7.532806,
  26.96924, 8.116384, -0.7147879, -2.624593, -2.045427, -1.958331, -3.891532, 
    -3.574209, 1.590985, 8.16889, 9.527815, 7.722002, 0.7398774, -2.990683, 
    -6.139617,
  32.80539, 14.70591, 1.940143, 1.230729, 0.5720527, -0.07222234, -2.137377, 
    -0.5339401, 2.18285, 7.709863, 10.18138, 6.817613, 1.579942, -2.351955, 
    -3.897361,
  31.49116, 21.23027, 6.259309, 4.348137, 3.749676, 1.076126, 3.012861, 
    4.741405, 5.852178, 16.61294, 13.89794, 7.886201, 0.9961908, -1.809693, 
    -4.685159 ;

 nv = 1, 2 ;

 pfull = 0.0252729048206747, 0.0885404738757409, 0.213072411383256, 
    0.41190537807884, 0.671080828691593, 0.987471468515016, 1.36790961365676, 
    1.82562112064242, 2.38097588033244, 3.06218961364243, 3.90121721567151, 
    4.9296281825995, 6.18008131929323, 7.68875807563375, 9.49537809361575, 
    11.643153995098, 14.1786857151188, 17.1517875598959, 20.6152476986609, 
    24.6245259348741, 29.237386591333, 34.5134757786445, 40.5138467378254, 
    47.3004421634272, 54.9355325495126, 63.4811392623337, 72.9984371159701, 
    83.5471442618119, 95.1849171805989, 107.966767294215, 121.944503506415, 
    137.166169497631, 153.675572970355, 171.511834307961, 190.708985325578, 
    211.295632932361, 233.294677858721, 256.723099608772, 281.591803639405, 
    307.905555737256, 335.66293113824, 364.856338389786, 395.47216160598, 
    427.490864234311, 460.887168786725, 495.630391513078, 531.761718445649, 
    569.289185351388, 607.768705103107, 646.445374671436, 684.792067788697, 
    722.468679913451, 759.124006783627, 794.401045766566, 827.769968639223, 
    858.597822486016, 886.389109609622, 910.841030891388, 931.860653469283, 
    949.549679924174, 964.159924710431, 976.012345333387, 985.470174132691, 
    992.77226220014, 997.948601287575 ;

 phalf = 0.01, 0.0513470268, 0.1404240036, 0.3072783852, 0.5379505539, 
    0.8245489502, 1.170559845, 1.5862843323, 2.0879000854, 2.700272522, 
    3.4550848389, 4.3841940308, 5.5185266113, 6.8925054932, 8.5440936279, 
    10.5147802734, 12.8495031738, 15.5965148926, 18.8071691895, 
    22.5356542969, 26.8386547852, 31.7749560547, 37.4049951172, 
    43.7903613281, 50.9932617188, 59.0759326172, 68.100078125, 78.1262353516, 
    89.2131933594, 101.4173632812, 114.7922466406, 129.3878501562, 
    145.2501478125, 162.4206823438, 180.9360560938, 200.8276451562, 
    222.1212074219, 244.8367185938, 268.9881007812, 294.5831945312, 
    321.6236510156, 350.1049399219, 380.0163883594, 411.3414303125, 
    444.0575547656, 478.1367280469, 513.5456339062, 550.403556875, 
    588.6019571094, 627.3470909766, 665.9273852344, 704.0097012891, 
    741.2475327734, 777.2856108203, 811.7659041211, 843.9830114648, 
    873.3803854492, 899.5263707422, 922.2501762402, 941.5376650684, 
    957.6070185254, 970.7426572876, 981.30107, 989.65107, 995.9000099865, 1000 ;

 pk = 1, 5.134703, 14.0424, 30.72784, 53.79506, 82.4549, 117.056, 158.6284, 
    208.79, 270.0273, 345.5085, 438.4194, 551.8527, 689.2505, 854.4094, 
    1051.478, 1284.95, 1559.651, 1880.717, 2253.565, 2683.865, 3177.496, 
    3740.5, 4379.036, 5099.326, 5907.593, 6810.008, 7812.624, 8921.319, 
    10141.74, 11285.93, 12188.79, 12884.3, 13400.12, 13758.85, 13979.1, 
    14076.26, 14063.13, 13950.46, 13747.31, 13461.45, 13099.54, 12667.38, 
    12170.08, 11612.19, 10997.8, 10330.65, 9611.055, 8843.304, 8045.85, 
    7236.312, 6424.557, 5606.509, 4778.059, 3944.972, 3146.775, 2416.634, 
    1778.226, 1246.215, 826.5195, 511.2139, 290.7407, 150, 68.893, 14.999, 0 ;

 scalar_axis = 0 ;

 time = 0.5, 1.5, 2.5, 3.5, 4.5, 5.5, 6.5, 7.5, 8.5, 9.5, 10.5, 11.5, 12.5, 
    13.5, 14.5, 15.5, 16.5, 17.5, 18.5, 19.5, 20.5, 21.5, 22.5, 23.5, 24.5, 
    25.5, 26.5, 27.5, 28.5, 29.5, 30.5, 31.5, 32.5, 33.5, 34.5, 35.5, 36.5, 
    37.5, 38.5, 39.5, 40.5, 41.5, 42.5, 43.5, 44.5, 45.5, 46.5, 47.5, 48.5, 
    49.5, 50.5, 51.5, 52.5, 53.5, 54.5, 55.5, 56.5, 57.5, 58.5, 59.5, 60.5, 
    61.5, 62.5, 63.5, 64.5, 65.5, 66.5, 67.5, 68.5, 69.5, 70.5, 71.5, 72.5, 
    73.5, 74.5, 75.5, 76.5, 77.5, 78.5, 79.5, 80.5, 81.5, 82.5, 83.5, 84.5, 
    85.5, 86.5, 87.5, 88.5, 89.5, 90.5, 91.5, 92.5, 93.5, 94.5, 95.5, 96.5, 
    97.5, 98.5, 99.5, 100.5, 101.5, 102.5, 103.5, 104.5, 105.5, 106.5, 107.5, 
    108.5, 109.5, 110.5, 111.5, 112.5, 113.5, 114.5, 115.5, 116.5, 117.5, 
    118.5, 119.5, 120.5, 121.5, 122.5, 123.5, 124.5, 125.5, 126.5, 127.5, 
    128.5, 129.5, 130.5, 131.5, 132.5, 133.5, 134.5, 135.5, 136.5, 137.5, 
    138.5, 139.5, 140.5, 141.5, 142.5, 143.5, 144.5, 145.5, 146.5, 147.5, 
    148.5, 149.5, 150.5, 151.5, 152.5, 153.5, 154.5, 155.5, 156.5, 157.5, 
    158.5, 159.5, 160.5, 161.5, 162.5, 163.5, 164.5, 165.5, 166.5, 167.5, 
    168.5, 169.5, 170.5, 171.5, 172.5, 173.5, 174.5, 175.5, 176.5, 177.5, 
    178.5, 179.5, 180.5, 181.5 ;

 time_bnds =
  0, 1,
  1, 2,
  2, 3,
  3, 4,
  4, 5,
  5, 6,
  6, 7,
  7, 8,
  8, 9,
  9, 10,
  10, 11,
  11, 12,
  12, 13,
  13, 14,
  14, 15,
  15, 16,
  16, 17,
  17, 18,
  18, 19,
  19, 20,
  20, 21,
  21, 22,
  22, 23,
  23, 24,
  24, 25,
  25, 26,
  26, 27,
  27, 28,
  28, 29,
  29, 30,
  30, 31,
  31, 32,
  32, 33,
  33, 34,
  34, 35,
  35, 36,
  36, 37,
  37, 38,
  38, 39,
  39, 40,
  40, 41,
  41, 42,
  42, 43,
  43, 44,
  44, 45,
  45, 46,
  46, 47,
  47, 48,
  48, 49,
  49, 50,
  50, 51,
  51, 52,
  52, 53,
  53, 54,
  54, 55,
  55, 56,
  56, 57,
  57, 58,
  58, 59,
  59, 60,
  60, 61,
  61, 62,
  62, 63,
  63, 64,
  64, 65,
  65, 66,
  66, 67,
  67, 68,
  68, 69,
  69, 70,
  70, 71,
  71, 72,
  72, 73,
  73, 74,
  74, 75,
  75, 76,
  76, 77,
  77, 78,
  78, 79,
  79, 80,
  80, 81,
  81, 82,
  82, 83,
  83, 84,
  84, 85,
  85, 86,
  86, 87,
  87, 88,
  88, 89,
  89, 90,
  90, 91,
  91, 92,
  92, 93,
  93, 94,
  94, 95,
  95, 96,
  96, 97,
  97, 98,
  98, 99,
  99, 100,
  100, 101,
  101, 102,
  102, 103,
  103, 104,
  104, 105,
  105, 106,
  106, 107,
  107, 108,
  108, 109,
  109, 110,
  110, 111,
  111, 112,
  112, 113,
  113, 114,
  114, 115,
  115, 116,
  116, 117,
  117, 118,
  118, 119,
  119, 120,
  120, 121,
  121, 122,
  122, 123,
  123, 124,
  124, 125,
  125, 126,
  126, 127,
  127, 128,
  128, 129,
  129, 130,
  130, 131,
  131, 132,
  132, 133,
  133, 134,
  134, 135,
  135, 136,
  136, 137,
  137, 138,
  138, 139,
  139, 140,
  140, 141,
  141, 142,
  142, 143,
  143, 144,
  144, 145,
  145, 146,
  146, 147,
  147, 148,
  148, 149,
  149, 150,
  150, 151,
  151, 152,
  152, 153,
  153, 154,
  154, 155,
  155, 156,
  156, 157,
  157, 158,
  158, 159,
  159, 160,
  160, 161,
  161, 162,
  162, 163,
  163, 164,
  164, 165,
  165, 166,
  166, 167,
  167, 168,
  168, 169,
  169, 170,
  170, 171,
  171, 172,
  172, 173,
  173, 174,
  174, 175,
  175, 176,
  176, 177,
  177, 178,
  178, 179,
  179, 180,
  180, 181,
  181, 182 ;
}
