netcdf \20030101.grid_spec.tile1 {
dimensions:
	grid_x = 97 ;
	grid_y = 97 ;
	time = UNLIMITED ; // (1 currently)
	grid_xt = 96 ;
	grid_yt = 96 ;
	phalf = 50 ;
variables:
	double grid_x(grid_x) ;
		grid_x:units = "degrees_E" ;
		grid_x:long_name = "cell corner longitude" ;
		grid_x:axis = "X" ;
	double grid_y(grid_y) ;
		grid_y:units = "degrees_N" ;
		grid_y:long_name = "cell corner latitude" ;
		grid_y:axis = "Y" ;
	double time(time) ;
		time:units = "days since 1870-01-01 00:00:00" ;
		time:long_name = "time" ;
		time:axis = "T" ;
		time:calendar_type = "JULIAN" ;
		time:calendar = "julian" ;
	double grid_xt(grid_xt) ;
		grid_xt:units = "degrees_E" ;
		grid_xt:long_name = "T-cell longitude" ;
		grid_xt:axis = "X" ;
	double grid_yt(grid_yt) ;
		grid_yt:units = "degrees_N" ;
		grid_yt:long_name = "T-cell latitude" ;
		grid_yt:axis = "Y" ;
	double phalf(phalf) ;
		phalf:units = "mb" ;
		phalf:long_name = "ref half pressure level" ;
		phalf:axis = "Z" ;
		phalf:positive = "down" ;
	float grid_lon(grid_y, grid_x) ;
		grid_lon:_FillValue = 1.e+20f ;
		grid_lon:missing_value = 1.e+20f ;
		grid_lon:units = "degrees_E" ;
		grid_lon:long_name = "longitude" ;
		grid_lon:cell_methods = "time: point" ;
	float grid_lat(grid_y, grid_x) ;
		grid_lat:_FillValue = 1.e+20f ;
		grid_lat:missing_value = 1.e+20f ;
		grid_lat:units = "degrees_N" ;
		grid_lat:long_name = "latitude" ;
		grid_lat:cell_methods = "time: point" ;
	float grid_lont(grid_yt, grid_xt) ;
		grid_lont:_FillValue = 1.e+20f ;
		grid_lont:missing_value = 1.e+20f ;
		grid_lont:units = "degrees_E" ;
		grid_lont:long_name = "longitude" ;
		grid_lont:cell_methods = "time: point" ;
	float grid_latt(grid_yt, grid_xt) ;
		grid_latt:_FillValue = 1.e+20f ;
		grid_latt:missing_value = 1.e+20f ;
		grid_latt:units = "degrees_N" ;
		grid_latt:long_name = "latitude" ;
		grid_latt:cell_methods = "time: point" ;
	float area(grid_yt, grid_xt) ;
		area:_FillValue = 1.e+20f ;
		area:missing_value = 1.e+20f ;
		area:units = "m**2" ;
		area:long_name = "cell area" ;
		area:cell_methods = "time: point" ;
	float bk(phalf) ;
		bk:_FillValue = 1.e+20f ;
		bk:missing_value = 1.e+20f ;
		bk:long_name = "vertical coordinate sigma value" ;
		bk:cell_methods = "time: point" ;
	float pk(phalf) ;
		pk:_FillValue = 1.e+20f ;
		pk:missing_value = 1.e+20f ;
		pk:units = "pascal" ;
		pk:long_name = "pressure part of the hybrid coordinate" ;
		pk:cell_methods = "time: point" ;
	float sftlf(grid_yt, grid_xt) ;
		sftlf:_FillValue = 1.e+20f ;
		sftlf:missing_value = 1.e+20f ;
		sftlf:units = "1.0" ;
		sftlf:long_name = "Fraction of the Grid Cell Occupied by Land" ;
		sftlf:cell_methods = "time: point" ;
		sftlf:cell_measures = "area: area" ;
		sftlf:standard_name = "land_area_fraction" ;
		sftlf:interp_method = "conserve_order1" ;
	float orog(grid_yt, grid_xt) ;
		orog:_FillValue = 1.e+20f ;
		orog:missing_value = 1.e+20f ;
		orog:units = "m" ;
		orog:long_name = "Surface Altitude" ;
		orog:cell_methods = "time: point" ;
		orog:cell_measures = "area: area" ;
		orog:standard_name = "surface_altitude" ;
		orog:interp_method = "conserve_order1" ;
	float land_mask(grid_yt, grid_xt) ;
		land_mask:_FillValue = 1.e+20f ;
		land_mask:missing_value = 1.e+20f ;
		land_mask:valid_range = -0.01f, 1.01f ;
		land_mask:long_name = "fractional amount of land" ;
		land_mask:cell_methods = "time: point" ;
		land_mask:interp_method = "conserve_order1" ;
	float zsurf(grid_yt, grid_xt) ;
		zsurf:_FillValue = 1.e+20f ;
		zsurf:missing_value = 1.e+20f ;
		zsurf:units = "m" ;
		zsurf:long_name = "surface height" ;
		zsurf:cell_methods = "time: point" ;

// global attributes:
		:title = "ESM4_longamip_D1_am4p2_proto7b_whiteCapsAlbedo_salt_SIS2" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
data:

 grid_x = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19, 
    20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 37, 
    38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 54, 55, 
    56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 72, 73, 
    74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 90, 91, 
    92, 93, 94, 95, 96, 97 ;

 grid_y = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19, 
    20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 37, 
    38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 54, 55, 
    56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 72, 73, 
    74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 90, 91, 
    92, 93, 94, 95, 96, 97 ;

 time = 0 ;

 grid_xt = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19, 
    20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 37, 
    38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 54, 55, 
    56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 72, 73, 
    74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 90, 91, 
    92, 93, 94, 95, 96 ;

 grid_yt = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19, 
    20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 37, 
    38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 54, 55, 
    56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 72, 73, 
    74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 90, 91, 
    92, 93, 94, 95, 96 ;

 phalf = 0.01, 0.0269722, 0.0517136, 0.0889455, 0.142479, 0.2207157, 
    0.3361283, 0.5048096, 0.7479993, 1.0940055, 1.580046, 2.2544108, 
    3.178956, 4.431935, 6.1111558, 8.3374392, 11.2583405, 15.0520759, 
    19.9315829, 26.1486254, 33.997842, 43.820624, 56.0087014, 71.0073115, 
    89.3178242, 111.4997021, 138.1716841, 170.012093, 207.7581856, 
    252.2033875, 304.1464563, 363.9522552, 430.6429622, 501.015122, 
    570.6113482, 635.806353, 694.8286462, 747.1992533, 793.0044191, 
    832.5750255, 866.4443202, 895.1917865, 919.4060705, 939.6860264, 
    956.4664631, 970.1833931, 981.1347983, 989.68, 995.9, 1000 ;

 grid_lon =
  305, 305.7828, 306.5727, 307.3698, 308.1741, 308.9857, 309.8047, 310.6309, 
    311.4646, 312.3057, 313.1541, 314.01, 314.8733, 315.744, 316.6221, 
    317.5075, 318.4002, 319.3002, 320.2073, 321.1216, 322.043, 322.9712, 
    323.9063, 324.8481, 325.7966, 326.7514, 327.7126, 328.6799, 329.6532, 
    330.6322, 331.6168, 332.6068, 333.6019, 334.6019, 335.6065, 336.6156, 
    337.6287, 338.6458, 339.6663, 340.6902, 341.717, 342.7465, 343.7783, 
    344.8122, 345.8477, 346.8846, 347.9225, 348.9611, 350, 351.0389, 
    352.0775, 353.1154, 354.1523, 355.1878, 356.2217, 357.2535, 358.283, 
    359.3098, 0.3336662, 1.354252, 2.371273, 3.384442, 4.393482, 5.398128, 
    6.39812, 7.393215, 8.383177, 9.367781, 10.34682, 11.32008, 12.28739, 
    13.24856, 14.20343, 15.15185, 16.09367, 17.02878, 17.95705, 18.87837, 
    19.79265, 20.69982, 21.59979, 22.49251, 23.37793, 24.256, 25.12669, 
    25.98999, 26.84588, 27.69435, 28.53541, 29.36907, 30.19535, 31.01428, 
    31.82589, 32.63021, 33.42731, 34.21722, 35,
  305, 305.7828, 306.5727, 307.3698, 308.1741, 308.9857, 309.8047, 310.6309, 
    311.4646, 312.3057, 313.1541, 314.01, 314.8733, 315.744, 316.6221, 
    317.5075, 318.4002, 319.3002, 320.2073, 321.1216, 322.043, 322.9712, 
    323.9063, 324.8481, 325.7966, 326.7514, 327.7126, 328.6799, 329.6532, 
    330.6322, 331.6168, 332.6068, 333.6019, 334.6019, 335.6065, 336.6156, 
    337.6287, 338.6458, 339.6663, 340.6902, 341.717, 342.7465, 343.7783, 
    344.8122, 345.8477, 346.8846, 347.9225, 348.9611, 350, 351.0389, 
    352.0775, 353.1154, 354.1523, 355.1878, 356.2217, 357.2535, 358.283, 
    359.3098, 0.3336662, 1.354252, 2.371273, 3.384442, 4.393482, 5.398128, 
    6.39812, 7.393215, 8.383177, 9.367781, 10.34682, 11.32008, 12.28739, 
    13.24856, 14.20343, 15.15185, 16.09367, 17.02878, 17.95705, 18.87837, 
    19.79265, 20.69982, 21.59979, 22.49251, 23.37793, 24.256, 25.12669, 
    25.98999, 26.84588, 27.69435, 28.53541, 29.36907, 30.19535, 31.01428, 
    31.82589, 32.63021, 33.42731, 34.21722, 35,
  305, 305.7828, 306.5727, 307.3698, 308.1741, 308.9857, 309.8047, 310.6309, 
    311.4646, 312.3057, 313.1541, 314.01, 314.8733, 315.744, 316.6221, 
    317.5075, 318.4002, 319.3002, 320.2073, 321.1216, 322.043, 322.9712, 
    323.9063, 324.8481, 325.7966, 326.7514, 327.7126, 328.6799, 329.6532, 
    330.6322, 331.6168, 332.6068, 333.6019, 334.6019, 335.6065, 336.6156, 
    337.6287, 338.6458, 339.6663, 340.6902, 341.717, 342.7465, 343.7783, 
    344.8122, 345.8477, 346.8846, 347.9225, 348.9611, 350, 351.0389, 
    352.0775, 353.1154, 354.1523, 355.1878, 356.2217, 357.2535, 358.283, 
    359.3098, 0.3336662, 1.354252, 2.371273, 3.384442, 4.393482, 5.398128, 
    6.39812, 7.393215, 8.383177, 9.367781, 10.34682, 11.32008, 12.28739, 
    13.24856, 14.20343, 15.15185, 16.09367, 17.02878, 17.95705, 18.87837, 
    19.79265, 20.69982, 21.59979, 22.49251, 23.37793, 24.256, 25.12669, 
    25.98999, 26.84588, 27.69435, 28.53541, 29.36907, 30.19535, 31.01428, 
    31.82589, 32.63021, 33.42731, 34.21722, 35,
  305, 305.7828, 306.5727, 307.3698, 308.1741, 308.9857, 309.8047, 310.6309, 
    311.4646, 312.3057, 313.1541, 314.01, 314.8733, 315.744, 316.6221, 
    317.5075, 318.4002, 319.3002, 320.2073, 321.1216, 322.043, 322.9712, 
    323.9063, 324.8481, 325.7966, 326.7514, 327.7126, 328.6799, 329.6532, 
    330.6322, 331.6168, 332.6068, 333.6019, 334.6019, 335.6065, 336.6156, 
    337.6287, 338.6458, 339.6663, 340.6902, 341.717, 342.7465, 343.7783, 
    344.8122, 345.8477, 346.8846, 347.9225, 348.9611, 350, 351.0389, 
    352.0775, 353.1154, 354.1523, 355.1878, 356.2217, 357.2535, 358.283, 
    359.3098, 0.3336662, 1.354252, 2.371273, 3.384442, 4.393482, 5.398128, 
    6.39812, 7.393215, 8.383177, 9.367781, 10.34682, 11.32008, 12.28739, 
    13.24856, 14.20343, 15.15185, 16.09367, 17.02878, 17.95705, 18.87837, 
    19.79265, 20.69982, 21.59979, 22.49251, 23.37793, 24.256, 25.12669, 
    25.98999, 26.84588, 27.69435, 28.53541, 29.36907, 30.19535, 31.01428, 
    31.82589, 32.63021, 33.42731, 34.21722, 35,
  305, 305.7828, 306.5727, 307.3698, 308.1741, 308.9857, 309.8047, 310.6309, 
    311.4646, 312.3057, 313.1541, 314.01, 314.8733, 315.744, 316.6221, 
    317.5075, 318.4002, 319.3002, 320.2073, 321.1216, 322.043, 322.9712, 
    323.9063, 324.8481, 325.7966, 326.7514, 327.7126, 328.6799, 329.6532, 
    330.6322, 331.6168, 332.6068, 333.6019, 334.6019, 335.6065, 336.6156, 
    337.6287, 338.6458, 339.6663, 340.6902, 341.717, 342.7465, 343.7783, 
    344.8122, 345.8477, 346.8846, 347.9225, 348.9611, 350, 351.0389, 
    352.0775, 353.1154, 354.1523, 355.1878, 356.2217, 357.2535, 358.283, 
    359.3098, 0.3336662, 1.354252, 2.371273, 3.384442, 4.393482, 5.398128, 
    6.39812, 7.393215, 8.383177, 9.367781, 10.34682, 11.32008, 12.28739, 
    13.24856, 14.20343, 15.15185, 16.09367, 17.02878, 17.95705, 18.87837, 
    19.79265, 20.69982, 21.59979, 22.49251, 23.37793, 24.256, 25.12669, 
    25.98999, 26.84588, 27.69435, 28.53541, 29.36907, 30.19535, 31.01428, 
    31.82589, 32.63021, 33.42731, 34.21722, 35,
  305, 305.7828, 306.5727, 307.3698, 308.1741, 308.9857, 309.8047, 310.6309, 
    311.4646, 312.3057, 313.1541, 314.01, 314.8733, 315.744, 316.6221, 
    317.5075, 318.4002, 319.3002, 320.2073, 321.1216, 322.043, 322.9712, 
    323.9063, 324.8481, 325.7966, 326.7514, 327.7126, 328.6799, 329.6532, 
    330.6322, 331.6168, 332.6068, 333.6019, 334.6019, 335.6065, 336.6156, 
    337.6287, 338.6458, 339.6663, 340.6902, 341.717, 342.7465, 343.7783, 
    344.8122, 345.8477, 346.8846, 347.9225, 348.9611, 350, 351.0389, 
    352.0775, 353.1154, 354.1523, 355.1878, 356.2217, 357.2535, 358.283, 
    359.3098, 0.3336662, 1.354252, 2.371273, 3.384442, 4.393482, 5.398128, 
    6.39812, 7.393215, 8.383177, 9.367781, 10.34682, 11.32008, 12.28739, 
    13.24856, 14.20343, 15.15185, 16.09367, 17.02878, 17.95705, 18.87837, 
    19.79265, 20.69982, 21.59979, 22.49251, 23.37793, 24.256, 25.12669, 
    25.98999, 26.84588, 27.69435, 28.53541, 29.36907, 30.19535, 31.01428, 
    31.82589, 32.63021, 33.42731, 34.21722, 35,
  305, 305.7828, 306.5727, 307.3698, 308.1741, 308.9857, 309.8047, 310.6309, 
    311.4646, 312.3057, 313.1541, 314.01, 314.8733, 315.744, 316.6221, 
    317.5075, 318.4002, 319.3002, 320.2073, 321.1216, 322.043, 322.9712, 
    323.9063, 324.8481, 325.7966, 326.7514, 327.7126, 328.6799, 329.6532, 
    330.6322, 331.6168, 332.6068, 333.6019, 334.6019, 335.6065, 336.6156, 
    337.6287, 338.6458, 339.6663, 340.6902, 341.717, 342.7465, 343.7783, 
    344.8122, 345.8477, 346.8846, 347.9225, 348.9611, 350, 351.0389, 
    352.0775, 353.1154, 354.1523, 355.1878, 356.2217, 357.2535, 358.283, 
    359.3098, 0.3336662, 1.354252, 2.371273, 3.384442, 4.393482, 5.398128, 
    6.39812, 7.393215, 8.383177, 9.367781, 10.34682, 11.32008, 12.28739, 
    13.24856, 14.20343, 15.15185, 16.09367, 17.02878, 17.95705, 18.87837, 
    19.79265, 20.69982, 21.59979, 22.49251, 23.37793, 24.256, 25.12669, 
    25.98999, 26.84588, 27.69435, 28.53541, 29.36907, 30.19535, 31.01428, 
    31.82589, 32.63021, 33.42731, 34.21722, 35,
  305, 305.7828, 306.5727, 307.3698, 308.1741, 308.9857, 309.8047, 310.6309, 
    311.4646, 312.3057, 313.1541, 314.01, 314.8733, 315.744, 316.6221, 
    317.5075, 318.4002, 319.3002, 320.2073, 321.1216, 322.043, 322.9712, 
    323.9063, 324.8481, 325.7966, 326.7514, 327.7126, 328.6799, 329.6532, 
    330.6322, 331.6168, 332.6068, 333.6019, 334.6019, 335.6065, 336.6156, 
    337.6287, 338.6458, 339.6663, 340.6902, 341.717, 342.7465, 343.7783, 
    344.8122, 345.8477, 346.8846, 347.9225, 348.9611, 350, 351.0389, 
    352.0775, 353.1154, 354.1523, 355.1878, 356.2217, 357.2535, 358.283, 
    359.3098, 0.3336662, 1.354252, 2.371273, 3.384442, 4.393482, 5.398128, 
    6.39812, 7.393215, 8.383177, 9.367781, 10.34682, 11.32008, 12.28739, 
    13.24856, 14.20343, 15.15185, 16.09367, 17.02878, 17.95705, 18.87837, 
    19.79265, 20.69982, 21.59979, 22.49251, 23.37793, 24.256, 25.12669, 
    25.98999, 26.84588, 27.69435, 28.53541, 29.36907, 30.19535, 31.01428, 
    31.82589, 32.63021, 33.42731, 34.21722, 35,
  305, 305.7828, 306.5727, 307.3698, 308.1741, 308.9857, 309.8047, 310.6309, 
    311.4646, 312.3057, 313.1541, 314.01, 314.8733, 315.744, 316.6221, 
    317.5075, 318.4002, 319.3002, 320.2073, 321.1216, 322.043, 322.9712, 
    323.9063, 324.8481, 325.7966, 326.7514, 327.7126, 328.6799, 329.6532, 
    330.6322, 331.6168, 332.6068, 333.6019, 334.6019, 335.6065, 336.6156, 
    337.6287, 338.6458, 339.6663, 340.6902, 341.717, 342.7465, 343.7783, 
    344.8122, 345.8477, 346.8846, 347.9225, 348.9611, 350, 351.0389, 
    352.0775, 353.1154, 354.1523, 355.1878, 356.2217, 357.2535, 358.283, 
    359.3098, 0.3336662, 1.354252, 2.371273, 3.384442, 4.393482, 5.398128, 
    6.39812, 7.393215, 8.383177, 9.367781, 10.34682, 11.32008, 12.28739, 
    13.24856, 14.20343, 15.15185, 16.09367, 17.02878, 17.95705, 18.87837, 
    19.79265, 20.69982, 21.59979, 22.49251, 23.37793, 24.256, 25.12669, 
    25.98999, 26.84588, 27.69435, 28.53541, 29.36907, 30.19535, 31.01428, 
    31.82589, 32.63021, 33.42731, 34.21722, 35,
  305, 305.7828, 306.5727, 307.3698, 308.1741, 308.9857, 309.8047, 310.6309, 
    311.4646, 312.3057, 313.1541, 314.01, 314.8733, 315.744, 316.6221, 
    317.5075, 318.4002, 319.3002, 320.2073, 321.1216, 322.043, 322.9712, 
    323.9063, 324.8481, 325.7966, 326.7514, 327.7126, 328.6799, 329.6532, 
    330.6322, 331.6168, 332.6068, 333.6019, 334.6019, 335.6065, 336.6156, 
    337.6287, 338.6458, 339.6663, 340.6902, 341.717, 342.7465, 343.7783, 
    344.8122, 345.8477, 346.8846, 347.9225, 348.9611, 350, 351.0389, 
    352.0775, 353.1154, 354.1523, 355.1878, 356.2217, 357.2535, 358.283, 
    359.3098, 0.3336662, 1.354252, 2.371273, 3.384442, 4.393482, 5.398128, 
    6.39812, 7.393215, 8.383177, 9.367781, 10.34682, 11.32008, 12.28739, 
    13.24856, 14.20343, 15.15185, 16.09367, 17.02878, 17.95705, 18.87837, 
    19.79265, 20.69982, 21.59979, 22.49251, 23.37793, 24.256, 25.12669, 
    25.98999, 26.84588, 27.69435, 28.53541, 29.36907, 30.19535, 31.01428, 
    31.82589, 32.63021, 33.42731, 34.21722, 35,
  305, 305.7828, 306.5727, 307.3698, 308.1741, 308.9857, 309.8047, 310.6309, 
    311.4646, 312.3057, 313.1541, 314.01, 314.8733, 315.744, 316.6221, 
    317.5075, 318.4002, 319.3002, 320.2073, 321.1216, 322.043, 322.9712, 
    323.9063, 324.8481, 325.7966, 326.7514, 327.7126, 328.6799, 329.6532, 
    330.6322, 331.6168, 332.6068, 333.6019, 334.6019, 335.6065, 336.6156, 
    337.6287, 338.6458, 339.6663, 340.6902, 341.717, 342.7465, 343.7783, 
    344.8122, 345.8477, 346.8846, 347.9225, 348.9611, 350, 351.0389, 
    352.0775, 353.1154, 354.1523, 355.1878, 356.2217, 357.2535, 358.283, 
    359.3098, 0.3336662, 1.354252, 2.371273, 3.384442, 4.393482, 5.398128, 
    6.39812, 7.393215, 8.383177, 9.367781, 10.34682, 11.32008, 12.28739, 
    13.24856, 14.20343, 15.15185, 16.09367, 17.02878, 17.95705, 18.87837, 
    19.79265, 20.69982, 21.59979, 22.49251, 23.37793, 24.256, 25.12669, 
    25.98999, 26.84588, 27.69435, 28.53541, 29.36907, 30.19535, 31.01428, 
    31.82589, 32.63021, 33.42731, 34.21722, 35,
  305, 305.7828, 306.5727, 307.3698, 308.1741, 308.9857, 309.8047, 310.6309, 
    311.4646, 312.3057, 313.1541, 314.01, 314.8733, 315.744, 316.6221, 
    317.5075, 318.4002, 319.3002, 320.2073, 321.1216, 322.043, 322.9712, 
    323.9063, 324.8481, 325.7966, 326.7514, 327.7126, 328.6799, 329.6532, 
    330.6322, 331.6168, 332.6068, 333.6019, 334.6019, 335.6065, 336.6156, 
    337.6287, 338.6458, 339.6663, 340.6902, 341.717, 342.7465, 343.7783, 
    344.8122, 345.8477, 346.8846, 347.9225, 348.9611, 350, 351.0389, 
    352.0775, 353.1154, 354.1523, 355.1878, 356.2217, 357.2535, 358.283, 
    359.3098, 0.3336662, 1.354252, 2.371273, 3.384442, 4.393482, 5.398128, 
    6.39812, 7.393215, 8.383177, 9.367781, 10.34682, 11.32008, 12.28739, 
    13.24856, 14.20343, 15.15185, 16.09367, 17.02878, 17.95705, 18.87837, 
    19.79265, 20.69982, 21.59979, 22.49251, 23.37793, 24.256, 25.12669, 
    25.98999, 26.84588, 27.69435, 28.53541, 29.36907, 30.19535, 31.01428, 
    31.82589, 32.63021, 33.42731, 34.21722, 35,
  305, 305.7828, 306.5727, 307.3698, 308.1741, 308.9857, 309.8047, 310.6309, 
    311.4646, 312.3057, 313.1541, 314.01, 314.8733, 315.744, 316.6221, 
    317.5075, 318.4002, 319.3002, 320.2073, 321.1216, 322.043, 322.9712, 
    323.9063, 324.8481, 325.7966, 326.7514, 327.7126, 328.6799, 329.6532, 
    330.6322, 331.6168, 332.6068, 333.6019, 334.6019, 335.6065, 336.6156, 
    337.6287, 338.6458, 339.6663, 340.6902, 341.717, 342.7465, 343.7783, 
    344.8122, 345.8477, 346.8846, 347.9225, 348.9611, 350, 351.0389, 
    352.0775, 353.1154, 354.1523, 355.1878, 356.2217, 357.2535, 358.283, 
    359.3098, 0.3336662, 1.354252, 2.371273, 3.384442, 4.393482, 5.398128, 
    6.39812, 7.393215, 8.383177, 9.367781, 10.34682, 11.32008, 12.28739, 
    13.24856, 14.20343, 15.15185, 16.09367, 17.02878, 17.95705, 18.87837, 
    19.79265, 20.69982, 21.59979, 22.49251, 23.37793, 24.256, 25.12669, 
    25.98999, 26.84588, 27.69435, 28.53541, 29.36907, 30.19535, 31.01428, 
    31.82589, 32.63021, 33.42731, 34.21722, 35,
  305, 305.7828, 306.5727, 307.3698, 308.1741, 308.9857, 309.8047, 310.6309, 
    311.4646, 312.3057, 313.1541, 314.01, 314.8733, 315.744, 316.6221, 
    317.5075, 318.4002, 319.3002, 320.2073, 321.1216, 322.043, 322.9712, 
    323.9063, 324.8481, 325.7966, 326.7514, 327.7126, 328.6799, 329.6532, 
    330.6322, 331.6168, 332.6068, 333.6019, 334.6019, 335.6065, 336.6156, 
    337.6287, 338.6458, 339.6663, 340.6902, 341.717, 342.7465, 343.7783, 
    344.8122, 345.8477, 346.8846, 347.9225, 348.9611, 350, 351.0389, 
    352.0775, 353.1154, 354.1523, 355.1878, 356.2217, 357.2535, 358.283, 
    359.3098, 0.3336662, 1.354252, 2.371273, 3.384442, 4.393482, 5.398128, 
    6.39812, 7.393215, 8.383177, 9.367781, 10.34682, 11.32008, 12.28739, 
    13.24856, 14.20343, 15.15185, 16.09367, 17.02878, 17.95705, 18.87837, 
    19.79265, 20.69982, 21.59979, 22.49251, 23.37793, 24.256, 25.12669, 
    25.98999, 26.84588, 27.69435, 28.53541, 29.36907, 30.19535, 31.01428, 
    31.82589, 32.63021, 33.42731, 34.21722, 35,
  305, 305.7828, 306.5727, 307.3698, 308.1741, 308.9857, 309.8047, 310.6309, 
    311.4646, 312.3057, 313.1541, 314.01, 314.8733, 315.744, 316.6221, 
    317.5075, 318.4002, 319.3002, 320.2073, 321.1216, 322.043, 322.9712, 
    323.9063, 324.8481, 325.7966, 326.7514, 327.7126, 328.6799, 329.6532, 
    330.6322, 331.6168, 332.6068, 333.6019, 334.6019, 335.6065, 336.6156, 
    337.6287, 338.6458, 339.6663, 340.6902, 341.717, 342.7465, 343.7783, 
    344.8122, 345.8477, 346.8846, 347.9225, 348.9611, 350, 351.0389, 
    352.0775, 353.1154, 354.1523, 355.1878, 356.2217, 357.2535, 358.283, 
    359.3098, 0.3336662, 1.354252, 2.371273, 3.384442, 4.393482, 5.398128, 
    6.39812, 7.393215, 8.383177, 9.367781, 10.34682, 11.32008, 12.28739, 
    13.24856, 14.20343, 15.15185, 16.09367, 17.02878, 17.95705, 18.87837, 
    19.79265, 20.69982, 21.59979, 22.49251, 23.37793, 24.256, 25.12669, 
    25.98999, 26.84588, 27.69435, 28.53541, 29.36907, 30.19535, 31.01428, 
    31.82589, 32.63021, 33.42731, 34.21722, 35,
  305, 305.7828, 306.5727, 307.3698, 308.1741, 308.9857, 309.8047, 310.6309, 
    311.4646, 312.3057, 313.1541, 314.01, 314.8733, 315.744, 316.6221, 
    317.5075, 318.4002, 319.3002, 320.2073, 321.1216, 322.043, 322.9712, 
    323.9063, 324.8481, 325.7966, 326.7514, 327.7126, 328.6799, 329.6532, 
    330.6322, 331.6168, 332.6068, 333.6019, 334.6019, 335.6065, 336.6156, 
    337.6287, 338.6458, 339.6663, 340.6902, 341.717, 342.7465, 343.7783, 
    344.8122, 345.8477, 346.8846, 347.9225, 348.9611, 350, 351.0389, 
    352.0775, 353.1154, 354.1523, 355.1878, 356.2217, 357.2535, 358.283, 
    359.3098, 0.3336662, 1.354252, 2.371273, 3.384442, 4.393482, 5.398128, 
    6.39812, 7.393215, 8.383177, 9.367781, 10.34682, 11.32008, 12.28739, 
    13.24856, 14.20343, 15.15185, 16.09367, 17.02878, 17.95705, 18.87837, 
    19.79265, 20.69982, 21.59979, 22.49251, 23.37793, 24.256, 25.12669, 
    25.98999, 26.84588, 27.69435, 28.53541, 29.36907, 30.19535, 31.01428, 
    31.82589, 32.63021, 33.42731, 34.21722, 35,
  305, 305.7828, 306.5727, 307.3698, 308.1741, 308.9857, 309.8047, 310.6309, 
    311.4646, 312.3057, 313.1541, 314.01, 314.8733, 315.744, 316.6221, 
    317.5075, 318.4002, 319.3002, 320.2073, 321.1216, 322.043, 322.9712, 
    323.9063, 324.8481, 325.7966, 326.7514, 327.7126, 328.6799, 329.6532, 
    330.6322, 331.6168, 332.6068, 333.6019, 334.6019, 335.6065, 336.6156, 
    337.6287, 338.6458, 339.6663, 340.6902, 341.717, 342.7465, 343.7783, 
    344.8122, 345.8477, 346.8846, 347.9225, 348.9611, 350, 351.0389, 
    352.0775, 353.1154, 354.1523, 355.1878, 356.2217, 357.2535, 358.283, 
    359.3098, 0.3336662, 1.354252, 2.371273, 3.384442, 4.393482, 5.398128, 
    6.39812, 7.393215, 8.383177, 9.367781, 10.34682, 11.32008, 12.28739, 
    13.24856, 14.20343, 15.15185, 16.09367, 17.02878, 17.95705, 18.87837, 
    19.79265, 20.69982, 21.59979, 22.49251, 23.37793, 24.256, 25.12669, 
    25.98999, 26.84588, 27.69435, 28.53541, 29.36907, 30.19535, 31.01428, 
    31.82589, 32.63021, 33.42731, 34.21722, 35,
  305, 305.7828, 306.5727, 307.3698, 308.1741, 308.9857, 309.8047, 310.6309, 
    311.4646, 312.3057, 313.1541, 314.01, 314.8733, 315.744, 316.6221, 
    317.5075, 318.4002, 319.3002, 320.2073, 321.1216, 322.043, 322.9712, 
    323.9063, 324.8481, 325.7966, 326.7514, 327.7126, 328.6799, 329.6532, 
    330.6322, 331.6168, 332.6068, 333.6019, 334.6019, 335.6065, 336.6156, 
    337.6287, 338.6458, 339.6663, 340.6902, 341.717, 342.7465, 343.7783, 
    344.8122, 345.8477, 346.8846, 347.9225, 348.9611, 350, 351.0389, 
    352.0775, 353.1154, 354.1523, 355.1878, 356.2217, 357.2535, 358.283, 
    359.3098, 0.3336662, 1.354252, 2.371273, 3.384442, 4.393482, 5.398128, 
    6.39812, 7.393215, 8.383177, 9.367781, 10.34682, 11.32008, 12.28739, 
    13.24856, 14.20343, 15.15185, 16.09367, 17.02878, 17.95705, 18.87837, 
    19.79265, 20.69982, 21.59979, 22.49251, 23.37793, 24.256, 25.12669, 
    25.98999, 26.84588, 27.69435, 28.53541, 29.36907, 30.19535, 31.01428, 
    31.82589, 32.63021, 33.42731, 34.21722, 35,
  305, 305.7828, 306.5727, 307.3698, 308.1741, 308.9857, 309.8047, 310.6309, 
    311.4646, 312.3057, 313.1541, 314.01, 314.8733, 315.744, 316.6221, 
    317.5075, 318.4002, 319.3002, 320.2073, 321.1216, 322.043, 322.9712, 
    323.9063, 324.8481, 325.7966, 326.7514, 327.7126, 328.6799, 329.6532, 
    330.6322, 331.6168, 332.6068, 333.6019, 334.6019, 335.6065, 336.6156, 
    337.6287, 338.6458, 339.6663, 340.6902, 341.717, 342.7465, 343.7783, 
    344.8122, 345.8477, 346.8846, 347.9225, 348.9611, 350, 351.0389, 
    352.0775, 353.1154, 354.1523, 355.1878, 356.2217, 357.2535, 358.283, 
    359.3098, 0.3336662, 1.354252, 2.371273, 3.384442, 4.393482, 5.398128, 
    6.39812, 7.393215, 8.383177, 9.367781, 10.34682, 11.32008, 12.28739, 
    13.24856, 14.20343, 15.15185, 16.09367, 17.02878, 17.95705, 18.87837, 
    19.79265, 20.69982, 21.59979, 22.49251, 23.37793, 24.256, 25.12669, 
    25.98999, 26.84588, 27.69435, 28.53541, 29.36907, 30.19535, 31.01428, 
    31.82589, 32.63021, 33.42731, 34.21722, 35,
  305, 305.7828, 306.5727, 307.3698, 308.1741, 308.9857, 309.8047, 310.6309, 
    311.4646, 312.3057, 313.1541, 314.01, 314.8733, 315.744, 316.6221, 
    317.5075, 318.4002, 319.3002, 320.2073, 321.1216, 322.043, 322.9712, 
    323.9063, 324.8481, 325.7966, 326.7514, 327.7126, 328.6799, 329.6532, 
    330.6322, 331.6168, 332.6068, 333.6019, 334.6019, 335.6065, 336.6156, 
    337.6287, 338.6458, 339.6663, 340.6902, 341.717, 342.7465, 343.7783, 
    344.8122, 345.8477, 346.8846, 347.9225, 348.9611, 350, 351.0389, 
    352.0775, 353.1154, 354.1523, 355.1878, 356.2217, 357.2535, 358.283, 
    359.3098, 0.3336662, 1.354252, 2.371273, 3.384442, 4.393482, 5.398128, 
    6.39812, 7.393215, 8.383177, 9.367781, 10.34682, 11.32008, 12.28739, 
    13.24856, 14.20343, 15.15185, 16.09367, 17.02878, 17.95705, 18.87837, 
    19.79265, 20.69982, 21.59979, 22.49251, 23.37793, 24.256, 25.12669, 
    25.98999, 26.84588, 27.69435, 28.53541, 29.36907, 30.19535, 31.01428, 
    31.82589, 32.63021, 33.42731, 34.21722, 35,
  305, 305.7828, 306.5727, 307.3698, 308.1741, 308.9857, 309.8047, 310.6309, 
    311.4646, 312.3057, 313.1541, 314.01, 314.8733, 315.744, 316.6221, 
    317.5075, 318.4002, 319.3002, 320.2073, 321.1216, 322.043, 322.9712, 
    323.9063, 324.8481, 325.7966, 326.7514, 327.7126, 328.6799, 329.6532, 
    330.6322, 331.6168, 332.6068, 333.6019, 334.6019, 335.6065, 336.6156, 
    337.6287, 338.6458, 339.6663, 340.6902, 341.717, 342.7465, 343.7783, 
    344.8122, 345.8477, 346.8846, 347.9225, 348.9611, 350, 351.0389, 
    352.0775, 353.1154, 354.1523, 355.1878, 356.2217, 357.2535, 358.283, 
    359.3098, 0.3336662, 1.354252, 2.371273, 3.384442, 4.393482, 5.398128, 
    6.39812, 7.393215, 8.383177, 9.367781, 10.34682, 11.32008, 12.28739, 
    13.24856, 14.20343, 15.15185, 16.09367, 17.02878, 17.95705, 18.87837, 
    19.79265, 20.69982, 21.59979, 22.49251, 23.37793, 24.256, 25.12669, 
    25.98999, 26.84588, 27.69435, 28.53541, 29.36907, 30.19535, 31.01428, 
    31.82589, 32.63021, 33.42731, 34.21722, 35,
  305, 305.7828, 306.5727, 307.3698, 308.1741, 308.9857, 309.8047, 310.6309, 
    311.4646, 312.3057, 313.1541, 314.01, 314.8733, 315.744, 316.6221, 
    317.5075, 318.4002, 319.3002, 320.2073, 321.1216, 322.043, 322.9712, 
    323.9063, 324.8481, 325.7966, 326.7514, 327.7126, 328.6799, 329.6532, 
    330.6322, 331.6168, 332.6068, 333.6019, 334.6019, 335.6065, 336.6156, 
    337.6287, 338.6458, 339.6663, 340.6902, 341.717, 342.7465, 343.7783, 
    344.8122, 345.8477, 346.8846, 347.9225, 348.9611, 350, 351.0389, 
    352.0775, 353.1154, 354.1523, 355.1878, 356.2217, 357.2535, 358.283, 
    359.3098, 0.3336662, 1.354252, 2.371273, 3.384442, 4.393482, 5.398128, 
    6.39812, 7.393215, 8.383177, 9.367781, 10.34682, 11.32008, 12.28739, 
    13.24856, 14.20343, 15.15185, 16.09367, 17.02878, 17.95705, 18.87837, 
    19.79265, 20.69982, 21.59979, 22.49251, 23.37793, 24.256, 25.12669, 
    25.98999, 26.84588, 27.69435, 28.53541, 29.36907, 30.19535, 31.01428, 
    31.82589, 32.63021, 33.42731, 34.21722, 35,
  305, 305.7828, 306.5727, 307.3698, 308.1741, 308.9857, 309.8047, 310.6309, 
    311.4646, 312.3057, 313.1541, 314.01, 314.8733, 315.744, 316.6221, 
    317.5075, 318.4002, 319.3002, 320.2073, 321.1216, 322.043, 322.9712, 
    323.9063, 324.8481, 325.7966, 326.7514, 327.7126, 328.6799, 329.6532, 
    330.6322, 331.6168, 332.6068, 333.6019, 334.6019, 335.6065, 336.6156, 
    337.6287, 338.6458, 339.6663, 340.6902, 341.717, 342.7465, 343.7783, 
    344.8122, 345.8477, 346.8846, 347.9225, 348.9611, 350, 351.0389, 
    352.0775, 353.1154, 354.1523, 355.1878, 356.2217, 357.2535, 358.283, 
    359.3098, 0.3336662, 1.354252, 2.371273, 3.384442, 4.393482, 5.398128, 
    6.39812, 7.393215, 8.383177, 9.367781, 10.34682, 11.32008, 12.28739, 
    13.24856, 14.20343, 15.15185, 16.09367, 17.02878, 17.95705, 18.87837, 
    19.79265, 20.69982, 21.59979, 22.49251, 23.37793, 24.256, 25.12669, 
    25.98999, 26.84588, 27.69435, 28.53541, 29.36907, 30.19535, 31.01428, 
    31.82589, 32.63021, 33.42731, 34.21722, 35,
  305, 305.7828, 306.5727, 307.3698, 308.1741, 308.9857, 309.8047, 310.6309, 
    311.4646, 312.3057, 313.1541, 314.01, 314.8733, 315.744, 316.6221, 
    317.5075, 318.4002, 319.3002, 320.2073, 321.1216, 322.043, 322.9712, 
    323.9063, 324.8481, 325.7966, 326.7514, 327.7126, 328.6799, 329.6532, 
    330.6322, 331.6168, 332.6068, 333.6019, 334.6019, 335.6065, 336.6156, 
    337.6287, 338.6458, 339.6663, 340.6902, 341.717, 342.7465, 343.7783, 
    344.8122, 345.8477, 346.8846, 347.9225, 348.9611, 350, 351.0389, 
    352.0775, 353.1154, 354.1523, 355.1878, 356.2217, 357.2535, 358.283, 
    359.3098, 0.3336662, 1.354252, 2.371273, 3.384442, 4.393482, 5.398128, 
    6.39812, 7.393215, 8.383177, 9.367781, 10.34682, 11.32008, 12.28739, 
    13.24856, 14.20343, 15.15185, 16.09367, 17.02878, 17.95705, 18.87837, 
    19.79265, 20.69982, 21.59979, 22.49251, 23.37793, 24.256, 25.12669, 
    25.98999, 26.84588, 27.69435, 28.53541, 29.36907, 30.19535, 31.01428, 
    31.82589, 32.63021, 33.42731, 34.21722, 35,
  305, 305.7828, 306.5727, 307.3698, 308.1741, 308.9857, 309.8047, 310.6309, 
    311.4646, 312.3057, 313.1541, 314.01, 314.8733, 315.744, 316.6221, 
    317.5075, 318.4002, 319.3002, 320.2073, 321.1216, 322.043, 322.9712, 
    323.9063, 324.8481, 325.7966, 326.7514, 327.7126, 328.6799, 329.6532, 
    330.6322, 331.6168, 332.6068, 333.6019, 334.6019, 335.6065, 336.6156, 
    337.6287, 338.6458, 339.6663, 340.6902, 341.717, 342.7465, 343.7783, 
    344.8122, 345.8477, 346.8846, 347.9225, 348.9611, 350, 351.0389, 
    352.0775, 353.1154, 354.1523, 355.1878, 356.2217, 357.2535, 358.283, 
    359.3098, 0.3336662, 1.354252, 2.371273, 3.384442, 4.393482, 5.398128, 
    6.39812, 7.393215, 8.383177, 9.367781, 10.34682, 11.32008, 12.28739, 
    13.24856, 14.20343, 15.15185, 16.09367, 17.02878, 17.95705, 18.87837, 
    19.79265, 20.69982, 21.59979, 22.49251, 23.37793, 24.256, 25.12669, 
    25.98999, 26.84588, 27.69435, 28.53541, 29.36907, 30.19535, 31.01428, 
    31.82589, 32.63021, 33.42731, 34.21722, 35,
  305, 305.7828, 306.5727, 307.3698, 308.1741, 308.9857, 309.8047, 310.6309, 
    311.4646, 312.3057, 313.1541, 314.01, 314.8733, 315.744, 316.6221, 
    317.5075, 318.4002, 319.3002, 320.2073, 321.1216, 322.043, 322.9712, 
    323.9063, 324.8481, 325.7966, 326.7514, 327.7126, 328.6799, 329.6532, 
    330.6322, 331.6168, 332.6068, 333.6019, 334.6019, 335.6065, 336.6156, 
    337.6287, 338.6458, 339.6663, 340.6902, 341.717, 342.7465, 343.7783, 
    344.8122, 345.8477, 346.8846, 347.9225, 348.9611, 350, 351.0389, 
    352.0775, 353.1154, 354.1523, 355.1878, 356.2217, 357.2535, 358.283, 
    359.3098, 0.3336662, 1.354252, 2.371273, 3.384442, 4.393482, 5.398128, 
    6.39812, 7.393215, 8.383177, 9.367781, 10.34682, 11.32008, 12.28739, 
    13.24856, 14.20343, 15.15185, 16.09367, 17.02878, 17.95705, 18.87837, 
    19.79265, 20.69982, 21.59979, 22.49251, 23.37793, 24.256, 25.12669, 
    25.98999, 26.84588, 27.69435, 28.53541, 29.36907, 30.19535, 31.01428, 
    31.82589, 32.63021, 33.42731, 34.21722, 35,
  305, 305.7828, 306.5727, 307.3698, 308.1741, 308.9857, 309.8047, 310.6309, 
    311.4646, 312.3057, 313.1541, 314.01, 314.8733, 315.744, 316.6221, 
    317.5075, 318.4002, 319.3002, 320.2073, 321.1216, 322.043, 322.9712, 
    323.9063, 324.8481, 325.7966, 326.7514, 327.7126, 328.6799, 329.6532, 
    330.6322, 331.6168, 332.6068, 333.6019, 334.6019, 335.6065, 336.6156, 
    337.6287, 338.6458, 339.6663, 340.6902, 341.717, 342.7465, 343.7783, 
    344.8122, 345.8477, 346.8846, 347.9225, 348.9611, 350, 351.0389, 
    352.0775, 353.1154, 354.1523, 355.1878, 356.2217, 357.2535, 358.283, 
    359.3098, 0.3336662, 1.354252, 2.371273, 3.384442, 4.393482, 5.398128, 
    6.39812, 7.393215, 8.383177, 9.367781, 10.34682, 11.32008, 12.28739, 
    13.24856, 14.20343, 15.15185, 16.09367, 17.02878, 17.95705, 18.87837, 
    19.79265, 20.69982, 21.59979, 22.49251, 23.37793, 24.256, 25.12669, 
    25.98999, 26.84588, 27.69435, 28.53541, 29.36907, 30.19535, 31.01428, 
    31.82589, 32.63021, 33.42731, 34.21722, 35,
  305, 305.7828, 306.5727, 307.3698, 308.1741, 308.9857, 309.8047, 310.6309, 
    311.4646, 312.3057, 313.1541, 314.01, 314.8733, 315.744, 316.6221, 
    317.5075, 318.4002, 319.3002, 320.2073, 321.1216, 322.043, 322.9712, 
    323.9063, 324.8481, 325.7966, 326.7514, 327.7126, 328.6799, 329.6532, 
    330.6322, 331.6168, 332.6068, 333.6019, 334.6019, 335.6065, 336.6156, 
    337.6287, 338.6458, 339.6663, 340.6902, 341.717, 342.7465, 343.7783, 
    344.8122, 345.8477, 346.8846, 347.9225, 348.9611, 350, 351.0389, 
    352.0775, 353.1154, 354.1523, 355.1878, 356.2217, 357.2535, 358.283, 
    359.3098, 0.3336662, 1.354252, 2.371273, 3.384442, 4.393482, 5.398128, 
    6.39812, 7.393215, 8.383177, 9.367781, 10.34682, 11.32008, 12.28739, 
    13.24856, 14.20343, 15.15185, 16.09367, 17.02878, 17.95705, 18.87837, 
    19.79265, 20.69982, 21.59979, 22.49251, 23.37793, 24.256, 25.12669, 
    25.98999, 26.84588, 27.69435, 28.53541, 29.36907, 30.19535, 31.01428, 
    31.82589, 32.63021, 33.42731, 34.21722, 35,
  305, 305.7828, 306.5727, 307.3698, 308.1741, 308.9857, 309.8047, 310.6309, 
    311.4646, 312.3057, 313.1541, 314.01, 314.8733, 315.744, 316.6221, 
    317.5075, 318.4002, 319.3002, 320.2073, 321.1216, 322.043, 322.9712, 
    323.9063, 324.8481, 325.7966, 326.7514, 327.7126, 328.6799, 329.6532, 
    330.6322, 331.6168, 332.6068, 333.6019, 334.6019, 335.6065, 336.6156, 
    337.6287, 338.6458, 339.6663, 340.6902, 341.717, 342.7465, 343.7783, 
    344.8122, 345.8477, 346.8846, 347.9225, 348.9611, 350, 351.0389, 
    352.0775, 353.1154, 354.1523, 355.1878, 356.2217, 357.2535, 358.283, 
    359.3098, 0.3336662, 1.354252, 2.371273, 3.384442, 4.393482, 5.398128, 
    6.39812, 7.393215, 8.383177, 9.367781, 10.34682, 11.32008, 12.28739, 
    13.24856, 14.20343, 15.15185, 16.09367, 17.02878, 17.95705, 18.87837, 
    19.79265, 20.69982, 21.59979, 22.49251, 23.37793, 24.256, 25.12669, 
    25.98999, 26.84588, 27.69435, 28.53541, 29.36907, 30.19535, 31.01428, 
    31.82589, 32.63021, 33.42731, 34.21722, 35,
  305, 305.7828, 306.5727, 307.3698, 308.1741, 308.9857, 309.8047, 310.6309, 
    311.4646, 312.3057, 313.1541, 314.01, 314.8733, 315.744, 316.6221, 
    317.5075, 318.4002, 319.3002, 320.2073, 321.1216, 322.043, 322.9712, 
    323.9063, 324.8481, 325.7966, 326.7514, 327.7126, 328.6799, 329.6532, 
    330.6322, 331.6168, 332.6068, 333.6019, 334.6019, 335.6065, 336.6156, 
    337.6287, 338.6458, 339.6663, 340.6902, 341.717, 342.7465, 343.7783, 
    344.8122, 345.8477, 346.8846, 347.9225, 348.9611, 350, 351.0389, 
    352.0775, 353.1154, 354.1523, 355.1878, 356.2217, 357.2535, 358.283, 
    359.3098, 0.3336662, 1.354252, 2.371273, 3.384442, 4.393482, 5.398128, 
    6.39812, 7.393215, 8.383177, 9.367781, 10.34682, 11.32008, 12.28739, 
    13.24856, 14.20343, 15.15185, 16.09367, 17.02878, 17.95705, 18.87837, 
    19.79265, 20.69982, 21.59979, 22.49251, 23.37793, 24.256, 25.12669, 
    25.98999, 26.84588, 27.69435, 28.53541, 29.36907, 30.19535, 31.01428, 
    31.82589, 32.63021, 33.42731, 34.21722, 35,
  305, 305.7828, 306.5727, 307.3698, 308.1741, 308.9857, 309.8047, 310.6309, 
    311.4646, 312.3057, 313.1541, 314.01, 314.8733, 315.744, 316.6221, 
    317.5075, 318.4002, 319.3002, 320.2073, 321.1216, 322.043, 322.9712, 
    323.9063, 324.8481, 325.7966, 326.7514, 327.7126, 328.6799, 329.6532, 
    330.6322, 331.6168, 332.6068, 333.6019, 334.6019, 335.6065, 336.6156, 
    337.6287, 338.6458, 339.6663, 340.6902, 341.717, 342.7465, 343.7783, 
    344.8122, 345.8477, 346.8846, 347.9225, 348.9611, 350, 351.0389, 
    352.0775, 353.1154, 354.1523, 355.1878, 356.2217, 357.2535, 358.283, 
    359.3098, 0.3336662, 1.354252, 2.371273, 3.384442, 4.393482, 5.398128, 
    6.39812, 7.393215, 8.383177, 9.367781, 10.34682, 11.32008, 12.28739, 
    13.24856, 14.20343, 15.15185, 16.09367, 17.02878, 17.95705, 18.87837, 
    19.79265, 20.69982, 21.59979, 22.49251, 23.37793, 24.256, 25.12669, 
    25.98999, 26.84588, 27.69435, 28.53541, 29.36907, 30.19535, 31.01428, 
    31.82589, 32.63021, 33.42731, 34.21722, 35,
  305, 305.7828, 306.5727, 307.3698, 308.1741, 308.9857, 309.8047, 310.6309, 
    311.4646, 312.3057, 313.1541, 314.01, 314.8733, 315.744, 316.6221, 
    317.5075, 318.4002, 319.3002, 320.2073, 321.1216, 322.043, 322.9712, 
    323.9063, 324.8481, 325.7966, 326.7514, 327.7126, 328.6799, 329.6532, 
    330.6322, 331.6168, 332.6068, 333.6019, 334.6019, 335.6065, 336.6156, 
    337.6287, 338.6458, 339.6663, 340.6902, 341.717, 342.7465, 343.7783, 
    344.8122, 345.8477, 346.8846, 347.9225, 348.9611, 350, 351.0389, 
    352.0775, 353.1154, 354.1523, 355.1878, 356.2217, 357.2535, 358.283, 
    359.3098, 0.3336662, 1.354252, 2.371273, 3.384442, 4.393482, 5.398128, 
    6.39812, 7.393215, 8.383177, 9.367781, 10.34682, 11.32008, 12.28739, 
    13.24856, 14.20343, 15.15185, 16.09367, 17.02878, 17.95705, 18.87837, 
    19.79265, 20.69982, 21.59979, 22.49251, 23.37793, 24.256, 25.12669, 
    25.98999, 26.84588, 27.69435, 28.53541, 29.36907, 30.19535, 31.01428, 
    31.82589, 32.63021, 33.42731, 34.21722, 35,
  305, 305.7828, 306.5727, 307.3698, 308.1741, 308.9857, 309.8047, 310.6309, 
    311.4646, 312.3057, 313.1541, 314.01, 314.8733, 315.744, 316.6221, 
    317.5075, 318.4002, 319.3002, 320.2073, 321.1216, 322.043, 322.9712, 
    323.9063, 324.8481, 325.7966, 326.7514, 327.7126, 328.6799, 329.6532, 
    330.6322, 331.6168, 332.6068, 333.6019, 334.6019, 335.6065, 336.6156, 
    337.6287, 338.6458, 339.6663, 340.6902, 341.717, 342.7465, 343.7783, 
    344.8122, 345.8477, 346.8846, 347.9225, 348.9611, 350, 351.0389, 
    352.0775, 353.1154, 354.1523, 355.1878, 356.2217, 357.2535, 358.283, 
    359.3098, 0.3336662, 1.354252, 2.371273, 3.384442, 4.393482, 5.398128, 
    6.39812, 7.393215, 8.383177, 9.367781, 10.34682, 11.32008, 12.28739, 
    13.24856, 14.20343, 15.15185, 16.09367, 17.02878, 17.95705, 18.87837, 
    19.79265, 20.69982, 21.59979, 22.49251, 23.37793, 24.256, 25.12669, 
    25.98999, 26.84588, 27.69435, 28.53541, 29.36907, 30.19535, 31.01428, 
    31.82589, 32.63021, 33.42731, 34.21722, 35,
  305, 305.7828, 306.5727, 307.3698, 308.1741, 308.9857, 309.8047, 310.6309, 
    311.4646, 312.3057, 313.1541, 314.01, 314.8733, 315.744, 316.6221, 
    317.5075, 318.4002, 319.3002, 320.2073, 321.1216, 322.043, 322.9712, 
    323.9063, 324.8481, 325.7966, 326.7514, 327.7126, 328.6799, 329.6532, 
    330.6322, 331.6168, 332.6068, 333.6019, 334.6019, 335.6065, 336.6156, 
    337.6287, 338.6458, 339.6663, 340.6902, 341.717, 342.7465, 343.7783, 
    344.8122, 345.8477, 346.8846, 347.9225, 348.9611, 350, 351.0389, 
    352.0775, 353.1154, 354.1523, 355.1878, 356.2217, 357.2535, 358.283, 
    359.3098, 0.3336662, 1.354252, 2.371273, 3.384442, 4.393482, 5.398128, 
    6.39812, 7.393215, 8.383177, 9.367781, 10.34682, 11.32008, 12.28739, 
    13.24856, 14.20343, 15.15185, 16.09367, 17.02878, 17.95705, 18.87837, 
    19.79265, 20.69982, 21.59979, 22.49251, 23.37793, 24.256, 25.12669, 
    25.98999, 26.84588, 27.69435, 28.53541, 29.36907, 30.19535, 31.01428, 
    31.82589, 32.63021, 33.42731, 34.21722, 35,
  305, 305.7828, 306.5727, 307.3698, 308.1741, 308.9857, 309.8047, 310.6309, 
    311.4646, 312.3057, 313.1541, 314.01, 314.8733, 315.744, 316.6221, 
    317.5075, 318.4002, 319.3002, 320.2073, 321.1216, 322.043, 322.9712, 
    323.9063, 324.8481, 325.7966, 326.7514, 327.7126, 328.6799, 329.6532, 
    330.6322, 331.6168, 332.6068, 333.6019, 334.6019, 335.6065, 336.6156, 
    337.6287, 338.6458, 339.6663, 340.6902, 341.717, 342.7465, 343.7783, 
    344.8122, 345.8477, 346.8846, 347.9225, 348.9611, 350, 351.0389, 
    352.0775, 353.1154, 354.1523, 355.1878, 356.2217, 357.2535, 358.283, 
    359.3098, 0.3336662, 1.354252, 2.371273, 3.384442, 4.393482, 5.398128, 
    6.39812, 7.393215, 8.383177, 9.367781, 10.34682, 11.32008, 12.28739, 
    13.24856, 14.20343, 15.15185, 16.09367, 17.02878, 17.95705, 18.87837, 
    19.79265, 20.69982, 21.59979, 22.49251, 23.37793, 24.256, 25.12669, 
    25.98999, 26.84588, 27.69435, 28.53541, 29.36907, 30.19535, 31.01428, 
    31.82589, 32.63021, 33.42731, 34.21722, 35,
  305, 305.7828, 306.5727, 307.3698, 308.1741, 308.9857, 309.8047, 310.6309, 
    311.4646, 312.3057, 313.1541, 314.01, 314.8733, 315.744, 316.6221, 
    317.5075, 318.4002, 319.3002, 320.2073, 321.1216, 322.043, 322.9712, 
    323.9063, 324.8481, 325.7966, 326.7514, 327.7126, 328.6799, 329.6532, 
    330.6322, 331.6168, 332.6068, 333.6019, 334.6019, 335.6065, 336.6156, 
    337.6287, 338.6458, 339.6663, 340.6902, 341.717, 342.7465, 343.7783, 
    344.8122, 345.8477, 346.8846, 347.9225, 348.9611, 350, 351.0389, 
    352.0775, 353.1154, 354.1523, 355.1878, 356.2217, 357.2535, 358.283, 
    359.3098, 0.3336662, 1.354252, 2.371273, 3.384442, 4.393482, 5.398128, 
    6.39812, 7.393215, 8.383177, 9.367781, 10.34682, 11.32008, 12.28739, 
    13.24856, 14.20343, 15.15185, 16.09367, 17.02878, 17.95705, 18.87837, 
    19.79265, 20.69982, 21.59979, 22.49251, 23.37793, 24.256, 25.12669, 
    25.98999, 26.84588, 27.69435, 28.53541, 29.36907, 30.19535, 31.01428, 
    31.82589, 32.63021, 33.42731, 34.21722, 35,
  305, 305.7828, 306.5727, 307.3698, 308.1741, 308.9857, 309.8047, 310.6309, 
    311.4646, 312.3057, 313.1541, 314.01, 314.8733, 315.744, 316.6221, 
    317.5075, 318.4002, 319.3002, 320.2073, 321.1216, 322.043, 322.9712, 
    323.9063, 324.8481, 325.7966, 326.7514, 327.7126, 328.6799, 329.6532, 
    330.6322, 331.6168, 332.6068, 333.6019, 334.6019, 335.6065, 336.6156, 
    337.6287, 338.6458, 339.6663, 340.6902, 341.717, 342.7465, 343.7783, 
    344.8122, 345.8477, 346.8846, 347.9225, 348.9611, 350, 351.0389, 
    352.0775, 353.1154, 354.1523, 355.1878, 356.2217, 357.2535, 358.283, 
    359.3098, 0.3336662, 1.354252, 2.371273, 3.384442, 4.393482, 5.398128, 
    6.39812, 7.393215, 8.383177, 9.367781, 10.34682, 11.32008, 12.28739, 
    13.24856, 14.20343, 15.15185, 16.09367, 17.02878, 17.95705, 18.87837, 
    19.79265, 20.69982, 21.59979, 22.49251, 23.37793, 24.256, 25.12669, 
    25.98999, 26.84588, 27.69435, 28.53541, 29.36907, 30.19535, 31.01428, 
    31.82589, 32.63021, 33.42731, 34.21722, 35,
  305, 305.7828, 306.5727, 307.3698, 308.1741, 308.9857, 309.8047, 310.6309, 
    311.4646, 312.3057, 313.1541, 314.01, 314.8733, 315.744, 316.6221, 
    317.5075, 318.4002, 319.3002, 320.2073, 321.1216, 322.043, 322.9712, 
    323.9063, 324.8481, 325.7966, 326.7514, 327.7126, 328.6799, 329.6532, 
    330.6322, 331.6168, 332.6068, 333.6019, 334.6019, 335.6065, 336.6156, 
    337.6287, 338.6458, 339.6663, 340.6902, 341.717, 342.7465, 343.7783, 
    344.8122, 345.8477, 346.8846, 347.9225, 348.9611, 350, 351.0389, 
    352.0775, 353.1154, 354.1523, 355.1878, 356.2217, 357.2535, 358.283, 
    359.3098, 0.3336662, 1.354252, 2.371273, 3.384442, 4.393482, 5.398128, 
    6.39812, 7.393215, 8.383177, 9.367781, 10.34682, 11.32008, 12.28739, 
    13.24856, 14.20343, 15.15185, 16.09367, 17.02878, 17.95705, 18.87837, 
    19.79265, 20.69982, 21.59979, 22.49251, 23.37793, 24.256, 25.12669, 
    25.98999, 26.84588, 27.69435, 28.53541, 29.36907, 30.19535, 31.01428, 
    31.82589, 32.63021, 33.42731, 34.21722, 35,
  305, 305.7828, 306.5727, 307.3698, 308.1741, 308.9857, 309.8047, 310.6309, 
    311.4646, 312.3057, 313.1541, 314.01, 314.8733, 315.744, 316.6221, 
    317.5075, 318.4002, 319.3002, 320.2073, 321.1216, 322.043, 322.9712, 
    323.9063, 324.8481, 325.7966, 326.7514, 327.7126, 328.6799, 329.6532, 
    330.6322, 331.6168, 332.6068, 333.6019, 334.6019, 335.6065, 336.6156, 
    337.6287, 338.6458, 339.6663, 340.6902, 341.717, 342.7465, 343.7783, 
    344.8122, 345.8477, 346.8846, 347.9225, 348.9611, 350, 351.0389, 
    352.0775, 353.1154, 354.1523, 355.1878, 356.2217, 357.2535, 358.283, 
    359.3098, 0.3336662, 1.354252, 2.371273, 3.384442, 4.393482, 5.398128, 
    6.39812, 7.393215, 8.383177, 9.367781, 10.34682, 11.32008, 12.28739, 
    13.24856, 14.20343, 15.15185, 16.09367, 17.02878, 17.95705, 18.87837, 
    19.79265, 20.69982, 21.59979, 22.49251, 23.37793, 24.256, 25.12669, 
    25.98999, 26.84588, 27.69435, 28.53541, 29.36907, 30.19535, 31.01428, 
    31.82589, 32.63021, 33.42731, 34.21722, 35,
  305, 305.7828, 306.5727, 307.3698, 308.1741, 308.9857, 309.8047, 310.6309, 
    311.4646, 312.3057, 313.1541, 314.01, 314.8733, 315.744, 316.6221, 
    317.5075, 318.4002, 319.3002, 320.2073, 321.1216, 322.043, 322.9712, 
    323.9063, 324.8481, 325.7966, 326.7514, 327.7126, 328.6799, 329.6532, 
    330.6322, 331.6168, 332.6068, 333.6019, 334.6019, 335.6065, 336.6156, 
    337.6287, 338.6458, 339.6663, 340.6902, 341.717, 342.7465, 343.7783, 
    344.8122, 345.8477, 346.8846, 347.9225, 348.9611, 350, 351.0389, 
    352.0775, 353.1154, 354.1523, 355.1878, 356.2217, 357.2535, 358.283, 
    359.3098, 0.3336662, 1.354252, 2.371273, 3.384442, 4.393482, 5.398128, 
    6.39812, 7.393215, 8.383177, 9.367781, 10.34682, 11.32008, 12.28739, 
    13.24856, 14.20343, 15.15185, 16.09367, 17.02878, 17.95705, 18.87837, 
    19.79265, 20.69982, 21.59979, 22.49251, 23.37793, 24.256, 25.12669, 
    25.98999, 26.84588, 27.69435, 28.53541, 29.36907, 30.19535, 31.01428, 
    31.82589, 32.63021, 33.42731, 34.21722, 35,
  305, 305.7828, 306.5727, 307.3698, 308.1741, 308.9857, 309.8047, 310.6309, 
    311.4646, 312.3057, 313.1541, 314.01, 314.8733, 315.744, 316.6221, 
    317.5075, 318.4002, 319.3002, 320.2073, 321.1216, 322.043, 322.9712, 
    323.9063, 324.8481, 325.7966, 326.7514, 327.7126, 328.6799, 329.6532, 
    330.6322, 331.6168, 332.6068, 333.6019, 334.6019, 335.6065, 336.6156, 
    337.6287, 338.6458, 339.6663, 340.6902, 341.717, 342.7465, 343.7783, 
    344.8122, 345.8477, 346.8846, 347.9225, 348.9611, 350, 351.0389, 
    352.0775, 353.1154, 354.1523, 355.1878, 356.2217, 357.2535, 358.283, 
    359.3098, 0.3336662, 1.354252, 2.371273, 3.384442, 4.393482, 5.398128, 
    6.39812, 7.393215, 8.383177, 9.367781, 10.34682, 11.32008, 12.28739, 
    13.24856, 14.20343, 15.15185, 16.09367, 17.02878, 17.95705, 18.87837, 
    19.79265, 20.69982, 21.59979, 22.49251, 23.37793, 24.256, 25.12669, 
    25.98999, 26.84588, 27.69435, 28.53541, 29.36907, 30.19535, 31.01428, 
    31.82589, 32.63021, 33.42731, 34.21722, 35,
  305, 305.7828, 306.5727, 307.3698, 308.1741, 308.9857, 309.8047, 310.6309, 
    311.4646, 312.3057, 313.1541, 314.01, 314.8733, 315.744, 316.6221, 
    317.5075, 318.4002, 319.3002, 320.2073, 321.1216, 322.043, 322.9712, 
    323.9063, 324.8481, 325.7966, 326.7514, 327.7126, 328.6799, 329.6532, 
    330.6322, 331.6168, 332.6068, 333.6019, 334.6019, 335.6065, 336.6156, 
    337.6287, 338.6458, 339.6663, 340.6902, 341.717, 342.7465, 343.7783, 
    344.8122, 345.8477, 346.8846, 347.9225, 348.9611, 350, 351.0389, 
    352.0775, 353.1154, 354.1523, 355.1878, 356.2217, 357.2535, 358.283, 
    359.3098, 0.3336662, 1.354252, 2.371273, 3.384442, 4.393482, 5.398128, 
    6.39812, 7.393215, 8.383177, 9.367781, 10.34682, 11.32008, 12.28739, 
    13.24856, 14.20343, 15.15185, 16.09367, 17.02878, 17.95705, 18.87837, 
    19.79265, 20.69982, 21.59979, 22.49251, 23.37793, 24.256, 25.12669, 
    25.98999, 26.84588, 27.69435, 28.53541, 29.36907, 30.19535, 31.01428, 
    31.82589, 32.63021, 33.42731, 34.21722, 35,
  305, 305.7828, 306.5727, 307.3698, 308.1741, 308.9857, 309.8047, 310.6309, 
    311.4646, 312.3057, 313.1541, 314.01, 314.8733, 315.744, 316.6221, 
    317.5075, 318.4002, 319.3002, 320.2073, 321.1216, 322.043, 322.9712, 
    323.9063, 324.8481, 325.7966, 326.7514, 327.7126, 328.6799, 329.6532, 
    330.6322, 331.6168, 332.6068, 333.6019, 334.6019, 335.6065, 336.6156, 
    337.6287, 338.6458, 339.6663, 340.6902, 341.717, 342.7465, 343.7783, 
    344.8122, 345.8477, 346.8846, 347.9225, 348.9611, 350, 351.0389, 
    352.0775, 353.1154, 354.1523, 355.1878, 356.2217, 357.2535, 358.283, 
    359.3098, 0.3336662, 1.354252, 2.371273, 3.384442, 4.393482, 5.398128, 
    6.39812, 7.393215, 8.383177, 9.367781, 10.34682, 11.32008, 12.28739, 
    13.24856, 14.20343, 15.15185, 16.09367, 17.02878, 17.95705, 18.87837, 
    19.79265, 20.69982, 21.59979, 22.49251, 23.37793, 24.256, 25.12669, 
    25.98999, 26.84588, 27.69435, 28.53541, 29.36907, 30.19535, 31.01428, 
    31.82589, 32.63021, 33.42731, 34.21722, 35,
  305, 305.7828, 306.5727, 307.3698, 308.1741, 308.9857, 309.8047, 310.6309, 
    311.4646, 312.3057, 313.1541, 314.01, 314.8733, 315.744, 316.6221, 
    317.5075, 318.4002, 319.3002, 320.2073, 321.1216, 322.043, 322.9712, 
    323.9063, 324.8481, 325.7966, 326.7514, 327.7126, 328.6799, 329.6532, 
    330.6322, 331.6168, 332.6068, 333.6019, 334.6019, 335.6065, 336.6156, 
    337.6287, 338.6458, 339.6663, 340.6902, 341.717, 342.7465, 343.7783, 
    344.8122, 345.8477, 346.8846, 347.9225, 348.9611, 350, 351.0389, 
    352.0775, 353.1154, 354.1523, 355.1878, 356.2217, 357.2535, 358.283, 
    359.3098, 0.3336662, 1.354252, 2.371273, 3.384442, 4.393482, 5.398128, 
    6.39812, 7.393215, 8.383177, 9.367781, 10.34682, 11.32008, 12.28739, 
    13.24856, 14.20343, 15.15185, 16.09367, 17.02878, 17.95705, 18.87837, 
    19.79265, 20.69982, 21.59979, 22.49251, 23.37793, 24.256, 25.12669, 
    25.98999, 26.84588, 27.69435, 28.53541, 29.36907, 30.19535, 31.01428, 
    31.82589, 32.63021, 33.42731, 34.21722, 35,
  305, 305.7828, 306.5727, 307.3698, 308.1741, 308.9857, 309.8047, 310.6309, 
    311.4646, 312.3057, 313.1541, 314.01, 314.8733, 315.744, 316.6221, 
    317.5075, 318.4002, 319.3002, 320.2073, 321.1216, 322.043, 322.9712, 
    323.9063, 324.8481, 325.7966, 326.7514, 327.7126, 328.6799, 329.6532, 
    330.6322, 331.6168, 332.6068, 333.6019, 334.6019, 335.6065, 336.6156, 
    337.6287, 338.6458, 339.6663, 340.6902, 341.717, 342.7465, 343.7783, 
    344.8122, 345.8477, 346.8846, 347.9225, 348.9611, 350, 351.0389, 
    352.0775, 353.1154, 354.1523, 355.1878, 356.2217, 357.2535, 358.283, 
    359.3098, 0.3336662, 1.354252, 2.371273, 3.384442, 4.393482, 5.398128, 
    6.39812, 7.393215, 8.383177, 9.367781, 10.34682, 11.32008, 12.28739, 
    13.24856, 14.20343, 15.15185, 16.09367, 17.02878, 17.95705, 18.87837, 
    19.79265, 20.69982, 21.59979, 22.49251, 23.37793, 24.256, 25.12669, 
    25.98999, 26.84588, 27.69435, 28.53541, 29.36907, 30.19535, 31.01428, 
    31.82589, 32.63021, 33.42731, 34.21722, 35,
  305, 305.7828, 306.5727, 307.3698, 308.1741, 308.9857, 309.8047, 310.6309, 
    311.4646, 312.3057, 313.1541, 314.01, 314.8733, 315.744, 316.6221, 
    317.5075, 318.4002, 319.3002, 320.2073, 321.1216, 322.043, 322.9712, 
    323.9063, 324.8481, 325.7966, 326.7514, 327.7126, 328.6799, 329.6532, 
    330.6322, 331.6168, 332.6068, 333.6019, 334.6019, 335.6065, 336.6156, 
    337.6287, 338.6458, 339.6663, 340.6902, 341.717, 342.7465, 343.7783, 
    344.8122, 345.8477, 346.8846, 347.9225, 348.9611, 350, 351.0389, 
    352.0775, 353.1154, 354.1523, 355.1878, 356.2217, 357.2535, 358.283, 
    359.3098, 0.3336662, 1.354252, 2.371273, 3.384442, 4.393482, 5.398128, 
    6.39812, 7.393215, 8.383177, 9.367781, 10.34682, 11.32008, 12.28739, 
    13.24856, 14.20343, 15.15185, 16.09367, 17.02878, 17.95705, 18.87837, 
    19.79265, 20.69982, 21.59979, 22.49251, 23.37793, 24.256, 25.12669, 
    25.98999, 26.84588, 27.69435, 28.53541, 29.36907, 30.19535, 31.01428, 
    31.82589, 32.63021, 33.42731, 34.21722, 35,
  305, 305.7828, 306.5727, 307.3698, 308.1741, 308.9857, 309.8047, 310.6309, 
    311.4646, 312.3057, 313.1541, 314.01, 314.8733, 315.744, 316.6221, 
    317.5075, 318.4002, 319.3002, 320.2073, 321.1216, 322.043, 322.9712, 
    323.9063, 324.8481, 325.7966, 326.7514, 327.7126, 328.6799, 329.6532, 
    330.6322, 331.6168, 332.6068, 333.6019, 334.6019, 335.6065, 336.6156, 
    337.6287, 338.6458, 339.6663, 340.6902, 341.717, 342.7465, 343.7783, 
    344.8122, 345.8477, 346.8846, 347.9225, 348.9611, 350, 351.0389, 
    352.0775, 353.1154, 354.1523, 355.1878, 356.2217, 357.2535, 358.283, 
    359.3098, 0.3336662, 1.354252, 2.371273, 3.384442, 4.393482, 5.398128, 
    6.39812, 7.393215, 8.383177, 9.367781, 10.34682, 11.32008, 12.28739, 
    13.24856, 14.20343, 15.15185, 16.09367, 17.02878, 17.95705, 18.87837, 
    19.79265, 20.69982, 21.59979, 22.49251, 23.37793, 24.256, 25.12669, 
    25.98999, 26.84588, 27.69435, 28.53541, 29.36907, 30.19535, 31.01428, 
    31.82589, 32.63021, 33.42731, 34.21722, 35,
  305, 305.7828, 306.5727, 307.3698, 308.1741, 308.9857, 309.8047, 310.6309, 
    311.4646, 312.3057, 313.1541, 314.01, 314.8733, 315.744, 316.6221, 
    317.5075, 318.4002, 319.3002, 320.2073, 321.1216, 322.043, 322.9712, 
    323.9063, 324.8481, 325.7966, 326.7514, 327.7126, 328.6799, 329.6532, 
    330.6322, 331.6168, 332.6068, 333.6019, 334.6019, 335.6065, 336.6156, 
    337.6287, 338.6458, 339.6663, 340.6902, 341.717, 342.7465, 343.7783, 
    344.8122, 345.8477, 346.8846, 347.9225, 348.9611, 350, 351.0389, 
    352.0775, 353.1154, 354.1523, 355.1878, 356.2217, 357.2535, 358.283, 
    359.3098, 0.3336662, 1.354252, 2.371273, 3.384442, 4.393482, 5.398128, 
    6.39812, 7.393215, 8.383177, 9.367781, 10.34682, 11.32008, 12.28739, 
    13.24856, 14.20343, 15.15185, 16.09367, 17.02878, 17.95705, 18.87837, 
    19.79265, 20.69982, 21.59979, 22.49251, 23.37793, 24.256, 25.12669, 
    25.98999, 26.84588, 27.69435, 28.53541, 29.36907, 30.19535, 31.01428, 
    31.82589, 32.63021, 33.42731, 34.21722, 35,
  305, 305.7828, 306.5727, 307.3698, 308.1741, 308.9857, 309.8047, 310.6309, 
    311.4646, 312.3057, 313.1541, 314.01, 314.8733, 315.744, 316.6221, 
    317.5075, 318.4002, 319.3002, 320.2073, 321.1216, 322.043, 322.9712, 
    323.9063, 324.8481, 325.7966, 326.7514, 327.7126, 328.6799, 329.6532, 
    330.6322, 331.6168, 332.6068, 333.6019, 334.6019, 335.6065, 336.6156, 
    337.6287, 338.6458, 339.6663, 340.6902, 341.717, 342.7465, 343.7783, 
    344.8122, 345.8477, 346.8846, 347.9225, 348.9611, 350, 351.0389, 
    352.0775, 353.1154, 354.1523, 355.1878, 356.2217, 357.2535, 358.283, 
    359.3098, 0.3336662, 1.354252, 2.371273, 3.384442, 4.393482, 5.398128, 
    6.39812, 7.393215, 8.383177, 9.367781, 10.34682, 11.32008, 12.28739, 
    13.24856, 14.20343, 15.15185, 16.09367, 17.02878, 17.95705, 18.87837, 
    19.79265, 20.69982, 21.59979, 22.49251, 23.37793, 24.256, 25.12669, 
    25.98999, 26.84588, 27.69435, 28.53541, 29.36907, 30.19535, 31.01428, 
    31.82589, 32.63021, 33.42731, 34.21722, 35,
  305, 305.7828, 306.5727, 307.3698, 308.1741, 308.9857, 309.8047, 310.6309, 
    311.4646, 312.3057, 313.1541, 314.01, 314.8733, 315.744, 316.6221, 
    317.5075, 318.4002, 319.3002, 320.2073, 321.1216, 322.043, 322.9712, 
    323.9063, 324.8481, 325.7966, 326.7514, 327.7126, 328.6799, 329.6532, 
    330.6322, 331.6168, 332.6068, 333.6019, 334.6019, 335.6065, 336.6156, 
    337.6287, 338.6458, 339.6663, 340.6902, 341.717, 342.7465, 343.7783, 
    344.8122, 345.8477, 346.8846, 347.9225, 348.9611, 350, 351.0389, 
    352.0775, 353.1154, 354.1523, 355.1878, 356.2217, 357.2535, 358.283, 
    359.3098, 0.3336662, 1.354252, 2.371273, 3.384442, 4.393482, 5.398128, 
    6.39812, 7.393215, 8.383177, 9.367781, 10.34682, 11.32008, 12.28739, 
    13.24856, 14.20343, 15.15185, 16.09367, 17.02878, 17.95705, 18.87837, 
    19.79265, 20.69982, 21.59979, 22.49251, 23.37793, 24.256, 25.12669, 
    25.98999, 26.84588, 27.69435, 28.53541, 29.36907, 30.19535, 31.01428, 
    31.82589, 32.63021, 33.42731, 34.21722, 35,
  305, 305.7828, 306.5727, 307.3698, 308.1741, 308.9857, 309.8047, 310.6309, 
    311.4646, 312.3057, 313.1541, 314.01, 314.8733, 315.744, 316.6221, 
    317.5075, 318.4002, 319.3002, 320.2073, 321.1216, 322.043, 322.9712, 
    323.9063, 324.8481, 325.7966, 326.7514, 327.7126, 328.6799, 329.6532, 
    330.6322, 331.6168, 332.6068, 333.6019, 334.6019, 335.6065, 336.6156, 
    337.6287, 338.6458, 339.6663, 340.6902, 341.717, 342.7465, 343.7783, 
    344.8122, 345.8477, 346.8846, 347.9225, 348.9611, 350, 351.0389, 
    352.0775, 353.1154, 354.1523, 355.1878, 356.2217, 357.2535, 358.283, 
    359.3098, 0.3336662, 1.354252, 2.371273, 3.384442, 4.393482, 5.398128, 
    6.39812, 7.393215, 8.383177, 9.367781, 10.34682, 11.32008, 12.28739, 
    13.24856, 14.20343, 15.15185, 16.09367, 17.02878, 17.95705, 18.87837, 
    19.79265, 20.69982, 21.59979, 22.49251, 23.37793, 24.256, 25.12669, 
    25.98999, 26.84588, 27.69435, 28.53541, 29.36907, 30.19535, 31.01428, 
    31.82589, 32.63021, 33.42731, 34.21722, 35,
  305, 305.7828, 306.5727, 307.3698, 308.1741, 308.9857, 309.8047, 310.6309, 
    311.4646, 312.3057, 313.1541, 314.01, 314.8733, 315.744, 316.6221, 
    317.5075, 318.4002, 319.3002, 320.2073, 321.1216, 322.043, 322.9712, 
    323.9063, 324.8481, 325.7966, 326.7514, 327.7126, 328.6799, 329.6532, 
    330.6322, 331.6168, 332.6068, 333.6019, 334.6019, 335.6065, 336.6156, 
    337.6287, 338.6458, 339.6663, 340.6902, 341.717, 342.7465, 343.7783, 
    344.8122, 345.8477, 346.8846, 347.9225, 348.9611, 350, 351.0389, 
    352.0775, 353.1154, 354.1523, 355.1878, 356.2217, 357.2535, 358.283, 
    359.3098, 0.3336662, 1.354252, 2.371273, 3.384442, 4.393482, 5.398128, 
    6.39812, 7.393215, 8.383177, 9.367781, 10.34682, 11.32008, 12.28739, 
    13.24856, 14.20343, 15.15185, 16.09367, 17.02878, 17.95705, 18.87837, 
    19.79265, 20.69982, 21.59979, 22.49251, 23.37793, 24.256, 25.12669, 
    25.98999, 26.84588, 27.69435, 28.53541, 29.36907, 30.19535, 31.01428, 
    31.82589, 32.63021, 33.42731, 34.21722, 35,
  305, 305.7828, 306.5727, 307.3698, 308.1741, 308.9857, 309.8047, 310.6309, 
    311.4646, 312.3057, 313.1541, 314.01, 314.8733, 315.744, 316.6221, 
    317.5075, 318.4002, 319.3002, 320.2073, 321.1216, 322.043, 322.9712, 
    323.9063, 324.8481, 325.7966, 326.7514, 327.7126, 328.6799, 329.6532, 
    330.6322, 331.6168, 332.6068, 333.6019, 334.6019, 335.6065, 336.6156, 
    337.6287, 338.6458, 339.6663, 340.6902, 341.717, 342.7465, 343.7783, 
    344.8122, 345.8477, 346.8846, 347.9225, 348.9611, 350, 351.0389, 
    352.0775, 353.1154, 354.1523, 355.1878, 356.2217, 357.2535, 358.283, 
    359.3098, 0.3336662, 1.354252, 2.371273, 3.384442, 4.393482, 5.398128, 
    6.39812, 7.393215, 8.383177, 9.367781, 10.34682, 11.32008, 12.28739, 
    13.24856, 14.20343, 15.15185, 16.09367, 17.02878, 17.95705, 18.87837, 
    19.79265, 20.69982, 21.59979, 22.49251, 23.37793, 24.256, 25.12669, 
    25.98999, 26.84588, 27.69435, 28.53541, 29.36907, 30.19535, 31.01428, 
    31.82589, 32.63021, 33.42731, 34.21722, 35,
  305, 305.7828, 306.5727, 307.3698, 308.1741, 308.9857, 309.8047, 310.6309, 
    311.4646, 312.3057, 313.1541, 314.01, 314.8733, 315.744, 316.6221, 
    317.5075, 318.4002, 319.3002, 320.2073, 321.1216, 322.043, 322.9712, 
    323.9063, 324.8481, 325.7966, 326.7514, 327.7126, 328.6799, 329.6532, 
    330.6322, 331.6168, 332.6068, 333.6019, 334.6019, 335.6065, 336.6156, 
    337.6287, 338.6458, 339.6663, 340.6902, 341.717, 342.7465, 343.7783, 
    344.8122, 345.8477, 346.8846, 347.9225, 348.9611, 350, 351.0389, 
    352.0775, 353.1154, 354.1523, 355.1878, 356.2217, 357.2535, 358.283, 
    359.3098, 0.3336662, 1.354252, 2.371273, 3.384442, 4.393482, 5.398128, 
    6.39812, 7.393215, 8.383177, 9.367781, 10.34682, 11.32008, 12.28739, 
    13.24856, 14.20343, 15.15185, 16.09367, 17.02878, 17.95705, 18.87837, 
    19.79265, 20.69982, 21.59979, 22.49251, 23.37793, 24.256, 25.12669, 
    25.98999, 26.84588, 27.69435, 28.53541, 29.36907, 30.19535, 31.01428, 
    31.82589, 32.63021, 33.42731, 34.21722, 35,
  305, 305.7828, 306.5727, 307.3698, 308.1741, 308.9857, 309.8047, 310.6309, 
    311.4646, 312.3057, 313.1541, 314.01, 314.8733, 315.744, 316.6221, 
    317.5075, 318.4002, 319.3002, 320.2073, 321.1216, 322.043, 322.9712, 
    323.9063, 324.8481, 325.7966, 326.7514, 327.7126, 328.6799, 329.6532, 
    330.6322, 331.6168, 332.6068, 333.6019, 334.6019, 335.6065, 336.6156, 
    337.6287, 338.6458, 339.6663, 340.6902, 341.717, 342.7465, 343.7783, 
    344.8122, 345.8477, 346.8846, 347.9225, 348.9611, 350, 351.0389, 
    352.0775, 353.1154, 354.1523, 355.1878, 356.2217, 357.2535, 358.283, 
    359.3098, 0.3336662, 1.354252, 2.371273, 3.384442, 4.393482, 5.398128, 
    6.39812, 7.393215, 8.383177, 9.367781, 10.34682, 11.32008, 12.28739, 
    13.24856, 14.20343, 15.15185, 16.09367, 17.02878, 17.95705, 18.87837, 
    19.79265, 20.69982, 21.59979, 22.49251, 23.37793, 24.256, 25.12669, 
    25.98999, 26.84588, 27.69435, 28.53541, 29.36907, 30.19535, 31.01428, 
    31.82589, 32.63021, 33.42731, 34.21722, 35,
  305, 305.7828, 306.5727, 307.3698, 308.1741, 308.9857, 309.8047, 310.6309, 
    311.4646, 312.3057, 313.1541, 314.01, 314.8733, 315.744, 316.6221, 
    317.5075, 318.4002, 319.3002, 320.2073, 321.1216, 322.043, 322.9712, 
    323.9063, 324.8481, 325.7966, 326.7514, 327.7126, 328.6799, 329.6532, 
    330.6322, 331.6168, 332.6068, 333.6019, 334.6019, 335.6065, 336.6156, 
    337.6287, 338.6458, 339.6663, 340.6902, 341.717, 342.7465, 343.7783, 
    344.8122, 345.8477, 346.8846, 347.9225, 348.9611, 350, 351.0389, 
    352.0775, 353.1154, 354.1523, 355.1878, 356.2217, 357.2535, 358.283, 
    359.3098, 0.3336662, 1.354252, 2.371273, 3.384442, 4.393482, 5.398128, 
    6.39812, 7.393215, 8.383177, 9.367781, 10.34682, 11.32008, 12.28739, 
    13.24856, 14.20343, 15.15185, 16.09367, 17.02878, 17.95705, 18.87837, 
    19.79265, 20.69982, 21.59979, 22.49251, 23.37793, 24.256, 25.12669, 
    25.98999, 26.84588, 27.69435, 28.53541, 29.36907, 30.19535, 31.01428, 
    31.82589, 32.63021, 33.42731, 34.21722, 35,
  305, 305.7828, 306.5727, 307.3698, 308.1741, 308.9857, 309.8047, 310.6309, 
    311.4646, 312.3057, 313.1541, 314.01, 314.8733, 315.744, 316.6221, 
    317.5075, 318.4002, 319.3002, 320.2073, 321.1216, 322.043, 322.9712, 
    323.9063, 324.8481, 325.7966, 326.7514, 327.7126, 328.6799, 329.6532, 
    330.6322, 331.6168, 332.6068, 333.6019, 334.6019, 335.6065, 336.6156, 
    337.6287, 338.6458, 339.6663, 340.6902, 341.717, 342.7465, 343.7783, 
    344.8122, 345.8477, 346.8846, 347.9225, 348.9611, 350, 351.0389, 
    352.0775, 353.1154, 354.1523, 355.1878, 356.2217, 357.2535, 358.283, 
    359.3098, 0.3336662, 1.354252, 2.371273, 3.384442, 4.393482, 5.398128, 
    6.39812, 7.393215, 8.383177, 9.367781, 10.34682, 11.32008, 12.28739, 
    13.24856, 14.20343, 15.15185, 16.09367, 17.02878, 17.95705, 18.87837, 
    19.79265, 20.69982, 21.59979, 22.49251, 23.37793, 24.256, 25.12669, 
    25.98999, 26.84588, 27.69435, 28.53541, 29.36907, 30.19535, 31.01428, 
    31.82589, 32.63021, 33.42731, 34.21722, 35,
  305, 305.7828, 306.5727, 307.3698, 308.1741, 308.9857, 309.8047, 310.6309, 
    311.4646, 312.3057, 313.1541, 314.01, 314.8733, 315.744, 316.6221, 
    317.5075, 318.4002, 319.3002, 320.2073, 321.1216, 322.043, 322.9712, 
    323.9063, 324.8481, 325.7966, 326.7514, 327.7126, 328.6799, 329.6532, 
    330.6322, 331.6168, 332.6068, 333.6019, 334.6019, 335.6065, 336.6156, 
    337.6287, 338.6458, 339.6663, 340.6902, 341.717, 342.7465, 343.7783, 
    344.8122, 345.8477, 346.8846, 347.9225, 348.9611, 350, 351.0389, 
    352.0775, 353.1154, 354.1523, 355.1878, 356.2217, 357.2535, 358.283, 
    359.3098, 0.3336662, 1.354252, 2.371273, 3.384442, 4.393482, 5.398128, 
    6.39812, 7.393215, 8.383177, 9.367781, 10.34682, 11.32008, 12.28739, 
    13.24856, 14.20343, 15.15185, 16.09367, 17.02878, 17.95705, 18.87837, 
    19.79265, 20.69982, 21.59979, 22.49251, 23.37793, 24.256, 25.12669, 
    25.98999, 26.84588, 27.69435, 28.53541, 29.36907, 30.19535, 31.01428, 
    31.82589, 32.63021, 33.42731, 34.21722, 35,
  305, 305.7828, 306.5727, 307.3698, 308.1741, 308.9857, 309.8047, 310.6309, 
    311.4646, 312.3057, 313.1541, 314.01, 314.8733, 315.744, 316.6221, 
    317.5075, 318.4002, 319.3002, 320.2073, 321.1216, 322.043, 322.9712, 
    323.9063, 324.8481, 325.7966, 326.7514, 327.7126, 328.6799, 329.6532, 
    330.6322, 331.6168, 332.6068, 333.6019, 334.6019, 335.6065, 336.6156, 
    337.6287, 338.6458, 339.6663, 340.6902, 341.717, 342.7465, 343.7783, 
    344.8122, 345.8477, 346.8846, 347.9225, 348.9611, 350, 351.0389, 
    352.0775, 353.1154, 354.1523, 355.1878, 356.2217, 357.2535, 358.283, 
    359.3098, 0.3336662, 1.354252, 2.371273, 3.384442, 4.393482, 5.398128, 
    6.39812, 7.393215, 8.383177, 9.367781, 10.34682, 11.32008, 12.28739, 
    13.24856, 14.20343, 15.15185, 16.09367, 17.02878, 17.95705, 18.87837, 
    19.79265, 20.69982, 21.59979, 22.49251, 23.37793, 24.256, 25.12669, 
    25.98999, 26.84588, 27.69435, 28.53541, 29.36907, 30.19535, 31.01428, 
    31.82589, 32.63021, 33.42731, 34.21722, 35,
  305, 305.7828, 306.5727, 307.3698, 308.1741, 308.9857, 309.8047, 310.6309, 
    311.4646, 312.3057, 313.1541, 314.01, 314.8733, 315.744, 316.6221, 
    317.5075, 318.4002, 319.3002, 320.2073, 321.1216, 322.043, 322.9712, 
    323.9063, 324.8481, 325.7966, 326.7514, 327.7126, 328.6799, 329.6532, 
    330.6322, 331.6168, 332.6068, 333.6019, 334.6019, 335.6065, 336.6156, 
    337.6287, 338.6458, 339.6663, 340.6902, 341.717, 342.7465, 343.7783, 
    344.8122, 345.8477, 346.8846, 347.9225, 348.9611, 350, 351.0389, 
    352.0775, 353.1154, 354.1523, 355.1878, 356.2217, 357.2535, 358.283, 
    359.3098, 0.3336662, 1.354252, 2.371273, 3.384442, 4.393482, 5.398128, 
    6.39812, 7.393215, 8.383177, 9.367781, 10.34682, 11.32008, 12.28739, 
    13.24856, 14.20343, 15.15185, 16.09367, 17.02878, 17.95705, 18.87837, 
    19.79265, 20.69982, 21.59979, 22.49251, 23.37793, 24.256, 25.12669, 
    25.98999, 26.84588, 27.69435, 28.53541, 29.36907, 30.19535, 31.01428, 
    31.82589, 32.63021, 33.42731, 34.21722, 35,
  305, 305.7828, 306.5727, 307.3698, 308.1741, 308.9857, 309.8047, 310.6309, 
    311.4646, 312.3057, 313.1541, 314.01, 314.8733, 315.744, 316.6221, 
    317.5075, 318.4002, 319.3002, 320.2073, 321.1216, 322.043, 322.9712, 
    323.9063, 324.8481, 325.7966, 326.7514, 327.7126, 328.6799, 329.6532, 
    330.6322, 331.6168, 332.6068, 333.6019, 334.6019, 335.6065, 336.6156, 
    337.6287, 338.6458, 339.6663, 340.6902, 341.717, 342.7465, 343.7783, 
    344.8122, 345.8477, 346.8846, 347.9225, 348.9611, 350, 351.0389, 
    352.0775, 353.1154, 354.1523, 355.1878, 356.2217, 357.2535, 358.283, 
    359.3098, 0.3336662, 1.354252, 2.371273, 3.384442, 4.393482, 5.398128, 
    6.39812, 7.393215, 8.383177, 9.367781, 10.34682, 11.32008, 12.28739, 
    13.24856, 14.20343, 15.15185, 16.09367, 17.02878, 17.95705, 18.87837, 
    19.79265, 20.69982, 21.59979, 22.49251, 23.37793, 24.256, 25.12669, 
    25.98999, 26.84588, 27.69435, 28.53541, 29.36907, 30.19535, 31.01428, 
    31.82589, 32.63021, 33.42731, 34.21722, 35,
  305, 305.7828, 306.5727, 307.3698, 308.1741, 308.9857, 309.8047, 310.6309, 
    311.4646, 312.3057, 313.1541, 314.01, 314.8733, 315.744, 316.6221, 
    317.5075, 318.4002, 319.3002, 320.2073, 321.1216, 322.043, 322.9712, 
    323.9063, 324.8481, 325.7966, 326.7514, 327.7126, 328.6799, 329.6532, 
    330.6322, 331.6168, 332.6068, 333.6019, 334.6019, 335.6065, 336.6156, 
    337.6287, 338.6458, 339.6663, 340.6902, 341.717, 342.7465, 343.7783, 
    344.8122, 345.8477, 346.8846, 347.9225, 348.9611, 350, 351.0389, 
    352.0775, 353.1154, 354.1523, 355.1878, 356.2217, 357.2535, 358.283, 
    359.3098, 0.3336662, 1.354252, 2.371273, 3.384442, 4.393482, 5.398128, 
    6.39812, 7.393215, 8.383177, 9.367781, 10.34682, 11.32008, 12.28739, 
    13.24856, 14.20343, 15.15185, 16.09367, 17.02878, 17.95705, 18.87837, 
    19.79265, 20.69982, 21.59979, 22.49251, 23.37793, 24.256, 25.12669, 
    25.98999, 26.84588, 27.69435, 28.53541, 29.36907, 30.19535, 31.01428, 
    31.82589, 32.63021, 33.42731, 34.21722, 35,
  305, 305.7828, 306.5727, 307.3698, 308.1741, 308.9857, 309.8047, 310.6309, 
    311.4646, 312.3057, 313.1541, 314.01, 314.8733, 315.744, 316.6221, 
    317.5075, 318.4002, 319.3002, 320.2073, 321.1216, 322.043, 322.9712, 
    323.9063, 324.8481, 325.7966, 326.7514, 327.7126, 328.6799, 329.6532, 
    330.6322, 331.6168, 332.6068, 333.6019, 334.6019, 335.6065, 336.6156, 
    337.6287, 338.6458, 339.6663, 340.6902, 341.717, 342.7465, 343.7783, 
    344.8122, 345.8477, 346.8846, 347.9225, 348.9611, 350, 351.0389, 
    352.0775, 353.1154, 354.1523, 355.1878, 356.2217, 357.2535, 358.283, 
    359.3098, 0.3336662, 1.354252, 2.371273, 3.384442, 4.393482, 5.398128, 
    6.39812, 7.393215, 8.383177, 9.367781, 10.34682, 11.32008, 12.28739, 
    13.24856, 14.20343, 15.15185, 16.09367, 17.02878, 17.95705, 18.87837, 
    19.79265, 20.69982, 21.59979, 22.49251, 23.37793, 24.256, 25.12669, 
    25.98999, 26.84588, 27.69435, 28.53541, 29.36907, 30.19535, 31.01428, 
    31.82589, 32.63021, 33.42731, 34.21722, 35,
  305, 305.7828, 306.5727, 307.3698, 308.1741, 308.9857, 309.8047, 310.6309, 
    311.4646, 312.3057, 313.1541, 314.01, 314.8733, 315.744, 316.6221, 
    317.5075, 318.4002, 319.3002, 320.2073, 321.1216, 322.043, 322.9712, 
    323.9063, 324.8481, 325.7966, 326.7514, 327.7126, 328.6799, 329.6532, 
    330.6322, 331.6168, 332.6068, 333.6019, 334.6019, 335.6065, 336.6156, 
    337.6287, 338.6458, 339.6663, 340.6902, 341.717, 342.7465, 343.7783, 
    344.8122, 345.8477, 346.8846, 347.9225, 348.9611, 350, 351.0389, 
    352.0775, 353.1154, 354.1523, 355.1878, 356.2217, 357.2535, 358.283, 
    359.3098, 0.3336662, 1.354252, 2.371273, 3.384442, 4.393482, 5.398128, 
    6.39812, 7.393215, 8.383177, 9.367781, 10.34682, 11.32008, 12.28739, 
    13.24856, 14.20343, 15.15185, 16.09367, 17.02878, 17.95705, 18.87837, 
    19.79265, 20.69982, 21.59979, 22.49251, 23.37793, 24.256, 25.12669, 
    25.98999, 26.84588, 27.69435, 28.53541, 29.36907, 30.19535, 31.01428, 
    31.82589, 32.63021, 33.42731, 34.21722, 35,
  305, 305.7828, 306.5727, 307.3698, 308.1741, 308.9857, 309.8047, 310.6309, 
    311.4646, 312.3057, 313.1541, 314.01, 314.8733, 315.744, 316.6221, 
    317.5075, 318.4002, 319.3002, 320.2073, 321.1216, 322.043, 322.9712, 
    323.9063, 324.8481, 325.7966, 326.7514, 327.7126, 328.6799, 329.6532, 
    330.6322, 331.6168, 332.6068, 333.6019, 334.6019, 335.6065, 336.6156, 
    337.6287, 338.6458, 339.6663, 340.6902, 341.717, 342.7465, 343.7783, 
    344.8122, 345.8477, 346.8846, 347.9225, 348.9611, 350, 351.0389, 
    352.0775, 353.1154, 354.1523, 355.1878, 356.2217, 357.2535, 358.283, 
    359.3098, 0.3336662, 1.354252, 2.371273, 3.384442, 4.393482, 5.398128, 
    6.39812, 7.393215, 8.383177, 9.367781, 10.34682, 11.32008, 12.28739, 
    13.24856, 14.20343, 15.15185, 16.09367, 17.02878, 17.95705, 18.87837, 
    19.79265, 20.69982, 21.59979, 22.49251, 23.37793, 24.256, 25.12669, 
    25.98999, 26.84588, 27.69435, 28.53541, 29.36907, 30.19535, 31.01428, 
    31.82589, 32.63021, 33.42731, 34.21722, 35,
  305, 305.7828, 306.5727, 307.3698, 308.1741, 308.9857, 309.8047, 310.6309, 
    311.4646, 312.3057, 313.1541, 314.01, 314.8733, 315.744, 316.6221, 
    317.5075, 318.4002, 319.3002, 320.2073, 321.1216, 322.043, 322.9712, 
    323.9063, 324.8481, 325.7966, 326.7514, 327.7126, 328.6799, 329.6532, 
    330.6322, 331.6168, 332.6068, 333.6019, 334.6019, 335.6065, 336.6156, 
    337.6287, 338.6458, 339.6663, 340.6902, 341.717, 342.7465, 343.7783, 
    344.8122, 345.8477, 346.8846, 347.9225, 348.9611, 350, 351.0389, 
    352.0775, 353.1154, 354.1523, 355.1878, 356.2217, 357.2535, 358.283, 
    359.3098, 0.3336662, 1.354252, 2.371273, 3.384442, 4.393482, 5.398128, 
    6.39812, 7.393215, 8.383177, 9.367781, 10.34682, 11.32008, 12.28739, 
    13.24856, 14.20343, 15.15185, 16.09367, 17.02878, 17.95705, 18.87837, 
    19.79265, 20.69982, 21.59979, 22.49251, 23.37793, 24.256, 25.12669, 
    25.98999, 26.84588, 27.69435, 28.53541, 29.36907, 30.19535, 31.01428, 
    31.82589, 32.63021, 33.42731, 34.21722, 35,
  305, 305.7828, 306.5727, 307.3698, 308.1741, 308.9857, 309.8047, 310.6309, 
    311.4646, 312.3057, 313.1541, 314.01, 314.8733, 315.744, 316.6221, 
    317.5075, 318.4002, 319.3002, 320.2073, 321.1216, 322.043, 322.9712, 
    323.9063, 324.8481, 325.7966, 326.7514, 327.7126, 328.6799, 329.6532, 
    330.6322, 331.6168, 332.6068, 333.6019, 334.6019, 335.6065, 336.6156, 
    337.6287, 338.6458, 339.6663, 340.6902, 341.717, 342.7465, 343.7783, 
    344.8122, 345.8477, 346.8846, 347.9225, 348.9611, 350, 351.0389, 
    352.0775, 353.1154, 354.1523, 355.1878, 356.2217, 357.2535, 358.283, 
    359.3098, 0.3336662, 1.354252, 2.371273, 3.384442, 4.393482, 5.398128, 
    6.39812, 7.393215, 8.383177, 9.367781, 10.34682, 11.32008, 12.28739, 
    13.24856, 14.20343, 15.15185, 16.09367, 17.02878, 17.95705, 18.87837, 
    19.79265, 20.69982, 21.59979, 22.49251, 23.37793, 24.256, 25.12669, 
    25.98999, 26.84588, 27.69435, 28.53541, 29.36907, 30.19535, 31.01428, 
    31.82589, 32.63021, 33.42731, 34.21722, 35,
  305, 305.7828, 306.5727, 307.3698, 308.1741, 308.9857, 309.8047, 310.6309, 
    311.4646, 312.3057, 313.1541, 314.01, 314.8733, 315.744, 316.6221, 
    317.5075, 318.4002, 319.3002, 320.2073, 321.1216, 322.043, 322.9712, 
    323.9063, 324.8481, 325.7966, 326.7514, 327.7126, 328.6799, 329.6532, 
    330.6322, 331.6168, 332.6068, 333.6019, 334.6019, 335.6065, 336.6156, 
    337.6287, 338.6458, 339.6663, 340.6902, 341.717, 342.7465, 343.7783, 
    344.8122, 345.8477, 346.8846, 347.9225, 348.9611, 350, 351.0389, 
    352.0775, 353.1154, 354.1523, 355.1878, 356.2217, 357.2535, 358.283, 
    359.3098, 0.3336662, 1.354252, 2.371273, 3.384442, 4.393482, 5.398128, 
    6.39812, 7.393215, 8.383177, 9.367781, 10.34682, 11.32008, 12.28739, 
    13.24856, 14.20343, 15.15185, 16.09367, 17.02878, 17.95705, 18.87837, 
    19.79265, 20.69982, 21.59979, 22.49251, 23.37793, 24.256, 25.12669, 
    25.98999, 26.84588, 27.69435, 28.53541, 29.36907, 30.19535, 31.01428, 
    31.82589, 32.63021, 33.42731, 34.21722, 35,
  305, 305.7828, 306.5727, 307.3698, 308.1741, 308.9857, 309.8047, 310.6309, 
    311.4646, 312.3057, 313.1541, 314.01, 314.8733, 315.744, 316.6221, 
    317.5075, 318.4002, 319.3002, 320.2073, 321.1216, 322.043, 322.9712, 
    323.9063, 324.8481, 325.7966, 326.7514, 327.7126, 328.6799, 329.6532, 
    330.6322, 331.6168, 332.6068, 333.6019, 334.6019, 335.6065, 336.6156, 
    337.6287, 338.6458, 339.6663, 340.6902, 341.717, 342.7465, 343.7783, 
    344.8122, 345.8477, 346.8846, 347.9225, 348.9611, 350, 351.0389, 
    352.0775, 353.1154, 354.1523, 355.1878, 356.2217, 357.2535, 358.283, 
    359.3098, 0.3336662, 1.354252, 2.371273, 3.384442, 4.393482, 5.398128, 
    6.39812, 7.393215, 8.383177, 9.367781, 10.34682, 11.32008, 12.28739, 
    13.24856, 14.20343, 15.15185, 16.09367, 17.02878, 17.95705, 18.87837, 
    19.79265, 20.69982, 21.59979, 22.49251, 23.37793, 24.256, 25.12669, 
    25.98999, 26.84588, 27.69435, 28.53541, 29.36907, 30.19535, 31.01428, 
    31.82589, 32.63021, 33.42731, 34.21722, 35,
  305, 305.7828, 306.5727, 307.3698, 308.1741, 308.9857, 309.8047, 310.6309, 
    311.4646, 312.3057, 313.1541, 314.01, 314.8733, 315.744, 316.6221, 
    317.5075, 318.4002, 319.3002, 320.2073, 321.1216, 322.043, 322.9712, 
    323.9063, 324.8481, 325.7966, 326.7514, 327.7126, 328.6799, 329.6532, 
    330.6322, 331.6168, 332.6068, 333.6019, 334.6019, 335.6065, 336.6156, 
    337.6287, 338.6458, 339.6663, 340.6902, 341.717, 342.7465, 343.7783, 
    344.8122, 345.8477, 346.8846, 347.9225, 348.9611, 350, 351.0389, 
    352.0775, 353.1154, 354.1523, 355.1878, 356.2217, 357.2535, 358.283, 
    359.3098, 0.3336662, 1.354252, 2.371273, 3.384442, 4.393482, 5.398128, 
    6.39812, 7.393215, 8.383177, 9.367781, 10.34682, 11.32008, 12.28739, 
    13.24856, 14.20343, 15.15185, 16.09367, 17.02878, 17.95705, 18.87837, 
    19.79265, 20.69982, 21.59979, 22.49251, 23.37793, 24.256, 25.12669, 
    25.98999, 26.84588, 27.69435, 28.53541, 29.36907, 30.19535, 31.01428, 
    31.82589, 32.63021, 33.42731, 34.21722, 35,
  305, 305.7828, 306.5727, 307.3698, 308.1741, 308.9857, 309.8047, 310.6309, 
    311.4646, 312.3057, 313.1541, 314.01, 314.8733, 315.744, 316.6221, 
    317.5075, 318.4002, 319.3002, 320.2073, 321.1216, 322.043, 322.9712, 
    323.9063, 324.8481, 325.7966, 326.7514, 327.7126, 328.6799, 329.6532, 
    330.6322, 331.6168, 332.6068, 333.6019, 334.6019, 335.6065, 336.6156, 
    337.6287, 338.6458, 339.6663, 340.6902, 341.717, 342.7465, 343.7783, 
    344.8122, 345.8477, 346.8846, 347.9225, 348.9611, 350, 351.0389, 
    352.0775, 353.1154, 354.1523, 355.1878, 356.2217, 357.2535, 358.283, 
    359.3098, 0.3336662, 1.354252, 2.371273, 3.384442, 4.393482, 5.398128, 
    6.39812, 7.393215, 8.383177, 9.367781, 10.34682, 11.32008, 12.28739, 
    13.24856, 14.20343, 15.15185, 16.09367, 17.02878, 17.95705, 18.87837, 
    19.79265, 20.69982, 21.59979, 22.49251, 23.37793, 24.256, 25.12669, 
    25.98999, 26.84588, 27.69435, 28.53541, 29.36907, 30.19535, 31.01428, 
    31.82589, 32.63021, 33.42731, 34.21722, 35,
  305, 305.7828, 306.5727, 307.3698, 308.1741, 308.9857, 309.8047, 310.6309, 
    311.4646, 312.3057, 313.1541, 314.01, 314.8733, 315.744, 316.6221, 
    317.5075, 318.4002, 319.3002, 320.2073, 321.1216, 322.043, 322.9712, 
    323.9063, 324.8481, 325.7966, 326.7514, 327.7126, 328.6799, 329.6532, 
    330.6322, 331.6168, 332.6068, 333.6019, 334.6019, 335.6065, 336.6156, 
    337.6287, 338.6458, 339.6663, 340.6902, 341.717, 342.7465, 343.7783, 
    344.8122, 345.8477, 346.8846, 347.9225, 348.9611, 350, 351.0389, 
    352.0775, 353.1154, 354.1523, 355.1878, 356.2217, 357.2535, 358.283, 
    359.3098, 0.3336662, 1.354252, 2.371273, 3.384442, 4.393482, 5.398128, 
    6.39812, 7.393215, 8.383177, 9.367781, 10.34682, 11.32008, 12.28739, 
    13.24856, 14.20343, 15.15185, 16.09367, 17.02878, 17.95705, 18.87837, 
    19.79265, 20.69982, 21.59979, 22.49251, 23.37793, 24.256, 25.12669, 
    25.98999, 26.84588, 27.69435, 28.53541, 29.36907, 30.19535, 31.01428, 
    31.82589, 32.63021, 33.42731, 34.21722, 35,
  305, 305.7828, 306.5727, 307.3698, 308.1741, 308.9857, 309.8047, 310.6309, 
    311.4646, 312.3057, 313.1541, 314.01, 314.8733, 315.744, 316.6221, 
    317.5075, 318.4002, 319.3002, 320.2073, 321.1216, 322.043, 322.9712, 
    323.9063, 324.8481, 325.7966, 326.7514, 327.7126, 328.6799, 329.6532, 
    330.6322, 331.6168, 332.6068, 333.6019, 334.6019, 335.6065, 336.6156, 
    337.6287, 338.6458, 339.6663, 340.6902, 341.717, 342.7465, 343.7783, 
    344.8122, 345.8477, 346.8846, 347.9225, 348.9611, 350, 351.0389, 
    352.0775, 353.1154, 354.1523, 355.1878, 356.2217, 357.2535, 358.283, 
    359.3098, 0.3336662, 1.354252, 2.371273, 3.384442, 4.393482, 5.398128, 
    6.39812, 7.393215, 8.383177, 9.367781, 10.34682, 11.32008, 12.28739, 
    13.24856, 14.20343, 15.15185, 16.09367, 17.02878, 17.95705, 18.87837, 
    19.79265, 20.69982, 21.59979, 22.49251, 23.37793, 24.256, 25.12669, 
    25.98999, 26.84588, 27.69435, 28.53541, 29.36907, 30.19535, 31.01428, 
    31.82589, 32.63021, 33.42731, 34.21722, 35,
  305, 305.7828, 306.5727, 307.3698, 308.1741, 308.9857, 309.8047, 310.6309, 
    311.4646, 312.3057, 313.1541, 314.01, 314.8733, 315.744, 316.6221, 
    317.5075, 318.4002, 319.3002, 320.2073, 321.1216, 322.043, 322.9712, 
    323.9063, 324.8481, 325.7966, 326.7514, 327.7126, 328.6799, 329.6532, 
    330.6322, 331.6168, 332.6068, 333.6019, 334.6019, 335.6065, 336.6156, 
    337.6287, 338.6458, 339.6663, 340.6902, 341.717, 342.7465, 343.7783, 
    344.8122, 345.8477, 346.8846, 347.9225, 348.9611, 350, 351.0389, 
    352.0775, 353.1154, 354.1523, 355.1878, 356.2217, 357.2535, 358.283, 
    359.3098, 0.3336662, 1.354252, 2.371273, 3.384442, 4.393482, 5.398128, 
    6.39812, 7.393215, 8.383177, 9.367781, 10.34682, 11.32008, 12.28739, 
    13.24856, 14.20343, 15.15185, 16.09367, 17.02878, 17.95705, 18.87837, 
    19.79265, 20.69982, 21.59979, 22.49251, 23.37793, 24.256, 25.12669, 
    25.98999, 26.84588, 27.69435, 28.53541, 29.36907, 30.19535, 31.01428, 
    31.82589, 32.63021, 33.42731, 34.21722, 35,
  305, 305.7828, 306.5727, 307.3698, 308.1741, 308.9857, 309.8047, 310.6309, 
    311.4646, 312.3057, 313.1541, 314.01, 314.8733, 315.744, 316.6221, 
    317.5075, 318.4002, 319.3002, 320.2073, 321.1216, 322.043, 322.9712, 
    323.9063, 324.8481, 325.7966, 326.7514, 327.7126, 328.6799, 329.6532, 
    330.6322, 331.6168, 332.6068, 333.6019, 334.6019, 335.6065, 336.6156, 
    337.6287, 338.6458, 339.6663, 340.6902, 341.717, 342.7465, 343.7783, 
    344.8122, 345.8477, 346.8846, 347.9225, 348.9611, 350, 351.0389, 
    352.0775, 353.1154, 354.1523, 355.1878, 356.2217, 357.2535, 358.283, 
    359.3098, 0.3336662, 1.354252, 2.371273, 3.384442, 4.393482, 5.398128, 
    6.39812, 7.393215, 8.383177, 9.367781, 10.34682, 11.32008, 12.28739, 
    13.24856, 14.20343, 15.15185, 16.09367, 17.02878, 17.95705, 18.87837, 
    19.79265, 20.69982, 21.59979, 22.49251, 23.37793, 24.256, 25.12669, 
    25.98999, 26.84588, 27.69435, 28.53541, 29.36907, 30.19535, 31.01428, 
    31.82589, 32.63021, 33.42731, 34.21722, 35,
  305, 305.7828, 306.5727, 307.3698, 308.1741, 308.9857, 309.8047, 310.6309, 
    311.4646, 312.3057, 313.1541, 314.01, 314.8733, 315.744, 316.6221, 
    317.5075, 318.4002, 319.3002, 320.2073, 321.1216, 322.043, 322.9712, 
    323.9063, 324.8481, 325.7966, 326.7514, 327.7126, 328.6799, 329.6532, 
    330.6322, 331.6168, 332.6068, 333.6019, 334.6019, 335.6065, 336.6156, 
    337.6287, 338.6458, 339.6663, 340.6902, 341.717, 342.7465, 343.7783, 
    344.8122, 345.8477, 346.8846, 347.9225, 348.9611, 350, 351.0389, 
    352.0775, 353.1154, 354.1523, 355.1878, 356.2217, 357.2535, 358.283, 
    359.3098, 0.3336662, 1.354252, 2.371273, 3.384442, 4.393482, 5.398128, 
    6.39812, 7.393215, 8.383177, 9.367781, 10.34682, 11.32008, 12.28739, 
    13.24856, 14.20343, 15.15185, 16.09367, 17.02878, 17.95705, 18.87837, 
    19.79265, 20.69982, 21.59979, 22.49251, 23.37793, 24.256, 25.12669, 
    25.98999, 26.84588, 27.69435, 28.53541, 29.36907, 30.19535, 31.01428, 
    31.82589, 32.63021, 33.42731, 34.21722, 35,
  305, 305.7828, 306.5727, 307.3698, 308.1741, 308.9857, 309.8047, 310.6309, 
    311.4646, 312.3057, 313.1541, 314.01, 314.8733, 315.744, 316.6221, 
    317.5075, 318.4002, 319.3002, 320.2073, 321.1216, 322.043, 322.9712, 
    323.9063, 324.8481, 325.7966, 326.7514, 327.7126, 328.6799, 329.6532, 
    330.6322, 331.6168, 332.6068, 333.6019, 334.6019, 335.6065, 336.6156, 
    337.6287, 338.6458, 339.6663, 340.6902, 341.717, 342.7465, 343.7783, 
    344.8122, 345.8477, 346.8846, 347.9225, 348.9611, 350, 351.0389, 
    352.0775, 353.1154, 354.1523, 355.1878, 356.2217, 357.2535, 358.283, 
    359.3098, 0.3336662, 1.354252, 2.371273, 3.384442, 4.393482, 5.398128, 
    6.39812, 7.393215, 8.383177, 9.367781, 10.34682, 11.32008, 12.28739, 
    13.24856, 14.20343, 15.15185, 16.09367, 17.02878, 17.95705, 18.87837, 
    19.79265, 20.69982, 21.59979, 22.49251, 23.37793, 24.256, 25.12669, 
    25.98999, 26.84588, 27.69435, 28.53541, 29.36907, 30.19535, 31.01428, 
    31.82589, 32.63021, 33.42731, 34.21722, 35,
  305, 305.7828, 306.5727, 307.3698, 308.1741, 308.9857, 309.8047, 310.6309, 
    311.4646, 312.3057, 313.1541, 314.01, 314.8733, 315.744, 316.6221, 
    317.5075, 318.4002, 319.3002, 320.2073, 321.1216, 322.043, 322.9712, 
    323.9063, 324.8481, 325.7966, 326.7514, 327.7126, 328.6799, 329.6532, 
    330.6322, 331.6168, 332.6068, 333.6019, 334.6019, 335.6065, 336.6156, 
    337.6287, 338.6458, 339.6663, 340.6902, 341.717, 342.7465, 343.7783, 
    344.8122, 345.8477, 346.8846, 347.9225, 348.9611, 350, 351.0389, 
    352.0775, 353.1154, 354.1523, 355.1878, 356.2217, 357.2535, 358.283, 
    359.3098, 0.3336662, 1.354252, 2.371273, 3.384442, 4.393482, 5.398128, 
    6.39812, 7.393215, 8.383177, 9.367781, 10.34682, 11.32008, 12.28739, 
    13.24856, 14.20343, 15.15185, 16.09367, 17.02878, 17.95705, 18.87837, 
    19.79265, 20.69982, 21.59979, 22.49251, 23.37793, 24.256, 25.12669, 
    25.98999, 26.84588, 27.69435, 28.53541, 29.36907, 30.19535, 31.01428, 
    31.82589, 32.63021, 33.42731, 34.21722, 35,
  305, 305.7828, 306.5727, 307.3698, 308.1741, 308.9857, 309.8047, 310.6309, 
    311.4646, 312.3057, 313.1541, 314.01, 314.8733, 315.744, 316.6221, 
    317.5075, 318.4002, 319.3002, 320.2073, 321.1216, 322.043, 322.9712, 
    323.9063, 324.8481, 325.7966, 326.7514, 327.7126, 328.6799, 329.6532, 
    330.6322, 331.6168, 332.6068, 333.6019, 334.6019, 335.6065, 336.6156, 
    337.6287, 338.6458, 339.6663, 340.6902, 341.717, 342.7465, 343.7783, 
    344.8122, 345.8477, 346.8846, 347.9225, 348.9611, 350, 351.0389, 
    352.0775, 353.1154, 354.1523, 355.1878, 356.2217, 357.2535, 358.283, 
    359.3098, 0.3336662, 1.354252, 2.371273, 3.384442, 4.393482, 5.398128, 
    6.39812, 7.393215, 8.383177, 9.367781, 10.34682, 11.32008, 12.28739, 
    13.24856, 14.20343, 15.15185, 16.09367, 17.02878, 17.95705, 18.87837, 
    19.79265, 20.69982, 21.59979, 22.49251, 23.37793, 24.256, 25.12669, 
    25.98999, 26.84588, 27.69435, 28.53541, 29.36907, 30.19535, 31.01428, 
    31.82589, 32.63021, 33.42731, 34.21722, 35,
  305, 305.7828, 306.5727, 307.3698, 308.1741, 308.9857, 309.8047, 310.6309, 
    311.4646, 312.3057, 313.1541, 314.01, 314.8733, 315.744, 316.6221, 
    317.5075, 318.4002, 319.3002, 320.2073, 321.1216, 322.043, 322.9712, 
    323.9063, 324.8481, 325.7966, 326.7514, 327.7126, 328.6799, 329.6532, 
    330.6322, 331.6168, 332.6068, 333.6019, 334.6019, 335.6065, 336.6156, 
    337.6287, 338.6458, 339.6663, 340.6902, 341.717, 342.7465, 343.7783, 
    344.8122, 345.8477, 346.8846, 347.9225, 348.9611, 350, 351.0389, 
    352.0775, 353.1154, 354.1523, 355.1878, 356.2217, 357.2535, 358.283, 
    359.3098, 0.3336662, 1.354252, 2.371273, 3.384442, 4.393482, 5.398128, 
    6.39812, 7.393215, 8.383177, 9.367781, 10.34682, 11.32008, 12.28739, 
    13.24856, 14.20343, 15.15185, 16.09367, 17.02878, 17.95705, 18.87837, 
    19.79265, 20.69982, 21.59979, 22.49251, 23.37793, 24.256, 25.12669, 
    25.98999, 26.84588, 27.69435, 28.53541, 29.36907, 30.19535, 31.01428, 
    31.82589, 32.63021, 33.42731, 34.21722, 35,
  305, 305.7828, 306.5727, 307.3698, 308.1741, 308.9857, 309.8047, 310.6309, 
    311.4646, 312.3057, 313.1541, 314.01, 314.8733, 315.744, 316.6221, 
    317.5075, 318.4002, 319.3002, 320.2073, 321.1216, 322.043, 322.9712, 
    323.9063, 324.8481, 325.7966, 326.7514, 327.7126, 328.6799, 329.6532, 
    330.6322, 331.6168, 332.6068, 333.6019, 334.6019, 335.6065, 336.6156, 
    337.6287, 338.6458, 339.6663, 340.6902, 341.717, 342.7465, 343.7783, 
    344.8122, 345.8477, 346.8846, 347.9225, 348.9611, 350, 351.0389, 
    352.0775, 353.1154, 354.1523, 355.1878, 356.2217, 357.2535, 358.283, 
    359.3098, 0.3336662, 1.354252, 2.371273, 3.384442, 4.393482, 5.398128, 
    6.39812, 7.393215, 8.383177, 9.367781, 10.34682, 11.32008, 12.28739, 
    13.24856, 14.20343, 15.15185, 16.09367, 17.02878, 17.95705, 18.87837, 
    19.79265, 20.69982, 21.59979, 22.49251, 23.37793, 24.256, 25.12669, 
    25.98999, 26.84588, 27.69435, 28.53541, 29.36907, 30.19535, 31.01428, 
    31.82589, 32.63021, 33.42731, 34.21722, 35,
  305, 305.7828, 306.5727, 307.3698, 308.1741, 308.9857, 309.8047, 310.6309, 
    311.4646, 312.3057, 313.1541, 314.01, 314.8733, 315.744, 316.6221, 
    317.5075, 318.4002, 319.3002, 320.2073, 321.1216, 322.043, 322.9712, 
    323.9063, 324.8481, 325.7966, 326.7514, 327.7126, 328.6799, 329.6532, 
    330.6322, 331.6168, 332.6068, 333.6019, 334.6019, 335.6065, 336.6156, 
    337.6287, 338.6458, 339.6663, 340.6902, 341.717, 342.7465, 343.7783, 
    344.8122, 345.8477, 346.8846, 347.9225, 348.9611, 350, 351.0389, 
    352.0775, 353.1154, 354.1523, 355.1878, 356.2217, 357.2535, 358.283, 
    359.3098, 0.3336662, 1.354252, 2.371273, 3.384442, 4.393482, 5.398128, 
    6.39812, 7.393215, 8.383177, 9.367781, 10.34682, 11.32008, 12.28739, 
    13.24856, 14.20343, 15.15185, 16.09367, 17.02878, 17.95705, 18.87837, 
    19.79265, 20.69982, 21.59979, 22.49251, 23.37793, 24.256, 25.12669, 
    25.98999, 26.84588, 27.69435, 28.53541, 29.36907, 30.19535, 31.01428, 
    31.82589, 32.63021, 33.42731, 34.21722, 35,
  305, 305.7828, 306.5727, 307.3698, 308.1741, 308.9857, 309.8047, 310.6309, 
    311.4646, 312.3057, 313.1541, 314.01, 314.8733, 315.744, 316.6221, 
    317.5075, 318.4002, 319.3002, 320.2073, 321.1216, 322.043, 322.9712, 
    323.9063, 324.8481, 325.7966, 326.7514, 327.7126, 328.6799, 329.6532, 
    330.6322, 331.6168, 332.6068, 333.6019, 334.6019, 335.6065, 336.6156, 
    337.6287, 338.6458, 339.6663, 340.6902, 341.717, 342.7465, 343.7783, 
    344.8122, 345.8477, 346.8846, 347.9225, 348.9611, 350, 351.0389, 
    352.0775, 353.1154, 354.1523, 355.1878, 356.2217, 357.2535, 358.283, 
    359.3098, 0.3336662, 1.354252, 2.371273, 3.384442, 4.393482, 5.398128, 
    6.39812, 7.393215, 8.383177, 9.367781, 10.34682, 11.32008, 12.28739, 
    13.24856, 14.20343, 15.15185, 16.09367, 17.02878, 17.95705, 18.87837, 
    19.79265, 20.69982, 21.59979, 22.49251, 23.37793, 24.256, 25.12669, 
    25.98999, 26.84588, 27.69435, 28.53541, 29.36907, 30.19535, 31.01428, 
    31.82589, 32.63021, 33.42731, 34.21722, 35,
  305, 305.7828, 306.5727, 307.3698, 308.1741, 308.9857, 309.8047, 310.6309, 
    311.4646, 312.3057, 313.1541, 314.01, 314.8733, 315.744, 316.6221, 
    317.5075, 318.4002, 319.3002, 320.2073, 321.1216, 322.043, 322.9712, 
    323.9063, 324.8481, 325.7966, 326.7514, 327.7126, 328.6799, 329.6532, 
    330.6322, 331.6168, 332.6068, 333.6019, 334.6019, 335.6065, 336.6156, 
    337.6287, 338.6458, 339.6663, 340.6902, 341.717, 342.7465, 343.7783, 
    344.8122, 345.8477, 346.8846, 347.9225, 348.9611, 350, 351.0389, 
    352.0775, 353.1154, 354.1523, 355.1878, 356.2217, 357.2535, 358.283, 
    359.3098, 0.3336662, 1.354252, 2.371273, 3.384442, 4.393482, 5.398128, 
    6.39812, 7.393215, 8.383177, 9.367781, 10.34682, 11.32008, 12.28739, 
    13.24856, 14.20343, 15.15185, 16.09367, 17.02878, 17.95705, 18.87837, 
    19.79265, 20.69982, 21.59979, 22.49251, 23.37793, 24.256, 25.12669, 
    25.98999, 26.84588, 27.69435, 28.53541, 29.36907, 30.19535, 31.01428, 
    31.82589, 32.63021, 33.42731, 34.21722, 35,
  305, 305.7828, 306.5727, 307.3698, 308.1741, 308.9857, 309.8047, 310.6309, 
    311.4646, 312.3057, 313.1541, 314.01, 314.8733, 315.744, 316.6221, 
    317.5075, 318.4002, 319.3002, 320.2073, 321.1216, 322.043, 322.9712, 
    323.9063, 324.8481, 325.7966, 326.7514, 327.7126, 328.6799, 329.6532, 
    330.6322, 331.6168, 332.6068, 333.6019, 334.6019, 335.6065, 336.6156, 
    337.6287, 338.6458, 339.6663, 340.6902, 341.717, 342.7465, 343.7783, 
    344.8122, 345.8477, 346.8846, 347.9225, 348.9611, 350, 351.0389, 
    352.0775, 353.1154, 354.1523, 355.1878, 356.2217, 357.2535, 358.283, 
    359.3098, 0.3336662, 1.354252, 2.371273, 3.384442, 4.393482, 5.398128, 
    6.39812, 7.393215, 8.383177, 9.367781, 10.34682, 11.32008, 12.28739, 
    13.24856, 14.20343, 15.15185, 16.09367, 17.02878, 17.95705, 18.87837, 
    19.79265, 20.69982, 21.59979, 22.49251, 23.37793, 24.256, 25.12669, 
    25.98999, 26.84588, 27.69435, 28.53541, 29.36907, 30.19535, 31.01428, 
    31.82589, 32.63021, 33.42731, 34.21722, 35,
  305, 305.7828, 306.5727, 307.3698, 308.1741, 308.9857, 309.8047, 310.6309, 
    311.4646, 312.3057, 313.1541, 314.01, 314.8733, 315.744, 316.6221, 
    317.5075, 318.4002, 319.3002, 320.2073, 321.1216, 322.043, 322.9712, 
    323.9063, 324.8481, 325.7966, 326.7514, 327.7126, 328.6799, 329.6532, 
    330.6322, 331.6168, 332.6068, 333.6019, 334.6019, 335.6065, 336.6156, 
    337.6287, 338.6458, 339.6663, 340.6902, 341.717, 342.7465, 343.7783, 
    344.8122, 345.8477, 346.8846, 347.9225, 348.9611, 350, 351.0389, 
    352.0775, 353.1154, 354.1523, 355.1878, 356.2217, 357.2535, 358.283, 
    359.3098, 0.3336662, 1.354252, 2.371273, 3.384442, 4.393482, 5.398128, 
    6.39812, 7.393215, 8.383177, 9.367781, 10.34682, 11.32008, 12.28739, 
    13.24856, 14.20343, 15.15185, 16.09367, 17.02878, 17.95705, 18.87837, 
    19.79265, 20.69982, 21.59979, 22.49251, 23.37793, 24.256, 25.12669, 
    25.98999, 26.84588, 27.69435, 28.53541, 29.36907, 30.19535, 31.01428, 
    31.82589, 32.63021, 33.42731, 34.21722, 35,
  305, 305.7828, 306.5727, 307.3698, 308.1741, 308.9857, 309.8047, 310.6309, 
    311.4646, 312.3057, 313.1541, 314.01, 314.8733, 315.744, 316.6221, 
    317.5075, 318.4002, 319.3002, 320.2073, 321.1216, 322.043, 322.9712, 
    323.9063, 324.8481, 325.7966, 326.7514, 327.7126, 328.6799, 329.6532, 
    330.6322, 331.6168, 332.6068, 333.6019, 334.6019, 335.6065, 336.6156, 
    337.6287, 338.6458, 339.6663, 340.6902, 341.717, 342.7465, 343.7783, 
    344.8122, 345.8477, 346.8846, 347.9225, 348.9611, 350, 351.0389, 
    352.0775, 353.1154, 354.1523, 355.1878, 356.2217, 357.2535, 358.283, 
    359.3098, 0.3336662, 1.354252, 2.371273, 3.384442, 4.393482, 5.398128, 
    6.39812, 7.393215, 8.383177, 9.367781, 10.34682, 11.32008, 12.28739, 
    13.24856, 14.20343, 15.15185, 16.09367, 17.02878, 17.95705, 18.87837, 
    19.79265, 20.69982, 21.59979, 22.49251, 23.37793, 24.256, 25.12669, 
    25.98999, 26.84588, 27.69435, 28.53541, 29.36907, 30.19535, 31.01428, 
    31.82589, 32.63021, 33.42731, 34.21722, 35,
  305, 305.7828, 306.5727, 307.3698, 308.1741, 308.9857, 309.8047, 310.6309, 
    311.4646, 312.3057, 313.1541, 314.01, 314.8733, 315.744, 316.6221, 
    317.5075, 318.4002, 319.3002, 320.2073, 321.1216, 322.043, 322.9712, 
    323.9063, 324.8481, 325.7966, 326.7514, 327.7126, 328.6799, 329.6532, 
    330.6322, 331.6168, 332.6068, 333.6019, 334.6019, 335.6065, 336.6156, 
    337.6287, 338.6458, 339.6663, 340.6902, 341.717, 342.7465, 343.7783, 
    344.8122, 345.8477, 346.8846, 347.9225, 348.9611, 350, 351.0389, 
    352.0775, 353.1154, 354.1523, 355.1878, 356.2217, 357.2535, 358.283, 
    359.3098, 0.3336662, 1.354252, 2.371273, 3.384442, 4.393482, 5.398128, 
    6.39812, 7.393215, 8.383177, 9.367781, 10.34682, 11.32008, 12.28739, 
    13.24856, 14.20343, 15.15185, 16.09367, 17.02878, 17.95705, 18.87837, 
    19.79265, 20.69982, 21.59979, 22.49251, 23.37793, 24.256, 25.12669, 
    25.98999, 26.84588, 27.69435, 28.53541, 29.36907, 30.19535, 31.01428, 
    31.82589, 32.63021, 33.42731, 34.21722, 35,
  305, 305.7828, 306.5727, 307.3698, 308.1741, 308.9857, 309.8047, 310.6309, 
    311.4646, 312.3057, 313.1541, 314.01, 314.8733, 315.744, 316.6221, 
    317.5075, 318.4002, 319.3002, 320.2073, 321.1216, 322.043, 322.9712, 
    323.9063, 324.8481, 325.7966, 326.7514, 327.7126, 328.6799, 329.6532, 
    330.6322, 331.6168, 332.6068, 333.6019, 334.6019, 335.6065, 336.6156, 
    337.6287, 338.6458, 339.6663, 340.6902, 341.717, 342.7465, 343.7783, 
    344.8122, 345.8477, 346.8846, 347.9225, 348.9611, 350, 351.0389, 
    352.0775, 353.1154, 354.1523, 355.1878, 356.2217, 357.2535, 358.283, 
    359.3098, 0.3336662, 1.354252, 2.371273, 3.384442, 4.393482, 5.398128, 
    6.39812, 7.393215, 8.383177, 9.367781, 10.34682, 11.32008, 12.28739, 
    13.24856, 14.20343, 15.15185, 16.09367, 17.02878, 17.95705, 18.87837, 
    19.79265, 20.69982, 21.59979, 22.49251, 23.37793, 24.256, 25.12669, 
    25.98999, 26.84588, 27.69435, 28.53541, 29.36907, 30.19535, 31.01428, 
    31.82589, 32.63021, 33.42731, 34.21722, 35,
  305, 305.7828, 306.5727, 307.3698, 308.1741, 308.9857, 309.8047, 310.6309, 
    311.4646, 312.3057, 313.1541, 314.01, 314.8733, 315.744, 316.6221, 
    317.5075, 318.4002, 319.3002, 320.2073, 321.1216, 322.043, 322.9712, 
    323.9063, 324.8481, 325.7966, 326.7514, 327.7126, 328.6799, 329.6532, 
    330.6322, 331.6168, 332.6068, 333.6019, 334.6019, 335.6065, 336.6156, 
    337.6287, 338.6458, 339.6663, 340.6902, 341.717, 342.7465, 343.7783, 
    344.8122, 345.8477, 346.8846, 347.9225, 348.9611, 350, 351.0389, 
    352.0775, 353.1154, 354.1523, 355.1878, 356.2217, 357.2535, 358.283, 
    359.3098, 0.3336662, 1.354252, 2.371273, 3.384442, 4.393482, 5.398128, 
    6.39812, 7.393215, 8.383177, 9.367781, 10.34682, 11.32008, 12.28739, 
    13.24856, 14.20343, 15.15185, 16.09367, 17.02878, 17.95705, 18.87837, 
    19.79265, 20.69982, 21.59979, 22.49251, 23.37793, 24.256, 25.12669, 
    25.98999, 26.84588, 27.69435, 28.53541, 29.36907, 30.19535, 31.01428, 
    31.82589, 32.63021, 33.42731, 34.21722, 35,
  305, 305.7828, 306.5727, 307.3698, 308.1741, 308.9857, 309.8047, 310.6309, 
    311.4646, 312.3057, 313.1541, 314.01, 314.8733, 315.744, 316.6221, 
    317.5075, 318.4002, 319.3002, 320.2073, 321.1216, 322.043, 322.9712, 
    323.9063, 324.8481, 325.7966, 326.7514, 327.7126, 328.6799, 329.6532, 
    330.6322, 331.6168, 332.6068, 333.6019, 334.6019, 335.6065, 336.6156, 
    337.6287, 338.6458, 339.6663, 340.6902, 341.717, 342.7465, 343.7783, 
    344.8122, 345.8477, 346.8846, 347.9225, 348.9611, 350, 351.0389, 
    352.0775, 353.1154, 354.1523, 355.1878, 356.2217, 357.2535, 358.283, 
    359.3098, 0.3336662, 1.354252, 2.371273, 3.384442, 4.393482, 5.398128, 
    6.39812, 7.393215, 8.383177, 9.367781, 10.34682, 11.32008, 12.28739, 
    13.24856, 14.20343, 15.15185, 16.09367, 17.02878, 17.95705, 18.87837, 
    19.79265, 20.69982, 21.59979, 22.49251, 23.37793, 24.256, 25.12669, 
    25.98999, 26.84588, 27.69435, 28.53541, 29.36907, 30.19535, 31.01428, 
    31.82589, 32.63021, 33.42731, 34.21722, 35,
  305, 305.7828, 306.5727, 307.3698, 308.1741, 308.9857, 309.8047, 310.6309, 
    311.4646, 312.3057, 313.1541, 314.01, 314.8733, 315.744, 316.6221, 
    317.5075, 318.4002, 319.3002, 320.2073, 321.1216, 322.043, 322.9712, 
    323.9063, 324.8481, 325.7966, 326.7514, 327.7126, 328.6799, 329.6532, 
    330.6322, 331.6168, 332.6068, 333.6019, 334.6019, 335.6065, 336.6156, 
    337.6287, 338.6458, 339.6663, 340.6902, 341.717, 342.7465, 343.7783, 
    344.8122, 345.8477, 346.8846, 347.9225, 348.9611, 350, 351.0389, 
    352.0775, 353.1154, 354.1523, 355.1878, 356.2217, 357.2535, 358.283, 
    359.3098, 0.3336662, 1.354252, 2.371273, 3.384442, 4.393482, 5.398128, 
    6.39812, 7.393215, 8.383177, 9.367781, 10.34682, 11.32008, 12.28739, 
    13.24856, 14.20343, 15.15185, 16.09367, 17.02878, 17.95705, 18.87837, 
    19.79265, 20.69982, 21.59979, 22.49251, 23.37793, 24.256, 25.12669, 
    25.98999, 26.84588, 27.69435, 28.53541, 29.36907, 30.19535, 31.01428, 
    31.82589, 32.63021, 33.42731, 34.21722, 35,
  305, 305.7828, 306.5727, 307.3698, 308.1741, 308.9857, 309.8047, 310.6309, 
    311.4646, 312.3057, 313.1541, 314.01, 314.8733, 315.744, 316.6221, 
    317.5075, 318.4002, 319.3002, 320.2073, 321.1216, 322.043, 322.9712, 
    323.9063, 324.8481, 325.7966, 326.7514, 327.7126, 328.6799, 329.6532, 
    330.6322, 331.6168, 332.6068, 333.6019, 334.6019, 335.6065, 336.6156, 
    337.6287, 338.6458, 339.6663, 340.6902, 341.717, 342.7465, 343.7783, 
    344.8122, 345.8477, 346.8846, 347.9225, 348.9611, 350, 351.0389, 
    352.0775, 353.1154, 354.1523, 355.1878, 356.2217, 357.2535, 358.283, 
    359.3098, 0.3336662, 1.354252, 2.371273, 3.384442, 4.393482, 5.398128, 
    6.39812, 7.393215, 8.383177, 9.367781, 10.34682, 11.32008, 12.28739, 
    13.24856, 14.20343, 15.15185, 16.09367, 17.02878, 17.95705, 18.87837, 
    19.79265, 20.69982, 21.59979, 22.49251, 23.37793, 24.256, 25.12669, 
    25.98999, 26.84588, 27.69435, 28.53541, 29.36907, 30.19535, 31.01428, 
    31.82589, 32.63021, 33.42731, 34.21722, 35,
  305, 305.7828, 306.5727, 307.3698, 308.1741, 308.9857, 309.8047, 310.6309, 
    311.4646, 312.3057, 313.1541, 314.01, 314.8733, 315.744, 316.6221, 
    317.5075, 318.4002, 319.3002, 320.2073, 321.1216, 322.043, 322.9712, 
    323.9063, 324.8481, 325.7966, 326.7514, 327.7126, 328.6799, 329.6532, 
    330.6322, 331.6168, 332.6068, 333.6019, 334.6019, 335.6065, 336.6156, 
    337.6287, 338.6458, 339.6663, 340.6902, 341.717, 342.7465, 343.7783, 
    344.8122, 345.8477, 346.8846, 347.9225, 348.9611, 350, 351.0389, 
    352.0775, 353.1154, 354.1523, 355.1878, 356.2217, 357.2535, 358.283, 
    359.3098, 0.3336662, 1.354252, 2.371273, 3.384442, 4.393482, 5.398128, 
    6.39812, 7.393215, 8.383177, 9.367781, 10.34682, 11.32008, 12.28739, 
    13.24856, 14.20343, 15.15185, 16.09367, 17.02878, 17.95705, 18.87837, 
    19.79265, 20.69982, 21.59979, 22.49251, 23.37793, 24.256, 25.12669, 
    25.98999, 26.84588, 27.69435, 28.53541, 29.36907, 30.19535, 31.01428, 
    31.82589, 32.63021, 33.42731, 34.21722, 35,
  305, 305.7828, 306.5727, 307.3698, 308.1741, 308.9857, 309.8047, 310.6309, 
    311.4646, 312.3057, 313.1541, 314.01, 314.8733, 315.744, 316.6221, 
    317.5075, 318.4002, 319.3002, 320.2073, 321.1216, 322.043, 322.9712, 
    323.9063, 324.8481, 325.7966, 326.7514, 327.7126, 328.6799, 329.6532, 
    330.6322, 331.6168, 332.6068, 333.6019, 334.6019, 335.6065, 336.6156, 
    337.6287, 338.6458, 339.6663, 340.6902, 341.717, 342.7465, 343.7783, 
    344.8122, 345.8477, 346.8846, 347.9225, 348.9611, 350, 351.0389, 
    352.0775, 353.1154, 354.1523, 355.1878, 356.2217, 357.2535, 358.283, 
    359.3098, 0.3336662, 1.354252, 2.371273, 3.384442, 4.393482, 5.398128, 
    6.39812, 7.393215, 8.383177, 9.367781, 10.34682, 11.32008, 12.28739, 
    13.24856, 14.20343, 15.15185, 16.09367, 17.02878, 17.95705, 18.87837, 
    19.79265, 20.69982, 21.59979, 22.49251, 23.37793, 24.256, 25.12669, 
    25.98999, 26.84588, 27.69435, 28.53541, 29.36907, 30.19535, 31.01428, 
    31.82589, 32.63021, 33.42731, 34.21722, 35,
  305, 305.7828, 306.5727, 307.3698, 308.1741, 308.9857, 309.8047, 310.6309, 
    311.4646, 312.3057, 313.1541, 314.01, 314.8733, 315.744, 316.6221, 
    317.5075, 318.4002, 319.3002, 320.2073, 321.1216, 322.043, 322.9712, 
    323.9063, 324.8481, 325.7966, 326.7514, 327.7126, 328.6799, 329.6532, 
    330.6322, 331.6168, 332.6068, 333.6019, 334.6019, 335.6065, 336.6156, 
    337.6287, 338.6458, 339.6663, 340.6902, 341.717, 342.7465, 343.7783, 
    344.8122, 345.8477, 346.8846, 347.9225, 348.9611, 350, 351.0389, 
    352.0775, 353.1154, 354.1523, 355.1878, 356.2217, 357.2535, 358.283, 
    359.3098, 0.3336662, 1.354252, 2.371273, 3.384442, 4.393482, 5.398128, 
    6.39812, 7.393215, 8.383177, 9.367781, 10.34682, 11.32008, 12.28739, 
    13.24856, 14.20343, 15.15185, 16.09367, 17.02878, 17.95705, 18.87837, 
    19.79265, 20.69982, 21.59979, 22.49251, 23.37793, 24.256, 25.12669, 
    25.98999, 26.84588, 27.69435, 28.53541, 29.36907, 30.19535, 31.01428, 
    31.82589, 32.63021, 33.42731, 34.21722, 35,
  305, 305.7828, 306.5727, 307.3698, 308.1741, 308.9857, 309.8047, 310.6309, 
    311.4646, 312.3057, 313.1541, 314.01, 314.8733, 315.744, 316.6221, 
    317.5075, 318.4002, 319.3002, 320.2073, 321.1216, 322.043, 322.9712, 
    323.9063, 324.8481, 325.7966, 326.7514, 327.7126, 328.6799, 329.6532, 
    330.6322, 331.6168, 332.6068, 333.6019, 334.6019, 335.6065, 336.6156, 
    337.6287, 338.6458, 339.6663, 340.6902, 341.717, 342.7465, 343.7783, 
    344.8122, 345.8477, 346.8846, 347.9225, 348.9611, 350, 351.0389, 
    352.0775, 353.1154, 354.1523, 355.1878, 356.2217, 357.2535, 358.283, 
    359.3098, 0.3336662, 1.354252, 2.371273, 3.384442, 4.393482, 5.398128, 
    6.39812, 7.393215, 8.383177, 9.367781, 10.34682, 11.32008, 12.28739, 
    13.24856, 14.20343, 15.15185, 16.09367, 17.02878, 17.95705, 18.87837, 
    19.79265, 20.69982, 21.59979, 22.49251, 23.37793, 24.256, 25.12669, 
    25.98999, 26.84588, 27.69435, 28.53541, 29.36907, 30.19535, 31.01428, 
    31.82589, 32.63021, 33.42731, 34.21722, 35 ;

 grid_lat =
  -35.26439, -35.62921, -35.98892, -36.34341, -36.69255, -37.03624, 
    -37.37434, -37.70675, -38.03334, -38.354, -38.66859, -38.977, -39.27911, 
    -39.57478, -39.8639, -40.14635, -40.42199, -40.69072, -40.9524, 
    -41.20691, -41.45414, -41.69396, -41.92625, -42.15091, -42.36781, 
    -42.57683, -42.77788, -42.97084, -43.1556, -43.33206, -43.50012, 
    -43.65969, -43.81068, -43.95298, -44.08652, -44.21122, -44.32701, 
    -44.4338, -44.53154, -44.62016, -44.6996, -44.76982, -44.83077, 
    -44.88241, -44.9247, -44.95763, -44.98116, -44.99529, -45, -44.99529, 
    -44.98116, -44.95763, -44.9247, -44.88241, -44.83077, -44.76982, 
    -44.6996, -44.62016, -44.53154, -44.4338, -44.32701, -44.21122, 
    -44.08652, -43.95298, -43.81068, -43.65969, -43.50012, -43.33206, 
    -43.1556, -42.97084, -42.77788, -42.57683, -42.36781, -42.15091, 
    -41.92625, -41.69396, -41.45414, -41.20691, -40.9524, -40.69072, 
    -40.42199, -40.14635, -39.8639, -39.57478, -39.27911, -38.977, -38.66859, 
    -38.354, -38.03334, -37.70675, -37.37434, -37.03624, -36.69255, 
    -36.34341, -35.98892, -35.62921, -35.26439,
  -34.52972, -34.89117, -35.24767, -35.59911, -35.94537, -36.28631, 
    -36.62183, -36.95179, -37.27608, -37.59457, -37.90713, -38.21363, 
    -38.51395, -38.80796, -39.09554, -39.37654, -39.65086, -39.91835, 
    -40.1789, -40.43238, -40.67865, -40.9176, -41.14911, -41.37305, -41.5893, 
    -41.79774, -41.99827, -42.19077, -42.37512, -42.55122, -42.71897, 
    -42.87827, -43.02901, -43.17111, -43.30448, -43.42903, -43.54469, 
    -43.65138, -43.74903, -43.83758, -43.91697, -43.98714, -44.04806, 
    -44.09967, -44.14195, -44.17486, -44.19839, -44.21251, -44.21722, 
    -44.21251, -44.19839, -44.17486, -44.14195, -44.09967, -44.04806, 
    -43.98714, -43.91697, -43.83758, -43.74903, -43.65138, -43.54469, 
    -43.42903, -43.30448, -43.17111, -43.02901, -42.87827, -42.71897, 
    -42.55122, -42.37512, -42.19077, -41.99827, -41.79774, -41.5893, 
    -41.37305, -41.14911, -40.9176, -40.67865, -40.43238, -40.1789, 
    -39.91835, -39.65086, -39.37654, -39.09554, -38.80796, -38.51395, 
    -38.21363, -37.90713, -37.59457, -37.27608, -36.95179, -36.62183, 
    -36.28631, -35.94537, -35.59911, -35.24767, -34.89117, -34.52972,
  -33.79504, -34.15289, -34.50594, -34.8541, -35.19722, -35.53519, -35.86789, 
    -36.19517, -36.51693, -36.83301, -37.14331, -37.44768, -37.746, 
    -38.03813, -38.32394, -38.6033, -38.87608, -39.14214, -39.40136, 
    -39.6536, -39.89874, -40.13664, -40.36718, -40.59023, -40.80568, 
    -41.01338, -41.21324, -41.40512, -41.58892, -41.76453, -41.93184, 
    -42.09073, -42.24112, -42.38291, -42.516, -42.64032, -42.75576, 
    -42.86227, -42.95976, -43.04817, -43.12745, -43.19752, -43.25835, 
    -43.3099, -43.35213, -43.385, -43.4085, -43.4226, -43.42731, -43.4226, 
    -43.4085, -43.385, -43.35213, -43.3099, -43.25835, -43.19752, -43.12745, 
    -43.04817, -42.95976, -42.86227, -42.75576, -42.64032, -42.516, 
    -42.38291, -42.24112, -42.09073, -41.93184, -41.76453, -41.58892, 
    -41.40512, -41.21324, -41.01338, -40.80568, -40.59023, -40.36718, 
    -40.13664, -39.89874, -39.6536, -39.40136, -39.14214, -38.87608, 
    -38.6033, -38.32394, -38.03813, -37.746, -37.44768, -37.14331, -36.83301, 
    -36.51693, -36.19517, -35.86789, -35.53519, -35.19722, -34.8541, 
    -34.50594, -34.15289, -33.79504,
  -33.06036, -33.41436, -33.76374, -34.10837, -34.44813, -34.78289, 
    -35.11252, -35.4369, -35.75588, -36.06934, -36.37715, -36.67916, 
    -36.97525, -37.26529, -37.54912, -37.82662, -38.09766, -38.36209, 
    -38.61978, -38.87059, -39.1144, -39.35107, -39.58046, -39.80246, 
    -40.01692, -40.22372, -40.42275, -40.61388, -40.79699, -40.97196, 
    -41.13869, -41.29707, -41.44698, -41.58834, -41.72106, -41.84503, 
    -41.96017, -42.06641, -42.16367, -42.25187, -42.33097, -42.40089, 
    -42.4616, -42.51304, -42.55518, -42.58799, -42.61144, -42.62552, 
    -42.63021, -42.62552, -42.61144, -42.58799, -42.55518, -42.51304, 
    -42.4616, -42.40089, -42.33097, -42.25187, -42.16367, -42.06641, 
    -41.96017, -41.84503, -41.72106, -41.58834, -41.44698, -41.29707, 
    -41.13869, -40.97196, -40.79699, -40.61388, -40.42275, -40.22372, 
    -40.01692, -39.80246, -39.58046, -39.35107, -39.1144, -38.87059, 
    -38.61978, -38.36209, -38.09766, -37.82662, -37.54912, -37.26529, 
    -36.97525, -36.67916, -36.37715, -36.06934, -35.75588, -35.4369, 
    -35.11252, -34.78289, -34.44813, -34.10837, -33.76374, -33.41436, 
    -33.06036,
  -32.32569, -32.67561, -33.02107, -33.36194, -33.6981, -34.02942, -34.35575, 
    -34.67698, -34.99296, -35.30357, -35.60866, -35.90809, -36.20173, 
    -36.48944, -36.77109, -37.04652, -37.3156, -37.57819, -37.83415, 
    -38.08334, -38.32563, -38.56088, -38.78895, -39.00971, -39.22302, 
    -39.42876, -39.6268, -39.81702, -39.99928, -40.17348, -40.3395, 
    -40.49723, -40.64656, -40.78738, -40.91961, -41.04314, -41.15789, 
    -41.26377, -41.36071, -41.44865, -41.5275, -41.59722, -41.65775, 
    -41.70904, -41.75106, -41.78378, -41.80717, -41.82121, -41.82589, 
    -41.82121, -41.80717, -41.78378, -41.75106, -41.70904, -41.65775, 
    -41.59722, -41.5275, -41.44865, -41.36071, -41.26377, -41.15789, 
    -41.04314, -40.91961, -40.78738, -40.64656, -40.49723, -40.3395, 
    -40.17348, -39.99928, -39.81702, -39.6268, -39.42876, -39.22302, 
    -39.00971, -38.78895, -38.56088, -38.32563, -38.08334, -37.83415, 
    -37.57819, -37.3156, -37.04652, -36.77109, -36.48944, -36.20173, 
    -35.90809, -35.60866, -35.30357, -34.99296, -34.67698, -34.35575, 
    -34.02942, -33.6981, -33.36194, -33.02107, -32.67561, -32.32569,
  -31.59101, -31.93662, -32.27793, -32.61481, -32.94714, -33.27477, 
    -33.59758, -33.91543, -34.22818, -34.5357, -34.83784, -35.13448, 
    -35.42545, -35.71062, -35.98985, -36.26299, -36.52991, -36.79046, 
    -37.04449, -37.29186, -37.53244, -37.76608, -37.99264, -38.21198, 
    -38.42397, -38.62848, -38.82537, -39.01452, -39.1958, -39.36908, 
    -39.53426, -39.69121, -39.83982, -39.97999, -40.11162, -40.23461, 
    -40.34887, -40.45432, -40.55087, -40.63845, -40.717, -40.78645, 
    -40.84675, -40.89785, -40.93972, -40.97232, -40.99562, -41.00961, 
    -41.01428, -41.00961, -40.99562, -40.97232, -40.93972, -40.89785, 
    -40.84675, -40.78645, -40.717, -40.63845, -40.55087, -40.45432, 
    -40.34887, -40.23461, -40.11162, -39.97999, -39.83982, -39.69121, 
    -39.53426, -39.36908, -39.1958, -39.01452, -38.82537, -38.62848, 
    -38.42397, -38.21198, -37.99264, -37.76608, -37.53244, -37.29186, 
    -37.04449, -36.79046, -36.52991, -36.26299, -35.98985, -35.71062, 
    -35.42545, -35.13448, -34.83784, -34.5357, -34.22818, -33.91543, 
    -33.59758, -33.27477, -32.94714, -32.61481, -32.27793, -31.93662, 
    -31.59101,
  -30.85634, -31.19741, -31.53433, -31.86699, -32.19525, -32.51897, 
    -32.83802, -33.15226, -33.46156, -33.76576, -34.06473, -34.35833, 
    -34.64641, -34.92882, -35.20542, -35.47607, -35.74061, -35.9989, 
    -36.2508, -36.49615, -36.73482, -36.96666, -37.19153, -37.40928, 
    -37.61977, -37.82288, -38.01846, -38.20639, -38.38652, -38.55875, 
    -38.72294, -38.87898, -39.02676, -39.16616, -39.29708, -39.41943, 
    -39.5331, -39.63801, -39.73409, -39.82125, -39.89942, -39.96855, 
    -40.02857, -40.07944, -40.12112, -40.15358, -40.17678, -40.1907, 
    -40.19535, -40.1907, -40.17678, -40.15358, -40.12112, -40.07944, 
    -40.02857, -39.96855, -39.89942, -39.82125, -39.73409, -39.63801, 
    -39.5331, -39.41943, -39.29708, -39.16616, -39.02676, -38.87898, 
    -38.72294, -38.55875, -38.38652, -38.20639, -38.01846, -37.82288, 
    -37.61977, -37.40928, -37.19153, -36.96666, -36.73482, -36.49615, 
    -36.2508, -35.9989, -35.74061, -35.47607, -35.20542, -34.92882, 
    -34.64641, -34.35833, -34.06473, -33.76576, -33.46156, -33.15226, 
    -32.83802, -32.51897, -32.19525, -31.86699, -31.53433, -31.19741, 
    -30.85634,
  -30.12167, -30.45796, -30.79028, -31.11849, -31.44245, -31.76203, -32.0771, 
    -32.3875, -32.6931, -32.99376, -33.28933, -33.57967, -33.86464, 
    -34.14407, -34.41782, -34.68575, -34.94771, -35.20354, -35.45309, 
    -35.69623, -35.9328, -36.16264, -36.38563, -36.6016, -36.81043, 
    -37.01196, -37.20607, -37.39261, -37.57145, -37.74247, -37.90554, 
    -38.06054, -38.20735, -38.34586, -38.47596, -38.59755, -38.71054, 
    -38.81484, -38.91036, -38.99702, -39.07475, -39.1435, -39.20319, 
    -39.25378, -39.29524, -39.32752, -39.3506, -39.36445, -39.36907, 
    -39.36445, -39.3506, -39.32752, -39.29524, -39.25378, -39.20319, 
    -39.1435, -39.07475, -38.99702, -38.91036, -38.81484, -38.71054, 
    -38.59755, -38.47596, -38.34586, -38.20735, -38.06054, -37.90554, 
    -37.74247, -37.57145, -37.39261, -37.20607, -37.01196, -36.81043, 
    -36.6016, -36.38563, -36.16264, -35.9328, -35.69623, -35.45309, 
    -35.20354, -34.94771, -34.68575, -34.41782, -34.14407, -33.86464, 
    -33.57967, -33.28933, -32.99376, -32.6931, -32.3875, -32.0771, -31.76203, 
    -31.44245, -31.11849, -30.79028, -30.45796, -30.12167,
  -29.38699, -29.7183, -30.04578, -30.36931, -30.68875, -31.00396, -31.31481, 
    -31.62114, -31.92283, -32.21972, -32.51167, -32.79853, -33.08015, 
    -33.35638, -33.62707, -33.89207, -34.15122, -34.40438, -34.6514, 
    -34.89211, -35.12637, -35.35404, -35.57495, -35.78897, -35.99594, 
    -36.19573, -36.38819, -36.57319, -36.75058, -36.92025, -37.08205, 
    -37.23587, -37.38158, -37.51908, -37.64825, -37.76899, -37.8812, 
    -37.98478, -38.07965, -38.16574, -38.24297, -38.31126, -38.37057, 
    -38.42085, -38.46204, -38.49412, -38.51705, -38.53082, -38.53541, 
    -38.53082, -38.51705, -38.49412, -38.46204, -38.42085, -38.37057, 
    -38.31126, -38.24297, -38.16574, -38.07965, -37.98478, -37.8812, 
    -37.76899, -37.64825, -37.51908, -37.38158, -37.23587, -37.08205, 
    -36.92025, -36.75058, -36.57319, -36.38819, -36.19573, -35.99594, 
    -35.78897, -35.57495, -35.35404, -35.12637, -34.89211, -34.6514, 
    -34.40438, -34.15122, -33.89207, -33.62707, -33.35638, -33.08015, 
    -32.79853, -32.51167, -32.21972, -31.92283, -31.62114, -31.31481, 
    -31.00396, -30.68875, -30.36931, -30.04578, -29.7183, -29.38699,
  -28.65232, -28.97841, -29.30084, -29.61947, -29.93416, -30.24478, 
    -30.55118, -30.85322, -31.15076, -31.44366, -31.73176, -32.01491, 
    -32.29297, -32.56578, -32.83318, -33.09504, -33.35118, -33.60146, 
    -33.84572, -34.08381, -34.31557, -34.54086, -34.75951, -34.97139, 
    -35.17633, -35.3742, -35.56485, -35.74813, -35.92393, -36.09208, 
    -36.25248, -36.40498, -36.54947, -36.68583, -36.81395, -36.93372, 
    -37.04504, -37.14782, -37.24197, -37.3274, -37.40405, -37.47184, 
    -37.53071, -37.58062, -37.62151, -37.65335, -37.67612, -37.68979, 
    -37.69435, -37.68979, -37.67612, -37.65335, -37.62151, -37.58062, 
    -37.53071, -37.47184, -37.40405, -37.3274, -37.24197, -37.14782, 
    -37.04504, -36.93372, -36.81395, -36.68583, -36.54947, -36.40498, 
    -36.25248, -36.09208, -35.92393, -35.74813, -35.56485, -35.3742, 
    -35.17633, -34.97139, -34.75951, -34.54086, -34.31557, -34.08381, 
    -33.84572, -33.60146, -33.35118, -33.09504, -32.83318, -32.56578, 
    -32.29297, -32.01491, -31.73176, -31.44366, -31.15076, -30.85322, 
    -30.55118, -30.24478, -29.93416, -29.61947, -29.30084, -28.97841, 
    -28.65232,
  -27.91764, -28.23831, -28.55546, -28.86897, -29.17869, -29.48449, 
    -29.78622, -30.08375, -30.37692, -30.6656, -30.94962, -31.22885, 
    -31.50312, -31.77229, -32.03619, -32.29469, -32.5476, -32.79479, 
    -33.03609, -33.27135, -33.50042, -33.72313, -33.93933, -34.14888, 
    -34.35161, -34.54738, -34.73605, -34.91746, -35.09149, -35.25799, 
    -35.41682, -35.56787, -35.71101, -35.8461, -35.97306, -36.09175, 
    -36.20208, -36.30396, -36.39729, -36.48199, -36.55799, -36.62521, 
    -36.68359, -36.73308, -36.77364, -36.80522, -36.8278, -36.84136, 
    -36.84588, -36.84136, -36.8278, -36.80522, -36.77364, -36.73308, 
    -36.68359, -36.62521, -36.55799, -36.48199, -36.39729, -36.30396, 
    -36.20208, -36.09175, -35.97306, -35.8461, -35.71101, -35.56787, 
    -35.41682, -35.25799, -35.09149, -34.91746, -34.73605, -34.54738, 
    -34.35161, -34.14888, -33.93933, -33.72313, -33.50042, -33.27135, 
    -33.03609, -32.79479, -32.5476, -32.29469, -32.03619, -31.77229, 
    -31.50312, -31.22885, -30.94962, -30.6656, -30.37692, -30.08375, 
    -29.78622, -29.48449, -29.17869, -28.86897, -28.55546, -28.23831, 
    -27.91764,
  -27.18297, -27.49799, -27.80966, -28.11782, -28.42235, -28.72311, 
    -29.01996, -29.31275, -29.60133, -29.88556, -30.16529, -30.44036, 
    -30.71063, -30.97594, -31.23613, -31.49104, -31.74052, -31.98441, 
    -32.22254, -32.45477, -32.68093, -32.90088, -33.11443, -33.32146, 
    -33.5218, -33.7153, -33.90181, -34.08119, -34.25329, -34.41798, 
    -34.57511, -34.72456, -34.8662, -34.99992, -35.12558, -35.24308, 
    -35.35233, -35.45321, -35.54563, -35.62952, -35.70479, -35.77137, 
    -35.8292, -35.87823, -35.91842, -35.94971, -35.97208, -35.98551, 
    -35.98999, -35.98551, -35.97208, -35.94971, -35.91842, -35.87823, 
    -35.8292, -35.77137, -35.70479, -35.62952, -35.54563, -35.45321, 
    -35.35233, -35.24308, -35.12558, -34.99992, -34.8662, -34.72456, 
    -34.57511, -34.41798, -34.25329, -34.08119, -33.90181, -33.7153, 
    -33.5218, -33.32146, -33.11443, -32.90088, -32.68093, -32.45477, 
    -32.22254, -31.98441, -31.74052, -31.49104, -31.23613, -30.97594, 
    -30.71063, -30.44036, -30.16529, -29.88556, -29.60133, -29.31275, 
    -29.01996, -28.72311, -28.42235, -28.11782, -27.80966, -27.49799, 
    -27.18297,
  -26.44829, -26.75747, -27.06343, -27.36604, -27.66517, -27.96067, 
    -28.25241, -28.54023, -28.82401, -29.10357, -29.37879, -29.64949, 
    -29.91554, -30.17676, -30.43301, -30.68413, -30.92996, -31.17034, 
    -31.4051, -31.63409, -31.85715, -32.07413, -32.28485, -32.48917, 
    -32.68693, -32.87798, -33.06216, -33.23934, -33.40936, -33.57207, 
    -33.72735, -33.87507, -34.01508, -34.14728, -34.27153, -34.38773, 
    -34.49578, -34.59556, -34.68699, -34.76999, -34.84446, -34.91034, 
    -34.96757, -35.01609, -35.05586, -35.08683, -35.10897, -35.12226, 
    -35.12669, -35.12226, -35.10897, -35.08683, -35.05586, -35.01609, 
    -34.96757, -34.91034, -34.84446, -34.76999, -34.68699, -34.59556, 
    -34.49578, -34.38773, -34.27153, -34.14728, -34.01508, -33.87507, 
    -33.72735, -33.57207, -33.40936, -33.23934, -33.06216, -32.87798, 
    -32.68693, -32.48917, -32.28485, -32.07413, -31.85715, -31.63409, 
    -31.4051, -31.17034, -30.92996, -30.68413, -30.43301, -30.17676, 
    -29.91554, -29.64949, -29.37879, -29.10357, -28.82401, -28.54023, 
    -28.25241, -27.96067, -27.66517, -27.36604, -27.06343, -26.75747, 
    -26.44829,
  -25.71362, -26.01674, -26.31679, -26.61363, -26.90714, -27.19717, 
    -27.48358, -27.76624, -28.04498, -28.31966, -28.59014, -28.85626, 
    -29.11786, -29.37479, -29.62689, -29.874, -30.11596, -30.35262, -30.5838, 
    -30.80936, -31.02912, -31.24292, -31.45062, -31.65205, -31.84704, 
    -32.03546, -32.21714, -32.39194, -32.55971, -32.7203, -32.87358, 
    -33.01942, -33.15767, -33.28822, -33.41094, -33.52573, -33.63246, 
    -33.73105, -33.8214, -33.90341, -33.97701, -34.04213, -34.0987, 
    -34.14666, -34.18597, -34.21658, -34.23848, -34.25162, -34.256, 
    -34.25162, -34.23848, -34.21658, -34.18597, -34.14666, -34.0987, 
    -34.04213, -33.97701, -33.90341, -33.8214, -33.73105, -33.63246, 
    -33.52573, -33.41094, -33.28822, -33.15767, -33.01942, -32.87358, 
    -32.7203, -32.55971, -32.39194, -32.21714, -32.03546, -31.84704, 
    -31.65205, -31.45062, -31.24292, -31.02912, -30.80936, -30.5838, 
    -30.35262, -30.11596, -29.874, -29.62689, -29.37479, -29.11786, 
    -28.85626, -28.59014, -28.31966, -28.04498, -27.76624, -27.48358, 
    -27.19717, -26.90714, -26.61363, -26.31679, -26.01674, -25.71362,
  -24.97894, -25.2758, -25.56974, -25.86061, -26.14829, -26.43264, -26.71351, 
    -26.99077, -27.26427, -27.53386, -27.79938, -28.0607, -28.31764, 
    -28.57006, -28.81779, -29.06068, -29.29857, -29.5313, -29.75869, 
    -29.9806, -30.19686, -30.4073, -30.61178, -30.81012, -31.00217, 
    -31.18778, -31.36679, -31.53904, -31.7044, -31.86271, -32.01384, 
    -32.15764, -32.29399, -32.42276, -32.54383, -32.65709, -32.76241, 
    -32.85971, -32.94887, -33.02983, -33.10248, -33.16676, -33.22261, 
    -33.26997, -33.30878, -33.33901, -33.36062, -33.3736, -33.37793, 
    -33.3736, -33.36062, -33.33901, -33.30878, -33.26997, -33.22261, 
    -33.16676, -33.10248, -33.02983, -32.94887, -32.85971, -32.76241, 
    -32.65709, -32.54383, -32.42276, -32.29399, -32.15764, -32.01384, 
    -31.86271, -31.7044, -31.53904, -31.36679, -31.18778, -31.00217, 
    -30.81012, -30.61178, -30.4073, -30.19686, -29.9806, -29.75869, -29.5313, 
    -29.29857, -29.06068, -28.81779, -28.57006, -28.31764, -28.0607, 
    -27.79938, -27.53386, -27.26427, -26.99077, -26.71351, -26.43264, 
    -26.14829, -25.86061, -25.56974, -25.2758, -24.97894,
  -24.24427, -24.53467, -24.82229, -25.10699, -25.38863, -25.66709, 
    -25.94222, -26.21387, -26.48191, -26.74619, -27.00655, -27.26284, 
    -27.51491, -27.76261, -28.00576, -28.24422, -28.47782, -28.70641, 
    -28.92981, -29.14787, -29.36043, -29.56732, -29.76838, -29.96344, 
    -30.15236, -30.33498, -30.51114, -30.68068, -30.84346, -30.99933, 
    -31.14815, -31.28979, -31.4241, -31.55096, -31.67025, -31.78186, 
    -31.88566, -31.98156, -32.06945, -32.14926, -32.22089, -32.28428, 
    -32.33934, -32.38604, -32.42432, -32.45413, -32.47544, -32.48825, 
    -32.49251, -32.48825, -32.47544, -32.45413, -32.42432, -32.38604, 
    -32.33934, -32.28428, -32.22089, -32.14926, -32.06945, -31.98156, 
    -31.88566, -31.78186, -31.67025, -31.55096, -31.4241, -31.28979, 
    -31.14815, -30.99933, -30.84346, -30.68068, -30.51114, -30.33498, 
    -30.15236, -29.96344, -29.76838, -29.56732, -29.36043, -29.14787, 
    -28.92981, -28.70641, -28.47782, -28.24422, -28.00576, -27.76261, 
    -27.51491, -27.26284, -27.00655, -26.74619, -26.48191, -26.21387, 
    -25.94222, -25.66709, -25.38863, -25.10699, -24.82229, -24.53467, 
    -24.24427,
  -23.50959, -23.79335, -24.07445, -24.35277, -24.62818, -24.90054, 
    -25.16972, -25.43556, -25.69794, -25.95669, -26.21167, -26.46273, 
    -26.70972, -26.95247, -27.19084, -27.42466, -27.65377, -27.87801, 
    -28.09721, -28.31122, -28.51988, -28.72301, -28.92046, -29.11207, 
    -29.29767, -29.47712, -29.65025, -29.8169, -29.97694, -30.13022, 
    -30.27658, -30.4159, -30.54803, -30.67286, -30.79025, -30.90008, 
    -31.00225, -31.09665, -31.18319, -31.26176, -31.33229, -31.39471, 
    -31.44894, -31.49493, -31.53263, -31.56199, -31.58298, -31.59559, 
    -31.59979, -31.59559, -31.58298, -31.56199, -31.53263, -31.49493, 
    -31.44894, -31.39471, -31.33229, -31.26176, -31.18319, -31.09665, 
    -31.00225, -30.90008, -30.79025, -30.67286, -30.54803, -30.4159, 
    -30.27658, -30.13022, -29.97694, -29.8169, -29.65025, -29.47712, 
    -29.29767, -29.11207, -28.92046, -28.72301, -28.51988, -28.31122, 
    -28.09721, -27.87801, -27.65377, -27.42466, -27.19084, -26.95247, 
    -26.70972, -26.46273, -26.21167, -25.95669, -25.69794, -25.43556, 
    -25.16972, -24.90054, -24.62818, -24.35277, -24.07445, -23.79335, 
    -23.50959,
  -22.77492, -23.05183, -23.32623, -23.59798, -23.86696, -24.13302, 
    -24.39604, -24.65587, -24.91236, -25.16539, -25.41478, -25.6604, 
    -25.9021, -26.13971, -26.37307, -26.60204, -26.82645, -27.04614, 
    -27.26094, -27.47071, -27.67526, -27.87444, -28.06809, -28.25605, 
    -28.43815, -28.61425, -28.78417, -28.94778, -29.10491, -29.25543, 
    -29.39919, -29.53604, -29.66586, -29.78851, -29.90387, -30.01182, 
    -30.11224, -30.20505, -30.29012, -30.36738, -30.43673, -30.49811, 
    -30.55145, -30.59668, -30.63375, -30.66263, -30.68328, -30.69568, 
    -30.69982, -30.69568, -30.68328, -30.66263, -30.63375, -30.59668, 
    -30.55145, -30.49811, -30.43673, -30.36738, -30.29012, -30.20505, 
    -30.11224, -30.01182, -29.90387, -29.78851, -29.66586, -29.53604, 
    -29.39919, -29.25543, -29.10491, -28.94778, -28.78417, -28.61425, 
    -28.43815, -28.25605, -28.06809, -27.87444, -27.67526, -27.47071, 
    -27.26094, -27.04614, -26.82645, -26.60204, -26.37307, -26.13971, 
    -25.9021, -25.6604, -25.41478, -25.16539, -24.91236, -24.65587, 
    -24.39604, -24.13302, -23.86696, -23.59798, -23.32623, -23.05183, 
    -22.77492,
  -22.04024, -22.31014, -22.57764, -22.84263, -23.10497, -23.36455, -23.6212, 
    -23.87482, -24.12524, -24.37232, -24.61593, -24.85591, -25.0921, 
    -25.32435, -25.55252, -25.77643, -25.99593, -26.21087, -26.42107, 
    -26.62638, -26.82663, -27.02167, -27.21133, -27.39545, -27.57387, 
    -27.74643, -27.91298, -28.07337, -28.22743, -28.37503, -28.51603, 
    -28.65027, -28.77763, -28.89797, -29.01118, -29.11712, -29.2157, 
    -29.3068, -29.39032, -29.46618, -29.53428, -29.59455, -29.64693, 
    -29.69135, -29.72776, -29.75613, -29.77641, -29.78859, -29.79265, 
    -29.78859, -29.77641, -29.75613, -29.72776, -29.69135, -29.64693, 
    -29.59455, -29.53428, -29.46618, -29.39032, -29.3068, -29.2157, 
    -29.11712, -29.01118, -28.89797, -28.77763, -28.65027, -28.51603, 
    -28.37503, -28.22743, -28.07337, -27.91298, -27.74643, -27.57387, 
    -27.39545, -27.21133, -27.02167, -26.82663, -26.62638, -26.42107, 
    -26.21087, -25.99593, -25.77643, -25.55252, -25.32435, -25.0921, 
    -24.85591, -24.61593, -24.37232, -24.12524, -23.87482, -23.6212, 
    -23.36455, -23.10497, -22.84263, -22.57764, -22.31014, -22.04024,
  -21.30557, -21.56826, -21.82868, -22.08672, -22.34225, -22.59513, 
    -22.84524, -23.09244, -23.33659, -23.57754, -23.81515, -24.04927, 
    -24.27976, -24.50646, -24.72922, -24.94787, -25.16227, -25.37224, 
    -25.57764, -25.77831, -25.97407, -26.16477, -26.35024, -26.53034, 
    -26.70489, -26.87375, -27.03675, -27.19374, -27.34457, -27.4891, 
    -27.62718, -27.75867, -27.88343, -28.00133, -28.11226, -28.21608, 
    -28.3127, -28.40199, -28.48387, -28.55823, -28.625, -28.6841, -28.73546, 
    -28.77902, -28.81473, -28.84255, -28.86244, -28.87439, -28.87837, 
    -28.87439, -28.86244, -28.84255, -28.81473, -28.77902, -28.73546, 
    -28.6841, -28.625, -28.55823, -28.48387, -28.40199, -28.3127, -28.21608, 
    -28.11226, -28.00133, -27.88343, -27.75867, -27.62718, -27.4891, 
    -27.34457, -27.19374, -27.03675, -26.87375, -26.70489, -26.53034, 
    -26.35024, -26.16477, -25.97407, -25.77831, -25.57764, -25.37224, 
    -25.16227, -24.94787, -24.72922, -24.50646, -24.27976, -24.04927, 
    -23.81515, -23.57754, -23.33659, -23.09244, -22.84524, -22.59513, 
    -22.34225, -22.08672, -21.82868, -21.56826, -21.30557,
  -20.57089, -20.8262, -21.07937, -21.33028, -21.5788, -21.82482, -22.06818, 
    -22.30877, -22.54645, -22.78106, -23.01249, -23.24056, -23.46515, 
    -23.68609, -23.90323, -24.11643, -24.32551, -24.53034, -24.73074, 
    -24.92656, -25.11763, -25.3038, -25.48491, -25.6608, -25.8313, -25.99627, 
    -26.15555, -26.30898, -26.45642, -26.59771, -26.73272, -26.86131, 
    -26.98333, -27.09867, -27.20719, -27.30877, -27.40331, -27.4907, 
    -27.57083, -27.64362, -27.70898, -27.76684, -27.81712, -27.85977, 
    -27.89473, -27.92197, -27.94145, -27.95315, -27.95705, -27.95315, 
    -27.94145, -27.92197, -27.89473, -27.85977, -27.81712, -27.76684, 
    -27.70898, -27.64362, -27.57083, -27.4907, -27.40331, -27.30877, 
    -27.20719, -27.09867, -26.98333, -26.86131, -26.73272, -26.59771, 
    -26.45642, -26.30898, -26.15555, -25.99627, -25.8313, -25.6608, 
    -25.48491, -25.3038, -25.11763, -24.92656, -24.73074, -24.53034, 
    -24.32551, -24.11643, -23.90323, -23.68609, -23.46515, -23.24056, 
    -23.01249, -22.78106, -22.54645, -22.30877, -22.06818, -21.82482, 
    -21.5788, -21.33028, -21.07937, -20.8262, -20.57089,
  -19.83622, -20.08398, -20.32972, -20.57332, -20.81466, -21.05361, 
    -21.29005, -21.52384, -21.75485, -21.98295, -22.20798, -22.42981, 
    -22.6483, -22.86328, -23.07462, -23.28216, -23.48574, -23.68522, 
    -23.88042, -24.0712, -24.2574, -24.43885, -24.6154, -24.7869, -24.95318, 
    -25.11408, -25.26947, -25.41917, -25.56305, -25.70096, -25.83275, 
    -25.95829, -26.07744, -26.19007, -26.29606, -26.39529, -26.48764, 
    -26.57302, -26.65132, -26.72244, -26.78632, -26.84286, -26.892, 
    -26.93369, -26.96786, -26.99449, -27.01353, -27.02497, -27.02878, 
    -27.02497, -27.01353, -26.99449, -26.96786, -26.93369, -26.892, 
    -26.84286, -26.78632, -26.72244, -26.65132, -26.57302, -26.48764, 
    -26.39529, -26.29606, -26.19007, -26.07744, -25.95829, -25.83275, 
    -25.70096, -25.56305, -25.41917, -25.26947, -25.11408, -24.95318, 
    -24.7869, -24.6154, -24.43885, -24.2574, -24.0712, -23.88042, -23.68522, 
    -23.48574, -23.28216, -23.07462, -22.86328, -22.6483, -22.42981, 
    -22.20798, -21.98295, -21.75485, -21.52384, -21.29005, -21.05361, 
    -20.81466, -20.57332, -20.32972, -20.08398, -19.83622,
  -19.10155, -19.34159, -19.57973, -19.81585, -20.04982, -20.28154, 
    -20.51087, -20.73768, -20.96184, -21.18322, -21.40168, -21.61708, 
    -21.82927, -22.03811, -22.24345, -22.44514, -22.64302, -22.83695, 
    -23.02677, -23.21232, -23.39345, -23.57, -23.74181, -23.90874, -24.07061, 
    -24.22728, -24.3786, -24.52441, -24.66457, -24.79893, -24.92736, 
    -25.0497, -25.16584, -25.27564, -25.37897, -25.47573, -25.56579, 
    -25.64905, -25.72542, -25.7948, -25.85711, -25.91227, -25.96022, 
    -26.00089, -26.03424, -26.06021, -26.0788, -26.08995, -26.09367, 
    -26.08995, -26.0788, -26.06021, -26.03424, -26.00089, -25.96022, 
    -25.91227, -25.85711, -25.7948, -25.72542, -25.64905, -25.56579, 
    -25.47573, -25.37897, -25.27564, -25.16584, -25.0497, -24.92736, 
    -24.79893, -24.66457, -24.52441, -24.3786, -24.22728, -24.07061, 
    -23.90874, -23.74181, -23.57, -23.39345, -23.21232, -23.02677, -22.83695, 
    -22.64302, -22.44514, -22.24345, -22.03811, -21.82927, -21.61708, 
    -21.40168, -21.18322, -20.96184, -20.73768, -20.51087, -20.28154, 
    -20.04982, -19.81585, -19.57973, -19.34159, -19.10155,
  -18.36687, -18.59904, -18.82941, -19.05788, -19.28433, -19.50863, 
    -19.73068, -19.95033, -20.16746, -20.38194, -20.59364, -20.80241, 
    -21.00812, -21.21062, -21.40977, -21.60542, -21.79742, -21.98561, 
    -22.16986, -22.35, -22.52588, -22.69734, -22.86423, -23.0264, -23.18369, 
    -23.33596, -23.48304, -23.6248, -23.76108, -23.89175, -24.01665, 
    -24.13567, -24.24865, -24.35549, -24.45604, -24.55021, -24.63787, 
    -24.71892, -24.79326, -24.86081, -24.92148, -24.97519, -25.02188, 
    -25.06149, -25.09396, -25.11926, -25.13736, -25.14822, -25.15185, 
    -25.14822, -25.13736, -25.11926, -25.09396, -25.06149, -25.02188, 
    -24.97519, -24.92148, -24.86081, -24.79326, -24.71892, -24.63787, 
    -24.55021, -24.45604, -24.35549, -24.24865, -24.13567, -24.01665, 
    -23.89175, -23.76108, -23.6248, -23.48304, -23.33596, -23.18369, 
    -23.0264, -22.86423, -22.69734, -22.52588, -22.35, -22.16986, -21.98561, 
    -21.79742, -21.60542, -21.40977, -21.21062, -21.00812, -20.80241, 
    -20.59364, -20.38194, -20.16746, -19.95033, -19.73068, -19.50863, 
    -19.28433, -19.05788, -18.82941, -18.59904, -18.36687,
  -17.63219, -17.85633, -18.07879, -18.29944, -18.51819, -18.73492, -18.9495, 
    -19.16182, -19.37174, -19.57915, -19.7839, -19.98587, -20.18491, 
    -20.38089, -20.57367, -20.76309, -20.94901, -21.13129, -21.30978, 
    -21.48432, -21.65476, -21.82095, -21.98275, -22.13999, -22.29253, 
    -22.44022, -22.5829, -22.72045, -22.85269, -22.97951, -23.10075, 
    -23.21629, -23.32599, -23.42973, -23.52739, -23.61885, -23.704, 
    -23.78273, -23.85496, -23.92059, -23.97954, -24.03174, -24.07711, 
    -24.1156, -24.14717, -24.17175, -24.18934, -24.19991, -24.20343, 
    -24.19991, -24.18934, -24.17175, -24.14717, -24.1156, -24.07711, 
    -24.03174, -23.97954, -23.92059, -23.85496, -23.78273, -23.704, 
    -23.61885, -23.52739, -23.42973, -23.32599, -23.21629, -23.10075, 
    -22.97951, -22.85269, -22.72045, -22.5829, -22.44022, -22.29253, 
    -22.13999, -21.98275, -21.82095, -21.65476, -21.48432, -21.30978, 
    -21.13129, -20.94901, -20.76309, -20.57367, -20.38089, -20.18491, 
    -19.98587, -19.7839, -19.57915, -19.37174, -19.16182, -18.9495, 
    -18.73492, -18.51819, -18.29944, -18.07879, -17.85633, -17.63219,
  -16.89752, -17.11348, -17.32786, -17.54054, -17.75143, -17.96042, 
    -18.16737, -18.37219, -18.57473, -18.77489, -18.97252, -19.16751, 
    -19.35971, -19.54898, -19.7352, -19.91821, -20.09789, -20.27407, 
    -20.44661, -20.61537, -20.7802, -20.94095, -21.09747, -21.24961, 
    -21.39723, -21.54018, -21.6783, -21.81147, -21.93953, -22.06234, 
    -22.17978, -22.2917, -22.39799, -22.49851, -22.59314, -22.68178, 
    -22.76431, -22.84064, -22.91066, -22.97429, -23.03145, -23.08206, 
    -23.12605, -23.16338, -23.19399, -23.21784, -23.2349, -23.24514, 
    -23.24856, -23.24514, -23.2349, -23.21784, -23.19399, -23.16338, 
    -23.12605, -23.08206, -23.03145, -22.97429, -22.91066, -22.84064, 
    -22.76431, -22.68178, -22.59314, -22.49851, -22.39799, -22.2917, 
    -22.17978, -22.06234, -21.93953, -21.81147, -21.6783, -21.54018, 
    -21.39723, -21.24961, -21.09747, -20.94095, -20.7802, -20.61537, 
    -20.44661, -20.27407, -20.09789, -19.91821, -19.7352, -19.54898, 
    -19.35971, -19.16751, -18.97252, -18.77489, -18.57473, -18.37219, 
    -18.16737, -17.96042, -17.75143, -17.54054, -17.32786, -17.11348, 
    -16.89752,
  -16.16285, -16.37048, -16.57663, -16.7812, -16.98408, -17.18516, -17.38433, 
    -17.58147, -17.77647, -17.96921, -18.15956, -18.34738, -18.53256, 
    -18.71496, -18.89445, -19.07088, -19.24412, -19.41402, -19.58045, 
    -19.74325, -19.9023, -20.05743, -20.20851, -20.35538, -20.49791, 
    -20.63595, -20.76936, -20.89799, -21.02171, -21.14038, -21.25386, 
    -21.36204, -21.46477, -21.56195, -21.65344, -21.73915, -21.81896, 
    -21.89278, -21.9605, -22.02205, -22.07734, -22.1263, -22.16886, 
    -22.20498, -22.23459, -22.25766, -22.27417, -22.28408, -22.28739, 
    -22.28408, -22.27417, -22.25766, -22.23459, -22.20498, -22.16886, 
    -22.1263, -22.07734, -22.02205, -21.9605, -21.89278, -21.81896, 
    -21.73915, -21.65344, -21.56195, -21.46477, -21.36204, -21.25386, 
    -21.14038, -21.02171, -20.89799, -20.76936, -20.63595, -20.49791, 
    -20.35538, -20.20851, -20.05743, -19.9023, -19.74325, -19.58045, 
    -19.41402, -19.24412, -19.07088, -18.89445, -18.71496, -18.53256, 
    -18.34738, -18.15956, -17.96921, -17.77647, -17.58147, -17.38433, 
    -17.18516, -16.98408, -16.7812, -16.57663, -16.37048, -16.16285,
  -15.42817, -15.62734, -15.82513, -16.02143, -16.21614, -16.40917, -16.6004, 
    -16.78971, -16.97701, -17.16216, -17.34505, -17.52556, -17.70355, 
    -17.8789, -18.05148, -18.22116, -18.38779, -18.55125, -18.71139, 
    -18.86807, -19.02115, -19.1705, -19.31597, -19.45741, -19.59469, 
    -19.72766, -19.85619, -19.98014, -20.09937, -20.21375, -20.32315, 
    -20.42744, -20.5265, -20.6202, -20.70844, -20.79111, -20.8681, -20.9393, 
    -21.00464, -21.06402, -21.11737, -21.16462, -21.20569, -21.24054, 
    -21.26912, -21.29139, -21.30732, -21.31689, -21.32008, -21.31689, 
    -21.30732, -21.29139, -21.26912, -21.24054, -21.20569, -21.16462, 
    -21.11737, -21.06402, -21.00464, -20.9393, -20.8681, -20.79111, 
    -20.70844, -20.6202, -20.5265, -20.42744, -20.32315, -20.21375, 
    -20.09937, -19.98014, -19.85619, -19.72766, -19.59469, -19.45741, 
    -19.31597, -19.1705, -19.02115, -18.86807, -18.71139, -18.55125, 
    -18.38779, -18.22116, -18.05148, -17.8789, -17.70355, -17.52556, 
    -17.34505, -17.16216, -16.97701, -16.78971, -16.6004, -16.40917, 
    -16.21614, -16.02143, -15.82513, -15.62734, -15.42817,
  -14.6935, -14.88407, -15.07335, -15.26124, -15.44765, -15.63248, -15.81561, 
    -15.99695, -16.17639, -16.3538, -16.52908, -16.7021, -16.87274, 
    -17.04088, -17.20639, -17.36914, -17.52901, -17.68585, -17.83953, 
    -17.98992, -18.13688, -18.28028, -18.41997, -18.55582, -18.68769, 
    -18.81544, -18.93895, -19.05806, -19.17266, -19.28261, -19.38778, 
    -19.48806, -19.58331, -19.67343, -19.7583, -19.83782, -19.91188, 
    -19.98038, -20.04325, -20.10039, -20.15172, -20.19719, -20.23672, 
    -20.27026, -20.29777, -20.3192, -20.33454, -20.34374, -20.34682, 
    -20.34374, -20.33454, -20.3192, -20.29777, -20.27026, -20.23672, 
    -20.19719, -20.15172, -20.10039, -20.04325, -19.98038, -19.91188, 
    -19.83782, -19.7583, -19.67343, -19.58331, -19.48806, -19.38778, 
    -19.28261, -19.17266, -19.05806, -18.93895, -18.81544, -18.68769, 
    -18.55582, -18.41997, -18.28028, -18.13688, -17.98992, -17.83953, 
    -17.68585, -17.52901, -17.36914, -17.20639, -17.04088, -16.87274, 
    -16.7021, -16.52908, -16.3538, -16.17639, -15.99695, -15.81561, 
    -15.63248, -15.44765, -15.26124, -15.07335, -14.88407, -14.6935,
  -13.95882, -14.14067, -14.32132, -14.50067, -14.67863, -14.85512, 
    -15.03002, -15.20323, -15.37465, -15.54417, -15.71168, -15.87706, 
    -16.0402, -16.20097, -16.35925, -16.51492, -16.66785, -16.81791, 
    -16.96498, -17.10892, -17.2496, -17.38689, -17.52065, -17.65075, 
    -17.77705, -17.89944, -18.01776, -18.1319, -18.24172, -18.34711, 
    -18.44792, -18.54405, -18.63538, -18.7218, -18.80319, -18.87945, 
    -18.95048, -19.0162, -19.0765, -19.13132, -19.18058, -19.2242, -19.26213, 
    -19.29432, -19.32071, -19.34128, -19.356, -19.36483, -19.36778, 
    -19.36483, -19.356, -19.34128, -19.32071, -19.29432, -19.26213, -19.2242, 
    -19.18058, -19.13132, -19.0765, -19.0162, -18.95048, -18.87945, 
    -18.80319, -18.7218, -18.63538, -18.54405, -18.44792, -18.34711, 
    -18.24172, -18.1319, -18.01776, -17.89944, -17.77705, -17.65075, 
    -17.52065, -17.38689, -17.2496, -17.10892, -16.96498, -16.81791, 
    -16.66785, -16.51492, -16.35925, -16.20097, -16.0402, -15.87706, 
    -15.71168, -15.54417, -15.37465, -15.20323, -15.03002, -14.85512, 
    -14.67863, -14.50067, -14.32132, -14.14067, -13.95882,
  -13.22415, -13.39715, -13.56903, -13.73972, -13.90911, -14.07711, 
    -14.24364, -14.40859, -14.57185, -14.73334, -14.89293, -15.05052, 
    -15.20599, -15.35924, -15.51014, -15.65857, -15.80442, -15.94755, 
    -16.08784, -16.22518, -16.35942, -16.49044, -16.61812, -16.74232, 
    -16.86292, -16.97978, -17.09279, -17.20181, -17.30672, -17.4074, 
    -17.50373, -17.5956, -17.68288, -17.76548, -17.84328, -17.91618, 
    -17.9841, -18.04693, -18.1046, -18.15702, -18.20412, -18.24584, 
    -18.28212, -18.31291, -18.33815, -18.35783, -18.3719, -18.38036, 
    -18.38318, -18.38036, -18.3719, -18.35783, -18.33815, -18.31291, 
    -18.28212, -18.24584, -18.20412, -18.15702, -18.1046, -18.04693, 
    -17.9841, -17.91618, -17.84328, -17.76548, -17.68288, -17.5956, 
    -17.50373, -17.4074, -17.30672, -17.20181, -17.09279, -16.97978, 
    -16.86292, -16.74232, -16.61812, -16.49044, -16.35942, -16.22518, 
    -16.08784, -15.94755, -15.80442, -15.65857, -15.51014, -15.35924, 
    -15.20599, -15.05052, -14.89293, -14.73334, -14.57185, -14.40859, 
    -14.24364, -14.07711, -13.90911, -13.73972, -13.56903, -13.39715, 
    -13.22415,
  -12.48947, -12.65351, -12.81652, -12.97841, -13.1391, -13.2985, -13.45652, 
    -13.61306, -13.76804, -13.92135, -14.07288, -14.22254, -14.37021, 
    -14.51579, -14.65916, -14.8002, -14.93881, -15.07486, -15.20823, 
    -15.33881, -15.46647, -15.59108, -15.71253, -15.83068, -15.94542, 
    -16.05663, -16.16418, -16.26795, -16.36782, -16.46367, -16.55539, 
    -16.64287, -16.72599, -16.80466, -16.87877, -16.94822, -17.01292, 
    -17.07278, -17.12773, -17.17768, -17.22256, -17.26232, -17.2969, 
    -17.32624, -17.3503, -17.36906, -17.38247, -17.39053, -17.39322, 
    -17.39053, -17.38247, -17.36906, -17.3503, -17.32624, -17.2969, 
    -17.26232, -17.22256, -17.17768, -17.12773, -17.07278, -17.01292, 
    -16.94822, -16.87877, -16.80466, -16.72599, -16.64287, -16.55539, 
    -16.46367, -16.36782, -16.26795, -16.16418, -16.05663, -15.94542, 
    -15.83068, -15.71253, -15.59108, -15.46647, -15.33881, -15.20823, 
    -15.07486, -14.93881, -14.8002, -14.65916, -14.51579, -14.37021, 
    -14.22254, -14.07288, -13.92135, -13.76804, -13.61306, -13.45652, 
    -13.2985, -13.1391, -12.97841, -12.81652, -12.65351, -12.48947,
  -11.7548, -11.90976, -12.06378, -12.21676, -12.36863, -12.5193, -12.66869, 
    -12.81671, -12.96326, -13.10826, -13.2516, -13.39319, -13.53292, 
    -13.67069, -13.80638, -13.9399, -14.07113, -14.19996, -14.32627, 
    -14.44994, -14.57087, -14.68893, -14.804, -14.91598, -15.02473, 
    -15.13014, -15.2321, -15.33048, -15.42518, -15.51608, -15.60307, 
    -15.68605, -15.7649, -15.83954, -15.90985, -15.97575, -16.03714, 
    -16.09396, -16.1461, -16.19351, -16.23612, -16.27386, -16.30668, 
    -16.33454, -16.35738, -16.37519, -16.38792, -16.39557, -16.39812, 
    -16.39557, -16.38792, -16.37519, -16.35738, -16.33454, -16.30668, 
    -16.27386, -16.23612, -16.19351, -16.1461, -16.09396, -16.03714, 
    -15.97575, -15.90985, -15.83954, -15.7649, -15.68605, -15.60307, 
    -15.51608, -15.42518, -15.33048, -15.2321, -15.13014, -15.02473, 
    -14.91598, -14.804, -14.68893, -14.57087, -14.44994, -14.32627, 
    -14.19996, -14.07113, -13.9399, -13.80638, -13.67069, -13.53292, 
    -13.39319, -13.2516, -13.10826, -12.96326, -12.81671, -12.66869, 
    -12.5193, -12.36863, -12.21676, -12.06378, -11.90976, -11.7548,
  -11.02012, -11.16591, -11.31083, -11.45479, -11.59772, -11.73955, 
    -11.88019, -12.01956, -12.15757, -12.29414, -12.42916, -12.56255, 
    -12.6942, -12.82403, -12.95192, -13.07777, -13.20149, -13.32295, 
    -13.44206, -13.5587, -13.67276, -13.78413, -13.8927, -13.99836, 
    -14.10098, -14.20047, -14.29671, -14.38959, -14.479, -14.56483, 
    -14.64697, -14.72534, -14.79981, -14.87031, -14.93673, -14.99899, 
    -15.05699, -15.11067, -15.15995, -15.20475, -15.24501, -15.28068, 
    -15.3117, -15.33803, -15.35962, -15.37645, -15.38849, -15.39572, 
    -15.39813, -15.39572, -15.38849, -15.37645, -15.35962, -15.33803, 
    -15.3117, -15.28068, -15.24501, -15.20475, -15.15995, -15.11067, 
    -15.05699, -14.99899, -14.93673, -14.87031, -14.79981, -14.72534, 
    -14.64697, -14.56483, -14.479, -14.38959, -14.29671, -14.20047, 
    -14.10098, -13.99836, -13.8927, -13.78413, -13.67276, -13.5587, 
    -13.44206, -13.32295, -13.20149, -13.07777, -12.95192, -12.82403, 
    -12.6942, -12.56255, -12.42916, -12.29414, -12.15757, -12.01956, 
    -11.88019, -11.73955, -11.59772, -11.45479, -11.31083, -11.16591, 
    -11.02012,
  -10.28545, -10.42197, -10.55768, -10.69252, -10.82641, -10.95929, 
    -11.09107, -11.22167, -11.35102, -11.47903, -11.60561, -11.73068, 
    -11.85414, -11.97589, -12.09585, -12.21391, -12.32998, -12.44396, 
    -12.55573, -12.66521, -12.77227, -12.87683, -12.97877, -13.07798, 
    -13.17436, -13.2678, -13.3582, -13.44545, -13.52945, -13.61009, 
    -13.68729, -13.76093, -13.83093, -13.89719, -13.95963, -14.01815, 
    -14.07269, -14.12316, -14.16949, -14.21162, -14.24948, -14.28303, 
    -14.3122, -14.33696, -14.35726, -14.37309, -14.38441, -14.39121, 
    -14.39348, -14.39121, -14.38441, -14.37309, -14.35726, -14.33696, 
    -14.3122, -14.28303, -14.24948, -14.21162, -14.16949, -14.12316, 
    -14.07269, -14.01815, -13.95963, -13.89719, -13.83093, -13.76093, 
    -13.68729, -13.61009, -13.52945, -13.44545, -13.3582, -13.2678, 
    -13.17436, -13.07798, -12.97877, -12.87683, -12.77227, -12.66521, 
    -12.55573, -12.44396, -12.32998, -12.21391, -12.09585, -11.97589, 
    -11.85414, -11.73068, -11.60561, -11.47903, -11.35102, -11.22167, 
    -11.09107, -10.95929, -10.82641, -10.69252, -10.55768, -10.42197, 
    -10.28545,
  -9.550773, -9.677926, -9.804344, -9.929964, -10.05472, -10.17854, 
    -10.30135, -10.42309, -10.54366, -10.66301, -10.78103, -10.89766, 
    -11.0128, -11.12637, -11.23828, -11.34843, -11.45673, -11.5631, 
    -11.66742, -11.7696, -11.86955, -11.96717, -12.06235, -12.155, -12.24501, 
    -12.33229, -12.41673, -12.49824, -12.57673, -12.65208, -12.72422, 
    -12.79304, -12.85847, -12.9204, -12.97877, -13.03348, -13.08447, 
    -13.13165, -13.17497, -13.21437, -13.24977, -13.28114, -13.30842, 
    -13.33158, -13.35057, -13.36537, -13.37596, -13.38232, -13.38444, 
    -13.38232, -13.37596, -13.36537, -13.35057, -13.33158, -13.30842, 
    -13.28114, -13.24977, -13.21437, -13.17497, -13.13165, -13.08447, 
    -13.03348, -12.97877, -12.9204, -12.85847, -12.79304, -12.72422, 
    -12.65208, -12.57673, -12.49824, -12.41673, -12.33229, -12.24501, 
    -12.155, -12.06235, -11.96717, -11.86955, -11.7696, -11.66742, -11.5631, 
    -11.45673, -11.34843, -11.23828, -11.12637, -11.0128, -10.89766, 
    -10.78103, -10.66301, -10.54366, -10.42309, -10.30135, -10.17854, 
    -10.05472, -9.929964, -9.804344, -9.677926, -9.550773,
  -8.816097, -8.933801, -9.050837, -9.167146, -9.282667, -9.397336, 
    -9.511086, -9.623848, -9.735553, -9.846126, -9.955491, -10.06357, 
    -10.17029, -10.27556, -10.3793, -10.48143, -10.58185, -10.68048, 
    -10.77724, -10.87202, -10.96474, -11.0553, -11.14361, -11.22959, 
    -11.31312, -11.39412, -11.47251, -11.54817, -11.62103, -11.691, 
    -11.75798, -11.82189, -11.88264, -11.94017, -11.99438, -12.0452, 
    -12.09256, -12.1364, -12.17664, -12.21324, -12.24614, -12.27528, 
    -12.30063, -12.32215, -12.3398, -12.35355, -12.36339, -12.3693, 
    -12.37127, -12.3693, -12.36339, -12.35355, -12.3398, -12.32215, 
    -12.30063, -12.27528, -12.24614, -12.21324, -12.17664, -12.1364, 
    -12.09256, -12.0452, -11.99438, -11.94017, -11.88264, -11.82189, 
    -11.75798, -11.691, -11.62103, -11.54817, -11.47251, -11.39412, 
    -11.31312, -11.22959, -11.14361, -11.0553, -10.96474, -10.87202, 
    -10.77724, -10.68048, -10.58185, -10.48143, -10.3793, -10.27556, 
    -10.17029, -10.06357, -9.955491, -9.846126, -9.735553, -9.623848, 
    -9.511086, -9.397336, -9.282667, -9.167146, -9.050837, -8.933801, 
    -8.816097,
  -8.081423, -8.189597, -8.297169, -8.404083, -8.510284, -8.615713, 
    -8.720308, -8.824006, -8.926742, -9.028447, -9.129053, -9.228487, 
    -9.326677, -9.423547, -9.519018, -9.613013, -9.705451, -9.79625, 
    -9.885328, -9.972599, -10.05798, -10.14138, -10.22272, -10.30191, 
    -10.37886, -10.45349, -10.52571, -10.59543, -10.66257, -10.72705, 
    -10.78878, -10.84769, -10.90369, -10.95672, -11.0067, -11.05355, 
    -11.09722, -11.13764, -11.17476, -11.2085, -11.23884, -11.26572, 
    -11.2891, -11.30894, -11.32522, -11.33791, -11.34698, -11.35243, 
    -11.35425, -11.35243, -11.34698, -11.33791, -11.32522, -11.30894, 
    -11.2891, -11.26572, -11.23884, -11.2085, -11.17476, -11.13764, 
    -11.09722, -11.05355, -11.0067, -10.95672, -10.90369, -10.84769, 
    -10.78878, -10.72705, -10.66257, -10.59543, -10.52571, -10.45349, 
    -10.37886, -10.30191, -10.22272, -10.14138, -10.05798, -9.972599, 
    -9.885328, -9.79625, -9.705451, -9.613013, -9.519018, -9.423547, 
    -9.326677, -9.228487, -9.129053, -9.028447, -8.926742, -8.824006, 
    -8.720308, -8.615713, -8.510284, -8.404083, -8.297169, -8.189597, 
    -8.081423,
  -7.346748, -7.445321, -7.543353, -7.640796, -7.737598, -7.833705, 
    -7.929061, -8.023608, -8.117288, -8.210036, -8.30179, -8.392486, 
    -8.482054, -8.570426, -8.657532, -8.743299, -8.827652, -8.910519, 
    -8.99182, -9.071482, -9.149424, -9.225567, -9.299832, -9.372141, 
    -9.442413, -9.510569, -9.576528, -9.640213, -9.701547, -9.760451, 
    -9.816853, -9.870676, -9.92185, -9.970306, -10.01598, -10.0588, 
    -10.09871, -10.13566, -10.16958, -10.20043, -10.22816, -10.25273, 
    -10.2741, -10.29224, -10.30712, -10.31872, -10.32702, -10.332, -10.33367, 
    -10.332, -10.32702, -10.31872, -10.30712, -10.29224, -10.2741, -10.25273, 
    -10.22816, -10.20043, -10.16958, -10.13566, -10.09871, -10.0588, 
    -10.01598, -9.970306, -9.92185, -9.870676, -9.816853, -9.760451, 
    -9.701547, -9.640213, -9.576528, -9.510569, -9.442413, -9.372141, 
    -9.299832, -9.225567, -9.149424, -9.071482, -8.99182, -8.910519, 
    -8.827652, -8.743299, -8.657532, -8.570426, -8.482054, -8.392486, 
    -8.30179, -8.210036, -8.117288, -8.023608, -7.929061, -7.833705, 
    -7.737598, -7.640796, -7.543353, -7.445321, -7.346748,
  -6.612073, -6.700978, -6.789403, -6.877304, -6.964634, -7.051345, 
    -7.137385, -7.222704, -7.307246, -7.390956, -7.473776, -7.555646, 
    -7.636507, -7.716295, -7.794946, -7.872395, -7.948575, -8.023417, 
    -8.096853, -8.168813, -8.239225, -8.308019, -8.375121, -8.44046, 
    -8.503963, -8.565559, -8.625175, -8.682739, -8.738181, -8.791431, 
    -8.842422, -8.891085, -8.937356, -8.981172, -9.02247, -9.061195, 
    -9.097291, -9.130703, -9.161384, -9.189286, -9.21437, -9.236594, 
    -9.255927, -9.272337, -9.285798, -9.29629, -9.303797, -9.308306, 
    -9.30981, -9.308306, -9.303797, -9.29629, -9.285798, -9.272337, 
    -9.255927, -9.236594, -9.21437, -9.189286, -9.161384, -9.130703, 
    -9.097291, -9.061195, -9.02247, -8.981172, -8.937356, -8.891085, 
    -8.842422, -8.791431, -8.738181, -8.682739, -8.625175, -8.565559, 
    -8.503963, -8.44046, -8.375121, -8.308019, -8.239225, -8.168813, 
    -8.096853, -8.023417, -7.948575, -7.872395, -7.794946, -7.716295, 
    -7.636507, -7.555646, -7.473776, -7.390956, -7.307246, -7.222704, 
    -7.137385, -7.051345, -6.964634, -6.877304, -6.789403, -6.700978, 
    -6.612073,
  -5.877398, -5.956575, -6.035332, -6.113627, -6.19142, -6.268667, -6.345323, 
    -6.421341, -6.496675, -6.571271, -6.645081, -6.718051, -6.790126, 
    -6.86125, -6.931367, -7.000417, -7.068341, -7.135077, -7.200565, 
    -7.26474, -7.327541, -7.388902, -7.448759, -7.507047, -7.563702, 
    -7.618658, -7.671851, -7.723217, -7.772693, -7.820215, -7.865723, 
    -7.909157, -7.950458, -7.989569, -8.026436, -8.061007, -8.09323, 
    -8.123061, -8.150454, -8.175366, -8.197762, -8.217607, -8.23487, 
    -8.249522, -8.261543, -8.270913, -8.277617, -8.281642, -8.282985, 
    -8.281642, -8.277617, -8.270913, -8.261543, -8.249522, -8.23487, 
    -8.217607, -8.197762, -8.175366, -8.150454, -8.123061, -8.09323, 
    -8.061007, -8.026436, -7.989569, -7.950458, -7.909157, -7.865723, 
    -7.820215, -7.772693, -7.723217, -7.671851, -7.618658, -7.563702, 
    -7.507047, -7.448759, -7.388902, -7.327541, -7.26474, -7.200565, 
    -7.135077, -7.068341, -7.000417, -6.931367, -6.86125, -6.790126, 
    -6.718051, -6.645081, -6.571271, -6.496675, -6.421341, -6.345323, 
    -6.268667, -6.19142, -6.113627, -6.035332, -5.956575, -5.877398,
  -5.142724, -5.21212, -5.281153, -5.349786, -5.417983, -5.485706, -5.552916, 
    -5.619571, -5.68563, -5.751048, -5.815781, -5.87978, -5.943, -6.00539, 
    -6.066901, -6.12748, -6.187074, -6.245632, -6.303097, -6.359414, 
    -6.414529, -6.468383, -6.520922, -6.572086, -6.621819, -6.670065, 
    -6.716765, -6.761864, -6.805305, -6.847034, -6.886996, -6.925138, 
    -6.96141, -6.995759, -7.02814, -7.058504, -7.086808, -7.113011, 
    -7.137073, -7.158958, -7.178632, -7.196066, -7.211231, -7.224104, 
    -7.234665, -7.242897, -7.248786, -7.252323, -7.253503, -7.252323, 
    -7.248786, -7.242897, -7.234665, -7.224104, -7.211231, -7.196066, 
    -7.178632, -7.158958, -7.137073, -7.113011, -7.086808, -7.058504, 
    -7.02814, -6.995759, -6.96141, -6.925138, -6.886996, -6.847034, 
    -6.805305, -6.761864, -6.716765, -6.670065, -6.621819, -6.572086, 
    -6.520922, -6.468383, -6.414529, -6.359414, -6.303097, -6.245632, 
    -6.187074, -6.12748, -6.066901, -6.00539, -5.943, -5.87978, -5.815781, 
    -5.751048, -5.68563, -5.619571, -5.552916, -5.485706, -5.417983, 
    -5.349786, -5.281153, -5.21212, -5.142724,
  -4.408049, -4.467618, -4.526879, -4.5858, -4.64435, -4.702497, -4.760206, 
    -4.817443, -4.874171, -4.930352, -4.985948, -5.040917, -5.095221, 
    -5.148814, -5.201655, -5.253699, -5.304901, -5.355214, -5.404592, 
    -5.452987, -5.50035, -5.546633, -5.591787, -5.635764, -5.678512, 
    -5.719984, -5.760129, -5.7989, -5.836247, -5.872125, -5.906484, 
    -5.939281, -5.970469, -6.000007, -6.027852, -6.053965, -6.078306, 
    -6.100842, -6.121536, -6.140359, -6.157281, -6.172276, -6.18532, 
    -6.196393, -6.205477, -6.212557, -6.217623, -6.220666, -6.221681, 
    -6.220666, -6.217623, -6.212557, -6.205477, -6.196393, -6.18532, 
    -6.172276, -6.157281, -6.140359, -6.121536, -6.100842, -6.078306, 
    -6.053965, -6.027852, -6.000007, -5.970469, -5.939281, -5.906484, 
    -5.872125, -5.836247, -5.7989, -5.760129, -5.719984, -5.678512, 
    -5.635764, -5.591787, -5.546633, -5.50035, -5.452987, -5.404592, 
    -5.355214, -5.304901, -5.253699, -5.201655, -5.148814, -5.095221, 
    -5.040917, -4.985948, -4.930352, -4.874171, -4.817443, -4.760206, 
    -4.702497, -4.64435, -4.5858, -4.526879, -4.467618, -4.408049,
  -3.673374, -3.723077, -3.772523, -3.82169, -3.870549, -3.919074, -3.967237, 
    -4.015007, -4.062356, -4.10925, -4.155657, -4.201545, -4.246879, 
    -4.291623, -4.335741, -4.379195, -4.421948, -4.463961, -4.505196, 
    -4.545611, -4.585167, -4.623823, -4.661538, -4.69827, -4.733978, 
    -4.768622, -4.802159, -4.834549, -4.865752, -4.895727, -4.924435, 
    -4.951838, -4.977899, -5.002581, -5.025849, -5.047671, -5.068013, 
    -5.086846, -5.104141, -5.119872, -5.134015, -5.146547, -5.15745, 
    -5.166705, -5.174297, -5.180215, -5.184449, -5.186993, -5.187841, 
    -5.186993, -5.184449, -5.180215, -5.174297, -5.166705, -5.15745, 
    -5.146547, -5.134015, -5.119872, -5.104141, -5.086846, -5.068013, 
    -5.047671, -5.025849, -5.002581, -4.977899, -4.951838, -4.924435, 
    -4.895727, -4.865752, -4.834549, -4.802159, -4.768622, -4.733978, 
    -4.69827, -4.661538, -4.623823, -4.585167, -4.545611, -4.505196, 
    -4.463961, -4.421948, -4.379195, -4.335741, -4.291623, -4.246879, 
    -4.201545, -4.155657, -4.10925, -4.062356, -4.015007, -3.967237, 
    -3.919074, -3.870549, -3.82169, -3.772523, -3.723077, -3.673374,
  -2.938699, -2.978501, -3.0181, -3.057476, -3.096608, -3.135473, -3.17405, 
    -3.212315, -3.250242, -3.287808, -3.324986, -3.361748, -3.398068, 
    -3.433917, -3.469266, -3.504085, -3.538343, -3.57201, -3.605054, 
    -3.637443, -3.669145, -3.700126, -3.730354, -3.759796, -3.788419, 
    -3.816189, -3.843073, -3.869038, -3.894052, -3.918083, -3.941099, 
    -3.963069, -3.983964, -4.003754, -4.022411, -4.039908, -4.05622, 
    -4.071321, -4.08519, -4.097805, -4.109146, -4.119196, -4.127939, 
    -4.135361, -4.14145, -4.146196, -4.149592, -4.151631, -4.152311, 
    -4.151631, -4.149592, -4.146196, -4.14145, -4.135361, -4.127939, 
    -4.119196, -4.109146, -4.097805, -4.08519, -4.071321, -4.05622, 
    -4.039908, -4.022411, -4.003754, -3.983964, -3.963069, -3.941099, 
    -3.918083, -3.894052, -3.869038, -3.843073, -3.816189, -3.788419, 
    -3.759796, -3.730354, -3.700126, -3.669145, -3.637443, -3.605054, 
    -3.57201, -3.538343, -3.504085, -3.469266, -3.433917, -3.398068, 
    -3.361748, -3.324986, -3.287808, -3.250242, -3.212315, -3.17405, 
    -3.135473, -3.096608, -3.057476, -3.0181, -2.978501, -2.938699,
  -2.204024, -2.233899, -2.263623, -2.29318, -2.322554, -2.35173, -2.38069, 
    -2.409416, -2.437891, -2.466094, -2.494007, -2.52161, -2.548881, 
    -2.575799, -2.602343, -2.628489, -2.654216, -2.679499, -2.704315, 
    -2.72864, -2.752449, -2.775718, -2.798423, -2.820537, -2.842036, 
    -2.862896, -2.883091, -2.902596, -2.921387, -2.93944, -2.956731, 
    -2.973237, -2.988935, -3.003803, -3.017821, -3.030967, -3.043222, 
    -3.054569, -3.06499, -3.074468, -3.08299, -3.090542, -3.097111, 
    -3.102689, -3.107264, -3.11083, -3.113382, -3.114914, -3.115426, 
    -3.114914, -3.113382, -3.11083, -3.107264, -3.102689, -3.097111, 
    -3.090542, -3.08299, -3.074468, -3.06499, -3.054569, -3.043222, 
    -3.030967, -3.017821, -3.003803, -2.988935, -2.973237, -2.956731, 
    -2.93944, -2.921387, -2.902596, -2.883091, -2.862896, -2.842036, 
    -2.820537, -2.798423, -2.775718, -2.752449, -2.72864, -2.704315, 
    -2.679499, -2.654216, -2.628489, -2.602343, -2.575799, -2.548881, 
    -2.52161, -2.494007, -2.466094, -2.437891, -2.409416, -2.38069, -2.35173, 
    -2.322554, -2.29318, -2.263623, -2.233899, -2.204024,
  -1.46935, -1.489277, -1.509105, -1.528821, -1.548416, -1.56788, -1.587199, 
    -1.606363, -1.62536, -1.644176, -1.662799, -1.681216, -1.699411, 
    -1.717372, -1.735083, -1.752529, -1.769696, -1.786567, -1.803126, 
    -1.819359, -1.835248, -1.850776, -1.865928, -1.880687, -1.895035, 
    -1.908957, -1.922435, -1.935454, -1.947996, -1.960045, -1.971586, 
    -1.982603, -1.993082, -2.003006, -2.012363, -2.021138, -2.029319, 
    -2.036894, -2.04385, -2.050177, -2.055866, -2.060907, -2.065293, 
    -2.069016, -2.07207, -2.074451, -2.076154, -2.077178, -2.077519, 
    -2.077178, -2.076154, -2.074451, -2.07207, -2.069016, -2.065293, 
    -2.060907, -2.055866, -2.050177, -2.04385, -2.036894, -2.029319, 
    -2.021138, -2.012363, -2.003006, -1.993082, -1.982603, -1.971586, 
    -1.960045, -1.947996, -1.935454, -1.922435, -1.908957, -1.895035, 
    -1.880687, -1.865928, -1.850776, -1.835248, -1.819359, -1.803126, 
    -1.786567, -1.769696, -1.752529, -1.735083, -1.717372, -1.699411, 
    -1.681216, -1.662799, -1.644176, -1.62536, -1.606363, -1.587199, 
    -1.56788, -1.548416, -1.528821, -1.509105, -1.489277, -1.46935,
  -0.7346748, -0.744642, -0.7545591, -0.7644209, -0.7742223, -0.7839577, 
    -0.7936214, -0.8032075, -0.8127099, -0.8221223, -0.8314381, -0.8406506, 
    -0.8497528, -0.8587376, -0.8675976, -0.8763254, -0.8849133, -0.8933536, 
    -0.9016382, -0.9097592, -0.9177083, -0.9254774, -0.9330581, -0.9404421, 
    -0.947621, -0.9545865, -0.9613302, -0.9678438, -0.9741191, -0.9801481, 
    -0.9859229, -0.9914355, -0.9966785, -1.001644, -1.006326, -1.010717, 
    -1.014811, -1.018601, -1.022082, -1.025248, -1.028095, -1.030618, 
    -1.032812, -1.034675, -1.036204, -1.037395, -1.038247, -1.038759, 
    -1.03893, -1.038759, -1.038247, -1.037395, -1.036204, -1.034675, 
    -1.032812, -1.030618, -1.028095, -1.025248, -1.022082, -1.018601, 
    -1.014811, -1.010717, -1.006326, -1.001644, -0.9966785, -0.9914355, 
    -0.9859229, -0.9801481, -0.9741191, -0.9678438, -0.9613302, -0.9545865, 
    -0.947621, -0.9404421, -0.9330581, -0.9254774, -0.9177083, -0.9097592, 
    -0.9016382, -0.8933536, -0.8849133, -0.8763254, -0.8675976, -0.8587376, 
    -0.8497528, -0.8406506, -0.8314381, -0.8221223, -0.8127099, -0.8032075, 
    -0.7936214, -0.7839577, -0.7742223, -0.7644209, -0.7545591, -0.744642, 
    -0.7346748,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0.7346748, 0.744642, 0.7545591, 0.7644209, 0.7742223, 0.7839577, 0.7936214, 
    0.8032075, 0.8127099, 0.8221223, 0.8314381, 0.8406506, 0.8497528, 
    0.8587376, 0.8675976, 0.8763254, 0.8849133, 0.8933536, 0.9016382, 
    0.9097592, 0.9177083, 0.9254774, 0.9330581, 0.9404421, 0.947621, 
    0.9545865, 0.9613302, 0.9678438, 0.9741191, 0.9801481, 0.9859229, 
    0.9914355, 0.9966785, 1.001644, 1.006326, 1.010717, 1.014811, 1.018601, 
    1.022082, 1.025248, 1.028095, 1.030618, 1.032812, 1.034675, 1.036204, 
    1.037395, 1.038247, 1.038759, 1.03893, 1.038759, 1.038247, 1.037395, 
    1.036204, 1.034675, 1.032812, 1.030618, 1.028095, 1.025248, 1.022082, 
    1.018601, 1.014811, 1.010717, 1.006326, 1.001644, 0.9966785, 0.9914355, 
    0.9859229, 0.9801481, 0.9741191, 0.9678438, 0.9613302, 0.9545865, 
    0.947621, 0.9404421, 0.9330581, 0.9254774, 0.9177083, 0.9097592, 
    0.9016382, 0.8933536, 0.8849133, 0.8763254, 0.8675976, 0.8587376, 
    0.8497528, 0.8406506, 0.8314381, 0.8221223, 0.8127099, 0.8032075, 
    0.7936214, 0.7839577, 0.7742223, 0.7644209, 0.7545591, 0.744642, 0.7346748,
  1.46935, 1.489277, 1.509105, 1.528821, 1.548416, 1.56788, 1.587199, 
    1.606363, 1.62536, 1.644176, 1.662799, 1.681216, 1.699411, 1.717372, 
    1.735083, 1.752529, 1.769696, 1.786567, 1.803126, 1.819359, 1.835248, 
    1.850776, 1.865928, 1.880687, 1.895035, 1.908957, 1.922435, 1.935454, 
    1.947996, 1.960045, 1.971586, 1.982603, 1.993082, 2.003006, 2.012363, 
    2.021138, 2.029319, 2.036894, 2.04385, 2.050177, 2.055866, 2.060907, 
    2.065293, 2.069016, 2.07207, 2.074451, 2.076154, 2.077178, 2.077519, 
    2.077178, 2.076154, 2.074451, 2.07207, 2.069016, 2.065293, 2.060907, 
    2.055866, 2.050177, 2.04385, 2.036894, 2.029319, 2.021138, 2.012363, 
    2.003006, 1.993082, 1.982603, 1.971586, 1.960045, 1.947996, 1.935454, 
    1.922435, 1.908957, 1.895035, 1.880687, 1.865928, 1.850776, 1.835248, 
    1.819359, 1.803126, 1.786567, 1.769696, 1.752529, 1.735083, 1.717372, 
    1.699411, 1.681216, 1.662799, 1.644176, 1.62536, 1.606363, 1.587199, 
    1.56788, 1.548416, 1.528821, 1.509105, 1.489277, 1.46935,
  2.204024, 2.233899, 2.263623, 2.29318, 2.322554, 2.35173, 2.38069, 
    2.409416, 2.437891, 2.466094, 2.494007, 2.52161, 2.548881, 2.575799, 
    2.602343, 2.628489, 2.654216, 2.679499, 2.704315, 2.72864, 2.752449, 
    2.775718, 2.798423, 2.820537, 2.842036, 2.862896, 2.883091, 2.902596, 
    2.921387, 2.93944, 2.956731, 2.973237, 2.988935, 3.003803, 3.017821, 
    3.030967, 3.043222, 3.054569, 3.06499, 3.074468, 3.08299, 3.090542, 
    3.097111, 3.102689, 3.107264, 3.11083, 3.113382, 3.114914, 3.115426, 
    3.114914, 3.113382, 3.11083, 3.107264, 3.102689, 3.097111, 3.090542, 
    3.08299, 3.074468, 3.06499, 3.054569, 3.043222, 3.030967, 3.017821, 
    3.003803, 2.988935, 2.973237, 2.956731, 2.93944, 2.921387, 2.902596, 
    2.883091, 2.862896, 2.842036, 2.820537, 2.798423, 2.775718, 2.752449, 
    2.72864, 2.704315, 2.679499, 2.654216, 2.628489, 2.602343, 2.575799, 
    2.548881, 2.52161, 2.494007, 2.466094, 2.437891, 2.409416, 2.38069, 
    2.35173, 2.322554, 2.29318, 2.263623, 2.233899, 2.204024,
  2.938699, 2.978501, 3.0181, 3.057476, 3.096608, 3.135473, 3.17405, 
    3.212315, 3.250242, 3.287808, 3.324986, 3.361748, 3.398068, 3.433917, 
    3.469266, 3.504085, 3.538343, 3.57201, 3.605054, 3.637443, 3.669145, 
    3.700126, 3.730354, 3.759796, 3.788419, 3.816189, 3.843073, 3.869038, 
    3.894052, 3.918083, 3.941099, 3.963069, 3.983964, 4.003754, 4.022411, 
    4.039908, 4.05622, 4.071321, 4.08519, 4.097805, 4.109146, 4.119196, 
    4.127939, 4.135361, 4.14145, 4.146196, 4.149592, 4.151631, 4.152311, 
    4.151631, 4.149592, 4.146196, 4.14145, 4.135361, 4.127939, 4.119196, 
    4.109146, 4.097805, 4.08519, 4.071321, 4.05622, 4.039908, 4.022411, 
    4.003754, 3.983964, 3.963069, 3.941099, 3.918083, 3.894052, 3.869038, 
    3.843073, 3.816189, 3.788419, 3.759796, 3.730354, 3.700126, 3.669145, 
    3.637443, 3.605054, 3.57201, 3.538343, 3.504085, 3.469266, 3.433917, 
    3.398068, 3.361748, 3.324986, 3.287808, 3.250242, 3.212315, 3.17405, 
    3.135473, 3.096608, 3.057476, 3.0181, 2.978501, 2.938699,
  3.673374, 3.723077, 3.772523, 3.82169, 3.870549, 3.919074, 3.967237, 
    4.015007, 4.062356, 4.10925, 4.155657, 4.201545, 4.246879, 4.291623, 
    4.335741, 4.379195, 4.421948, 4.463961, 4.505196, 4.545611, 4.585167, 
    4.623823, 4.661538, 4.69827, 4.733978, 4.768622, 4.802159, 4.834549, 
    4.865752, 4.895727, 4.924435, 4.951838, 4.977899, 5.002581, 5.025849, 
    5.047671, 5.068013, 5.086846, 5.104141, 5.119872, 5.134015, 5.146547, 
    5.15745, 5.166705, 5.174297, 5.180215, 5.184449, 5.186993, 5.187841, 
    5.186993, 5.184449, 5.180215, 5.174297, 5.166705, 5.15745, 5.146547, 
    5.134015, 5.119872, 5.104141, 5.086846, 5.068013, 5.047671, 5.025849, 
    5.002581, 4.977899, 4.951838, 4.924435, 4.895727, 4.865752, 4.834549, 
    4.802159, 4.768622, 4.733978, 4.69827, 4.661538, 4.623823, 4.585167, 
    4.545611, 4.505196, 4.463961, 4.421948, 4.379195, 4.335741, 4.291623, 
    4.246879, 4.201545, 4.155657, 4.10925, 4.062356, 4.015007, 3.967237, 
    3.919074, 3.870549, 3.82169, 3.772523, 3.723077, 3.673374,
  4.408049, 4.467618, 4.526879, 4.5858, 4.64435, 4.702497, 4.760206, 
    4.817443, 4.874171, 4.930352, 4.985948, 5.040917, 5.095221, 5.148814, 
    5.201655, 5.253699, 5.304901, 5.355214, 5.404592, 5.452987, 5.50035, 
    5.546633, 5.591787, 5.635764, 5.678512, 5.719984, 5.760129, 5.7989, 
    5.836247, 5.872125, 5.906484, 5.939281, 5.970469, 6.000007, 6.027852, 
    6.053965, 6.078306, 6.100842, 6.121536, 6.140359, 6.157281, 6.172276, 
    6.18532, 6.196393, 6.205477, 6.212557, 6.217623, 6.220666, 6.221681, 
    6.220666, 6.217623, 6.212557, 6.205477, 6.196393, 6.18532, 6.172276, 
    6.157281, 6.140359, 6.121536, 6.100842, 6.078306, 6.053965, 6.027852, 
    6.000007, 5.970469, 5.939281, 5.906484, 5.872125, 5.836247, 5.7989, 
    5.760129, 5.719984, 5.678512, 5.635764, 5.591787, 5.546633, 5.50035, 
    5.452987, 5.404592, 5.355214, 5.304901, 5.253699, 5.201655, 5.148814, 
    5.095221, 5.040917, 4.985948, 4.930352, 4.874171, 4.817443, 4.760206, 
    4.702497, 4.64435, 4.5858, 4.526879, 4.467618, 4.408049,
  5.142724, 5.21212, 5.281153, 5.349786, 5.417983, 5.485706, 5.552916, 
    5.619571, 5.68563, 5.751048, 5.815781, 5.87978, 5.943, 6.00539, 6.066901, 
    6.12748, 6.187074, 6.245632, 6.303097, 6.359414, 6.414529, 6.468383, 
    6.520922, 6.572086, 6.621819, 6.670065, 6.716765, 6.761864, 6.805305, 
    6.847034, 6.886996, 6.925138, 6.96141, 6.995759, 7.02814, 7.058504, 
    7.086808, 7.113011, 7.137073, 7.158958, 7.178632, 7.196066, 7.211231, 
    7.224104, 7.234665, 7.242897, 7.248786, 7.252323, 7.253503, 7.252323, 
    7.248786, 7.242897, 7.234665, 7.224104, 7.211231, 7.196066, 7.178632, 
    7.158958, 7.137073, 7.113011, 7.086808, 7.058504, 7.02814, 6.995759, 
    6.96141, 6.925138, 6.886996, 6.847034, 6.805305, 6.761864, 6.716765, 
    6.670065, 6.621819, 6.572086, 6.520922, 6.468383, 6.414529, 6.359414, 
    6.303097, 6.245632, 6.187074, 6.12748, 6.066901, 6.00539, 5.943, 5.87978, 
    5.815781, 5.751048, 5.68563, 5.619571, 5.552916, 5.485706, 5.417983, 
    5.349786, 5.281153, 5.21212, 5.142724,
  5.877398, 5.956575, 6.035332, 6.113627, 6.19142, 6.268667, 6.345323, 
    6.421341, 6.496675, 6.571271, 6.645081, 6.718051, 6.790126, 6.86125, 
    6.931367, 7.000417, 7.068341, 7.135077, 7.200565, 7.26474, 7.327541, 
    7.388902, 7.448759, 7.507047, 7.563702, 7.618658, 7.671851, 7.723217, 
    7.772693, 7.820215, 7.865723, 7.909157, 7.950458, 7.989569, 8.026436, 
    8.061007, 8.09323, 8.123061, 8.150454, 8.175366, 8.197762, 8.217607, 
    8.23487, 8.249522, 8.261543, 8.270913, 8.277617, 8.281642, 8.282985, 
    8.281642, 8.277617, 8.270913, 8.261543, 8.249522, 8.23487, 8.217607, 
    8.197762, 8.175366, 8.150454, 8.123061, 8.09323, 8.061007, 8.026436, 
    7.989569, 7.950458, 7.909157, 7.865723, 7.820215, 7.772693, 7.723217, 
    7.671851, 7.618658, 7.563702, 7.507047, 7.448759, 7.388902, 7.327541, 
    7.26474, 7.200565, 7.135077, 7.068341, 7.000417, 6.931367, 6.86125, 
    6.790126, 6.718051, 6.645081, 6.571271, 6.496675, 6.421341, 6.345323, 
    6.268667, 6.19142, 6.113627, 6.035332, 5.956575, 5.877398,
  6.612073, 6.700978, 6.789403, 6.877304, 6.964634, 7.051345, 7.137385, 
    7.222704, 7.307246, 7.390956, 7.473776, 7.555646, 7.636507, 7.716295, 
    7.794946, 7.872395, 7.948575, 8.023417, 8.096853, 8.168813, 8.239225, 
    8.308019, 8.375121, 8.44046, 8.503963, 8.565559, 8.625175, 8.682739, 
    8.738181, 8.791431, 8.842422, 8.891085, 8.937356, 8.981172, 9.02247, 
    9.061195, 9.097291, 9.130703, 9.161384, 9.189286, 9.21437, 9.236594, 
    9.255927, 9.272337, 9.285798, 9.29629, 9.303797, 9.308306, 9.30981, 
    9.308306, 9.303797, 9.29629, 9.285798, 9.272337, 9.255927, 9.236594, 
    9.21437, 9.189286, 9.161384, 9.130703, 9.097291, 9.061195, 9.02247, 
    8.981172, 8.937356, 8.891085, 8.842422, 8.791431, 8.738181, 8.682739, 
    8.625175, 8.565559, 8.503963, 8.44046, 8.375121, 8.308019, 8.239225, 
    8.168813, 8.096853, 8.023417, 7.948575, 7.872395, 7.794946, 7.716295, 
    7.636507, 7.555646, 7.473776, 7.390956, 7.307246, 7.222704, 7.137385, 
    7.051345, 6.964634, 6.877304, 6.789403, 6.700978, 6.612073,
  7.346748, 7.445321, 7.543353, 7.640796, 7.737598, 7.833705, 7.929061, 
    8.023608, 8.117288, 8.210036, 8.30179, 8.392486, 8.482054, 8.570426, 
    8.657532, 8.743299, 8.827652, 8.910519, 8.99182, 9.071482, 9.149424, 
    9.225567, 9.299832, 9.372141, 9.442413, 9.510569, 9.576528, 9.640213, 
    9.701547, 9.760451, 9.816853, 9.870676, 9.92185, 9.970306, 10.01598, 
    10.0588, 10.09871, 10.13566, 10.16958, 10.20043, 10.22816, 10.25273, 
    10.2741, 10.29224, 10.30712, 10.31872, 10.32702, 10.332, 10.33367, 
    10.332, 10.32702, 10.31872, 10.30712, 10.29224, 10.2741, 10.25273, 
    10.22816, 10.20043, 10.16958, 10.13566, 10.09871, 10.0588, 10.01598, 
    9.970306, 9.92185, 9.870676, 9.816853, 9.760451, 9.701547, 9.640213, 
    9.576528, 9.510569, 9.442413, 9.372141, 9.299832, 9.225567, 9.149424, 
    9.071482, 8.99182, 8.910519, 8.827652, 8.743299, 8.657532, 8.570426, 
    8.482054, 8.392486, 8.30179, 8.210036, 8.117288, 8.023608, 7.929061, 
    7.833705, 7.737598, 7.640796, 7.543353, 7.445321, 7.346748,
  8.081423, 8.189597, 8.297169, 8.404083, 8.510284, 8.615713, 8.720308, 
    8.824006, 8.926742, 9.028447, 9.129053, 9.228487, 9.326677, 9.423547, 
    9.519018, 9.613013, 9.705451, 9.79625, 9.885328, 9.972599, 10.05798, 
    10.14138, 10.22272, 10.30191, 10.37886, 10.45349, 10.52571, 10.59543, 
    10.66257, 10.72705, 10.78878, 10.84769, 10.90369, 10.95672, 11.0067, 
    11.05355, 11.09722, 11.13764, 11.17476, 11.2085, 11.23884, 11.26572, 
    11.2891, 11.30894, 11.32522, 11.33791, 11.34698, 11.35243, 11.35425, 
    11.35243, 11.34698, 11.33791, 11.32522, 11.30894, 11.2891, 11.26572, 
    11.23884, 11.2085, 11.17476, 11.13764, 11.09722, 11.05355, 11.0067, 
    10.95672, 10.90369, 10.84769, 10.78878, 10.72705, 10.66257, 10.59543, 
    10.52571, 10.45349, 10.37886, 10.30191, 10.22272, 10.14138, 10.05798, 
    9.972599, 9.885328, 9.79625, 9.705451, 9.613013, 9.519018, 9.423547, 
    9.326677, 9.228487, 9.129053, 9.028447, 8.926742, 8.824006, 8.720308, 
    8.615713, 8.510284, 8.404083, 8.297169, 8.189597, 8.081423,
  8.816097, 8.933801, 9.050837, 9.167146, 9.282667, 9.397336, 9.511086, 
    9.623848, 9.735553, 9.846126, 9.955491, 10.06357, 10.17029, 10.27556, 
    10.3793, 10.48143, 10.58185, 10.68048, 10.77724, 10.87202, 10.96474, 
    11.0553, 11.14361, 11.22959, 11.31312, 11.39412, 11.47251, 11.54817, 
    11.62103, 11.691, 11.75798, 11.82189, 11.88264, 11.94017, 11.99438, 
    12.0452, 12.09256, 12.1364, 12.17664, 12.21324, 12.24614, 12.27528, 
    12.30063, 12.32215, 12.3398, 12.35355, 12.36339, 12.3693, 12.37127, 
    12.3693, 12.36339, 12.35355, 12.3398, 12.32215, 12.30063, 12.27528, 
    12.24614, 12.21324, 12.17664, 12.1364, 12.09256, 12.0452, 11.99438, 
    11.94017, 11.88264, 11.82189, 11.75798, 11.691, 11.62103, 11.54817, 
    11.47251, 11.39412, 11.31312, 11.22959, 11.14361, 11.0553, 10.96474, 
    10.87202, 10.77724, 10.68048, 10.58185, 10.48143, 10.3793, 10.27556, 
    10.17029, 10.06357, 9.955491, 9.846126, 9.735553, 9.623848, 9.511086, 
    9.397336, 9.282667, 9.167146, 9.050837, 8.933801, 8.816097,
  9.550773, 9.677926, 9.804344, 9.929964, 10.05472, 10.17854, 10.30135, 
    10.42309, 10.54366, 10.66301, 10.78103, 10.89766, 11.0128, 11.12637, 
    11.23828, 11.34843, 11.45673, 11.5631, 11.66742, 11.7696, 11.86955, 
    11.96717, 12.06235, 12.155, 12.24501, 12.33229, 12.41673, 12.49824, 
    12.57673, 12.65208, 12.72422, 12.79304, 12.85847, 12.9204, 12.97877, 
    13.03348, 13.08447, 13.13165, 13.17497, 13.21437, 13.24977, 13.28114, 
    13.30842, 13.33158, 13.35057, 13.36537, 13.37596, 13.38232, 13.38444, 
    13.38232, 13.37596, 13.36537, 13.35057, 13.33158, 13.30842, 13.28114, 
    13.24977, 13.21437, 13.17497, 13.13165, 13.08447, 13.03348, 12.97877, 
    12.9204, 12.85847, 12.79304, 12.72422, 12.65208, 12.57673, 12.49824, 
    12.41673, 12.33229, 12.24501, 12.155, 12.06235, 11.96717, 11.86955, 
    11.7696, 11.66742, 11.5631, 11.45673, 11.34843, 11.23828, 11.12637, 
    11.0128, 10.89766, 10.78103, 10.66301, 10.54366, 10.42309, 10.30135, 
    10.17854, 10.05472, 9.929964, 9.804344, 9.677926, 9.550773,
  10.28545, 10.42197, 10.55768, 10.69252, 10.82641, 10.95929, 11.09107, 
    11.22167, 11.35102, 11.47903, 11.60561, 11.73068, 11.85414, 11.97589, 
    12.09585, 12.21391, 12.32998, 12.44396, 12.55573, 12.66521, 12.77227, 
    12.87683, 12.97877, 13.07798, 13.17436, 13.2678, 13.3582, 13.44545, 
    13.52945, 13.61009, 13.68729, 13.76093, 13.83093, 13.89719, 13.95963, 
    14.01815, 14.07269, 14.12316, 14.16949, 14.21162, 14.24948, 14.28303, 
    14.3122, 14.33696, 14.35726, 14.37309, 14.38441, 14.39121, 14.39348, 
    14.39121, 14.38441, 14.37309, 14.35726, 14.33696, 14.3122, 14.28303, 
    14.24948, 14.21162, 14.16949, 14.12316, 14.07269, 14.01815, 13.95963, 
    13.89719, 13.83093, 13.76093, 13.68729, 13.61009, 13.52945, 13.44545, 
    13.3582, 13.2678, 13.17436, 13.07798, 12.97877, 12.87683, 12.77227, 
    12.66521, 12.55573, 12.44396, 12.32998, 12.21391, 12.09585, 11.97589, 
    11.85414, 11.73068, 11.60561, 11.47903, 11.35102, 11.22167, 11.09107, 
    10.95929, 10.82641, 10.69252, 10.55768, 10.42197, 10.28545,
  11.02012, 11.16591, 11.31083, 11.45479, 11.59772, 11.73955, 11.88019, 
    12.01956, 12.15757, 12.29414, 12.42916, 12.56255, 12.6942, 12.82403, 
    12.95192, 13.07777, 13.20149, 13.32295, 13.44206, 13.5587, 13.67276, 
    13.78413, 13.8927, 13.99836, 14.10098, 14.20047, 14.29671, 14.38959, 
    14.479, 14.56483, 14.64697, 14.72534, 14.79981, 14.87031, 14.93673, 
    14.99899, 15.05699, 15.11067, 15.15995, 15.20475, 15.24501, 15.28068, 
    15.3117, 15.33803, 15.35962, 15.37645, 15.38849, 15.39572, 15.39813, 
    15.39572, 15.38849, 15.37645, 15.35962, 15.33803, 15.3117, 15.28068, 
    15.24501, 15.20475, 15.15995, 15.11067, 15.05699, 14.99899, 14.93673, 
    14.87031, 14.79981, 14.72534, 14.64697, 14.56483, 14.479, 14.38959, 
    14.29671, 14.20047, 14.10098, 13.99836, 13.8927, 13.78413, 13.67276, 
    13.5587, 13.44206, 13.32295, 13.20149, 13.07777, 12.95192, 12.82403, 
    12.6942, 12.56255, 12.42916, 12.29414, 12.15757, 12.01956, 11.88019, 
    11.73955, 11.59772, 11.45479, 11.31083, 11.16591, 11.02012,
  11.7548, 11.90976, 12.06378, 12.21676, 12.36863, 12.5193, 12.66869, 
    12.81671, 12.96326, 13.10826, 13.2516, 13.39319, 13.53292, 13.67069, 
    13.80638, 13.9399, 14.07113, 14.19996, 14.32627, 14.44994, 14.57087, 
    14.68893, 14.804, 14.91598, 15.02473, 15.13014, 15.2321, 15.33048, 
    15.42518, 15.51608, 15.60307, 15.68605, 15.7649, 15.83954, 15.90985, 
    15.97575, 16.03714, 16.09396, 16.1461, 16.19351, 16.23612, 16.27386, 
    16.30668, 16.33454, 16.35738, 16.37519, 16.38792, 16.39557, 16.39812, 
    16.39557, 16.38792, 16.37519, 16.35738, 16.33454, 16.30668, 16.27386, 
    16.23612, 16.19351, 16.1461, 16.09396, 16.03714, 15.97575, 15.90985, 
    15.83954, 15.7649, 15.68605, 15.60307, 15.51608, 15.42518, 15.33048, 
    15.2321, 15.13014, 15.02473, 14.91598, 14.804, 14.68893, 14.57087, 
    14.44994, 14.32627, 14.19996, 14.07113, 13.9399, 13.80638, 13.67069, 
    13.53292, 13.39319, 13.2516, 13.10826, 12.96326, 12.81671, 12.66869, 
    12.5193, 12.36863, 12.21676, 12.06378, 11.90976, 11.7548,
  12.48947, 12.65351, 12.81652, 12.97841, 13.1391, 13.2985, 13.45652, 
    13.61306, 13.76804, 13.92135, 14.07288, 14.22254, 14.37021, 14.51579, 
    14.65916, 14.8002, 14.93881, 15.07486, 15.20823, 15.33881, 15.46647, 
    15.59108, 15.71253, 15.83068, 15.94542, 16.05663, 16.16418, 16.26795, 
    16.36782, 16.46367, 16.55539, 16.64287, 16.72599, 16.80466, 16.87877, 
    16.94822, 17.01292, 17.07278, 17.12773, 17.17768, 17.22256, 17.26232, 
    17.2969, 17.32624, 17.3503, 17.36906, 17.38247, 17.39053, 17.39322, 
    17.39053, 17.38247, 17.36906, 17.3503, 17.32624, 17.2969, 17.26232, 
    17.22256, 17.17768, 17.12773, 17.07278, 17.01292, 16.94822, 16.87877, 
    16.80466, 16.72599, 16.64287, 16.55539, 16.46367, 16.36782, 16.26795, 
    16.16418, 16.05663, 15.94542, 15.83068, 15.71253, 15.59108, 15.46647, 
    15.33881, 15.20823, 15.07486, 14.93881, 14.8002, 14.65916, 14.51579, 
    14.37021, 14.22254, 14.07288, 13.92135, 13.76804, 13.61306, 13.45652, 
    13.2985, 13.1391, 12.97841, 12.81652, 12.65351, 12.48947,
  13.22415, 13.39715, 13.56903, 13.73972, 13.90911, 14.07711, 14.24364, 
    14.40859, 14.57185, 14.73334, 14.89293, 15.05052, 15.20599, 15.35924, 
    15.51014, 15.65857, 15.80442, 15.94755, 16.08784, 16.22518, 16.35942, 
    16.49044, 16.61812, 16.74232, 16.86292, 16.97978, 17.09279, 17.20181, 
    17.30672, 17.4074, 17.50373, 17.5956, 17.68288, 17.76548, 17.84328, 
    17.91618, 17.9841, 18.04693, 18.1046, 18.15702, 18.20412, 18.24584, 
    18.28212, 18.31291, 18.33815, 18.35783, 18.3719, 18.38036, 18.38318, 
    18.38036, 18.3719, 18.35783, 18.33815, 18.31291, 18.28212, 18.24584, 
    18.20412, 18.15702, 18.1046, 18.04693, 17.9841, 17.91618, 17.84328, 
    17.76548, 17.68288, 17.5956, 17.50373, 17.4074, 17.30672, 17.20181, 
    17.09279, 16.97978, 16.86292, 16.74232, 16.61812, 16.49044, 16.35942, 
    16.22518, 16.08784, 15.94755, 15.80442, 15.65857, 15.51014, 15.35924, 
    15.20599, 15.05052, 14.89293, 14.73334, 14.57185, 14.40859, 14.24364, 
    14.07711, 13.90911, 13.73972, 13.56903, 13.39715, 13.22415,
  13.95882, 14.14067, 14.32132, 14.50067, 14.67863, 14.85512, 15.03002, 
    15.20323, 15.37465, 15.54417, 15.71168, 15.87706, 16.0402, 16.20097, 
    16.35925, 16.51492, 16.66785, 16.81791, 16.96498, 17.10892, 17.2496, 
    17.38689, 17.52065, 17.65075, 17.77705, 17.89944, 18.01776, 18.1319, 
    18.24172, 18.34711, 18.44792, 18.54405, 18.63538, 18.7218, 18.80319, 
    18.87945, 18.95048, 19.0162, 19.0765, 19.13132, 19.18058, 19.2242, 
    19.26213, 19.29432, 19.32071, 19.34128, 19.356, 19.36483, 19.36778, 
    19.36483, 19.356, 19.34128, 19.32071, 19.29432, 19.26213, 19.2242, 
    19.18058, 19.13132, 19.0765, 19.0162, 18.95048, 18.87945, 18.80319, 
    18.7218, 18.63538, 18.54405, 18.44792, 18.34711, 18.24172, 18.1319, 
    18.01776, 17.89944, 17.77705, 17.65075, 17.52065, 17.38689, 17.2496, 
    17.10892, 16.96498, 16.81791, 16.66785, 16.51492, 16.35925, 16.20097, 
    16.0402, 15.87706, 15.71168, 15.54417, 15.37465, 15.20323, 15.03002, 
    14.85512, 14.67863, 14.50067, 14.32132, 14.14067, 13.95882,
  14.6935, 14.88407, 15.07335, 15.26124, 15.44765, 15.63248, 15.81561, 
    15.99695, 16.17639, 16.3538, 16.52908, 16.7021, 16.87274, 17.04088, 
    17.20639, 17.36914, 17.52901, 17.68585, 17.83953, 17.98992, 18.13688, 
    18.28028, 18.41997, 18.55582, 18.68769, 18.81544, 18.93895, 19.05806, 
    19.17266, 19.28261, 19.38778, 19.48806, 19.58331, 19.67343, 19.7583, 
    19.83782, 19.91188, 19.98038, 20.04325, 20.10039, 20.15172, 20.19719, 
    20.23672, 20.27026, 20.29777, 20.3192, 20.33454, 20.34374, 20.34682, 
    20.34374, 20.33454, 20.3192, 20.29777, 20.27026, 20.23672, 20.19719, 
    20.15172, 20.10039, 20.04325, 19.98038, 19.91188, 19.83782, 19.7583, 
    19.67343, 19.58331, 19.48806, 19.38778, 19.28261, 19.17266, 19.05806, 
    18.93895, 18.81544, 18.68769, 18.55582, 18.41997, 18.28028, 18.13688, 
    17.98992, 17.83953, 17.68585, 17.52901, 17.36914, 17.20639, 17.04088, 
    16.87274, 16.7021, 16.52908, 16.3538, 16.17639, 15.99695, 15.81561, 
    15.63248, 15.44765, 15.26124, 15.07335, 14.88407, 14.6935,
  15.42817, 15.62734, 15.82513, 16.02143, 16.21614, 16.40917, 16.6004, 
    16.78971, 16.97701, 17.16216, 17.34505, 17.52556, 17.70355, 17.8789, 
    18.05148, 18.22116, 18.38779, 18.55125, 18.71139, 18.86807, 19.02115, 
    19.1705, 19.31597, 19.45741, 19.59469, 19.72766, 19.85619, 19.98014, 
    20.09937, 20.21375, 20.32315, 20.42744, 20.5265, 20.6202, 20.70844, 
    20.79111, 20.8681, 20.9393, 21.00464, 21.06402, 21.11737, 21.16462, 
    21.20569, 21.24054, 21.26912, 21.29139, 21.30732, 21.31689, 21.32008, 
    21.31689, 21.30732, 21.29139, 21.26912, 21.24054, 21.20569, 21.16462, 
    21.11737, 21.06402, 21.00464, 20.9393, 20.8681, 20.79111, 20.70844, 
    20.6202, 20.5265, 20.42744, 20.32315, 20.21375, 20.09937, 19.98014, 
    19.85619, 19.72766, 19.59469, 19.45741, 19.31597, 19.1705, 19.02115, 
    18.86807, 18.71139, 18.55125, 18.38779, 18.22116, 18.05148, 17.8789, 
    17.70355, 17.52556, 17.34505, 17.16216, 16.97701, 16.78971, 16.6004, 
    16.40917, 16.21614, 16.02143, 15.82513, 15.62734, 15.42817,
  16.16285, 16.37048, 16.57663, 16.7812, 16.98408, 17.18516, 17.38433, 
    17.58147, 17.77647, 17.96921, 18.15956, 18.34738, 18.53256, 18.71496, 
    18.89445, 19.07088, 19.24412, 19.41402, 19.58045, 19.74325, 19.9023, 
    20.05743, 20.20851, 20.35538, 20.49791, 20.63595, 20.76936, 20.89799, 
    21.02171, 21.14038, 21.25386, 21.36204, 21.46477, 21.56195, 21.65344, 
    21.73915, 21.81896, 21.89278, 21.9605, 22.02205, 22.07734, 22.1263, 
    22.16886, 22.20498, 22.23459, 22.25766, 22.27417, 22.28408, 22.28739, 
    22.28408, 22.27417, 22.25766, 22.23459, 22.20498, 22.16886, 22.1263, 
    22.07734, 22.02205, 21.9605, 21.89278, 21.81896, 21.73915, 21.65344, 
    21.56195, 21.46477, 21.36204, 21.25386, 21.14038, 21.02171, 20.89799, 
    20.76936, 20.63595, 20.49791, 20.35538, 20.20851, 20.05743, 19.9023, 
    19.74325, 19.58045, 19.41402, 19.24412, 19.07088, 18.89445, 18.71496, 
    18.53256, 18.34738, 18.15956, 17.96921, 17.77647, 17.58147, 17.38433, 
    17.18516, 16.98408, 16.7812, 16.57663, 16.37048, 16.16285,
  16.89752, 17.11348, 17.32786, 17.54054, 17.75143, 17.96042, 18.16737, 
    18.37219, 18.57473, 18.77489, 18.97252, 19.16751, 19.35971, 19.54898, 
    19.7352, 19.91821, 20.09789, 20.27407, 20.44661, 20.61537, 20.7802, 
    20.94095, 21.09747, 21.24961, 21.39723, 21.54018, 21.6783, 21.81147, 
    21.93953, 22.06234, 22.17978, 22.2917, 22.39799, 22.49851, 22.59314, 
    22.68178, 22.76431, 22.84064, 22.91066, 22.97429, 23.03145, 23.08206, 
    23.12605, 23.16338, 23.19399, 23.21784, 23.2349, 23.24514, 23.24856, 
    23.24514, 23.2349, 23.21784, 23.19399, 23.16338, 23.12605, 23.08206, 
    23.03145, 22.97429, 22.91066, 22.84064, 22.76431, 22.68178, 22.59314, 
    22.49851, 22.39799, 22.2917, 22.17978, 22.06234, 21.93953, 21.81147, 
    21.6783, 21.54018, 21.39723, 21.24961, 21.09747, 20.94095, 20.7802, 
    20.61537, 20.44661, 20.27407, 20.09789, 19.91821, 19.7352, 19.54898, 
    19.35971, 19.16751, 18.97252, 18.77489, 18.57473, 18.37219, 18.16737, 
    17.96042, 17.75143, 17.54054, 17.32786, 17.11348, 16.89752,
  17.63219, 17.85633, 18.07879, 18.29944, 18.51819, 18.73492, 18.9495, 
    19.16182, 19.37174, 19.57915, 19.7839, 19.98587, 20.18491, 20.38089, 
    20.57367, 20.76309, 20.94901, 21.13129, 21.30978, 21.48432, 21.65476, 
    21.82095, 21.98275, 22.13999, 22.29253, 22.44022, 22.5829, 22.72045, 
    22.85269, 22.97951, 23.10075, 23.21629, 23.32599, 23.42973, 23.52739, 
    23.61885, 23.704, 23.78273, 23.85496, 23.92059, 23.97954, 24.03174, 
    24.07711, 24.1156, 24.14717, 24.17175, 24.18934, 24.19991, 24.20343, 
    24.19991, 24.18934, 24.17175, 24.14717, 24.1156, 24.07711, 24.03174, 
    23.97954, 23.92059, 23.85496, 23.78273, 23.704, 23.61885, 23.52739, 
    23.42973, 23.32599, 23.21629, 23.10075, 22.97951, 22.85269, 22.72045, 
    22.5829, 22.44022, 22.29253, 22.13999, 21.98275, 21.82095, 21.65476, 
    21.48432, 21.30978, 21.13129, 20.94901, 20.76309, 20.57367, 20.38089, 
    20.18491, 19.98587, 19.7839, 19.57915, 19.37174, 19.16182, 18.9495, 
    18.73492, 18.51819, 18.29944, 18.07879, 17.85633, 17.63219,
  18.36687, 18.59904, 18.82941, 19.05788, 19.28433, 19.50863, 19.73068, 
    19.95033, 20.16746, 20.38194, 20.59364, 20.80241, 21.00812, 21.21062, 
    21.40977, 21.60542, 21.79742, 21.98561, 22.16986, 22.35, 22.52588, 
    22.69734, 22.86423, 23.0264, 23.18369, 23.33596, 23.48304, 23.6248, 
    23.76108, 23.89175, 24.01665, 24.13567, 24.24865, 24.35549, 24.45604, 
    24.55021, 24.63787, 24.71892, 24.79326, 24.86081, 24.92148, 24.97519, 
    25.02188, 25.06149, 25.09396, 25.11926, 25.13736, 25.14822, 25.15185, 
    25.14822, 25.13736, 25.11926, 25.09396, 25.06149, 25.02188, 24.97519, 
    24.92148, 24.86081, 24.79326, 24.71892, 24.63787, 24.55021, 24.45604, 
    24.35549, 24.24865, 24.13567, 24.01665, 23.89175, 23.76108, 23.6248, 
    23.48304, 23.33596, 23.18369, 23.0264, 22.86423, 22.69734, 22.52588, 
    22.35, 22.16986, 21.98561, 21.79742, 21.60542, 21.40977, 21.21062, 
    21.00812, 20.80241, 20.59364, 20.38194, 20.16746, 19.95033, 19.73068, 
    19.50863, 19.28433, 19.05788, 18.82941, 18.59904, 18.36687,
  19.10155, 19.34159, 19.57973, 19.81585, 20.04982, 20.28154, 20.51087, 
    20.73768, 20.96184, 21.18322, 21.40168, 21.61708, 21.82927, 22.03811, 
    22.24345, 22.44514, 22.64302, 22.83695, 23.02677, 23.21232, 23.39345, 
    23.57, 23.74181, 23.90874, 24.07061, 24.22728, 24.3786, 24.52441, 
    24.66457, 24.79893, 24.92736, 25.0497, 25.16584, 25.27564, 25.37897, 
    25.47573, 25.56579, 25.64905, 25.72542, 25.7948, 25.85711, 25.91227, 
    25.96022, 26.00089, 26.03424, 26.06021, 26.0788, 26.08995, 26.09367, 
    26.08995, 26.0788, 26.06021, 26.03424, 26.00089, 25.96022, 25.91227, 
    25.85711, 25.7948, 25.72542, 25.64905, 25.56579, 25.47573, 25.37897, 
    25.27564, 25.16584, 25.0497, 24.92736, 24.79893, 24.66457, 24.52441, 
    24.3786, 24.22728, 24.07061, 23.90874, 23.74181, 23.57, 23.39345, 
    23.21232, 23.02677, 22.83695, 22.64302, 22.44514, 22.24345, 22.03811, 
    21.82927, 21.61708, 21.40168, 21.18322, 20.96184, 20.73768, 20.51087, 
    20.28154, 20.04982, 19.81585, 19.57973, 19.34159, 19.10155,
  19.83622, 20.08398, 20.32972, 20.57332, 20.81466, 21.05361, 21.29005, 
    21.52384, 21.75485, 21.98295, 22.20798, 22.42981, 22.6483, 22.86328, 
    23.07462, 23.28216, 23.48574, 23.68522, 23.88042, 24.0712, 24.2574, 
    24.43885, 24.6154, 24.7869, 24.95318, 25.11408, 25.26947, 25.41917, 
    25.56305, 25.70096, 25.83275, 25.95829, 26.07744, 26.19007, 26.29606, 
    26.39529, 26.48764, 26.57302, 26.65132, 26.72244, 26.78632, 26.84286, 
    26.892, 26.93369, 26.96786, 26.99449, 27.01353, 27.02497, 27.02878, 
    27.02497, 27.01353, 26.99449, 26.96786, 26.93369, 26.892, 26.84286, 
    26.78632, 26.72244, 26.65132, 26.57302, 26.48764, 26.39529, 26.29606, 
    26.19007, 26.07744, 25.95829, 25.83275, 25.70096, 25.56305, 25.41917, 
    25.26947, 25.11408, 24.95318, 24.7869, 24.6154, 24.43885, 24.2574, 
    24.0712, 23.88042, 23.68522, 23.48574, 23.28216, 23.07462, 22.86328, 
    22.6483, 22.42981, 22.20798, 21.98295, 21.75485, 21.52384, 21.29005, 
    21.05361, 20.81466, 20.57332, 20.32972, 20.08398, 19.83622,
  20.57089, 20.8262, 21.07937, 21.33028, 21.5788, 21.82482, 22.06818, 
    22.30877, 22.54645, 22.78106, 23.01249, 23.24056, 23.46515, 23.68609, 
    23.90323, 24.11643, 24.32551, 24.53034, 24.73074, 24.92656, 25.11763, 
    25.3038, 25.48491, 25.6608, 25.8313, 25.99627, 26.15555, 26.30898, 
    26.45642, 26.59771, 26.73272, 26.86131, 26.98333, 27.09867, 27.20719, 
    27.30877, 27.40331, 27.4907, 27.57083, 27.64362, 27.70898, 27.76684, 
    27.81712, 27.85977, 27.89473, 27.92197, 27.94145, 27.95315, 27.95705, 
    27.95315, 27.94145, 27.92197, 27.89473, 27.85977, 27.81712, 27.76684, 
    27.70898, 27.64362, 27.57083, 27.4907, 27.40331, 27.30877, 27.20719, 
    27.09867, 26.98333, 26.86131, 26.73272, 26.59771, 26.45642, 26.30898, 
    26.15555, 25.99627, 25.8313, 25.6608, 25.48491, 25.3038, 25.11763, 
    24.92656, 24.73074, 24.53034, 24.32551, 24.11643, 23.90323, 23.68609, 
    23.46515, 23.24056, 23.01249, 22.78106, 22.54645, 22.30877, 22.06818, 
    21.82482, 21.5788, 21.33028, 21.07937, 20.8262, 20.57089,
  21.30557, 21.56826, 21.82868, 22.08672, 22.34225, 22.59513, 22.84524, 
    23.09244, 23.33659, 23.57754, 23.81515, 24.04927, 24.27976, 24.50646, 
    24.72922, 24.94787, 25.16227, 25.37224, 25.57764, 25.77831, 25.97407, 
    26.16477, 26.35024, 26.53034, 26.70489, 26.87375, 27.03675, 27.19374, 
    27.34457, 27.4891, 27.62718, 27.75867, 27.88343, 28.00133, 28.11226, 
    28.21608, 28.3127, 28.40199, 28.48387, 28.55823, 28.625, 28.6841, 
    28.73546, 28.77902, 28.81473, 28.84255, 28.86244, 28.87439, 28.87837, 
    28.87439, 28.86244, 28.84255, 28.81473, 28.77902, 28.73546, 28.6841, 
    28.625, 28.55823, 28.48387, 28.40199, 28.3127, 28.21608, 28.11226, 
    28.00133, 27.88343, 27.75867, 27.62718, 27.4891, 27.34457, 27.19374, 
    27.03675, 26.87375, 26.70489, 26.53034, 26.35024, 26.16477, 25.97407, 
    25.77831, 25.57764, 25.37224, 25.16227, 24.94787, 24.72922, 24.50646, 
    24.27976, 24.04927, 23.81515, 23.57754, 23.33659, 23.09244, 22.84524, 
    22.59513, 22.34225, 22.08672, 21.82868, 21.56826, 21.30557,
  22.04024, 22.31014, 22.57764, 22.84263, 23.10497, 23.36455, 23.6212, 
    23.87482, 24.12524, 24.37232, 24.61593, 24.85591, 25.0921, 25.32435, 
    25.55252, 25.77643, 25.99593, 26.21087, 26.42107, 26.62638, 26.82663, 
    27.02167, 27.21133, 27.39545, 27.57387, 27.74643, 27.91298, 28.07337, 
    28.22743, 28.37503, 28.51603, 28.65027, 28.77763, 28.89797, 29.01118, 
    29.11712, 29.2157, 29.3068, 29.39032, 29.46618, 29.53428, 29.59455, 
    29.64693, 29.69135, 29.72776, 29.75613, 29.77641, 29.78859, 29.79265, 
    29.78859, 29.77641, 29.75613, 29.72776, 29.69135, 29.64693, 29.59455, 
    29.53428, 29.46618, 29.39032, 29.3068, 29.2157, 29.11712, 29.01118, 
    28.89797, 28.77763, 28.65027, 28.51603, 28.37503, 28.22743, 28.07337, 
    27.91298, 27.74643, 27.57387, 27.39545, 27.21133, 27.02167, 26.82663, 
    26.62638, 26.42107, 26.21087, 25.99593, 25.77643, 25.55252, 25.32435, 
    25.0921, 24.85591, 24.61593, 24.37232, 24.12524, 23.87482, 23.6212, 
    23.36455, 23.10497, 22.84263, 22.57764, 22.31014, 22.04024,
  22.77492, 23.05183, 23.32623, 23.59798, 23.86696, 24.13302, 24.39604, 
    24.65587, 24.91236, 25.16539, 25.41478, 25.6604, 25.9021, 26.13971, 
    26.37307, 26.60204, 26.82645, 27.04614, 27.26094, 27.47071, 27.67526, 
    27.87444, 28.06809, 28.25605, 28.43815, 28.61425, 28.78417, 28.94778, 
    29.10491, 29.25543, 29.39919, 29.53604, 29.66586, 29.78851, 29.90387, 
    30.01182, 30.11224, 30.20505, 30.29012, 30.36738, 30.43673, 30.49811, 
    30.55145, 30.59668, 30.63375, 30.66263, 30.68328, 30.69568, 30.69982, 
    30.69568, 30.68328, 30.66263, 30.63375, 30.59668, 30.55145, 30.49811, 
    30.43673, 30.36738, 30.29012, 30.20505, 30.11224, 30.01182, 29.90387, 
    29.78851, 29.66586, 29.53604, 29.39919, 29.25543, 29.10491, 28.94778, 
    28.78417, 28.61425, 28.43815, 28.25605, 28.06809, 27.87444, 27.67526, 
    27.47071, 27.26094, 27.04614, 26.82645, 26.60204, 26.37307, 26.13971, 
    25.9021, 25.6604, 25.41478, 25.16539, 24.91236, 24.65587, 24.39604, 
    24.13302, 23.86696, 23.59798, 23.32623, 23.05183, 22.77492,
  23.50959, 23.79335, 24.07445, 24.35277, 24.62818, 24.90054, 25.16972, 
    25.43556, 25.69794, 25.95669, 26.21167, 26.46273, 26.70972, 26.95247, 
    27.19084, 27.42466, 27.65377, 27.87801, 28.09721, 28.31122, 28.51988, 
    28.72301, 28.92046, 29.11207, 29.29767, 29.47712, 29.65025, 29.8169, 
    29.97694, 30.13022, 30.27658, 30.4159, 30.54803, 30.67286, 30.79025, 
    30.90008, 31.00225, 31.09665, 31.18319, 31.26176, 31.33229, 31.39471, 
    31.44894, 31.49493, 31.53263, 31.56199, 31.58298, 31.59559, 31.59979, 
    31.59559, 31.58298, 31.56199, 31.53263, 31.49493, 31.44894, 31.39471, 
    31.33229, 31.26176, 31.18319, 31.09665, 31.00225, 30.90008, 30.79025, 
    30.67286, 30.54803, 30.4159, 30.27658, 30.13022, 29.97694, 29.8169, 
    29.65025, 29.47712, 29.29767, 29.11207, 28.92046, 28.72301, 28.51988, 
    28.31122, 28.09721, 27.87801, 27.65377, 27.42466, 27.19084, 26.95247, 
    26.70972, 26.46273, 26.21167, 25.95669, 25.69794, 25.43556, 25.16972, 
    24.90054, 24.62818, 24.35277, 24.07445, 23.79335, 23.50959,
  24.24427, 24.53467, 24.82229, 25.10699, 25.38863, 25.66709, 25.94222, 
    26.21387, 26.48191, 26.74619, 27.00655, 27.26284, 27.51491, 27.76261, 
    28.00576, 28.24422, 28.47782, 28.70641, 28.92981, 29.14787, 29.36043, 
    29.56732, 29.76838, 29.96344, 30.15236, 30.33498, 30.51114, 30.68068, 
    30.84346, 30.99933, 31.14815, 31.28979, 31.4241, 31.55096, 31.67025, 
    31.78186, 31.88566, 31.98156, 32.06945, 32.14926, 32.22089, 32.28428, 
    32.33934, 32.38604, 32.42432, 32.45413, 32.47544, 32.48825, 32.49251, 
    32.48825, 32.47544, 32.45413, 32.42432, 32.38604, 32.33934, 32.28428, 
    32.22089, 32.14926, 32.06945, 31.98156, 31.88566, 31.78186, 31.67025, 
    31.55096, 31.4241, 31.28979, 31.14815, 30.99933, 30.84346, 30.68068, 
    30.51114, 30.33498, 30.15236, 29.96344, 29.76838, 29.56732, 29.36043, 
    29.14787, 28.92981, 28.70641, 28.47782, 28.24422, 28.00576, 27.76261, 
    27.51491, 27.26284, 27.00655, 26.74619, 26.48191, 26.21387, 25.94222, 
    25.66709, 25.38863, 25.10699, 24.82229, 24.53467, 24.24427,
  24.97894, 25.2758, 25.56974, 25.86061, 26.14829, 26.43264, 26.71351, 
    26.99077, 27.26427, 27.53386, 27.79938, 28.0607, 28.31764, 28.57006, 
    28.81779, 29.06068, 29.29857, 29.5313, 29.75869, 29.9806, 30.19686, 
    30.4073, 30.61178, 30.81012, 31.00217, 31.18778, 31.36679, 31.53904, 
    31.7044, 31.86271, 32.01384, 32.15764, 32.29399, 32.42276, 32.54383, 
    32.65709, 32.76241, 32.85971, 32.94887, 33.02983, 33.10248, 33.16676, 
    33.22261, 33.26997, 33.30878, 33.33901, 33.36062, 33.3736, 33.37793, 
    33.3736, 33.36062, 33.33901, 33.30878, 33.26997, 33.22261, 33.16676, 
    33.10248, 33.02983, 32.94887, 32.85971, 32.76241, 32.65709, 32.54383, 
    32.42276, 32.29399, 32.15764, 32.01384, 31.86271, 31.7044, 31.53904, 
    31.36679, 31.18778, 31.00217, 30.81012, 30.61178, 30.4073, 30.19686, 
    29.9806, 29.75869, 29.5313, 29.29857, 29.06068, 28.81779, 28.57006, 
    28.31764, 28.0607, 27.79938, 27.53386, 27.26427, 26.99077, 26.71351, 
    26.43264, 26.14829, 25.86061, 25.56974, 25.2758, 24.97894,
  25.71362, 26.01674, 26.31679, 26.61363, 26.90714, 27.19717, 27.48358, 
    27.76624, 28.04498, 28.31966, 28.59014, 28.85626, 29.11786, 29.37479, 
    29.62689, 29.874, 30.11596, 30.35262, 30.5838, 30.80936, 31.02912, 
    31.24292, 31.45062, 31.65205, 31.84704, 32.03546, 32.21714, 32.39194, 
    32.55971, 32.7203, 32.87358, 33.01942, 33.15767, 33.28822, 33.41094, 
    33.52573, 33.63246, 33.73105, 33.8214, 33.90341, 33.97701, 34.04213, 
    34.0987, 34.14666, 34.18597, 34.21658, 34.23848, 34.25162, 34.256, 
    34.25162, 34.23848, 34.21658, 34.18597, 34.14666, 34.0987, 34.04213, 
    33.97701, 33.90341, 33.8214, 33.73105, 33.63246, 33.52573, 33.41094, 
    33.28822, 33.15767, 33.01942, 32.87358, 32.7203, 32.55971, 32.39194, 
    32.21714, 32.03546, 31.84704, 31.65205, 31.45062, 31.24292, 31.02912, 
    30.80936, 30.5838, 30.35262, 30.11596, 29.874, 29.62689, 29.37479, 
    29.11786, 28.85626, 28.59014, 28.31966, 28.04498, 27.76624, 27.48358, 
    27.19717, 26.90714, 26.61363, 26.31679, 26.01674, 25.71362,
  26.44829, 26.75747, 27.06343, 27.36604, 27.66517, 27.96067, 28.25241, 
    28.54023, 28.82401, 29.10357, 29.37879, 29.64949, 29.91554, 30.17676, 
    30.43301, 30.68413, 30.92996, 31.17034, 31.4051, 31.63409, 31.85715, 
    32.07413, 32.28485, 32.48917, 32.68693, 32.87798, 33.06216, 33.23934, 
    33.40936, 33.57207, 33.72735, 33.87507, 34.01508, 34.14728, 34.27153, 
    34.38773, 34.49578, 34.59556, 34.68699, 34.76999, 34.84446, 34.91034, 
    34.96757, 35.01609, 35.05586, 35.08683, 35.10897, 35.12226, 35.12669, 
    35.12226, 35.10897, 35.08683, 35.05586, 35.01609, 34.96757, 34.91034, 
    34.84446, 34.76999, 34.68699, 34.59556, 34.49578, 34.38773, 34.27153, 
    34.14728, 34.01508, 33.87507, 33.72735, 33.57207, 33.40936, 33.23934, 
    33.06216, 32.87798, 32.68693, 32.48917, 32.28485, 32.07413, 31.85715, 
    31.63409, 31.4051, 31.17034, 30.92996, 30.68413, 30.43301, 30.17676, 
    29.91554, 29.64949, 29.37879, 29.10357, 28.82401, 28.54023, 28.25241, 
    27.96067, 27.66517, 27.36604, 27.06343, 26.75747, 26.44829,
  27.18297, 27.49799, 27.80966, 28.11782, 28.42235, 28.72311, 29.01996, 
    29.31275, 29.60133, 29.88556, 30.16529, 30.44036, 30.71063, 30.97594, 
    31.23613, 31.49104, 31.74052, 31.98441, 32.22254, 32.45477, 32.68093, 
    32.90088, 33.11443, 33.32146, 33.5218, 33.7153, 33.90181, 34.08119, 
    34.25329, 34.41798, 34.57511, 34.72456, 34.8662, 34.99992, 35.12558, 
    35.24308, 35.35233, 35.45321, 35.54563, 35.62952, 35.70479, 35.77137, 
    35.8292, 35.87823, 35.91842, 35.94971, 35.97208, 35.98551, 35.98999, 
    35.98551, 35.97208, 35.94971, 35.91842, 35.87823, 35.8292, 35.77137, 
    35.70479, 35.62952, 35.54563, 35.45321, 35.35233, 35.24308, 35.12558, 
    34.99992, 34.8662, 34.72456, 34.57511, 34.41798, 34.25329, 34.08119, 
    33.90181, 33.7153, 33.5218, 33.32146, 33.11443, 32.90088, 32.68093, 
    32.45477, 32.22254, 31.98441, 31.74052, 31.49104, 31.23613, 30.97594, 
    30.71063, 30.44036, 30.16529, 29.88556, 29.60133, 29.31275, 29.01996, 
    28.72311, 28.42235, 28.11782, 27.80966, 27.49799, 27.18297,
  27.91764, 28.23831, 28.55546, 28.86897, 29.17869, 29.48449, 29.78622, 
    30.08375, 30.37692, 30.6656, 30.94962, 31.22885, 31.50312, 31.77229, 
    32.03619, 32.29469, 32.5476, 32.79479, 33.03609, 33.27135, 33.50042, 
    33.72313, 33.93933, 34.14888, 34.35161, 34.54738, 34.73605, 34.91746, 
    35.09149, 35.25799, 35.41682, 35.56787, 35.71101, 35.8461, 35.97306, 
    36.09175, 36.20208, 36.30396, 36.39729, 36.48199, 36.55799, 36.62521, 
    36.68359, 36.73308, 36.77364, 36.80522, 36.8278, 36.84136, 36.84588, 
    36.84136, 36.8278, 36.80522, 36.77364, 36.73308, 36.68359, 36.62521, 
    36.55799, 36.48199, 36.39729, 36.30396, 36.20208, 36.09175, 35.97306, 
    35.8461, 35.71101, 35.56787, 35.41682, 35.25799, 35.09149, 34.91746, 
    34.73605, 34.54738, 34.35161, 34.14888, 33.93933, 33.72313, 33.50042, 
    33.27135, 33.03609, 32.79479, 32.5476, 32.29469, 32.03619, 31.77229, 
    31.50312, 31.22885, 30.94962, 30.6656, 30.37692, 30.08375, 29.78622, 
    29.48449, 29.17869, 28.86897, 28.55546, 28.23831, 27.91764,
  28.65232, 28.97841, 29.30084, 29.61947, 29.93416, 30.24478, 30.55118, 
    30.85322, 31.15076, 31.44366, 31.73176, 32.01491, 32.29297, 32.56578, 
    32.83318, 33.09504, 33.35118, 33.60146, 33.84572, 34.08381, 34.31557, 
    34.54086, 34.75951, 34.97139, 35.17633, 35.3742, 35.56485, 35.74813, 
    35.92393, 36.09208, 36.25248, 36.40498, 36.54947, 36.68583, 36.81395, 
    36.93372, 37.04504, 37.14782, 37.24197, 37.3274, 37.40405, 37.47184, 
    37.53071, 37.58062, 37.62151, 37.65335, 37.67612, 37.68979, 37.69435, 
    37.68979, 37.67612, 37.65335, 37.62151, 37.58062, 37.53071, 37.47184, 
    37.40405, 37.3274, 37.24197, 37.14782, 37.04504, 36.93372, 36.81395, 
    36.68583, 36.54947, 36.40498, 36.25248, 36.09208, 35.92393, 35.74813, 
    35.56485, 35.3742, 35.17633, 34.97139, 34.75951, 34.54086, 34.31557, 
    34.08381, 33.84572, 33.60146, 33.35118, 33.09504, 32.83318, 32.56578, 
    32.29297, 32.01491, 31.73176, 31.44366, 31.15076, 30.85322, 30.55118, 
    30.24478, 29.93416, 29.61947, 29.30084, 28.97841, 28.65232,
  29.38699, 29.7183, 30.04578, 30.36931, 30.68875, 31.00396, 31.31481, 
    31.62114, 31.92283, 32.21972, 32.51167, 32.79853, 33.08015, 33.35638, 
    33.62707, 33.89207, 34.15122, 34.40438, 34.6514, 34.89211, 35.12637, 
    35.35404, 35.57495, 35.78897, 35.99594, 36.19573, 36.38819, 36.57319, 
    36.75058, 36.92025, 37.08205, 37.23587, 37.38158, 37.51908, 37.64825, 
    37.76899, 37.8812, 37.98478, 38.07965, 38.16574, 38.24297, 38.31126, 
    38.37057, 38.42085, 38.46204, 38.49412, 38.51705, 38.53082, 38.53541, 
    38.53082, 38.51705, 38.49412, 38.46204, 38.42085, 38.37057, 38.31126, 
    38.24297, 38.16574, 38.07965, 37.98478, 37.8812, 37.76899, 37.64825, 
    37.51908, 37.38158, 37.23587, 37.08205, 36.92025, 36.75058, 36.57319, 
    36.38819, 36.19573, 35.99594, 35.78897, 35.57495, 35.35404, 35.12637, 
    34.89211, 34.6514, 34.40438, 34.15122, 33.89207, 33.62707, 33.35638, 
    33.08015, 32.79853, 32.51167, 32.21972, 31.92283, 31.62114, 31.31481, 
    31.00396, 30.68875, 30.36931, 30.04578, 29.7183, 29.38699,
  30.12167, 30.45796, 30.79028, 31.11849, 31.44245, 31.76203, 32.0771, 
    32.3875, 32.6931, 32.99376, 33.28933, 33.57967, 33.86464, 34.14407, 
    34.41782, 34.68575, 34.94771, 35.20354, 35.45309, 35.69623, 35.9328, 
    36.16264, 36.38563, 36.6016, 36.81043, 37.01196, 37.20607, 37.39261, 
    37.57145, 37.74247, 37.90554, 38.06054, 38.20735, 38.34586, 38.47596, 
    38.59755, 38.71054, 38.81484, 38.91036, 38.99702, 39.07475, 39.1435, 
    39.20319, 39.25378, 39.29524, 39.32752, 39.3506, 39.36445, 39.36907, 
    39.36445, 39.3506, 39.32752, 39.29524, 39.25378, 39.20319, 39.1435, 
    39.07475, 38.99702, 38.91036, 38.81484, 38.71054, 38.59755, 38.47596, 
    38.34586, 38.20735, 38.06054, 37.90554, 37.74247, 37.57145, 37.39261, 
    37.20607, 37.01196, 36.81043, 36.6016, 36.38563, 36.16264, 35.9328, 
    35.69623, 35.45309, 35.20354, 34.94771, 34.68575, 34.41782, 34.14407, 
    33.86464, 33.57967, 33.28933, 32.99376, 32.6931, 32.3875, 32.0771, 
    31.76203, 31.44245, 31.11849, 30.79028, 30.45796, 30.12167,
  30.85634, 31.19741, 31.53433, 31.86699, 32.19525, 32.51897, 32.83802, 
    33.15226, 33.46156, 33.76576, 34.06473, 34.35833, 34.64641, 34.92882, 
    35.20542, 35.47607, 35.74061, 35.9989, 36.2508, 36.49615, 36.73482, 
    36.96666, 37.19153, 37.40928, 37.61977, 37.82288, 38.01846, 38.20639, 
    38.38652, 38.55875, 38.72294, 38.87898, 39.02676, 39.16616, 39.29708, 
    39.41943, 39.5331, 39.63801, 39.73409, 39.82125, 39.89942, 39.96855, 
    40.02857, 40.07944, 40.12112, 40.15358, 40.17678, 40.1907, 40.19535, 
    40.1907, 40.17678, 40.15358, 40.12112, 40.07944, 40.02857, 39.96855, 
    39.89942, 39.82125, 39.73409, 39.63801, 39.5331, 39.41943, 39.29708, 
    39.16616, 39.02676, 38.87898, 38.72294, 38.55875, 38.38652, 38.20639, 
    38.01846, 37.82288, 37.61977, 37.40928, 37.19153, 36.96666, 36.73482, 
    36.49615, 36.2508, 35.9989, 35.74061, 35.47607, 35.20542, 34.92882, 
    34.64641, 34.35833, 34.06473, 33.76576, 33.46156, 33.15226, 32.83802, 
    32.51897, 32.19525, 31.86699, 31.53433, 31.19741, 30.85634,
  31.59101, 31.93662, 32.27793, 32.61481, 32.94714, 33.27477, 33.59758, 
    33.91543, 34.22818, 34.5357, 34.83784, 35.13448, 35.42545, 35.71062, 
    35.98985, 36.26299, 36.52991, 36.79046, 37.04449, 37.29186, 37.53244, 
    37.76608, 37.99264, 38.21198, 38.42397, 38.62848, 38.82537, 39.01452, 
    39.1958, 39.36908, 39.53426, 39.69121, 39.83982, 39.97999, 40.11162, 
    40.23461, 40.34887, 40.45432, 40.55087, 40.63845, 40.717, 40.78645, 
    40.84675, 40.89785, 40.93972, 40.97232, 40.99562, 41.00961, 41.01428, 
    41.00961, 40.99562, 40.97232, 40.93972, 40.89785, 40.84675, 40.78645, 
    40.717, 40.63845, 40.55087, 40.45432, 40.34887, 40.23461, 40.11162, 
    39.97999, 39.83982, 39.69121, 39.53426, 39.36908, 39.1958, 39.01452, 
    38.82537, 38.62848, 38.42397, 38.21198, 37.99264, 37.76608, 37.53244, 
    37.29186, 37.04449, 36.79046, 36.52991, 36.26299, 35.98985, 35.71062, 
    35.42545, 35.13448, 34.83784, 34.5357, 34.22818, 33.91543, 33.59758, 
    33.27477, 32.94714, 32.61481, 32.27793, 31.93662, 31.59101,
  32.32569, 32.67561, 33.02107, 33.36194, 33.6981, 34.02942, 34.35575, 
    34.67698, 34.99296, 35.30357, 35.60866, 35.90809, 36.20173, 36.48944, 
    36.77109, 37.04652, 37.3156, 37.57819, 37.83415, 38.08334, 38.32563, 
    38.56088, 38.78895, 39.00971, 39.22302, 39.42876, 39.6268, 39.81702, 
    39.99928, 40.17348, 40.3395, 40.49723, 40.64656, 40.78738, 40.91961, 
    41.04314, 41.15789, 41.26377, 41.36071, 41.44865, 41.5275, 41.59722, 
    41.65775, 41.70904, 41.75106, 41.78378, 41.80717, 41.82121, 41.82589, 
    41.82121, 41.80717, 41.78378, 41.75106, 41.70904, 41.65775, 41.59722, 
    41.5275, 41.44865, 41.36071, 41.26377, 41.15789, 41.04314, 40.91961, 
    40.78738, 40.64656, 40.49723, 40.3395, 40.17348, 39.99928, 39.81702, 
    39.6268, 39.42876, 39.22302, 39.00971, 38.78895, 38.56088, 38.32563, 
    38.08334, 37.83415, 37.57819, 37.3156, 37.04652, 36.77109, 36.48944, 
    36.20173, 35.90809, 35.60866, 35.30357, 34.99296, 34.67698, 34.35575, 
    34.02942, 33.6981, 33.36194, 33.02107, 32.67561, 32.32569,
  33.06036, 33.41436, 33.76374, 34.10837, 34.44813, 34.78289, 35.11252, 
    35.4369, 35.75588, 36.06934, 36.37715, 36.67916, 36.97525, 37.26529, 
    37.54912, 37.82662, 38.09766, 38.36209, 38.61978, 38.87059, 39.1144, 
    39.35107, 39.58046, 39.80246, 40.01692, 40.22372, 40.42275, 40.61388, 
    40.79699, 40.97196, 41.13869, 41.29707, 41.44698, 41.58834, 41.72106, 
    41.84503, 41.96017, 42.06641, 42.16367, 42.25187, 42.33097, 42.40089, 
    42.4616, 42.51304, 42.55518, 42.58799, 42.61144, 42.62552, 42.63021, 
    42.62552, 42.61144, 42.58799, 42.55518, 42.51304, 42.4616, 42.40089, 
    42.33097, 42.25187, 42.16367, 42.06641, 41.96017, 41.84503, 41.72106, 
    41.58834, 41.44698, 41.29707, 41.13869, 40.97196, 40.79699, 40.61388, 
    40.42275, 40.22372, 40.01692, 39.80246, 39.58046, 39.35107, 39.1144, 
    38.87059, 38.61978, 38.36209, 38.09766, 37.82662, 37.54912, 37.26529, 
    36.97525, 36.67916, 36.37715, 36.06934, 35.75588, 35.4369, 35.11252, 
    34.78289, 34.44813, 34.10837, 33.76374, 33.41436, 33.06036,
  33.79504, 34.15289, 34.50594, 34.8541, 35.19722, 35.53519, 35.86789, 
    36.19517, 36.51693, 36.83301, 37.14331, 37.44768, 37.746, 38.03813, 
    38.32394, 38.6033, 38.87608, 39.14214, 39.40136, 39.6536, 39.89874, 
    40.13664, 40.36718, 40.59023, 40.80568, 41.01338, 41.21324, 41.40512, 
    41.58892, 41.76453, 41.93184, 42.09073, 42.24112, 42.38291, 42.516, 
    42.64032, 42.75576, 42.86227, 42.95976, 43.04817, 43.12745, 43.19752, 
    43.25835, 43.3099, 43.35213, 43.385, 43.4085, 43.4226, 43.42731, 43.4226, 
    43.4085, 43.385, 43.35213, 43.3099, 43.25835, 43.19752, 43.12745, 
    43.04817, 42.95976, 42.86227, 42.75576, 42.64032, 42.516, 42.38291, 
    42.24112, 42.09073, 41.93184, 41.76453, 41.58892, 41.40512, 41.21324, 
    41.01338, 40.80568, 40.59023, 40.36718, 40.13664, 39.89874, 39.6536, 
    39.40136, 39.14214, 38.87608, 38.6033, 38.32394, 38.03813, 37.746, 
    37.44768, 37.14331, 36.83301, 36.51693, 36.19517, 35.86789, 35.53519, 
    35.19722, 34.8541, 34.50594, 34.15289, 33.79504,
  34.52972, 34.89117, 35.24767, 35.59911, 35.94537, 36.28631, 36.62183, 
    36.95179, 37.27608, 37.59457, 37.90713, 38.21363, 38.51395, 38.80796, 
    39.09554, 39.37654, 39.65086, 39.91835, 40.1789, 40.43238, 40.67865, 
    40.9176, 41.14911, 41.37305, 41.5893, 41.79774, 41.99827, 42.19077, 
    42.37512, 42.55122, 42.71897, 42.87827, 43.02901, 43.17111, 43.30448, 
    43.42903, 43.54469, 43.65138, 43.74903, 43.83758, 43.91697, 43.98714, 
    44.04806, 44.09967, 44.14195, 44.17486, 44.19839, 44.21251, 44.21722, 
    44.21251, 44.19839, 44.17486, 44.14195, 44.09967, 44.04806, 43.98714, 
    43.91697, 43.83758, 43.74903, 43.65138, 43.54469, 43.42903, 43.30448, 
    43.17111, 43.02901, 42.87827, 42.71897, 42.55122, 42.37512, 42.19077, 
    41.99827, 41.79774, 41.5893, 41.37305, 41.14911, 40.9176, 40.67865, 
    40.43238, 40.1789, 39.91835, 39.65086, 39.37654, 39.09554, 38.80796, 
    38.51395, 38.21363, 37.90713, 37.59457, 37.27608, 36.95179, 36.62183, 
    36.28631, 35.94537, 35.59911, 35.24767, 34.89117, 34.52972,
  35.26439, 35.62921, 35.98892, 36.34341, 36.69255, 37.03624, 37.37434, 
    37.70675, 38.03334, 38.354, 38.66859, 38.977, 39.27911, 39.57478, 
    39.8639, 40.14635, 40.42199, 40.69072, 40.9524, 41.20691, 41.45414, 
    41.69396, 41.92625, 42.15091, 42.36781, 42.57683, 42.77788, 42.97084, 
    43.1556, 43.33206, 43.50012, 43.65969, 43.81068, 43.95298, 44.08652, 
    44.21122, 44.32701, 44.4338, 44.53154, 44.62016, 44.6996, 44.76982, 
    44.83077, 44.88241, 44.9247, 44.95763, 44.98116, 44.99529, 45, 44.99529, 
    44.98116, 44.95763, 44.9247, 44.88241, 44.83077, 44.76982, 44.6996, 
    44.62016, 44.53154, 44.4338, 44.32701, 44.21122, 44.08652, 43.95298, 
    43.81068, 43.65969, 43.50012, 43.33206, 43.1556, 42.97084, 42.77788, 
    42.57683, 42.36781, 42.15091, 41.92625, 41.69396, 41.45414, 41.20691, 
    40.9524, 40.69072, 40.42199, 40.14635, 39.8639, 39.57478, 39.27911, 
    38.977, 38.66859, 38.354, 38.03334, 37.70675, 37.37434, 37.03624, 
    36.69255, 36.34341, 35.98892, 35.62921, 35.26439 ;

 grid_lont =
  305.3905, 306.1768, 306.9704, 307.7711, 308.579, 309.3943, 310.2169, 
    311.0468, 311.8842, 312.729, 313.5811, 314.4407, 315.3077, 316.1821, 
    317.0639, 317.9529, 318.8493, 319.7529, 320.6636, 321.5814, 322.5062, 
    323.4379, 324.3764, 325.3216, 326.2732, 327.2313, 328.1955, 329.1658, 
    330.142, 331.1238, 332.1111, 333.1037, 334.1013, 335.1036, 336.1105, 
    337.1216, 338.1368, 339.1556, 340.1779, 341.2032, 342.2314, 343.2621, 
    344.295, 345.3297, 346.366, 347.4034, 348.4417, 349.4805, 350.5195, 
    351.5583, 352.5966, 353.634, 354.6703, 355.705, 356.7379, 357.7686, 
    358.7968, 359.8221, 0.8443806, 1.86322, 2.878349, 3.889488, 4.896363, 
    5.898713, 6.896286, 7.888842, 8.876152, 9.857996, 10.83417, 11.80448, 
    12.76874, 13.72678, 14.67844, 15.62358, 16.56206, 17.49376, 18.41857, 
    19.33638, 20.24712, 21.1507, 22.04705, 22.93612, 23.81787, 24.69226, 
    25.55925, 26.41885, 27.27102, 28.11579, 28.95315, 29.78312, 30.60571, 
    31.42098, 32.22894, 33.02964, 33.82314, 34.60948,
  305.3906, 306.1769, 306.9704, 307.7711, 308.579, 309.3943, 310.2169, 
    311.0469, 311.8842, 312.729, 313.5812, 314.4408, 315.3078, 316.1822, 
    317.0639, 317.953, 318.8493, 319.7529, 320.6636, 321.5815, 322.5063, 
    323.438, 324.3764, 325.3216, 326.2733, 327.2313, 328.1956, 329.1659, 
    330.142, 331.1239, 332.1112, 333.1037, 334.1013, 335.1037, 336.1105, 
    337.1217, 338.1368, 339.1556, 340.1779, 341.2033, 342.2314, 343.2621, 
    344.295, 345.3297, 346.366, 347.4034, 348.4417, 349.4805, 350.5195, 
    351.5583, 352.5966, 353.634, 354.6703, 355.705, 356.7379, 357.7686, 
    358.7967, 359.8221, 0.8443687, 1.863207, 2.878335, 3.889472, 4.896347, 
    5.898695, 6.896268, 7.888824, 8.876132, 9.857976, 10.83415, 11.80446, 
    12.76871, 13.72675, 14.67842, 15.62356, 16.56204, 17.49373, 18.41854, 
    19.33636, 20.24709, 21.15067, 22.04702, 22.93609, 23.81784, 24.69223, 
    25.55922, 26.41882, 27.27099, 28.11576, 28.95312, 29.78308, 30.60568, 
    31.42095, 32.22891, 33.02961, 33.82311, 34.60945,
  305.3906, 306.1769, 306.9704, 307.7711, 308.5791, 309.3943, 310.2169, 
    311.0469, 311.8843, 312.729, 313.5812, 314.4408, 315.3078, 316.1822, 
    317.0639, 317.953, 318.8494, 319.7529, 320.6637, 321.5815, 322.5063, 
    323.438, 324.3765, 325.3216, 326.2733, 327.2313, 328.1956, 329.1659, 
    330.1421, 331.1239, 332.1112, 333.1038, 334.1013, 335.1037, 336.1105, 
    337.1217, 338.1368, 339.1556, 340.1779, 341.2033, 342.2315, 343.2621, 
    344.295, 345.3297, 346.366, 347.4034, 348.4417, 349.4805, 350.5195, 
    351.5583, 352.5966, 353.634, 354.6703, 355.705, 356.7379, 357.7685, 
    358.7967, 359.8221, 0.8443567, 1.863194, 2.878321, 3.889457, 4.89633, 
    5.898679, 6.89625, 7.888804, 8.876112, 9.857955, 10.83413, 11.80443, 
    12.76869, 13.72673, 14.67839, 15.62353, 16.56201, 17.49371, 18.41851, 
    19.33633, 20.24706, 21.15064, 22.04699, 22.93606, 23.81781, 24.6922, 
    25.55919, 26.41879, 27.27096, 28.11573, 28.95308, 29.78305, 30.60565, 
    31.42092, 32.22888, 33.02958, 33.82308, 34.60942,
  305.3906, 306.1769, 306.9705, 307.7711, 308.5791, 309.3944, 310.217, 
    311.0469, 311.8843, 312.7291, 313.5812, 314.4408, 315.3078, 316.1822, 
    317.064, 317.953, 318.8494, 319.753, 320.6637, 321.5815, 322.5063, 
    323.438, 324.3765, 325.3216, 326.2733, 327.2313, 328.1956, 329.1659, 
    330.1421, 331.1239, 332.1112, 333.1038, 334.1013, 335.1037, 336.1106, 
    337.1217, 338.1368, 339.1557, 340.1779, 341.2033, 342.2315, 343.2622, 
    344.295, 345.3297, 346.366, 347.4034, 348.4417, 349.4805, 350.5195, 
    351.5583, 352.5966, 353.634, 354.6703, 355.705, 356.7378, 357.7685, 
    358.7967, 359.8221, 0.8443446, 1.863181, 2.878307, 3.889442, 4.896314, 
    5.898661, 6.896232, 7.888785, 8.876092, 9.857934, 10.83411, 11.80441, 
    12.76867, 13.72671, 14.67837, 15.62351, 16.56199, 17.49368, 18.41849, 
    19.3363, 20.24703, 21.15061, 22.04696, 22.93604, 23.81778, 24.69217, 
    25.55916, 26.41875, 27.27093, 28.1157, 28.95305, 29.78302, 30.60562, 
    31.42089, 32.22885, 33.02955, 33.82305, 34.60939,
  305.3907, 306.177, 306.9705, 307.7712, 308.5791, 309.3944, 310.217, 
    311.047, 311.8843, 312.7291, 313.5813, 314.4409, 315.3079, 316.1823, 
    317.064, 317.9531, 318.8494, 319.753, 320.6637, 321.5815, 322.5063, 
    323.438, 324.3765, 325.3217, 326.2733, 327.2314, 328.1956, 329.1659, 
    330.1421, 331.1239, 332.1112, 333.1038, 334.1013, 335.1037, 336.1106, 
    337.1217, 338.1368, 339.1557, 340.1779, 341.2033, 342.2315, 343.2622, 
    344.295, 345.3297, 346.366, 347.4034, 348.4417, 349.4805, 350.5195, 
    351.5583, 352.5966, 353.634, 354.6703, 355.705, 356.7378, 357.7685, 
    358.7967, 359.8221, 0.8443325, 1.863167, 2.878293, 3.889427, 4.896298, 
    5.898644, 6.896214, 7.888766, 8.876072, 9.857914, 10.83408, 11.80439, 
    12.76865, 13.72668, 14.67834, 15.62348, 16.56196, 17.49366, 18.41846, 
    19.33627, 20.24701, 21.15058, 22.04693, 22.93601, 23.81775, 24.69214, 
    25.55913, 26.41872, 27.2709, 28.11567, 28.95302, 29.78299, 30.60559, 
    31.42085, 32.22882, 33.02952, 33.82301, 34.60936,
  305.3907, 306.177, 306.9705, 307.7712, 308.5792, 309.3944, 310.217, 
    311.047, 311.8844, 312.7291, 313.5813, 314.4409, 315.3079, 316.1823, 
    317.064, 317.9531, 318.8495, 319.753, 320.6638, 321.5816, 322.5064, 
    323.4381, 324.3766, 325.3217, 326.2733, 327.2314, 328.1956, 329.1659, 
    330.1421, 331.124, 332.1113, 333.1038, 334.1014, 335.1037, 336.1106, 
    337.1217, 338.1368, 339.1557, 340.1779, 341.2033, 342.2315, 343.2622, 
    344.295, 345.3298, 346.366, 347.4034, 348.4417, 349.4805, 350.5195, 
    351.5583, 352.5966, 353.634, 354.6702, 355.705, 356.7378, 357.7685, 
    358.7967, 359.8221, 0.8443203, 1.863154, 2.878278, 3.889411, 4.896282, 
    5.898627, 6.896195, 7.888747, 8.876052, 9.857893, 10.83406, 11.80437, 
    12.76862, 13.72666, 14.67832, 15.62346, 16.56193, 17.49363, 18.41843, 
    19.33625, 20.24698, 21.15055, 22.04691, 22.93598, 23.81772, 24.69211, 
    25.5591, 26.4187, 27.27087, 28.11563, 28.95299, 29.78296, 30.60556, 
    31.42082, 32.22879, 33.02949, 33.82298, 34.60933,
  305.3907, 306.177, 306.9706, 307.7712, 308.5792, 309.3945, 310.2171, 
    311.047, 311.8844, 312.7292, 313.5813, 314.4409, 315.3079, 316.1823, 
    317.0641, 317.9531, 318.8495, 319.7531, 320.6638, 321.5816, 322.5064, 
    323.4381, 324.3766, 325.3217, 326.2734, 327.2314, 328.1956, 329.166, 
    330.1421, 331.124, 332.1113, 333.1038, 334.1014, 335.1037, 336.1106, 
    337.1217, 338.1369, 339.1557, 340.1779, 341.2033, 342.2315, 343.2622, 
    344.295, 345.3298, 346.366, 347.4034, 348.4417, 349.4805, 350.5195, 
    351.5583, 352.5966, 353.634, 354.6702, 355.705, 356.7378, 357.7685, 
    358.7967, 359.8221, 0.844308, 1.863141, 2.878264, 3.889396, 4.896265, 
    5.89861, 6.896177, 7.888728, 8.876032, 9.857872, 10.83404, 11.80434, 
    12.7686, 13.72663, 14.67829, 15.62343, 16.56191, 17.4936, 18.41841, 
    19.33622, 20.24695, 21.15053, 22.04688, 22.93595, 23.81769, 24.69208, 
    25.55907, 26.41866, 27.27084, 28.1156, 28.95296, 29.78293, 30.60553, 
    31.42079, 32.22876, 33.02946, 33.82296, 34.60929,
  305.3907, 306.1771, 306.9706, 307.7713, 308.5792, 309.3945, 310.2171, 
    311.0471, 311.8844, 312.7292, 313.5814, 314.4409, 315.308, 316.1823, 
    317.0641, 317.9532, 318.8495, 319.7531, 320.6638, 321.5816, 322.5064, 
    323.4381, 324.3766, 325.3217, 326.2734, 327.2314, 328.1957, 329.166, 
    330.1422, 331.124, 332.1113, 333.1039, 334.1014, 335.1038, 336.1106, 
    337.1218, 338.1369, 339.1557, 340.1779, 341.2033, 342.2315, 343.2622, 
    344.295, 345.3298, 346.366, 347.4034, 348.4417, 349.4805, 350.5195, 
    351.5583, 352.5966, 353.634, 354.6702, 355.705, 356.7378, 357.7685, 
    358.7967, 359.8221, 0.8442957, 1.863127, 2.878249, 3.889381, 4.896249, 
    5.898592, 6.896159, 7.888709, 8.876012, 9.857851, 10.83402, 11.80432, 
    12.76858, 13.72661, 14.67827, 15.6234, 16.56188, 17.49358, 18.41838, 
    19.33619, 20.24692, 21.1505, 22.04685, 22.93592, 23.81767, 24.69205, 
    25.55904, 26.41864, 27.27081, 28.11558, 28.95293, 29.7829, 30.6055, 
    31.42076, 32.22873, 33.02943, 33.82293, 34.60926,
  305.3908, 306.1771, 306.9706, 307.7713, 308.5793, 309.3945, 310.2171, 
    311.0471, 311.8845, 312.7292, 313.5814, 314.441, 315.308, 316.1824, 
    317.0641, 317.9532, 318.8495, 319.7531, 320.6638, 321.5816, 322.5064, 
    323.4381, 324.3766, 325.3217, 326.2734, 327.2314, 328.1957, 329.166, 
    330.1422, 331.124, 332.1113, 333.1039, 334.1014, 335.1038, 336.1106, 
    337.1218, 338.1369, 339.1557, 340.178, 341.2033, 342.2315, 343.2622, 
    344.2951, 345.3298, 346.366, 347.4034, 348.4417, 349.4805, 350.5195, 
    351.5583, 352.5966, 353.634, 354.6702, 355.7049, 356.7378, 357.7685, 
    358.7967, 359.822, 0.8442835, 1.863114, 2.878235, 3.889365, 4.896233, 
    5.898575, 6.896141, 7.88869, 8.875992, 9.85783, 10.834, 11.8043, 
    12.76855, 13.72659, 14.67825, 15.62338, 16.56186, 17.49355, 18.41835, 
    19.33616, 20.2469, 21.15047, 22.04682, 22.93589, 23.81764, 24.69202, 
    25.55902, 26.41861, 27.27078, 28.11555, 28.9529, 29.78287, 30.60547, 
    31.42073, 32.22869, 33.0294, 33.8229, 34.60923,
  305.3908, 306.1771, 306.9706, 307.7713, 308.5793, 309.3946, 310.2172, 
    311.0471, 311.8845, 312.7292, 313.5814, 314.441, 315.308, 316.1824, 
    317.0641, 317.9532, 318.8495, 319.7531, 320.6638, 321.5817, 322.5065, 
    323.4382, 324.3766, 325.3218, 326.2734, 327.2315, 328.1957, 329.166, 
    330.1422, 331.124, 332.1113, 333.1039, 334.1014, 335.1038, 336.1107, 
    337.1218, 338.1369, 339.1557, 340.178, 341.2033, 342.2315, 343.2622, 
    344.2951, 345.3298, 346.366, 347.4034, 348.4417, 349.4805, 350.5195, 
    351.5583, 352.5966, 353.634, 354.6702, 355.7049, 356.7378, 357.7685, 
    358.7967, 359.822, 0.8442712, 1.863101, 2.878221, 3.88935, 4.896216, 
    5.898557, 6.896122, 7.88867, 8.875972, 9.857809, 10.83398, 11.80428, 
    12.76853, 13.72656, 14.67822, 15.62335, 16.56183, 17.49352, 18.41833, 
    19.33614, 20.24687, 21.15044, 22.04679, 22.93586, 23.81761, 24.69199, 
    25.55899, 26.41858, 27.27075, 28.11552, 28.95288, 29.78284, 30.60544, 
    31.4207, 32.22867, 33.02937, 33.82287, 34.60921,
  305.3908, 306.1772, 306.9706, 307.7714, 308.5793, 309.3946, 310.2172, 
    311.0471, 311.8845, 312.7293, 313.5815, 314.441, 315.308, 316.1824, 
    317.0642, 317.9532, 318.8496, 319.7531, 320.6639, 321.5817, 322.5065, 
    323.4382, 324.3767, 325.3218, 326.2735, 327.2315, 328.1957, 329.166, 
    330.1422, 331.1241, 332.1114, 333.1039, 334.1015, 335.1038, 336.1107, 
    337.1218, 338.1369, 339.1557, 340.178, 341.2034, 342.2315, 343.2622, 
    344.2951, 345.3298, 346.366, 347.4034, 348.4417, 349.4805, 350.5195, 
    351.5583, 352.5966, 353.634, 354.6702, 355.7049, 356.7378, 357.7685, 
    358.7966, 359.822, 0.8442588, 1.863087, 2.878206, 3.889334, 4.8962, 
    5.89854, 6.896104, 7.888651, 8.875953, 9.857789, 10.83395, 11.80425, 
    12.76851, 13.72654, 14.6782, 15.62333, 16.56181, 17.4935, 18.4183, 
    19.33611, 20.24684, 21.15042, 22.04676, 22.93583, 23.81758, 24.69196, 
    25.55896, 26.41855, 27.27073, 28.11549, 28.95284, 29.78281, 30.60541, 
    31.42068, 32.22864, 33.02934, 33.82284, 34.60918,
  305.3908, 306.1772, 306.9707, 307.7714, 308.5793, 309.3946, 310.2172, 
    311.0472, 311.8846, 312.7293, 313.5815, 314.4411, 315.3081, 316.1824, 
    317.0642, 317.9532, 318.8496, 319.7532, 320.6639, 321.5817, 322.5065, 
    323.4382, 324.3767, 325.3218, 326.2735, 327.2315, 328.1958, 329.1661, 
    330.1422, 331.1241, 332.1114, 333.1039, 334.1015, 335.1038, 336.1107, 
    337.1218, 338.1369, 339.1558, 340.178, 341.2034, 342.2315, 343.2622, 
    344.2951, 345.3298, 346.366, 347.4034, 348.4417, 349.4805, 350.5195, 
    351.5583, 352.5966, 353.634, 354.6702, 355.7049, 356.7378, 357.7685, 
    358.7966, 359.822, 0.8442466, 1.863074, 2.878192, 3.889319, 4.896183, 
    5.898523, 6.896086, 7.888632, 8.875933, 9.857768, 10.83393, 11.80423, 
    12.76848, 13.72652, 14.67817, 15.62331, 16.56178, 17.49347, 18.41828, 
    19.33608, 20.24681, 21.15039, 22.04674, 22.93581, 23.81755, 24.69193, 
    25.55893, 26.41852, 27.2707, 28.11546, 28.95282, 29.78278, 30.60538, 
    31.42065, 32.22861, 33.02932, 33.82281, 34.60915,
  305.3909, 306.1772, 306.9707, 307.7714, 308.5794, 309.3947, 310.2173, 
    311.0472, 311.8846, 312.7293, 313.5815, 314.4411, 315.3081, 316.1825, 
    317.0642, 317.9533, 318.8496, 319.7532, 320.6639, 321.5818, 322.5066, 
    323.4382, 324.3767, 325.3218, 326.2735, 327.2315, 328.1958, 329.1661, 
    330.1422, 331.1241, 332.1114, 333.1039, 334.1015, 335.1038, 336.1107, 
    337.1218, 338.1369, 339.1558, 340.178, 341.2034, 342.2316, 343.2622, 
    344.2951, 345.3298, 346.366, 347.4035, 348.4417, 349.4805, 350.5195, 
    351.5583, 352.5965, 353.634, 354.6702, 355.7049, 356.7378, 357.7684, 
    358.7966, 359.822, 0.8442343, 1.863061, 2.878178, 3.889304, 4.896167, 
    5.898506, 6.896068, 7.888614, 8.875913, 9.857747, 10.83391, 11.80421, 
    12.76846, 13.72649, 14.67815, 15.62328, 16.56175, 17.49345, 18.41825, 
    19.33606, 20.24679, 21.15036, 22.04671, 22.93578, 23.81752, 24.69191, 
    25.5589, 26.41849, 27.27067, 28.11543, 28.95279, 29.78276, 30.60536, 
    31.42062, 32.22858, 33.02929, 33.82278, 34.60912,
  305.3909, 306.1772, 306.9707, 307.7715, 308.5794, 309.3947, 310.2173, 
    311.0472, 311.8846, 312.7294, 313.5815, 314.4411, 315.3081, 316.1825, 
    317.0642, 317.9533, 318.8497, 319.7532, 320.664, 321.5818, 322.5066, 
    323.4383, 324.3767, 325.3219, 326.2735, 327.2316, 328.1958, 329.1661, 
    330.1423, 331.1241, 332.1114, 333.1039, 334.1015, 335.1039, 336.1107, 
    337.1218, 338.137, 339.1558, 340.178, 341.2034, 342.2316, 343.2622, 
    344.2951, 345.3298, 346.366, 347.4035, 348.4417, 349.4805, 350.5195, 
    351.5583, 352.5965, 353.634, 354.6702, 355.7049, 356.7378, 357.7684, 
    358.7966, 359.822, 0.8442221, 1.863047, 2.878163, 3.889288, 4.896151, 
    5.898489, 6.89605, 7.888595, 8.875893, 9.857727, 10.83389, 11.80419, 
    12.76844, 13.72647, 14.67813, 15.62326, 16.56173, 17.49342, 18.41822, 
    19.33603, 20.24676, 21.15034, 22.04668, 22.93575, 23.8175, 24.69188, 
    25.55888, 26.41846, 27.27064, 28.1154, 28.95276, 29.78273, 30.60533, 
    31.42059, 32.22855, 33.02926, 33.82276, 34.6091,
  305.3909, 306.1773, 306.9708, 307.7715, 308.5794, 309.3947, 310.2173, 
    311.0473, 311.8846, 312.7294, 313.5816, 314.4412, 315.3081, 316.1825, 
    317.0643, 317.9533, 318.8497, 319.7533, 320.664, 321.5818, 322.5066, 
    323.4383, 324.3768, 325.3219, 326.2736, 327.2316, 328.1958, 329.1661, 
    330.1423, 331.1241, 332.1114, 333.104, 334.1015, 335.1039, 336.1107, 
    337.1219, 338.137, 339.1558, 340.178, 341.2034, 342.2316, 343.2622, 
    344.2951, 345.3298, 346.3661, 347.4035, 348.4417, 349.4805, 350.5195, 
    351.5583, 352.5965, 353.6339, 354.6702, 355.7049, 356.7378, 357.7684, 
    358.7966, 359.822, 0.84421, 1.863034, 2.878149, 3.889273, 4.896135, 
    5.898471, 6.896032, 7.888576, 8.875874, 9.857707, 10.83387, 11.80417, 
    12.76842, 13.72645, 14.6781, 15.62323, 16.56171, 17.4934, 18.4182, 
    19.33601, 20.24674, 21.15031, 22.04666, 22.93573, 23.81747, 24.69185, 
    25.55885, 26.41844, 27.27061, 28.11538, 28.95273, 29.7827, 30.6053, 
    31.42057, 32.22853, 33.02924, 33.82273, 34.60907,
  305.391, 306.1773, 306.9708, 307.7715, 308.5795, 309.3947, 310.2173, 
    311.0473, 311.8846, 312.7294, 313.5816, 314.4412, 315.3082, 316.1826, 
    317.0643, 317.9534, 318.8497, 319.7533, 320.664, 321.5818, 322.5066, 
    323.4383, 324.3768, 325.3219, 326.2736, 327.2316, 328.1959, 329.1661, 
    330.1423, 331.1241, 332.1115, 333.104, 334.1015, 335.1039, 336.1107, 
    337.1219, 338.137, 339.1558, 340.178, 341.2034, 342.2316, 343.2623, 
    344.2951, 345.3298, 346.3661, 347.4035, 348.4417, 349.4805, 350.5195, 
    351.5583, 352.5965, 353.6339, 354.6702, 355.7049, 356.7377, 357.7684, 
    358.7966, 359.822, 0.844198, 1.863021, 2.878135, 3.889258, 4.896119, 
    5.898455, 6.896014, 7.888557, 8.875854, 9.857687, 10.83385, 11.80414, 
    12.76839, 13.72643, 14.67808, 15.62321, 16.56168, 17.49337, 18.41817, 
    19.33598, 20.24671, 21.15028, 22.04663, 22.9357, 23.81744, 24.69183, 
    25.55882, 26.41841, 27.27059, 28.11535, 28.95271, 29.78267, 30.60528, 
    31.42054, 32.2285, 33.02921, 33.8227, 34.60905,
  305.391, 306.1773, 306.9708, 307.7715, 308.5795, 309.3947, 310.2173, 
    311.0473, 311.8847, 312.7294, 313.5816, 314.4412, 315.3082, 316.1826, 
    317.0643, 317.9534, 318.8497, 319.7533, 320.664, 321.5818, 322.5067, 
    323.4384, 324.3768, 325.3219, 326.2736, 327.2316, 328.1959, 329.1662, 
    330.1423, 331.1242, 332.1115, 333.104, 334.1016, 335.1039, 336.1107, 
    337.1219, 338.137, 339.1558, 340.1781, 341.2034, 342.2316, 343.2623, 
    344.2951, 345.3298, 346.3661, 347.4035, 348.4417, 349.4805, 350.5195, 
    351.5583, 352.5965, 353.6339, 354.6702, 355.7049, 356.7377, 357.7684, 
    358.7966, 359.8219, 0.844186, 1.863008, 2.878121, 3.889243, 4.896103, 
    5.898438, 6.895997, 7.888539, 8.875834, 9.857667, 10.83383, 11.80412, 
    12.76837, 13.7264, 14.67806, 15.62319, 16.56166, 17.49335, 18.41815, 
    19.33596, 20.24669, 21.15026, 22.04661, 22.93567, 23.81742, 24.6918, 
    25.5588, 26.41838, 27.27056, 28.11532, 28.95268, 29.78265, 30.60525, 
    31.42051, 32.22848, 33.02918, 33.82268, 34.60902,
  305.391, 306.1773, 306.9709, 307.7715, 308.5795, 309.3948, 310.2174, 
    311.0473, 311.8847, 312.7295, 313.5816, 314.4412, 315.3082, 316.1826, 
    317.0644, 317.9534, 318.8498, 319.7533, 320.6641, 321.5819, 322.5067, 
    323.4384, 324.3768, 325.322, 326.2736, 327.2317, 328.1959, 329.1662, 
    330.1424, 331.1242, 332.1115, 333.104, 334.1016, 335.1039, 336.1108, 
    337.1219, 338.137, 339.1558, 340.1781, 341.2034, 342.2316, 343.2623, 
    344.2951, 345.3298, 346.3661, 347.4035, 348.4417, 349.4805, 350.5195, 
    351.5583, 352.5965, 353.6339, 354.6702, 355.7049, 356.7377, 357.7684, 
    358.7966, 359.8219, 0.8441741, 1.862995, 2.878107, 3.889229, 4.896087, 
    5.898421, 6.895979, 7.888521, 8.875816, 9.857647, 10.83381, 11.8041, 
    12.76835, 13.72638, 14.67803, 15.62316, 16.56163, 17.49333, 18.41813, 
    19.33593, 20.24666, 21.15023, 22.04658, 22.93565, 23.81739, 24.69177, 
    25.55877, 26.41836, 27.27054, 28.1153, 28.95266, 29.78262, 30.60522, 
    31.42049, 32.22845, 33.02916, 33.82265, 34.609,
  305.391, 306.1774, 306.9709, 307.7716, 308.5795, 309.3948, 310.2174, 
    311.0474, 311.8847, 312.7295, 313.5817, 314.4413, 315.3083, 316.1826, 
    317.0644, 317.9534, 318.8498, 319.7534, 320.6641, 321.5819, 322.5067, 
    323.4384, 324.3769, 325.322, 326.2737, 327.2317, 328.1959, 329.1662, 
    330.1424, 331.1242, 332.1115, 333.104, 334.1016, 335.1039, 336.1108, 
    337.1219, 338.137, 339.1558, 340.1781, 341.2034, 342.2316, 343.2623, 
    344.2951, 345.3298, 346.3661, 347.4035, 348.4417, 349.4805, 350.5195, 
    351.5583, 352.5965, 353.6339, 354.6702, 355.7049, 356.7377, 357.7684, 
    358.7966, 359.8219, 0.8441625, 1.862983, 2.878093, 3.889214, 4.896072, 
    5.898405, 6.895962, 7.888503, 8.875797, 9.857628, 10.83379, 11.80408, 
    12.76833, 13.72636, 14.67801, 15.62314, 16.56161, 17.4933, 18.4181, 
    19.33591, 20.24664, 21.15021, 22.04656, 22.93563, 23.81737, 24.69175, 
    25.55874, 26.41833, 27.27051, 28.11527, 28.95263, 29.7826, 30.6052, 
    31.42046, 32.22843, 33.02913, 33.82263, 34.60897,
  305.3911, 306.1774, 306.9709, 307.7716, 308.5796, 309.3948, 310.2174, 
    311.0474, 311.8847, 312.7295, 313.5817, 314.4413, 315.3083, 316.1826, 
    317.0644, 317.9535, 318.8498, 319.7534, 320.6641, 321.5819, 322.5067, 
    323.4384, 324.3769, 325.322, 326.2737, 327.2317, 328.1959, 329.1662, 
    330.1424, 331.1242, 332.1115, 333.1041, 334.1016, 335.1039, 336.1108, 
    337.1219, 338.137, 339.1559, 340.1781, 341.2034, 342.2316, 343.2623, 
    344.2951, 345.3298, 346.3661, 347.4035, 348.4417, 349.4805, 350.5195, 
    351.5583, 352.5965, 353.6339, 354.6702, 355.7049, 356.7377, 357.7684, 
    358.7966, 359.8219, 0.8441509, 1.86297, 2.87808, 3.889199, 4.896057, 
    5.898389, 6.895945, 7.888485, 8.875779, 9.857609, 10.83377, 11.80406, 
    12.76831, 13.72634, 14.67799, 15.62312, 16.56159, 17.49328, 18.41808, 
    19.33588, 20.24661, 21.15018, 22.04653, 22.9356, 23.81734, 24.69172, 
    25.55872, 26.41831, 27.27049, 28.11525, 28.95261, 29.78258, 30.60518, 
    31.42044, 32.2284, 33.02911, 33.82261, 34.60895,
  305.3911, 306.1774, 306.9709, 307.7716, 308.5796, 309.3948, 310.2174, 
    311.0474, 311.8848, 312.7295, 313.5817, 314.4413, 315.3083, 316.1827, 
    317.0644, 317.9535, 318.8499, 319.7534, 320.6641, 321.5819, 322.5067, 
    323.4384, 324.3769, 325.322, 326.2737, 327.2317, 328.196, 329.1663, 
    330.1424, 331.1242, 332.1115, 333.1041, 334.1016, 335.104, 336.1108, 
    337.1219, 338.1371, 339.1559, 340.1781, 341.2035, 342.2316, 343.2623, 
    344.2951, 345.3298, 346.3661, 347.4035, 348.4417, 349.4805, 350.5195, 
    351.5583, 352.5965, 353.6339, 354.6702, 355.7049, 356.7377, 357.7684, 
    358.7965, 359.8219, 0.8441395, 1.862958, 2.878067, 3.889185, 4.896041, 
    5.898373, 6.895928, 7.888468, 8.875761, 9.85759, 10.83375, 11.80404, 
    12.76829, 13.72632, 14.67797, 15.6231, 16.56157, 17.49326, 18.41805, 
    19.33586, 20.24659, 21.15016, 22.04651, 22.93558, 23.81732, 24.6917, 
    25.5587, 26.41829, 27.27046, 28.11522, 28.95258, 29.78255, 30.60515, 
    31.42042, 32.22838, 33.02909, 33.82259, 34.60892,
  305.3911, 306.1774, 306.9709, 307.7716, 308.5796, 309.3949, 310.2175, 
    311.0475, 311.8848, 312.7296, 313.5817, 314.4413, 315.3083, 316.1827, 
    317.0645, 317.9535, 318.8499, 319.7534, 320.6642, 321.582, 322.5068, 
    323.4384, 324.3769, 325.3221, 326.2737, 327.2317, 328.196, 329.1663, 
    330.1424, 331.1243, 332.1115, 333.1041, 334.1017, 335.104, 336.1108, 
    337.1219, 338.1371, 339.1559, 340.1781, 341.2035, 342.2316, 343.2623, 
    344.2951, 345.3298, 346.3661, 347.4035, 348.4417, 349.4805, 350.5195, 
    351.5583, 352.5965, 353.6339, 354.6702, 355.7049, 356.7377, 357.7684, 
    358.7965, 359.8219, 0.8441283, 1.862946, 2.878054, 3.889171, 4.896027, 
    5.898357, 6.895912, 7.888451, 8.875743, 9.857572, 10.83373, 11.80402, 
    12.76827, 13.7263, 14.67795, 15.62307, 16.56154, 17.49323, 18.41803, 
    19.33584, 20.24657, 21.15014, 22.04648, 22.93555, 23.8173, 24.69168, 
    25.55867, 26.41826, 27.27044, 28.1152, 28.95256, 29.78253, 30.60513, 
    31.42039, 32.22836, 33.02906, 33.82256, 34.60891,
  305.3911, 306.1775, 306.9709, 307.7717, 308.5796, 309.3949, 310.2175, 
    311.0475, 311.8848, 312.7296, 313.5818, 314.4413, 315.3083, 316.1827, 
    317.0645, 317.9536, 318.8499, 319.7534, 320.6642, 321.582, 322.5068, 
    323.4385, 324.377, 325.3221, 326.2737, 327.2318, 328.196, 329.1663, 
    330.1425, 331.1243, 332.1116, 333.1041, 334.1017, 335.104, 336.1108, 
    337.1219, 338.1371, 339.1559, 340.1781, 341.2035, 342.2316, 343.2623, 
    344.2952, 345.3299, 346.3661, 347.4035, 348.4417, 349.4805, 350.5195, 
    351.5583, 352.5965, 353.6339, 354.6701, 355.7048, 356.7377, 357.7684, 
    358.7965, 359.8219, 0.8441173, 1.862934, 2.878041, 3.889158, 4.896012, 
    5.898342, 6.895896, 7.888434, 8.875726, 9.857553, 10.83371, 11.804, 
    12.76825, 13.72628, 14.67793, 15.62305, 16.56152, 17.49321, 18.41801, 
    19.33582, 20.24654, 21.15011, 22.04646, 22.93553, 23.81727, 24.69166, 
    25.55865, 26.41824, 27.27042, 28.11518, 28.95254, 29.78251, 30.60511, 
    31.42037, 32.22834, 33.02905, 33.82254, 34.60888,
  305.3911, 306.1775, 306.971, 307.7717, 308.5797, 309.3949, 310.2175, 
    311.0475, 311.8849, 312.7296, 313.5818, 314.4414, 315.3084, 316.1827, 
    317.0645, 317.9536, 318.8499, 319.7535, 320.6642, 321.582, 322.5068, 
    323.4385, 324.377, 325.3221, 326.2737, 327.2318, 328.196, 329.1663, 
    330.1425, 331.1243, 332.1116, 333.1041, 334.1017, 335.104, 336.1109, 
    337.122, 338.1371, 339.1559, 340.1781, 341.2035, 342.2317, 343.2623, 
    344.2952, 345.3299, 346.3661, 347.4035, 348.4417, 349.4805, 350.5195, 
    351.5583, 352.5965, 353.6339, 354.6701, 355.7048, 356.7377, 357.7683, 
    358.7965, 359.8219, 0.8441065, 1.862922, 2.878028, 3.889144, 4.895998, 
    5.898327, 6.89588, 7.888417, 8.875709, 9.857535, 10.83369, 11.80398, 
    12.76823, 13.72626, 14.67791, 15.62303, 16.5615, 17.49319, 18.41799, 
    19.33579, 20.24652, 21.15009, 22.04644, 22.93551, 23.81725, 24.69163, 
    25.55863, 26.41822, 27.2704, 28.11516, 28.95252, 29.78248, 30.60509, 
    31.42035, 32.22832, 33.02902, 33.82252, 34.60886,
  305.3911, 306.1775, 306.971, 307.7717, 308.5797, 309.3949, 310.2175, 
    311.0475, 311.8849, 312.7296, 313.5818, 314.4414, 315.3084, 316.1828, 
    317.0645, 317.9536, 318.8499, 319.7535, 320.6642, 321.582, 322.5068, 
    323.4385, 324.377, 325.3221, 326.2738, 327.2318, 328.196, 329.1663, 
    330.1425, 331.1243, 332.1116, 333.1041, 334.1017, 335.104, 336.1109, 
    337.122, 338.1371, 339.1559, 340.1781, 341.2035, 342.2317, 343.2623, 
    344.2952, 345.3299, 346.3661, 347.4035, 348.4417, 349.4805, 350.5195, 
    351.5583, 352.5965, 353.6339, 354.6701, 355.7048, 356.7377, 357.7683, 
    358.7965, 359.8219, 0.8440959, 1.86291, 2.878016, 3.889131, 4.895984, 
    5.898313, 6.895865, 7.888402, 8.875691, 9.857518, 10.83367, 11.80397, 
    12.76821, 13.72624, 14.67789, 15.62301, 16.56148, 17.49317, 18.41797, 
    19.33577, 20.2465, 21.15007, 22.04642, 22.93549, 23.81723, 24.69161, 
    25.55861, 26.4182, 27.27037, 28.11514, 28.9525, 29.78246, 30.60506, 
    31.42033, 32.22829, 33.029, 33.8225, 34.60884,
  305.3912, 306.1775, 306.971, 307.7717, 308.5797, 309.395, 310.2176, 
    311.0475, 311.8849, 312.7296, 313.5818, 314.4414, 315.3084, 316.1828, 
    317.0645, 317.9536, 318.8499, 319.7535, 320.6642, 321.5821, 322.5068, 
    323.4385, 324.377, 325.3221, 326.2738, 327.2318, 328.196, 329.1664, 
    330.1425, 331.1243, 332.1116, 333.1042, 334.1017, 335.104, 336.1109, 
    337.122, 338.1371, 339.1559, 340.1782, 341.2035, 342.2317, 343.2623, 
    344.2952, 345.3299, 346.3661, 347.4035, 348.4417, 349.4805, 350.5195, 
    351.5583, 352.5965, 353.6339, 354.6701, 355.7048, 356.7377, 357.7683, 
    358.7965, 359.8218, 0.8440856, 1.862899, 2.878004, 3.889118, 4.89597, 
    5.898298, 6.89585, 7.888386, 8.875675, 9.857501, 10.83366, 11.80395, 
    12.76819, 13.72622, 14.67787, 15.62299, 16.56146, 17.49315, 18.41795, 
    19.33575, 20.24648, 21.15005, 22.0464, 22.93546, 23.81721, 24.69159, 
    25.55859, 26.41818, 27.27035, 28.11512, 28.95247, 29.78244, 30.60505, 
    31.42031, 32.22828, 33.02898, 33.82248, 34.60883,
  305.3912, 306.1776, 306.971, 307.7717, 308.5797, 309.395, 310.2176, 
    311.0475, 311.8849, 312.7297, 313.5818, 314.4414, 315.3084, 316.1828, 
    317.0645, 317.9536, 318.85, 319.7535, 320.6643, 321.5821, 322.5069, 
    323.4386, 324.377, 325.3221, 326.2738, 327.2318, 328.1961, 329.1664, 
    330.1425, 331.1243, 332.1116, 333.1042, 334.1017, 335.104, 336.1109, 
    337.122, 338.1371, 339.1559, 340.1782, 341.2035, 342.2317, 343.2623, 
    344.2952, 345.3299, 346.3661, 347.4035, 348.4418, 349.4805, 350.5195, 
    351.5582, 352.5965, 353.6339, 354.6701, 355.7048, 356.7377, 357.7683, 
    358.7965, 359.8218, 0.8440756, 1.862888, 2.877992, 3.889106, 4.895957, 
    5.898284, 6.895835, 7.888371, 8.87566, 9.857485, 10.83364, 11.80393, 
    12.76817, 13.7262, 14.67785, 15.62297, 16.56144, 17.49313, 18.41793, 
    19.33573, 20.24646, 21.15003, 22.04638, 22.93545, 23.81719, 24.69157, 
    25.55857, 26.41816, 27.27033, 28.1151, 28.95246, 29.78242, 30.60503, 
    31.42029, 32.22826, 33.02896, 33.82246, 34.60881,
  305.3912, 306.1776, 306.971, 307.7718, 308.5797, 309.395, 310.2176, 
    311.0476, 311.8849, 312.7297, 313.5819, 314.4415, 315.3084, 316.1828, 
    317.0646, 317.9536, 318.85, 319.7536, 320.6643, 321.5821, 322.5069, 
    323.4386, 324.377, 325.3222, 326.2738, 327.2318, 328.1961, 329.1664, 
    330.1425, 331.1244, 332.1116, 333.1042, 334.1017, 335.1041, 336.1109, 
    337.122, 338.1371, 339.1559, 340.1782, 341.2035, 342.2317, 343.2623, 
    344.2952, 345.3299, 346.3661, 347.4035, 348.4418, 349.4805, 350.5195, 
    351.5582, 352.5965, 353.6339, 354.6701, 355.7048, 356.7377, 357.7683, 
    358.7965, 359.8218, 0.8440659, 1.862878, 2.877981, 3.889094, 4.895945, 
    5.898271, 6.895822, 7.888356, 8.875645, 9.85747, 10.83362, 11.80391, 
    12.76816, 13.72618, 14.67783, 15.62296, 16.56142, 17.49311, 18.41791, 
    19.33571, 20.24644, 21.15001, 22.04636, 22.93543, 23.81717, 24.69155, 
    25.55855, 26.41814, 27.27031, 28.11508, 28.95244, 29.7824, 30.60501, 
    31.42027, 32.22824, 33.02895, 33.82244, 34.60879,
  305.3912, 306.1776, 306.9711, 307.7718, 308.5797, 309.395, 310.2176, 
    311.0476, 311.8849, 312.7297, 313.5819, 314.4415, 315.3085, 316.1829, 
    317.0646, 317.9537, 318.85, 319.7536, 320.6643, 321.5821, 322.5069, 
    323.4386, 324.3771, 325.3222, 326.2738, 327.2319, 328.1961, 329.1664, 
    330.1425, 331.1244, 332.1117, 333.1042, 334.1017, 335.1041, 336.1109, 
    337.122, 338.1371, 339.1559, 340.1782, 341.2035, 342.2317, 343.2624, 
    344.2952, 345.3299, 346.3661, 347.4035, 348.4418, 349.4805, 350.5195, 
    351.5582, 352.5965, 353.6339, 354.6701, 355.7048, 356.7376, 357.7683, 
    358.7965, 359.8218, 0.8440565, 1.862868, 2.87797, 3.889082, 4.895932, 
    5.898258, 6.895808, 7.888342, 8.875629, 9.857454, 10.83361, 11.8039, 
    12.76814, 13.72616, 14.67781, 15.62294, 16.56141, 17.4931, 18.41789, 
    19.3357, 20.24642, 21.14999, 22.04634, 22.93541, 23.81715, 24.69153, 
    25.55853, 26.41812, 27.27029, 28.11506, 28.95242, 29.78239, 30.60499, 
    31.42026, 32.22822, 33.02893, 33.82243, 34.60877,
  305.3912, 306.1776, 306.9711, 307.7718, 308.5798, 309.395, 310.2176, 
    311.0476, 311.8849, 312.7297, 313.5819, 314.4415, 315.3085, 316.1829, 
    317.0646, 317.9537, 318.85, 319.7536, 320.6643, 321.5821, 322.5069, 
    323.4386, 324.3771, 325.3222, 326.2739, 327.2319, 328.1961, 329.1664, 
    330.1425, 331.1244, 332.1117, 333.1042, 334.1017, 335.1041, 336.1109, 
    337.122, 338.1371, 339.1559, 340.1782, 341.2035, 342.2317, 343.2624, 
    344.2952, 345.3299, 346.3661, 347.4035, 348.4418, 349.4805, 350.5195, 
    351.5582, 352.5965, 353.6339, 354.6701, 355.7048, 356.7376, 357.7683, 
    358.7965, 359.8218, 0.8440474, 1.862858, 2.877959, 3.889071, 4.89592, 
    5.898245, 6.895795, 7.888328, 8.875615, 9.857439, 10.83359, 11.80388, 
    12.76812, 13.72615, 14.6778, 15.62292, 16.56139, 17.49308, 18.41787, 
    19.33568, 20.2464, 21.14997, 22.04632, 22.93539, 23.81713, 24.69151, 
    25.55851, 26.4181, 27.27028, 28.11504, 28.9524, 29.78237, 30.60497, 
    31.42024, 32.2282, 33.02891, 33.82241, 34.60876,
  305.3913, 306.1776, 306.9711, 307.7718, 308.5798, 309.3951, 310.2177, 
    311.0476, 311.885, 312.7297, 313.5819, 314.4415, 315.3085, 316.1829, 
    317.0646, 317.9537, 318.85, 319.7536, 320.6643, 321.5822, 322.5069, 
    323.4386, 324.3771, 325.3222, 326.2739, 327.2319, 328.1961, 329.1664, 
    330.1426, 331.1244, 332.1117, 333.1042, 334.1018, 335.1041, 336.1109, 
    337.122, 338.1371, 339.156, 340.1782, 341.2035, 342.2317, 343.2624, 
    344.2952, 345.3299, 346.3661, 347.4035, 348.4418, 349.4805, 350.5195, 
    351.5582, 352.5965, 353.6339, 354.6701, 355.7048, 356.7376, 357.7683, 
    358.7965, 359.8218, 0.8440387, 1.862849, 2.877949, 3.88906, 4.895909, 
    5.898233, 6.895782, 7.888315, 8.875602, 9.857426, 10.83358, 11.80387, 
    12.76811, 13.72613, 14.67778, 15.62291, 16.56137, 17.49306, 18.41786, 
    19.33566, 20.24639, 21.14996, 22.0463, 22.93537, 23.81712, 24.6915, 
    25.55849, 26.41808, 27.27026, 28.11502, 28.95238, 29.78235, 30.60496, 
    31.42022, 32.22819, 33.0289, 33.8224, 34.60874,
  305.3913, 306.1776, 306.9711, 307.7718, 308.5798, 309.3951, 310.2177, 
    311.0476, 311.885, 312.7298, 313.5819, 314.4415, 315.3085, 316.1829, 
    317.0646, 317.9537, 318.8501, 319.7536, 320.6644, 321.5822, 322.507, 
    323.4386, 324.3771, 325.3222, 326.2739, 327.2319, 328.1961, 329.1664, 
    330.1426, 331.1244, 332.1117, 333.1042, 334.1018, 335.1041, 336.111, 
    337.1221, 338.1371, 339.156, 340.1782, 341.2036, 342.2317, 343.2624, 
    344.2952, 345.3299, 346.3661, 347.4035, 348.4418, 349.4805, 350.5195, 
    351.5582, 352.5965, 353.6339, 354.6701, 355.7048, 356.7376, 357.7683, 
    358.7964, 359.8218, 0.8440303, 1.862839, 2.87794, 3.88905, 4.895898, 
    5.898222, 6.89577, 7.888302, 8.875588, 9.857411, 10.83356, 11.80385, 
    12.7681, 13.72612, 14.67777, 15.62289, 16.56136, 17.49305, 18.41784, 
    19.33565, 20.24637, 21.14994, 22.04629, 22.93536, 23.8171, 24.69148, 
    25.55848, 26.41807, 27.27024, 28.11501, 28.95237, 29.78234, 30.60494, 
    31.42021, 32.22817, 33.02888, 33.82238, 34.60873,
  305.3913, 306.1776, 306.9711, 307.7719, 308.5798, 309.3951, 310.2177, 
    311.0476, 311.885, 312.7298, 313.5819, 314.4415, 315.3085, 316.1829, 
    317.0647, 317.9537, 318.8501, 319.7536, 320.6644, 321.5822, 322.507, 
    323.4387, 324.3771, 325.3222, 326.2739, 327.2319, 328.1962, 329.1664, 
    330.1426, 331.1244, 332.1117, 333.1042, 334.1018, 335.1041, 336.111, 
    337.1221, 338.1372, 339.156, 340.1782, 341.2036, 342.2317, 343.2624, 
    344.2952, 345.3299, 346.3661, 347.4035, 348.4418, 349.4805, 350.5195, 
    351.5582, 352.5965, 353.6339, 354.6701, 355.7048, 356.7376, 357.7683, 
    358.7964, 359.8218, 0.8440224, 1.862831, 2.87793, 3.88904, 4.895887, 
    5.898211, 6.895759, 7.88829, 8.875576, 9.857399, 10.83355, 11.80384, 
    12.76808, 13.7261, 14.67775, 15.62288, 16.56134, 17.49303, 18.41783, 
    19.33563, 20.24636, 21.14993, 22.04627, 22.93534, 23.81708, 24.69147, 
    25.55846, 26.41805, 27.27023, 28.11499, 28.95235, 29.78232, 30.60493, 
    31.42019, 32.22816, 33.02887, 33.82237, 34.60871,
  305.3913, 306.1776, 306.9711, 307.7719, 308.5798, 309.3951, 310.2177, 
    311.0477, 311.885, 312.7298, 313.582, 314.4416, 315.3086, 316.1829, 
    317.0647, 317.9537, 318.8501, 319.7537, 320.6644, 321.5822, 322.507, 
    323.4387, 324.3771, 325.3223, 326.2739, 327.2319, 328.1962, 329.1665, 
    330.1426, 331.1244, 332.1117, 333.1042, 334.1018, 335.1041, 336.111, 
    337.1221, 338.1372, 339.156, 340.1782, 341.2036, 342.2317, 343.2624, 
    344.2952, 345.3299, 346.3661, 347.4035, 348.4418, 349.4805, 350.5195, 
    351.5582, 352.5965, 353.6339, 354.6701, 355.7048, 356.7376, 357.7683, 
    358.7964, 359.8218, 0.8440148, 1.862823, 2.877922, 3.889031, 4.895877, 
    5.898201, 6.895748, 7.888279, 8.875565, 9.857387, 10.83354, 11.80383, 
    12.76807, 13.72609, 14.67774, 15.62286, 16.56133, 17.49302, 18.41781, 
    19.33562, 20.24634, 21.14991, 22.04626, 22.93533, 23.81707, 24.69145, 
    25.55845, 26.41804, 27.27022, 28.11498, 28.95234, 29.78231, 30.60491, 
    31.42018, 32.22815, 33.02885, 33.82235, 34.6087,
  305.3913, 306.1776, 306.9712, 307.7719, 308.5798, 309.3951, 310.2177, 
    311.0477, 311.885, 312.7298, 313.582, 314.4416, 315.3086, 316.183, 
    317.0647, 317.9538, 318.8501, 319.7537, 320.6644, 321.5822, 322.507, 
    323.4387, 324.3771, 325.3223, 326.2739, 327.2319, 328.1962, 329.1665, 
    330.1426, 331.1245, 332.1117, 333.1042, 334.1018, 335.1041, 336.111, 
    337.1221, 338.1372, 339.156, 340.1782, 341.2036, 342.2317, 343.2624, 
    344.2952, 345.3299, 346.3661, 347.4035, 348.4418, 349.4805, 350.5195, 
    351.5582, 352.5965, 353.6339, 354.6701, 355.7048, 356.7376, 357.7683, 
    358.7964, 359.8218, 0.8440077, 1.862815, 2.877913, 3.889022, 4.895868, 
    5.89819, 6.895738, 7.888268, 8.875554, 9.857375, 10.83353, 11.80381, 
    12.76805, 13.72608, 14.67772, 15.62285, 16.56132, 17.493, 18.4178, 
    19.3356, 20.24633, 21.1499, 22.04625, 22.93531, 23.81706, 24.69144, 
    25.55843, 26.41802, 27.2702, 28.11497, 28.95233, 29.7823, 30.6049, 
    31.42017, 32.22813, 33.02884, 33.82234, 34.60869,
  305.3913, 306.1777, 306.9712, 307.7719, 308.5798, 309.3951, 310.2177, 
    311.0477, 311.885, 312.7298, 313.582, 314.4416, 315.3086, 316.183, 
    317.0647, 317.9538, 318.8501, 319.7537, 320.6644, 321.5822, 322.507, 
    323.4387, 324.3772, 325.3223, 326.2739, 327.232, 328.1962, 329.1665, 
    330.1426, 331.1245, 332.1118, 333.1043, 334.1018, 335.1041, 336.111, 
    337.1221, 338.1372, 339.156, 340.1782, 341.2036, 342.2317, 343.2624, 
    344.2952, 345.3299, 346.3661, 347.4035, 348.4418, 349.4805, 350.5195, 
    351.5582, 352.5965, 353.6339, 354.6701, 355.7048, 356.7376, 357.7683, 
    358.7964, 359.8218, 0.844001, 1.862808, 2.877906, 3.889014, 4.895859, 
    5.898181, 6.895728, 7.888258, 8.875544, 9.857365, 10.83352, 11.8038, 
    12.76804, 13.72607, 14.67771, 15.62284, 16.5613, 17.49299, 18.41779, 
    19.33559, 20.24632, 21.14989, 22.04623, 22.9353, 23.81704, 24.69143, 
    25.55842, 26.41801, 27.27019, 28.11495, 28.95231, 29.78228, 30.60489, 
    31.42015, 32.22812, 33.02883, 33.82233, 34.60868,
  305.3913, 306.1777, 306.9712, 307.7719, 308.5799, 309.3951, 310.2177, 
    311.0477, 311.8851, 312.7298, 313.582, 314.4416, 315.3086, 316.183, 
    317.0647, 317.9538, 318.8501, 319.7537, 320.6644, 321.5822, 322.507, 
    323.4387, 324.3772, 325.3223, 326.274, 327.232, 328.1962, 329.1665, 
    330.1426, 331.1245, 332.1118, 333.1043, 334.1018, 335.1042, 336.111, 
    337.1221, 338.1372, 339.156, 340.1782, 341.2036, 342.2317, 343.2624, 
    344.2952, 345.3299, 346.3661, 347.4035, 348.4418, 349.4805, 350.5195, 
    351.5582, 352.5965, 353.6339, 354.6701, 355.7048, 356.7376, 357.7683, 
    358.7964, 359.8218, 0.8439947, 1.862801, 2.877898, 3.889006, 4.895851, 
    5.898173, 6.895719, 7.888249, 8.875533, 9.857354, 10.83351, 11.80379, 
    12.76803, 13.72606, 14.6777, 15.62283, 16.56129, 17.49298, 18.41777, 
    19.33558, 20.2463, 21.14987, 22.04622, 22.93529, 23.81703, 24.69141, 
    25.55841, 26.418, 27.27018, 28.11494, 28.9523, 29.78227, 30.60488, 
    31.42014, 32.22811, 33.02882, 33.82232, 34.60867,
  305.3914, 306.1777, 306.9712, 307.7719, 308.5799, 309.3951, 310.2177, 
    311.0477, 311.8851, 312.7298, 313.582, 314.4416, 315.3086, 316.183, 
    317.0647, 317.9538, 318.8501, 319.7537, 320.6644, 321.5822, 322.507, 
    323.4387, 324.3772, 325.3223, 326.274, 327.232, 328.1962, 329.1665, 
    330.1427, 331.1245, 332.1118, 333.1043, 334.1018, 335.1042, 336.111, 
    337.1221, 338.1372, 339.156, 340.1782, 341.2036, 342.2317, 343.2624, 
    344.2952, 345.3299, 346.3661, 347.4035, 348.4418, 349.4805, 350.5195, 
    351.5582, 352.5965, 353.6339, 354.6701, 355.7048, 356.7376, 357.7683, 
    358.7964, 359.8218, 0.843989, 1.862795, 2.877892, 3.888999, 4.895844, 
    5.898165, 6.89571, 7.88824, 8.875525, 9.857346, 10.8335, 11.80378, 
    12.76802, 13.72604, 14.67769, 15.62282, 16.56128, 17.49297, 18.41776, 
    19.33557, 20.24629, 21.14986, 22.04621, 22.93528, 23.81702, 24.6914, 
    25.5584, 26.41799, 27.27017, 28.11493, 28.95229, 29.78226, 30.60487, 
    31.42013, 32.2281, 33.02881, 33.82231, 34.60866,
  305.3914, 306.1777, 306.9712, 307.7719, 308.5799, 309.3951, 310.2177, 
    311.0477, 311.8851, 312.7298, 313.582, 314.4416, 315.3086, 316.183, 
    317.0647, 317.9538, 318.8502, 319.7537, 320.6644, 321.5822, 322.507, 
    323.4387, 324.3772, 325.3223, 326.274, 327.232, 328.1962, 329.1665, 
    330.1427, 331.1245, 332.1118, 333.1043, 334.1018, 335.1042, 336.111, 
    337.1221, 338.1372, 339.156, 340.1783, 341.2036, 342.2318, 343.2624, 
    344.2952, 345.3299, 346.3661, 347.4035, 348.4418, 349.4805, 350.5195, 
    351.5582, 352.5965, 353.6339, 354.6701, 355.7048, 356.7376, 357.7682, 
    358.7964, 359.8217, 0.8439837, 1.862789, 2.877886, 3.888992, 4.895837, 
    5.898158, 6.895703, 7.888232, 8.875516, 9.857337, 10.83349, 11.80377, 
    12.76801, 13.72604, 14.67768, 15.6228, 16.56127, 17.49296, 18.41775, 
    19.33556, 20.24628, 21.14985, 22.0462, 22.93527, 23.81701, 24.69139, 
    25.55839, 26.41798, 27.27016, 28.11492, 28.95228, 29.78225, 30.60486, 
    31.42012, 32.22809, 33.0288, 33.8223, 34.60865,
  305.3914, 306.1777, 306.9712, 307.7719, 308.5799, 309.3951, 310.2177, 
    311.0477, 311.8851, 312.7299, 313.582, 314.4416, 315.3086, 316.183, 
    317.0647, 317.9538, 318.8502, 319.7537, 320.6645, 321.5822, 322.507, 
    323.4388, 324.3772, 325.3223, 326.274, 327.232, 328.1962, 329.1665, 
    330.1427, 331.1245, 332.1118, 333.1043, 334.1018, 335.1042, 336.111, 
    337.1221, 338.1372, 339.156, 340.1783, 341.2036, 342.2318, 343.2624, 
    344.2952, 345.3299, 346.3661, 347.4035, 348.4418, 349.4805, 350.5195, 
    351.5582, 352.5965, 353.6339, 354.6701, 355.7048, 356.7376, 357.7682, 
    358.7964, 359.8217, 0.8439789, 1.862784, 2.87788, 3.888986, 4.895831, 
    5.898151, 6.895696, 7.888225, 8.875509, 9.857329, 10.83348, 11.80377, 
    12.76801, 13.72603, 14.67767, 15.6228, 16.56126, 17.49295, 18.41774, 
    19.33555, 20.24627, 21.14984, 22.04619, 22.93526, 23.817, 24.69138, 
    25.55838, 26.41797, 27.27015, 28.11491, 28.95227, 29.78224, 30.60485, 
    31.42012, 32.22808, 33.02879, 33.82229, 34.60864,
  305.3914, 306.1777, 306.9712, 307.7719, 308.5799, 309.3952, 310.2178, 
    311.0477, 311.8851, 312.7299, 313.582, 314.4416, 315.3086, 316.183, 
    317.0648, 317.9538, 318.8502, 319.7537, 320.6645, 321.5823, 322.507, 
    323.4388, 324.3772, 325.3223, 326.274, 327.232, 328.1962, 329.1665, 
    330.1427, 331.1245, 332.1118, 333.1043, 334.1019, 335.1042, 336.111, 
    337.1221, 338.1372, 339.156, 340.1783, 341.2036, 342.2318, 343.2624, 
    344.2952, 345.3299, 346.3661, 347.4035, 348.4418, 349.4805, 350.5195, 
    351.5582, 352.5965, 353.6339, 354.6701, 355.7048, 356.7376, 357.7682, 
    358.7964, 359.8217, 0.8439746, 1.862779, 2.877875, 3.888981, 4.895825, 
    5.898145, 6.89569, 7.888219, 8.875503, 9.857323, 10.83347, 11.80376, 
    12.768, 13.72602, 14.67767, 15.62279, 16.56125, 17.49294, 18.41774, 
    19.33554, 20.24627, 21.14984, 22.04618, 22.93525, 23.81699, 24.69138, 
    25.55837, 26.41796, 27.27014, 28.11491, 28.95227, 29.78224, 30.60484, 
    31.42011, 32.22808, 33.02879, 33.82229, 34.60863,
  305.3914, 306.1777, 306.9712, 307.7719, 308.5799, 309.3952, 310.2178, 
    311.0477, 311.8851, 312.7299, 313.582, 314.4417, 315.3086, 316.183, 
    317.0648, 317.9538, 318.8502, 319.7538, 320.6645, 321.5823, 322.5071, 
    323.4388, 324.3772, 325.3223, 326.274, 327.232, 328.1963, 329.1665, 
    330.1427, 331.1245, 332.1118, 333.1043, 334.1019, 335.1042, 336.111, 
    337.1221, 338.1372, 339.156, 340.1783, 341.2036, 342.2318, 343.2624, 
    344.2952, 345.3299, 346.3661, 347.4035, 348.4418, 349.4805, 350.5195, 
    351.5582, 352.5965, 353.6339, 354.6701, 355.7048, 356.7376, 357.7682, 
    358.7964, 359.8217, 0.8439708, 1.862775, 2.877871, 3.888976, 4.89582, 
    5.89814, 6.895684, 7.888213, 8.875497, 9.857316, 10.83347, 11.80375, 
    12.76799, 13.72601, 14.67766, 15.62278, 16.56125, 17.49293, 18.41773, 
    19.33553, 20.24626, 21.14983, 22.04618, 22.93524, 23.81699, 24.69137, 
    25.55836, 26.41796, 27.27013, 28.1149, 28.95226, 29.78223, 30.60483, 
    31.4201, 32.22807, 33.02878, 33.82228, 34.60863,
  305.3914, 306.1777, 306.9712, 307.7719, 308.5799, 309.3952, 310.2178, 
    311.0478, 311.8851, 312.7299, 313.5821, 314.4417, 315.3086, 316.183, 
    317.0648, 317.9538, 318.8502, 319.7538, 320.6645, 321.5823, 322.5071, 
    323.4388, 324.3772, 325.3224, 326.274, 327.232, 328.1963, 329.1665, 
    330.1427, 331.1245, 332.1118, 333.1043, 334.1019, 335.1042, 336.111, 
    337.1221, 338.1372, 339.156, 340.1783, 341.2036, 342.2318, 343.2624, 
    344.2952, 345.3299, 346.3661, 347.4035, 348.4418, 349.4805, 350.5195, 
    351.5582, 352.5965, 353.6339, 354.6701, 355.7048, 356.7376, 357.7682, 
    358.7964, 359.8217, 0.8439676, 1.862772, 2.877867, 3.888972, 4.895816, 
    5.898136, 6.89568, 7.888208, 8.875491, 9.857311, 10.83346, 11.80375, 
    12.76799, 13.72601, 14.67765, 15.62278, 16.56124, 17.49293, 18.41772, 
    19.33553, 20.24625, 21.14982, 22.04617, 22.93524, 23.81698, 24.69136, 
    25.55836, 26.41795, 27.27013, 28.11489, 28.95225, 29.78222, 30.60483, 
    31.4201, 32.22807, 33.02877, 33.82228, 34.60862,
  305.3914, 306.1777, 306.9712, 307.7719, 308.5799, 309.3952, 310.2178, 
    311.0478, 311.8851, 312.7299, 313.5821, 314.4417, 315.3087, 316.183, 
    317.0648, 317.9538, 318.8502, 319.7538, 320.6645, 321.5823, 322.5071, 
    323.4388, 324.3772, 325.3224, 326.274, 327.232, 328.1963, 329.1665, 
    330.1427, 331.1245, 332.1118, 333.1043, 334.1019, 335.1042, 336.111, 
    337.1221, 338.1372, 339.156, 340.1783, 341.2036, 342.2318, 343.2624, 
    344.2952, 345.3299, 346.3661, 347.4035, 348.4418, 349.4805, 350.5195, 
    351.5582, 352.5965, 353.6339, 354.6701, 355.7048, 356.7376, 357.7682, 
    358.7964, 359.8217, 0.8439648, 1.862769, 2.877864, 3.888969, 4.895812, 
    5.898132, 6.895676, 7.888204, 8.875487, 9.857306, 10.83346, 11.80374, 
    12.76798, 13.726, 14.67765, 15.62277, 16.56124, 17.49292, 18.41772, 
    19.33552, 20.24625, 21.14982, 22.04616, 22.93523, 23.81697, 24.69136, 
    25.55835, 26.41794, 27.27012, 28.11489, 28.95225, 29.78222, 30.60482, 
    31.42009, 32.22806, 33.02877, 33.82227, 34.60862,
  305.3914, 306.1777, 306.9712, 307.7719, 308.5799, 309.3952, 310.2178, 
    311.0478, 311.8851, 312.7299, 313.5821, 314.4417, 315.3087, 316.183, 
    317.0648, 317.9538, 318.8502, 319.7538, 320.6645, 321.5823, 322.5071, 
    323.4388, 324.3772, 325.3224, 326.274, 327.232, 328.1963, 329.1665, 
    330.1427, 331.1245, 332.1118, 333.1043, 334.1019, 335.1042, 336.111, 
    337.1221, 338.1372, 339.156, 340.1783, 341.2036, 342.2318, 343.2624, 
    344.2952, 345.3299, 346.3661, 347.4035, 348.4418, 349.4805, 350.5195, 
    351.5582, 352.5965, 353.6339, 354.6701, 355.7048, 356.7376, 357.7682, 
    358.7964, 359.8217, 0.8439626, 1.862766, 2.877861, 3.888966, 4.895809, 
    5.898129, 6.895673, 7.888201, 8.875484, 9.857304, 10.83345, 11.80374, 
    12.76798, 13.726, 14.67764, 15.62277, 16.56123, 17.49292, 18.41771, 
    19.33552, 20.24624, 21.14981, 22.04616, 22.93523, 23.81697, 24.69135, 
    25.55835, 26.41794, 27.27012, 28.11488, 28.95224, 29.78222, 30.60482, 
    31.42009, 32.22805, 33.02877, 33.82227, 34.60861,
  305.3914, 306.1777, 306.9712, 307.7719, 308.5799, 309.3952, 310.2178, 
    311.0478, 311.8851, 312.7299, 313.5821, 314.4417, 315.3087, 316.183, 
    317.0648, 317.9539, 318.8502, 319.7538, 320.6645, 321.5823, 322.5071, 
    323.4388, 324.3772, 325.3224, 326.274, 327.232, 328.1963, 329.1665, 
    330.1427, 331.1245, 332.1118, 333.1043, 334.1019, 335.1042, 336.111, 
    337.1221, 338.1372, 339.156, 340.1783, 341.2036, 342.2318, 343.2624, 
    344.2952, 345.3299, 346.3661, 347.4035, 348.4418, 349.4805, 350.5195, 
    351.5582, 352.5965, 353.6339, 354.6701, 355.7048, 356.7376, 357.7682, 
    358.7964, 359.8217, 0.8439609, 1.862764, 2.877859, 3.888964, 4.895807, 
    5.898127, 6.89567, 7.888198, 8.875482, 9.857301, 10.83345, 11.80374, 
    12.76797, 13.726, 14.67764, 15.62276, 16.56123, 17.49292, 18.41771, 
    19.33552, 20.24624, 21.14981, 22.04616, 22.93522, 23.81697, 24.69135, 
    25.55835, 26.41794, 27.27012, 28.11488, 28.95224, 29.78221, 30.60482, 
    31.42008, 32.22805, 33.02876, 33.82227, 34.60861,
  305.3914, 306.1777, 306.9713, 307.7719, 308.5799, 309.3952, 310.2178, 
    311.0478, 311.8851, 312.7299, 313.5821, 314.4417, 315.3087, 316.183, 
    317.0648, 317.9539, 318.8502, 319.7538, 320.6645, 321.5823, 322.5071, 
    323.4388, 324.3772, 325.3224, 326.274, 327.232, 328.1963, 329.1666, 
    330.1427, 331.1245, 332.1118, 333.1043, 334.1019, 335.1042, 336.111, 
    337.1221, 338.1372, 339.156, 340.1783, 341.2036, 342.2318, 343.2624, 
    344.2952, 345.3299, 346.3661, 347.4035, 348.4418, 349.4805, 350.5195, 
    351.5582, 352.5965, 353.6339, 354.6701, 355.7048, 356.7376, 357.7682, 
    358.7964, 359.8217, 0.8439599, 1.862763, 2.877858, 3.888963, 4.895806, 
    5.898125, 6.895669, 7.888197, 8.87548, 9.857299, 10.83345, 11.80373, 
    12.76797, 13.72599, 14.67764, 15.62276, 16.56123, 17.49291, 18.41771, 
    19.33551, 20.24624, 21.14981, 22.04615, 22.93522, 23.81697, 24.69135, 
    25.55834, 26.41794, 27.27011, 28.11488, 28.95224, 29.78221, 30.60481, 
    31.42008, 32.22805, 33.02876, 33.82226, 34.60861,
  305.3914, 306.1777, 306.9713, 307.7719, 308.5799, 309.3952, 310.2178, 
    311.0478, 311.8851, 312.7299, 313.5821, 314.4417, 315.3087, 316.183, 
    317.0648, 317.9539, 318.8502, 319.7538, 320.6645, 321.5823, 322.5071, 
    323.4388, 324.3772, 325.3224, 326.274, 327.232, 328.1963, 329.1666, 
    330.1427, 331.1245, 332.1118, 333.1043, 334.1019, 335.1042, 336.111, 
    337.1221, 338.1372, 339.156, 340.1783, 341.2036, 342.2318, 343.2624, 
    344.2952, 345.3299, 346.3661, 347.4035, 348.4418, 349.4805, 350.5195, 
    351.5582, 352.5965, 353.6339, 354.6701, 355.7048, 356.7376, 357.7682, 
    358.7964, 359.8217, 0.8439593, 1.862763, 2.877857, 3.888962, 4.895805, 
    5.898124, 6.895668, 7.888196, 8.875479, 9.857298, 10.83345, 11.80373, 
    12.76797, 13.72599, 14.67764, 15.62276, 16.56123, 17.49291, 18.41771, 
    19.33551, 20.24624, 21.14981, 22.04615, 22.93522, 23.81697, 24.69135, 
    25.55834, 26.41793, 27.27011, 28.11488, 28.95224, 29.78221, 30.60481, 
    31.42008, 32.22805, 33.02876, 33.82226, 34.60861,
  305.3914, 306.1777, 306.9713, 307.7719, 308.5799, 309.3952, 310.2178, 
    311.0478, 311.8851, 312.7299, 313.5821, 314.4417, 315.3087, 316.183, 
    317.0648, 317.9539, 318.8502, 319.7538, 320.6645, 321.5823, 322.5071, 
    323.4388, 324.3772, 325.3224, 326.274, 327.232, 328.1963, 329.1666, 
    330.1427, 331.1245, 332.1118, 333.1043, 334.1019, 335.1042, 336.111, 
    337.1221, 338.1372, 339.156, 340.1783, 341.2036, 342.2318, 343.2624, 
    344.2952, 345.3299, 346.3661, 347.4035, 348.4418, 349.4805, 350.5195, 
    351.5582, 352.5965, 353.6339, 354.6701, 355.7048, 356.7376, 357.7682, 
    358.7964, 359.8217, 0.8439593, 1.862763, 2.877857, 3.888962, 4.895805, 
    5.898124, 6.895668, 7.888196, 8.875479, 9.857298, 10.83345, 11.80373, 
    12.76797, 13.72599, 14.67764, 15.62276, 16.56123, 17.49291, 18.41771, 
    19.33551, 20.24624, 21.14981, 22.04615, 22.93522, 23.81697, 24.69135, 
    25.55834, 26.41793, 27.27011, 28.11488, 28.95224, 29.78221, 30.60481, 
    31.42008, 32.22805, 33.02876, 33.82226, 34.60861,
  305.3914, 306.1777, 306.9713, 307.7719, 308.5799, 309.3952, 310.2178, 
    311.0478, 311.8851, 312.7299, 313.5821, 314.4417, 315.3087, 316.183, 
    317.0648, 317.9539, 318.8502, 319.7538, 320.6645, 321.5823, 322.5071, 
    323.4388, 324.3772, 325.3224, 326.274, 327.232, 328.1963, 329.1666, 
    330.1427, 331.1245, 332.1118, 333.1043, 334.1019, 335.1042, 336.111, 
    337.1221, 338.1372, 339.156, 340.1783, 341.2036, 342.2318, 343.2624, 
    344.2952, 345.3299, 346.3661, 347.4035, 348.4418, 349.4805, 350.5195, 
    351.5582, 352.5965, 353.6339, 354.6701, 355.7048, 356.7376, 357.7682, 
    358.7964, 359.8217, 0.8439599, 1.862763, 2.877858, 3.888963, 4.895806, 
    5.898125, 6.895669, 7.888197, 8.87548, 9.857299, 10.83345, 11.80373, 
    12.76797, 13.72599, 14.67764, 15.62276, 16.56123, 17.49291, 18.41771, 
    19.33551, 20.24624, 21.14981, 22.04615, 22.93522, 23.81697, 24.69135, 
    25.55834, 26.41794, 27.27011, 28.11488, 28.95224, 29.78221, 30.60481, 
    31.42008, 32.22805, 33.02876, 33.82226, 34.60861,
  305.3914, 306.1777, 306.9712, 307.7719, 308.5799, 309.3952, 310.2178, 
    311.0478, 311.8851, 312.7299, 313.5821, 314.4417, 315.3087, 316.183, 
    317.0648, 317.9539, 318.8502, 319.7538, 320.6645, 321.5823, 322.5071, 
    323.4388, 324.3772, 325.3224, 326.274, 327.232, 328.1963, 329.1665, 
    330.1427, 331.1245, 332.1118, 333.1043, 334.1019, 335.1042, 336.111, 
    337.1221, 338.1372, 339.156, 340.1783, 341.2036, 342.2318, 343.2624, 
    344.2952, 345.3299, 346.3661, 347.4035, 348.4418, 349.4805, 350.5195, 
    351.5582, 352.5965, 353.6339, 354.6701, 355.7048, 356.7376, 357.7682, 
    358.7964, 359.8217, 0.8439609, 1.862764, 2.877859, 3.888964, 4.895807, 
    5.898127, 6.89567, 7.888198, 8.875482, 9.857301, 10.83345, 11.80374, 
    12.76797, 13.726, 14.67764, 15.62276, 16.56123, 17.49292, 18.41771, 
    19.33552, 20.24624, 21.14981, 22.04616, 22.93522, 23.81697, 24.69135, 
    25.55835, 26.41794, 27.27012, 28.11488, 28.95224, 29.78221, 30.60482, 
    31.42008, 32.22805, 33.02876, 33.82227, 34.60861,
  305.3914, 306.1777, 306.9712, 307.7719, 308.5799, 309.3952, 310.2178, 
    311.0478, 311.8851, 312.7299, 313.5821, 314.4417, 315.3087, 316.183, 
    317.0648, 317.9538, 318.8502, 319.7538, 320.6645, 321.5823, 322.5071, 
    323.4388, 324.3772, 325.3224, 326.274, 327.232, 328.1963, 329.1665, 
    330.1427, 331.1245, 332.1118, 333.1043, 334.1019, 335.1042, 336.111, 
    337.1221, 338.1372, 339.156, 340.1783, 341.2036, 342.2318, 343.2624, 
    344.2952, 345.3299, 346.3661, 347.4035, 348.4418, 349.4805, 350.5195, 
    351.5582, 352.5965, 353.6339, 354.6701, 355.7048, 356.7376, 357.7682, 
    358.7964, 359.8217, 0.8439626, 1.862766, 2.877861, 3.888966, 4.895809, 
    5.898129, 6.895673, 7.888201, 8.875484, 9.857304, 10.83345, 11.80374, 
    12.76798, 13.726, 14.67764, 15.62277, 16.56123, 17.49292, 18.41771, 
    19.33552, 20.24624, 21.14981, 22.04616, 22.93523, 23.81697, 24.69135, 
    25.55835, 26.41794, 27.27012, 28.11488, 28.95224, 29.78222, 30.60482, 
    31.42009, 32.22805, 33.02877, 33.82227, 34.60861,
  305.3914, 306.1777, 306.9712, 307.7719, 308.5799, 309.3952, 310.2178, 
    311.0478, 311.8851, 312.7299, 313.5821, 314.4417, 315.3087, 316.183, 
    317.0648, 317.9538, 318.8502, 319.7538, 320.6645, 321.5823, 322.5071, 
    323.4388, 324.3772, 325.3224, 326.274, 327.232, 328.1963, 329.1665, 
    330.1427, 331.1245, 332.1118, 333.1043, 334.1019, 335.1042, 336.111, 
    337.1221, 338.1372, 339.156, 340.1783, 341.2036, 342.2318, 343.2624, 
    344.2952, 345.3299, 346.3661, 347.4035, 348.4418, 349.4805, 350.5195, 
    351.5582, 352.5965, 353.6339, 354.6701, 355.7048, 356.7376, 357.7682, 
    358.7964, 359.8217, 0.8439648, 1.862769, 2.877864, 3.888969, 4.895812, 
    5.898132, 6.895676, 7.888204, 8.875487, 9.857306, 10.83346, 11.80374, 
    12.76798, 13.726, 14.67765, 15.62277, 16.56124, 17.49292, 18.41772, 
    19.33552, 20.24625, 21.14982, 22.04616, 22.93523, 23.81697, 24.69136, 
    25.55835, 26.41794, 27.27012, 28.11489, 28.95225, 29.78222, 30.60482, 
    31.42009, 32.22806, 33.02877, 33.82227, 34.60862,
  305.3914, 306.1777, 306.9712, 307.7719, 308.5799, 309.3952, 310.2178, 
    311.0478, 311.8851, 312.7299, 313.5821, 314.4417, 315.3086, 316.183, 
    317.0648, 317.9538, 318.8502, 319.7538, 320.6645, 321.5823, 322.5071, 
    323.4388, 324.3772, 325.3224, 326.274, 327.232, 328.1963, 329.1665, 
    330.1427, 331.1245, 332.1118, 333.1043, 334.1019, 335.1042, 336.111, 
    337.1221, 338.1372, 339.156, 340.1783, 341.2036, 342.2318, 343.2624, 
    344.2952, 345.3299, 346.3661, 347.4035, 348.4418, 349.4805, 350.5195, 
    351.5582, 352.5965, 353.6339, 354.6701, 355.7048, 356.7376, 357.7682, 
    358.7964, 359.8217, 0.8439676, 1.862772, 2.877867, 3.888972, 4.895816, 
    5.898136, 6.89568, 7.888208, 8.875491, 9.857311, 10.83346, 11.80375, 
    12.76799, 13.72601, 14.67765, 15.62278, 16.56124, 17.49293, 18.41772, 
    19.33553, 20.24625, 21.14982, 22.04617, 22.93524, 23.81698, 24.69136, 
    25.55836, 26.41795, 27.27013, 28.11489, 28.95225, 29.78222, 30.60483, 
    31.4201, 32.22807, 33.02877, 33.82228, 34.60862,
  305.3914, 306.1777, 306.9712, 307.7719, 308.5799, 309.3952, 310.2178, 
    311.0477, 311.8851, 312.7299, 313.582, 314.4417, 315.3086, 316.183, 
    317.0648, 317.9538, 318.8502, 319.7538, 320.6645, 321.5823, 322.5071, 
    323.4388, 324.3772, 325.3223, 326.274, 327.232, 328.1963, 329.1665, 
    330.1427, 331.1245, 332.1118, 333.1043, 334.1019, 335.1042, 336.111, 
    337.1221, 338.1372, 339.156, 340.1783, 341.2036, 342.2318, 343.2624, 
    344.2952, 345.3299, 346.3661, 347.4035, 348.4418, 349.4805, 350.5195, 
    351.5582, 352.5965, 353.6339, 354.6701, 355.7048, 356.7376, 357.7682, 
    358.7964, 359.8217, 0.8439708, 1.862775, 2.877871, 3.888976, 4.89582, 
    5.89814, 6.895684, 7.888213, 8.875497, 9.857316, 10.83347, 11.80375, 
    12.76799, 13.72601, 14.67766, 15.62278, 16.56125, 17.49293, 18.41773, 
    19.33553, 20.24626, 21.14983, 22.04618, 22.93524, 23.81699, 24.69137, 
    25.55836, 26.41796, 27.27013, 28.1149, 28.95226, 29.78223, 30.60483, 
    31.4201, 32.22807, 33.02878, 33.82228, 34.60863,
  305.3914, 306.1777, 306.9712, 307.7719, 308.5799, 309.3952, 310.2178, 
    311.0477, 311.8851, 312.7299, 313.582, 314.4416, 315.3086, 316.183, 
    317.0648, 317.9538, 318.8502, 319.7537, 320.6645, 321.5823, 322.507, 
    323.4388, 324.3772, 325.3223, 326.274, 327.232, 328.1962, 329.1665, 
    330.1427, 331.1245, 332.1118, 333.1043, 334.1019, 335.1042, 336.111, 
    337.1221, 338.1372, 339.156, 340.1783, 341.2036, 342.2318, 343.2624, 
    344.2952, 345.3299, 346.3661, 347.4035, 348.4418, 349.4805, 350.5195, 
    351.5582, 352.5965, 353.6339, 354.6701, 355.7048, 356.7376, 357.7682, 
    358.7964, 359.8217, 0.8439746, 1.862779, 2.877875, 3.888981, 4.895825, 
    5.898145, 6.89569, 7.888219, 8.875503, 9.857323, 10.83347, 11.80376, 
    12.768, 13.72602, 14.67767, 15.62279, 16.56125, 17.49294, 18.41774, 
    19.33554, 20.24627, 21.14984, 22.04618, 22.93525, 23.81699, 24.69138, 
    25.55837, 26.41796, 27.27014, 28.11491, 28.95227, 29.78224, 30.60484, 
    31.42011, 32.22808, 33.02879, 33.82229, 34.60863,
  305.3914, 306.1777, 306.9712, 307.7719, 308.5799, 309.3951, 310.2177, 
    311.0477, 311.8851, 312.7299, 313.582, 314.4416, 315.3086, 316.183, 
    317.0647, 317.9538, 318.8502, 319.7537, 320.6645, 321.5822, 322.507, 
    323.4388, 324.3772, 325.3223, 326.274, 327.232, 328.1962, 329.1665, 
    330.1427, 331.1245, 332.1118, 333.1043, 334.1018, 335.1042, 336.111, 
    337.1221, 338.1372, 339.156, 340.1783, 341.2036, 342.2318, 343.2624, 
    344.2952, 345.3299, 346.3661, 347.4035, 348.4418, 349.4805, 350.5195, 
    351.5582, 352.5965, 353.6339, 354.6701, 355.7048, 356.7376, 357.7682, 
    358.7964, 359.8217, 0.8439789, 1.862784, 2.87788, 3.888986, 4.895831, 
    5.898151, 6.895696, 7.888225, 8.875509, 9.857329, 10.83348, 11.80377, 
    12.76801, 13.72603, 14.67767, 15.6228, 16.56126, 17.49295, 18.41774, 
    19.33555, 20.24627, 21.14984, 22.04619, 22.93526, 23.817, 24.69138, 
    25.55838, 26.41797, 27.27015, 28.11491, 28.95227, 29.78224, 30.60485, 
    31.42012, 32.22808, 33.02879, 33.82229, 34.60864,
  305.3914, 306.1777, 306.9712, 307.7719, 308.5799, 309.3951, 310.2177, 
    311.0477, 311.8851, 312.7298, 313.582, 314.4416, 315.3086, 316.183, 
    317.0647, 317.9538, 318.8502, 319.7537, 320.6644, 321.5822, 322.507, 
    323.4387, 324.3772, 325.3223, 326.274, 327.232, 328.1962, 329.1665, 
    330.1427, 331.1245, 332.1118, 333.1043, 334.1018, 335.1042, 336.111, 
    337.1221, 338.1372, 339.156, 340.1783, 341.2036, 342.2318, 343.2624, 
    344.2952, 345.3299, 346.3661, 347.4035, 348.4418, 349.4805, 350.5195, 
    351.5582, 352.5965, 353.6339, 354.6701, 355.7048, 356.7376, 357.7682, 
    358.7964, 359.8217, 0.8439837, 1.862789, 2.877886, 3.888992, 4.895837, 
    5.898158, 6.895703, 7.888232, 8.875516, 9.857337, 10.83349, 11.80377, 
    12.76801, 13.72604, 14.67768, 15.6228, 16.56127, 17.49296, 18.41775, 
    19.33556, 20.24628, 21.14985, 22.0462, 22.93527, 23.81701, 24.69139, 
    25.55839, 26.41798, 27.27016, 28.11492, 28.95228, 29.78225, 30.60486, 
    31.42012, 32.22809, 33.0288, 33.8223, 34.60865,
  305.3914, 306.1777, 306.9712, 307.7719, 308.5799, 309.3951, 310.2177, 
    311.0477, 311.8851, 312.7298, 313.582, 314.4416, 315.3086, 316.183, 
    317.0647, 317.9538, 318.8501, 319.7537, 320.6644, 321.5822, 322.507, 
    323.4387, 324.3772, 325.3223, 326.274, 327.232, 328.1962, 329.1665, 
    330.1427, 331.1245, 332.1118, 333.1043, 334.1018, 335.1042, 336.111, 
    337.1221, 338.1372, 339.156, 340.1782, 341.2036, 342.2317, 343.2624, 
    344.2952, 345.3299, 346.3661, 347.4035, 348.4418, 349.4805, 350.5195, 
    351.5582, 352.5965, 353.6339, 354.6701, 355.7048, 356.7376, 357.7683, 
    358.7964, 359.8218, 0.843989, 1.862795, 2.877892, 3.888999, 4.895844, 
    5.898165, 6.89571, 7.88824, 8.875525, 9.857346, 10.8335, 11.80378, 
    12.76802, 13.72604, 14.67769, 15.62282, 16.56128, 17.49297, 18.41776, 
    19.33557, 20.24629, 21.14986, 22.04621, 22.93528, 23.81702, 24.6914, 
    25.5584, 26.41799, 27.27017, 28.11493, 28.95229, 29.78226, 30.60487, 
    31.42013, 32.2281, 33.02881, 33.82231, 34.60866,
  305.3913, 306.1777, 306.9712, 307.7719, 308.5799, 309.3951, 310.2177, 
    311.0477, 311.8851, 312.7298, 313.582, 314.4416, 315.3086, 316.183, 
    317.0647, 317.9538, 318.8501, 319.7537, 320.6644, 321.5822, 322.507, 
    323.4387, 324.3772, 325.3223, 326.274, 327.232, 328.1962, 329.1665, 
    330.1426, 331.1245, 332.1118, 333.1043, 334.1018, 335.1042, 336.111, 
    337.1221, 338.1372, 339.156, 340.1782, 341.2036, 342.2317, 343.2624, 
    344.2952, 345.3299, 346.3661, 347.4035, 348.4418, 349.4805, 350.5195, 
    351.5582, 352.5965, 353.6339, 354.6701, 355.7048, 356.7376, 357.7683, 
    358.7964, 359.8218, 0.8439947, 1.862801, 2.877898, 3.889006, 4.895851, 
    5.898173, 6.895719, 7.888249, 8.875533, 9.857354, 10.83351, 11.80379, 
    12.76803, 13.72606, 14.6777, 15.62283, 16.56129, 17.49298, 18.41777, 
    19.33558, 20.2463, 21.14987, 22.04622, 22.93529, 23.81703, 24.69141, 
    25.55841, 26.418, 27.27018, 28.11494, 28.9523, 29.78227, 30.60488, 
    31.42014, 32.22811, 33.02882, 33.82232, 34.60867,
  305.3913, 306.1777, 306.9712, 307.7719, 308.5798, 309.3951, 310.2177, 
    311.0477, 311.885, 312.7298, 313.582, 314.4416, 315.3086, 316.183, 
    317.0647, 317.9538, 318.8501, 319.7537, 320.6644, 321.5822, 322.507, 
    323.4387, 324.3772, 325.3223, 326.2739, 327.232, 328.1962, 329.1665, 
    330.1426, 331.1245, 332.1118, 333.1043, 334.1018, 335.1041, 336.111, 
    337.1221, 338.1372, 339.156, 340.1782, 341.2036, 342.2317, 343.2624, 
    344.2952, 345.3299, 346.3661, 347.4035, 348.4418, 349.4805, 350.5195, 
    351.5582, 352.5965, 353.6339, 354.6701, 355.7048, 356.7376, 357.7683, 
    358.7964, 359.8218, 0.844001, 1.862808, 2.877906, 3.889014, 4.895859, 
    5.898181, 6.895728, 7.888258, 8.875544, 9.857365, 10.83352, 11.8038, 
    12.76804, 13.72607, 14.67771, 15.62284, 16.5613, 17.49299, 18.41779, 
    19.33559, 20.24632, 21.14989, 22.04623, 22.9353, 23.81704, 24.69143, 
    25.55842, 26.41801, 27.27019, 28.11495, 28.95231, 29.78228, 30.60489, 
    31.42015, 32.22812, 33.02883, 33.82233, 34.60868,
  305.3913, 306.1776, 306.9712, 307.7719, 308.5798, 309.3951, 310.2177, 
    311.0477, 311.885, 312.7298, 313.582, 314.4416, 315.3086, 316.183, 
    317.0647, 317.9538, 318.8501, 319.7537, 320.6644, 321.5822, 322.507, 
    323.4387, 324.3771, 325.3223, 326.2739, 327.2319, 328.1962, 329.1665, 
    330.1426, 331.1245, 332.1117, 333.1042, 334.1018, 335.1041, 336.111, 
    337.1221, 338.1372, 339.156, 340.1782, 341.2036, 342.2317, 343.2624, 
    344.2952, 345.3299, 346.3661, 347.4035, 348.4418, 349.4805, 350.5195, 
    351.5582, 352.5965, 353.6339, 354.6701, 355.7048, 356.7376, 357.7683, 
    358.7964, 359.8218, 0.8440077, 1.862815, 2.877913, 3.889022, 4.895868, 
    5.89819, 6.895738, 7.888268, 8.875554, 9.857375, 10.83353, 11.80381, 
    12.76805, 13.72608, 14.67772, 15.62285, 16.56132, 17.493, 18.4178, 
    19.3356, 20.24633, 21.1499, 22.04625, 22.93531, 23.81706, 24.69144, 
    25.55843, 26.41802, 27.2702, 28.11497, 28.95233, 29.7823, 30.6049, 
    31.42017, 32.22813, 33.02884, 33.82234, 34.60869,
  305.3913, 306.1776, 306.9711, 307.7719, 308.5798, 309.3951, 310.2177, 
    311.0477, 311.885, 312.7298, 313.582, 314.4416, 315.3086, 316.1829, 
    317.0647, 317.9537, 318.8501, 319.7537, 320.6644, 321.5822, 322.507, 
    323.4387, 324.3771, 325.3223, 326.2739, 327.2319, 328.1962, 329.1665, 
    330.1426, 331.1244, 332.1117, 333.1042, 334.1018, 335.1041, 336.111, 
    337.1221, 338.1372, 339.156, 340.1782, 341.2036, 342.2317, 343.2624, 
    344.2952, 345.3299, 346.3661, 347.4035, 348.4418, 349.4805, 350.5195, 
    351.5582, 352.5965, 353.6339, 354.6701, 355.7048, 356.7376, 357.7683, 
    358.7964, 359.8218, 0.8440148, 1.862823, 2.877922, 3.889031, 4.895877, 
    5.898201, 6.895748, 7.888279, 8.875565, 9.857387, 10.83354, 11.80383, 
    12.76807, 13.72609, 14.67774, 15.62286, 16.56133, 17.49302, 18.41781, 
    19.33562, 20.24634, 21.14991, 22.04626, 22.93533, 23.81707, 24.69145, 
    25.55845, 26.41804, 27.27022, 28.11498, 28.95234, 29.78231, 30.60491, 
    31.42018, 32.22815, 33.02885, 33.82235, 34.6087,
  305.3913, 306.1776, 306.9711, 307.7719, 308.5798, 309.3951, 310.2177, 
    311.0476, 311.885, 312.7298, 313.5819, 314.4415, 315.3085, 316.1829, 
    317.0647, 317.9537, 318.8501, 319.7536, 320.6644, 321.5822, 322.507, 
    323.4387, 324.3771, 325.3222, 326.2739, 327.2319, 328.1962, 329.1664, 
    330.1426, 331.1244, 332.1117, 333.1042, 334.1018, 335.1041, 336.111, 
    337.1221, 338.1372, 339.156, 340.1782, 341.2036, 342.2317, 343.2624, 
    344.2952, 345.3299, 346.3661, 347.4035, 348.4418, 349.4805, 350.5195, 
    351.5582, 352.5965, 353.6339, 354.6701, 355.7048, 356.7376, 357.7683, 
    358.7964, 359.8218, 0.8440224, 1.862831, 2.87793, 3.88904, 4.895887, 
    5.898211, 6.895759, 7.88829, 8.875576, 9.857399, 10.83355, 11.80384, 
    12.76808, 13.7261, 14.67775, 15.62288, 16.56134, 17.49303, 18.41783, 
    19.33563, 20.24636, 21.14993, 22.04627, 22.93534, 23.81708, 24.69147, 
    25.55846, 26.41805, 27.27023, 28.11499, 28.95235, 29.78232, 30.60493, 
    31.42019, 32.22816, 33.02887, 33.82237, 34.60871,
  305.3913, 306.1776, 306.9711, 307.7718, 308.5798, 309.3951, 310.2177, 
    311.0476, 311.885, 312.7298, 313.5819, 314.4415, 315.3085, 316.1829, 
    317.0646, 317.9537, 318.8501, 319.7536, 320.6644, 321.5822, 322.507, 
    323.4386, 324.3771, 325.3222, 326.2739, 327.2319, 328.1961, 329.1664, 
    330.1426, 331.1244, 332.1117, 333.1042, 334.1018, 335.1041, 336.111, 
    337.1221, 338.1371, 339.156, 340.1782, 341.2036, 342.2317, 343.2624, 
    344.2952, 345.3299, 346.3661, 347.4035, 348.4418, 349.4805, 350.5195, 
    351.5582, 352.5965, 353.6339, 354.6701, 355.7048, 356.7376, 357.7683, 
    358.7964, 359.8218, 0.8440303, 1.862839, 2.87794, 3.88905, 4.895898, 
    5.898222, 6.89577, 7.888302, 8.875588, 9.857411, 10.83356, 11.80385, 
    12.7681, 13.72612, 14.67777, 15.62289, 16.56136, 17.49305, 18.41784, 
    19.33565, 20.24637, 21.14994, 22.04629, 22.93536, 23.8171, 24.69148, 
    25.55848, 26.41807, 27.27024, 28.11501, 28.95237, 29.78234, 30.60494, 
    31.42021, 32.22817, 33.02888, 33.82238, 34.60873,
  305.3913, 306.1776, 306.9711, 307.7718, 308.5798, 309.3951, 310.2177, 
    311.0476, 311.885, 312.7297, 313.5819, 314.4415, 315.3085, 316.1829, 
    317.0646, 317.9537, 318.85, 319.7536, 320.6643, 321.5822, 322.5069, 
    323.4386, 324.3771, 325.3222, 326.2739, 327.2319, 328.1961, 329.1664, 
    330.1426, 331.1244, 332.1117, 333.1042, 334.1018, 335.1041, 336.1109, 
    337.122, 338.1371, 339.156, 340.1782, 341.2035, 342.2317, 343.2624, 
    344.2952, 345.3299, 346.3661, 347.4035, 348.4418, 349.4805, 350.5195, 
    351.5582, 352.5965, 353.6339, 354.6701, 355.7048, 356.7376, 357.7683, 
    358.7965, 359.8218, 0.8440387, 1.862849, 2.877949, 3.88906, 4.895909, 
    5.898233, 6.895782, 7.888315, 8.875602, 9.857426, 10.83358, 11.80387, 
    12.76811, 13.72613, 14.67778, 15.62291, 16.56137, 17.49306, 18.41786, 
    19.33566, 20.24639, 21.14996, 22.0463, 22.93537, 23.81712, 24.6915, 
    25.55849, 26.41808, 27.27026, 28.11502, 28.95238, 29.78235, 30.60496, 
    31.42022, 32.22819, 33.0289, 33.8224, 34.60874,
  305.3912, 306.1776, 306.9711, 307.7718, 308.5798, 309.395, 310.2176, 
    311.0476, 311.8849, 312.7297, 313.5819, 314.4415, 315.3085, 316.1829, 
    317.0646, 317.9537, 318.85, 319.7536, 320.6643, 321.5821, 322.5069, 
    323.4386, 324.3771, 325.3222, 326.2739, 327.2319, 328.1961, 329.1664, 
    330.1425, 331.1244, 332.1117, 333.1042, 334.1017, 335.1041, 336.1109, 
    337.122, 338.1371, 339.1559, 340.1782, 341.2035, 342.2317, 343.2624, 
    344.2952, 345.3299, 346.3661, 347.4035, 348.4418, 349.4805, 350.5195, 
    351.5582, 352.5965, 353.6339, 354.6701, 355.7048, 356.7376, 357.7683, 
    358.7965, 359.8218, 0.8440474, 1.862858, 2.877959, 3.889071, 4.89592, 
    5.898245, 6.895795, 7.888328, 8.875615, 9.857439, 10.83359, 11.80388, 
    12.76812, 13.72615, 14.6778, 15.62292, 16.56139, 17.49308, 18.41787, 
    19.33568, 20.2464, 21.14997, 22.04632, 22.93539, 23.81713, 24.69151, 
    25.55851, 26.4181, 27.27028, 28.11504, 28.9524, 29.78237, 30.60497, 
    31.42024, 32.2282, 33.02891, 33.82241, 34.60876,
  305.3912, 306.1776, 306.9711, 307.7718, 308.5797, 309.395, 310.2176, 
    311.0476, 311.8849, 312.7297, 313.5819, 314.4415, 315.3085, 316.1829, 
    317.0646, 317.9537, 318.85, 319.7536, 320.6643, 321.5821, 322.5069, 
    323.4386, 324.3771, 325.3222, 326.2738, 327.2319, 328.1961, 329.1664, 
    330.1425, 331.1244, 332.1117, 333.1042, 334.1017, 335.1041, 336.1109, 
    337.122, 338.1371, 339.1559, 340.1782, 341.2035, 342.2317, 343.2624, 
    344.2952, 345.3299, 346.3661, 347.4035, 348.4418, 349.4805, 350.5195, 
    351.5582, 352.5965, 353.6339, 354.6701, 355.7048, 356.7376, 357.7683, 
    358.7965, 359.8218, 0.8440565, 1.862868, 2.87797, 3.889082, 4.895932, 
    5.898258, 6.895808, 7.888342, 8.875629, 9.857454, 10.83361, 11.8039, 
    12.76814, 13.72616, 14.67781, 15.62294, 16.56141, 17.4931, 18.41789, 
    19.3357, 20.24642, 21.14999, 22.04634, 22.93541, 23.81715, 24.69153, 
    25.55853, 26.41812, 27.27029, 28.11506, 28.95242, 29.78239, 30.60499, 
    31.42026, 32.22822, 33.02893, 33.82243, 34.60877,
  305.3912, 306.1776, 306.971, 307.7718, 308.5797, 309.395, 310.2176, 
    311.0476, 311.8849, 312.7297, 313.5819, 314.4415, 315.3084, 316.1828, 
    317.0646, 317.9536, 318.85, 319.7536, 320.6643, 321.5821, 322.5069, 
    323.4386, 324.377, 325.3222, 326.2738, 327.2318, 328.1961, 329.1664, 
    330.1425, 331.1244, 332.1116, 333.1042, 334.1017, 335.1041, 336.1109, 
    337.122, 338.1371, 339.1559, 340.1782, 341.2035, 342.2317, 343.2623, 
    344.2952, 345.3299, 346.3661, 347.4035, 348.4418, 349.4805, 350.5195, 
    351.5582, 352.5965, 353.6339, 354.6701, 355.7048, 356.7377, 357.7683, 
    358.7965, 359.8218, 0.8440659, 1.862878, 2.877981, 3.889094, 4.895945, 
    5.898271, 6.895822, 7.888356, 8.875645, 9.85747, 10.83362, 11.80391, 
    12.76816, 13.72618, 14.67783, 15.62296, 16.56142, 17.49311, 18.41791, 
    19.33571, 20.24644, 21.15001, 22.04636, 22.93543, 23.81717, 24.69155, 
    25.55855, 26.41814, 27.27031, 28.11508, 28.95244, 29.7824, 30.60501, 
    31.42027, 32.22824, 33.02895, 33.82244, 34.60879,
  305.3912, 306.1776, 306.971, 307.7717, 308.5797, 309.395, 310.2176, 
    311.0475, 311.8849, 312.7297, 313.5818, 314.4414, 315.3084, 316.1828, 
    317.0645, 317.9536, 318.85, 319.7535, 320.6643, 321.5821, 322.5069, 
    323.4386, 324.377, 325.3221, 326.2738, 327.2318, 328.1961, 329.1664, 
    330.1425, 331.1243, 332.1116, 333.1042, 334.1017, 335.104, 336.1109, 
    337.122, 338.1371, 339.1559, 340.1782, 341.2035, 342.2317, 343.2623, 
    344.2952, 345.3299, 346.3661, 347.4035, 348.4418, 349.4805, 350.5195, 
    351.5582, 352.5965, 353.6339, 354.6701, 355.7048, 356.7377, 357.7683, 
    358.7965, 359.8218, 0.8440756, 1.862888, 2.877992, 3.889106, 4.895957, 
    5.898284, 6.895835, 7.888371, 8.87566, 9.857485, 10.83364, 11.80393, 
    12.76817, 13.7262, 14.67785, 15.62297, 16.56144, 17.49313, 18.41793, 
    19.33573, 20.24646, 21.15003, 22.04638, 22.93545, 23.81719, 24.69157, 
    25.55857, 26.41816, 27.27033, 28.1151, 28.95246, 29.78242, 30.60503, 
    31.42029, 32.22826, 33.02896, 33.82246, 34.60881,
  305.3912, 306.1775, 306.971, 307.7717, 308.5797, 309.395, 310.2176, 
    311.0475, 311.8849, 312.7296, 313.5818, 314.4414, 315.3084, 316.1828, 
    317.0645, 317.9536, 318.8499, 319.7535, 320.6642, 321.5821, 322.5068, 
    323.4385, 324.377, 325.3221, 326.2738, 327.2318, 328.196, 329.1664, 
    330.1425, 331.1243, 332.1116, 333.1042, 334.1017, 335.104, 336.1109, 
    337.122, 338.1371, 339.1559, 340.1782, 341.2035, 342.2317, 343.2623, 
    344.2952, 345.3299, 346.3661, 347.4035, 348.4417, 349.4805, 350.5195, 
    351.5583, 352.5965, 353.6339, 354.6701, 355.7048, 356.7377, 357.7683, 
    358.7965, 359.8218, 0.8440856, 1.862899, 2.878004, 3.889118, 4.89597, 
    5.898298, 6.89585, 7.888386, 8.875675, 9.857501, 10.83366, 11.80395, 
    12.76819, 13.72622, 14.67787, 15.62299, 16.56146, 17.49315, 18.41795, 
    19.33575, 20.24648, 21.15005, 22.0464, 22.93546, 23.81721, 24.69159, 
    25.55859, 26.41818, 27.27035, 28.11512, 28.95247, 29.78244, 30.60505, 
    31.42031, 32.22828, 33.02898, 33.82248, 34.60883,
  305.3911, 306.1775, 306.971, 307.7717, 308.5797, 309.3949, 310.2175, 
    311.0475, 311.8849, 312.7296, 313.5818, 314.4414, 315.3084, 316.1828, 
    317.0645, 317.9536, 318.8499, 319.7535, 320.6642, 321.582, 322.5068, 
    323.4385, 324.377, 325.3221, 326.2738, 327.2318, 328.196, 329.1663, 
    330.1425, 331.1243, 332.1116, 333.1041, 334.1017, 335.104, 336.1109, 
    337.122, 338.1371, 339.1559, 340.1781, 341.2035, 342.2317, 343.2623, 
    344.2952, 345.3299, 346.3661, 347.4035, 348.4417, 349.4805, 350.5195, 
    351.5583, 352.5965, 353.6339, 354.6701, 355.7048, 356.7377, 357.7683, 
    358.7965, 359.8219, 0.8440959, 1.86291, 2.878016, 3.889131, 4.895984, 
    5.898313, 6.895865, 7.888402, 8.875691, 9.857518, 10.83367, 11.80397, 
    12.76821, 13.72624, 14.67789, 15.62301, 16.56148, 17.49317, 18.41797, 
    19.33577, 20.2465, 21.15007, 22.04642, 22.93549, 23.81723, 24.69161, 
    25.55861, 26.4182, 27.27037, 28.11514, 28.9525, 29.78246, 30.60506, 
    31.42033, 32.22829, 33.029, 33.8225, 34.60884,
  305.3911, 306.1775, 306.971, 307.7717, 308.5797, 309.3949, 310.2175, 
    311.0475, 311.8849, 312.7296, 313.5818, 314.4414, 315.3084, 316.1827, 
    317.0645, 317.9536, 318.8499, 319.7535, 320.6642, 321.582, 322.5068, 
    323.4385, 324.377, 325.3221, 326.2737, 327.2318, 328.196, 329.1663, 
    330.1425, 331.1243, 332.1116, 333.1041, 334.1017, 335.104, 336.1109, 
    337.122, 338.1371, 339.1559, 340.1781, 341.2035, 342.2317, 343.2623, 
    344.2952, 345.3299, 346.3661, 347.4035, 348.4417, 349.4805, 350.5195, 
    351.5583, 352.5965, 353.6339, 354.6701, 355.7048, 356.7377, 357.7683, 
    358.7965, 359.8219, 0.8441065, 1.862922, 2.878028, 3.889144, 4.895998, 
    5.898327, 6.89588, 7.888417, 8.875709, 9.857535, 10.83369, 11.80398, 
    12.76823, 13.72626, 14.67791, 15.62303, 16.5615, 17.49319, 18.41799, 
    19.33579, 20.24652, 21.15009, 22.04644, 22.93551, 23.81725, 24.69163, 
    25.55863, 26.41822, 27.2704, 28.11516, 28.95252, 29.78248, 30.60509, 
    31.42035, 32.22832, 33.02902, 33.82252, 34.60886,
  305.3911, 306.1775, 306.9709, 307.7717, 308.5796, 309.3949, 310.2175, 
    311.0475, 311.8848, 312.7296, 313.5818, 314.4413, 315.3083, 316.1827, 
    317.0645, 317.9536, 318.8499, 319.7534, 320.6642, 321.582, 322.5068, 
    323.4385, 324.377, 325.3221, 326.2737, 327.2318, 328.196, 329.1663, 
    330.1425, 331.1243, 332.1116, 333.1041, 334.1017, 335.104, 336.1108, 
    337.1219, 338.1371, 339.1559, 340.1781, 341.2035, 342.2316, 343.2623, 
    344.2952, 345.3299, 346.3661, 347.4035, 348.4417, 349.4805, 350.5195, 
    351.5583, 352.5965, 353.6339, 354.6701, 355.7048, 356.7377, 357.7684, 
    358.7965, 359.8219, 0.8441173, 1.862934, 2.878041, 3.889158, 4.896012, 
    5.898342, 6.895896, 7.888434, 8.875726, 9.857553, 10.83371, 11.804, 
    12.76825, 13.72628, 14.67793, 15.62305, 16.56152, 17.49321, 18.41801, 
    19.33582, 20.24654, 21.15011, 22.04646, 22.93553, 23.81727, 24.69166, 
    25.55865, 26.41824, 27.27042, 28.11518, 28.95254, 29.78251, 30.60511, 
    31.42037, 32.22834, 33.02905, 33.82254, 34.60888,
  305.3911, 306.1774, 306.9709, 307.7716, 308.5796, 309.3949, 310.2175, 
    311.0475, 311.8848, 312.7296, 313.5817, 314.4413, 315.3083, 316.1827, 
    317.0645, 317.9535, 318.8499, 319.7534, 320.6642, 321.582, 322.5068, 
    323.4384, 324.3769, 325.3221, 326.2737, 327.2317, 328.196, 329.1663, 
    330.1424, 331.1243, 332.1115, 333.1041, 334.1017, 335.104, 336.1108, 
    337.1219, 338.1371, 339.1559, 340.1781, 341.2035, 342.2316, 343.2623, 
    344.2951, 345.3298, 346.3661, 347.4035, 348.4417, 349.4805, 350.5195, 
    351.5583, 352.5965, 353.6339, 354.6702, 355.7049, 356.7377, 357.7684, 
    358.7965, 359.8219, 0.8441283, 1.862946, 2.878054, 3.889171, 4.896027, 
    5.898357, 6.895912, 7.888451, 8.875743, 9.857572, 10.83373, 11.80402, 
    12.76827, 13.7263, 14.67795, 15.62307, 16.56154, 17.49323, 18.41803, 
    19.33584, 20.24657, 21.15014, 22.04648, 22.93555, 23.8173, 24.69168, 
    25.55867, 26.41826, 27.27044, 28.1152, 28.95256, 29.78253, 30.60513, 
    31.42039, 32.22836, 33.02906, 33.82256, 34.60891,
  305.3911, 306.1774, 306.9709, 307.7716, 308.5796, 309.3948, 310.2174, 
    311.0474, 311.8848, 312.7295, 313.5817, 314.4413, 315.3083, 316.1827, 
    317.0644, 317.9535, 318.8499, 319.7534, 320.6641, 321.5819, 322.5067, 
    323.4384, 324.3769, 325.322, 326.2737, 327.2317, 328.196, 329.1663, 
    330.1424, 331.1242, 332.1115, 333.1041, 334.1016, 335.104, 336.1108, 
    337.1219, 338.1371, 339.1559, 340.1781, 341.2035, 342.2316, 343.2623, 
    344.2951, 345.3298, 346.3661, 347.4035, 348.4417, 349.4805, 350.5195, 
    351.5583, 352.5965, 353.6339, 354.6702, 355.7049, 356.7377, 357.7684, 
    358.7965, 359.8219, 0.8441395, 1.862958, 2.878067, 3.889185, 4.896041, 
    5.898373, 6.895928, 7.888468, 8.875761, 9.85759, 10.83375, 11.80404, 
    12.76829, 13.72632, 14.67797, 15.6231, 16.56157, 17.49326, 18.41805, 
    19.33586, 20.24659, 21.15016, 22.04651, 22.93558, 23.81732, 24.6917, 
    25.5587, 26.41829, 27.27046, 28.11522, 28.95258, 29.78255, 30.60515, 
    31.42042, 32.22838, 33.02909, 33.82259, 34.60892,
  305.3911, 306.1774, 306.9709, 307.7716, 308.5796, 309.3948, 310.2174, 
    311.0474, 311.8847, 312.7295, 313.5817, 314.4413, 315.3083, 316.1826, 
    317.0644, 317.9535, 318.8498, 319.7534, 320.6641, 321.5819, 322.5067, 
    323.4384, 324.3769, 325.322, 326.2737, 327.2317, 328.1959, 329.1662, 
    330.1424, 331.1242, 332.1115, 333.1041, 334.1016, 335.1039, 336.1108, 
    337.1219, 338.137, 339.1559, 340.1781, 341.2034, 342.2316, 343.2623, 
    344.2951, 345.3298, 346.3661, 347.4035, 348.4417, 349.4805, 350.5195, 
    351.5583, 352.5965, 353.6339, 354.6702, 355.7049, 356.7377, 357.7684, 
    358.7966, 359.8219, 0.8441509, 1.86297, 2.87808, 3.889199, 4.896057, 
    5.898389, 6.895945, 7.888485, 8.875779, 9.857609, 10.83377, 11.80406, 
    12.76831, 13.72634, 14.67799, 15.62312, 16.56159, 17.49328, 18.41808, 
    19.33588, 20.24661, 21.15018, 22.04653, 22.9356, 23.81734, 24.69172, 
    25.55872, 26.41831, 27.27049, 28.11525, 28.95261, 29.78258, 30.60518, 
    31.42044, 32.2284, 33.02911, 33.82261, 34.60895,
  305.391, 306.1774, 306.9709, 307.7716, 308.5795, 309.3948, 310.2174, 
    311.0474, 311.8847, 312.7295, 313.5817, 314.4413, 315.3083, 316.1826, 
    317.0644, 317.9534, 318.8498, 319.7534, 320.6641, 321.5819, 322.5067, 
    323.4384, 324.3769, 325.322, 326.2737, 327.2317, 328.1959, 329.1662, 
    330.1424, 331.1242, 332.1115, 333.104, 334.1016, 335.1039, 336.1108, 
    337.1219, 338.137, 339.1558, 340.1781, 341.2034, 342.2316, 343.2623, 
    344.2951, 345.3298, 346.3661, 347.4035, 348.4417, 349.4805, 350.5195, 
    351.5583, 352.5965, 353.6339, 354.6702, 355.7049, 356.7377, 357.7684, 
    358.7966, 359.8219, 0.8441625, 1.862983, 2.878093, 3.889214, 4.896072, 
    5.898405, 6.895962, 7.888503, 8.875797, 9.857628, 10.83379, 11.80408, 
    12.76833, 13.72636, 14.67801, 15.62314, 16.56161, 17.4933, 18.4181, 
    19.33591, 20.24664, 21.15021, 22.04656, 22.93563, 23.81737, 24.69175, 
    25.55874, 26.41833, 27.27051, 28.11527, 28.95263, 29.7826, 30.6052, 
    31.42046, 32.22843, 33.02913, 33.82263, 34.60897,
  305.391, 306.1773, 306.9709, 307.7715, 308.5795, 309.3948, 310.2174, 
    311.0473, 311.8847, 312.7295, 313.5816, 314.4412, 315.3082, 316.1826, 
    317.0644, 317.9534, 318.8498, 319.7533, 320.6641, 321.5819, 322.5067, 
    323.4384, 324.3768, 325.322, 326.2736, 327.2317, 328.1959, 329.1662, 
    330.1424, 331.1242, 332.1115, 333.104, 334.1016, 335.1039, 336.1108, 
    337.1219, 338.137, 339.1558, 340.1781, 341.2034, 342.2316, 343.2623, 
    344.2951, 345.3298, 346.3661, 347.4035, 348.4417, 349.4805, 350.5195, 
    351.5583, 352.5965, 353.6339, 354.6702, 355.7049, 356.7377, 357.7684, 
    358.7966, 359.8219, 0.8441741, 1.862995, 2.878107, 3.889229, 4.896087, 
    5.898421, 6.895979, 7.888521, 8.875816, 9.857647, 10.83381, 11.8041, 
    12.76835, 13.72638, 14.67803, 15.62316, 16.56163, 17.49333, 18.41813, 
    19.33593, 20.24666, 21.15023, 22.04658, 22.93565, 23.81739, 24.69177, 
    25.55877, 26.41836, 27.27054, 28.1153, 28.95266, 29.78262, 30.60522, 
    31.42049, 32.22845, 33.02916, 33.82265, 34.609,
  305.391, 306.1773, 306.9708, 307.7715, 308.5795, 309.3947, 310.2173, 
    311.0473, 311.8847, 312.7294, 313.5816, 314.4412, 315.3082, 316.1826, 
    317.0643, 317.9534, 318.8497, 319.7533, 320.664, 321.5818, 322.5067, 
    323.4384, 324.3768, 325.3219, 326.2736, 327.2316, 328.1959, 329.1662, 
    330.1423, 331.1242, 332.1115, 333.104, 334.1016, 335.1039, 336.1107, 
    337.1219, 338.137, 339.1558, 340.1781, 341.2034, 342.2316, 343.2623, 
    344.2951, 345.3298, 346.3661, 347.4035, 348.4417, 349.4805, 350.5195, 
    351.5583, 352.5965, 353.6339, 354.6702, 355.7049, 356.7377, 357.7684, 
    358.7966, 359.8219, 0.844186, 1.863008, 2.878121, 3.889243, 4.896103, 
    5.898438, 6.895997, 7.888539, 8.875834, 9.857667, 10.83383, 11.80412, 
    12.76837, 13.7264, 14.67806, 15.62319, 16.56166, 17.49335, 18.41815, 
    19.33596, 20.24669, 21.15026, 22.04661, 22.93567, 23.81742, 24.6918, 
    25.5588, 26.41838, 27.27056, 28.11532, 28.95268, 29.78265, 30.60525, 
    31.42051, 32.22848, 33.02918, 33.82268, 34.60902,
  305.391, 306.1773, 306.9708, 307.7715, 308.5795, 309.3947, 310.2173, 
    311.0473, 311.8846, 312.7294, 313.5816, 314.4412, 315.3082, 316.1826, 
    317.0643, 317.9534, 318.8497, 319.7533, 320.664, 321.5818, 322.5066, 
    323.4383, 324.3768, 325.3219, 326.2736, 327.2316, 328.1959, 329.1661, 
    330.1423, 331.1241, 332.1115, 333.104, 334.1015, 335.1039, 336.1107, 
    337.1219, 338.137, 339.1558, 340.178, 341.2034, 342.2316, 343.2623, 
    344.2951, 345.3298, 346.3661, 347.4035, 348.4417, 349.4805, 350.5195, 
    351.5583, 352.5965, 353.6339, 354.6702, 355.7049, 356.7377, 357.7684, 
    358.7966, 359.822, 0.844198, 1.863021, 2.878135, 3.889258, 4.896119, 
    5.898455, 6.896014, 7.888557, 8.875854, 9.857687, 10.83385, 11.80414, 
    12.76839, 13.72643, 14.67808, 15.62321, 16.56168, 17.49337, 18.41817, 
    19.33598, 20.24671, 21.15028, 22.04663, 22.9357, 23.81744, 24.69183, 
    25.55882, 26.41841, 27.27059, 28.11535, 28.95271, 29.78267, 30.60528, 
    31.42054, 32.2285, 33.02921, 33.8227, 34.60905,
  305.3909, 306.1773, 306.9708, 307.7715, 308.5794, 309.3947, 310.2173, 
    311.0473, 311.8846, 312.7294, 313.5816, 314.4412, 315.3081, 316.1825, 
    317.0643, 317.9533, 318.8497, 319.7533, 320.664, 321.5818, 322.5066, 
    323.4383, 324.3768, 325.3219, 326.2736, 327.2316, 328.1958, 329.1661, 
    330.1423, 331.1241, 332.1114, 333.104, 334.1015, 335.1039, 336.1107, 
    337.1219, 338.137, 339.1558, 340.178, 341.2034, 342.2316, 343.2622, 
    344.2951, 345.3298, 346.3661, 347.4035, 348.4417, 349.4805, 350.5195, 
    351.5583, 352.5965, 353.6339, 354.6702, 355.7049, 356.7378, 357.7684, 
    358.7966, 359.822, 0.84421, 1.863034, 2.878149, 3.889273, 4.896135, 
    5.898471, 6.896032, 7.888576, 8.875874, 9.857707, 10.83387, 11.80417, 
    12.76842, 13.72645, 14.6781, 15.62323, 16.56171, 17.4934, 18.4182, 
    19.33601, 20.24674, 21.15031, 22.04666, 22.93573, 23.81747, 24.69185, 
    25.55885, 26.41844, 27.27061, 28.11538, 28.95273, 29.7827, 30.6053, 
    31.42057, 32.22853, 33.02924, 33.82273, 34.60907,
  305.3909, 306.1772, 306.9707, 307.7715, 308.5794, 309.3947, 310.2173, 
    311.0472, 311.8846, 312.7294, 313.5815, 314.4411, 315.3081, 316.1825, 
    317.0642, 317.9533, 318.8497, 319.7532, 320.664, 321.5818, 322.5066, 
    323.4383, 324.3767, 325.3219, 326.2735, 327.2316, 328.1958, 329.1661, 
    330.1423, 331.1241, 332.1114, 333.1039, 334.1015, 335.1039, 336.1107, 
    337.1218, 338.137, 339.1558, 340.178, 341.2034, 342.2316, 343.2622, 
    344.2951, 345.3298, 346.366, 347.4035, 348.4417, 349.4805, 350.5195, 
    351.5583, 352.5965, 353.634, 354.6702, 355.7049, 356.7378, 357.7684, 
    358.7966, 359.822, 0.8442221, 1.863047, 2.878163, 3.889288, 4.896151, 
    5.898489, 6.89605, 7.888595, 8.875893, 9.857727, 10.83389, 11.80419, 
    12.76844, 13.72647, 14.67813, 15.62326, 16.56173, 17.49342, 18.41822, 
    19.33603, 20.24676, 21.15034, 22.04668, 22.93575, 23.8175, 24.69188, 
    25.55888, 26.41846, 27.27064, 28.1154, 28.95276, 29.78273, 30.60533, 
    31.42059, 32.22855, 33.02926, 33.82276, 34.6091,
  305.3909, 306.1772, 306.9707, 307.7714, 308.5794, 309.3947, 310.2173, 
    311.0472, 311.8846, 312.7293, 313.5815, 314.4411, 315.3081, 316.1825, 
    317.0642, 317.9533, 318.8496, 319.7532, 320.6639, 321.5818, 322.5066, 
    323.4382, 324.3767, 325.3218, 326.2735, 327.2315, 328.1958, 329.1661, 
    330.1422, 331.1241, 332.1114, 333.1039, 334.1015, 335.1038, 336.1107, 
    337.1218, 338.1369, 339.1558, 340.178, 341.2034, 342.2316, 343.2622, 
    344.2951, 345.3298, 346.366, 347.4035, 348.4417, 349.4805, 350.5195, 
    351.5583, 352.5965, 353.634, 354.6702, 355.7049, 356.7378, 357.7684, 
    358.7966, 359.822, 0.8442343, 1.863061, 2.878178, 3.889304, 4.896167, 
    5.898506, 6.896068, 7.888614, 8.875913, 9.857747, 10.83391, 11.80421, 
    12.76846, 13.72649, 14.67815, 15.62328, 16.56175, 17.49345, 18.41825, 
    19.33606, 20.24679, 21.15036, 22.04671, 22.93578, 23.81752, 24.69191, 
    25.5589, 26.41849, 27.27067, 28.11543, 28.95279, 29.78276, 30.60536, 
    31.42062, 32.22858, 33.02929, 33.82278, 34.60912,
  305.3908, 306.1772, 306.9707, 307.7714, 308.5793, 309.3946, 310.2172, 
    311.0472, 311.8846, 312.7293, 313.5815, 314.4411, 315.3081, 316.1824, 
    317.0642, 317.9532, 318.8496, 319.7532, 320.6639, 321.5817, 322.5065, 
    323.4382, 324.3767, 325.3218, 326.2735, 327.2315, 328.1958, 329.1661, 
    330.1422, 331.1241, 332.1114, 333.1039, 334.1015, 335.1038, 336.1107, 
    337.1218, 338.1369, 339.1558, 340.178, 341.2034, 342.2315, 343.2622, 
    344.2951, 345.3298, 346.366, 347.4034, 348.4417, 349.4805, 350.5195, 
    351.5583, 352.5966, 353.634, 354.6702, 355.7049, 356.7378, 357.7685, 
    358.7966, 359.822, 0.8442466, 1.863074, 2.878192, 3.889319, 4.896183, 
    5.898523, 6.896086, 7.888632, 8.875933, 9.857768, 10.83393, 11.80423, 
    12.76848, 13.72652, 14.67817, 15.62331, 16.56178, 17.49347, 18.41828, 
    19.33608, 20.24681, 21.15039, 22.04674, 22.93581, 23.81755, 24.69193, 
    25.55893, 26.41852, 27.2707, 28.11546, 28.95282, 29.78278, 30.60538, 
    31.42065, 32.22861, 33.02932, 33.82281, 34.60915,
  305.3908, 306.1772, 306.9706, 307.7714, 308.5793, 309.3946, 310.2172, 
    311.0471, 311.8845, 312.7293, 313.5815, 314.441, 315.308, 316.1824, 
    317.0642, 317.9532, 318.8496, 319.7531, 320.6639, 321.5817, 322.5065, 
    323.4382, 324.3767, 325.3218, 326.2735, 327.2315, 328.1957, 329.166, 
    330.1422, 331.1241, 332.1114, 333.1039, 334.1015, 335.1038, 336.1107, 
    337.1218, 338.1369, 339.1557, 340.178, 341.2034, 342.2315, 343.2622, 
    344.2951, 345.3298, 346.366, 347.4034, 348.4417, 349.4805, 350.5195, 
    351.5583, 352.5966, 353.634, 354.6702, 355.7049, 356.7378, 357.7685, 
    358.7966, 359.822, 0.8442588, 1.863087, 2.878206, 3.889334, 4.8962, 
    5.89854, 6.896104, 7.888651, 8.875953, 9.857789, 10.83395, 11.80425, 
    12.76851, 13.72654, 14.6782, 15.62333, 16.56181, 17.4935, 18.4183, 
    19.33611, 20.24684, 21.15042, 22.04676, 22.93583, 23.81758, 24.69196, 
    25.55896, 26.41855, 27.27073, 28.11549, 28.95284, 29.78281, 30.60541, 
    31.42068, 32.22864, 33.02934, 33.82284, 34.60918,
  305.3908, 306.1771, 306.9706, 307.7713, 308.5793, 309.3946, 310.2172, 
    311.0471, 311.8845, 312.7292, 313.5814, 314.441, 315.308, 316.1824, 
    317.0641, 317.9532, 318.8495, 319.7531, 320.6638, 321.5817, 322.5065, 
    323.4382, 324.3766, 325.3218, 326.2734, 327.2315, 328.1957, 329.166, 
    330.1422, 331.124, 332.1113, 333.1039, 334.1014, 335.1038, 336.1107, 
    337.1218, 338.1369, 339.1557, 340.178, 341.2033, 342.2315, 343.2622, 
    344.2951, 345.3298, 346.366, 347.4034, 348.4417, 349.4805, 350.5195, 
    351.5583, 352.5966, 353.634, 354.6702, 355.7049, 356.7378, 357.7685, 
    358.7967, 359.822, 0.8442712, 1.863101, 2.878221, 3.88935, 4.896216, 
    5.898557, 6.896122, 7.88867, 8.875972, 9.857809, 10.83398, 11.80428, 
    12.76853, 13.72656, 14.67822, 15.62335, 16.56183, 17.49352, 18.41833, 
    19.33614, 20.24687, 21.15044, 22.04679, 22.93586, 23.81761, 24.69199, 
    25.55899, 26.41858, 27.27075, 28.11552, 28.95288, 29.78284, 30.60544, 
    31.4207, 32.22867, 33.02937, 33.82287, 34.60921,
  305.3908, 306.1771, 306.9706, 307.7713, 308.5793, 309.3945, 310.2171, 
    311.0471, 311.8845, 312.7292, 313.5814, 314.441, 315.308, 316.1824, 
    317.0641, 317.9532, 318.8495, 319.7531, 320.6638, 321.5816, 322.5064, 
    323.4381, 324.3766, 325.3217, 326.2734, 327.2314, 328.1957, 329.166, 
    330.1422, 331.124, 332.1113, 333.1039, 334.1014, 335.1038, 336.1106, 
    337.1218, 338.1369, 339.1557, 340.178, 341.2033, 342.2315, 343.2622, 
    344.2951, 345.3298, 346.366, 347.4034, 348.4417, 349.4805, 350.5195, 
    351.5583, 352.5966, 353.634, 354.6702, 355.7049, 356.7378, 357.7685, 
    358.7967, 359.822, 0.8442835, 1.863114, 2.878235, 3.889365, 4.896233, 
    5.898575, 6.896141, 7.88869, 8.875992, 9.85783, 10.834, 11.8043, 
    12.76855, 13.72659, 14.67825, 15.62338, 16.56186, 17.49355, 18.41835, 
    19.33616, 20.2469, 21.15047, 22.04682, 22.93589, 23.81764, 24.69202, 
    25.55902, 26.41861, 27.27078, 28.11555, 28.9529, 29.78287, 30.60547, 
    31.42073, 32.22869, 33.0294, 33.8229, 34.60923,
  305.3907, 306.1771, 306.9706, 307.7713, 308.5792, 309.3945, 310.2171, 
    311.0471, 311.8844, 312.7292, 313.5814, 314.4409, 315.308, 316.1823, 
    317.0641, 317.9532, 318.8495, 319.7531, 320.6638, 321.5816, 322.5064, 
    323.4381, 324.3766, 325.3217, 326.2734, 327.2314, 328.1957, 329.166, 
    330.1422, 331.124, 332.1113, 333.1039, 334.1014, 335.1038, 336.1106, 
    337.1218, 338.1369, 339.1557, 340.1779, 341.2033, 342.2315, 343.2622, 
    344.295, 345.3298, 346.366, 347.4034, 348.4417, 349.4805, 350.5195, 
    351.5583, 352.5966, 353.634, 354.6702, 355.705, 356.7378, 357.7685, 
    358.7967, 359.8221, 0.8442957, 1.863127, 2.878249, 3.889381, 4.896249, 
    5.898592, 6.896159, 7.888709, 8.876012, 9.857851, 10.83402, 11.80432, 
    12.76858, 13.72661, 14.67827, 15.6234, 16.56188, 17.49358, 18.41838, 
    19.33619, 20.24692, 21.1505, 22.04685, 22.93592, 23.81767, 24.69205, 
    25.55904, 26.41864, 27.27081, 28.11558, 28.95293, 29.7829, 30.6055, 
    31.42076, 32.22873, 33.02943, 33.82293, 34.60926,
  305.3907, 306.177, 306.9706, 307.7712, 308.5792, 309.3945, 310.2171, 
    311.047, 311.8844, 312.7292, 313.5813, 314.4409, 315.3079, 316.1823, 
    317.0641, 317.9531, 318.8495, 319.7531, 320.6638, 321.5816, 322.5064, 
    323.4381, 324.3766, 325.3217, 326.2734, 327.2314, 328.1956, 329.166, 
    330.1421, 331.124, 332.1113, 333.1038, 334.1014, 335.1037, 336.1106, 
    337.1217, 338.1369, 339.1557, 340.1779, 341.2033, 342.2315, 343.2622, 
    344.295, 345.3298, 346.366, 347.4034, 348.4417, 349.4805, 350.5195, 
    351.5583, 352.5966, 353.634, 354.6702, 355.705, 356.7378, 357.7685, 
    358.7967, 359.8221, 0.844308, 1.863141, 2.878264, 3.889396, 4.896265, 
    5.89861, 6.896177, 7.888728, 8.876032, 9.857872, 10.83404, 11.80434, 
    12.7686, 13.72663, 14.67829, 15.62343, 16.56191, 17.4936, 18.41841, 
    19.33622, 20.24695, 21.15053, 22.04688, 22.93595, 23.81769, 24.69208, 
    25.55907, 26.41866, 27.27084, 28.1156, 28.95296, 29.78293, 30.60553, 
    31.42079, 32.22876, 33.02946, 33.82296, 34.60929,
  305.3907, 306.177, 306.9705, 307.7712, 308.5792, 309.3944, 310.217, 
    311.047, 311.8844, 312.7291, 313.5813, 314.4409, 315.3079, 316.1823, 
    317.064, 317.9531, 318.8495, 319.753, 320.6638, 321.5816, 322.5064, 
    323.4381, 324.3766, 325.3217, 326.2733, 327.2314, 328.1956, 329.1659, 
    330.1421, 331.124, 332.1113, 333.1038, 334.1014, 335.1037, 336.1106, 
    337.1217, 338.1368, 339.1557, 340.1779, 341.2033, 342.2315, 343.2622, 
    344.295, 345.3298, 346.366, 347.4034, 348.4417, 349.4805, 350.5195, 
    351.5583, 352.5966, 353.634, 354.6702, 355.705, 356.7378, 357.7685, 
    358.7967, 359.8221, 0.8443203, 1.863154, 2.878278, 3.889411, 4.896282, 
    5.898627, 6.896195, 7.888747, 8.876052, 9.857893, 10.83406, 11.80437, 
    12.76862, 13.72666, 14.67832, 15.62346, 16.56193, 17.49363, 18.41843, 
    19.33625, 20.24698, 21.15055, 22.04691, 22.93598, 23.81772, 24.69211, 
    25.5591, 26.4187, 27.27087, 28.11563, 28.95299, 29.78296, 30.60556, 
    31.42082, 32.22879, 33.02949, 33.82298, 34.60933,
  305.3907, 306.177, 306.9705, 307.7712, 308.5791, 309.3944, 310.217, 
    311.047, 311.8843, 312.7291, 313.5813, 314.4409, 315.3079, 316.1823, 
    317.064, 317.9531, 318.8494, 319.753, 320.6637, 321.5815, 322.5063, 
    323.438, 324.3765, 325.3217, 326.2733, 327.2314, 328.1956, 329.1659, 
    330.1421, 331.1239, 332.1112, 333.1038, 334.1013, 335.1037, 336.1106, 
    337.1217, 338.1368, 339.1557, 340.1779, 341.2033, 342.2315, 343.2622, 
    344.295, 345.3297, 346.366, 347.4034, 348.4417, 349.4805, 350.5195, 
    351.5583, 352.5966, 353.634, 354.6703, 355.705, 356.7378, 357.7685, 
    358.7967, 359.8221, 0.8443325, 1.863167, 2.878293, 3.889427, 4.896298, 
    5.898644, 6.896214, 7.888766, 8.876072, 9.857914, 10.83408, 11.80439, 
    12.76865, 13.72668, 14.67834, 15.62348, 16.56196, 17.49366, 18.41846, 
    19.33627, 20.24701, 21.15058, 22.04693, 22.93601, 23.81775, 24.69214, 
    25.55913, 26.41872, 27.2709, 28.11567, 28.95302, 29.78299, 30.60559, 
    31.42085, 32.22882, 33.02952, 33.82301, 34.60936,
  305.3906, 306.1769, 306.9705, 307.7711, 308.5791, 309.3944, 310.217, 
    311.0469, 311.8843, 312.7291, 313.5812, 314.4408, 315.3078, 316.1822, 
    317.064, 317.953, 318.8494, 319.753, 320.6637, 321.5815, 322.5063, 
    323.438, 324.3765, 325.3216, 326.2733, 327.2313, 328.1956, 329.1659, 
    330.1421, 331.1239, 332.1112, 333.1038, 334.1013, 335.1037, 336.1106, 
    337.1217, 338.1368, 339.1557, 340.1779, 341.2033, 342.2315, 343.2622, 
    344.295, 345.3297, 346.366, 347.4034, 348.4417, 349.4805, 350.5195, 
    351.5583, 352.5966, 353.634, 354.6703, 355.705, 356.7378, 357.7685, 
    358.7967, 359.8221, 0.8443446, 1.863181, 2.878307, 3.889442, 4.896314, 
    5.898661, 6.896232, 7.888785, 8.876092, 9.857934, 10.83411, 11.80441, 
    12.76867, 13.72671, 14.67837, 15.62351, 16.56199, 17.49368, 18.41849, 
    19.3363, 20.24703, 21.15061, 22.04696, 22.93604, 23.81778, 24.69217, 
    25.55916, 26.41875, 27.27093, 28.1157, 28.95305, 29.78302, 30.60562, 
    31.42089, 32.22885, 33.02955, 33.82305, 34.60939,
  305.3906, 306.1769, 306.9704, 307.7711, 308.5791, 309.3943, 310.2169, 
    311.0469, 311.8843, 312.729, 313.5812, 314.4408, 315.3078, 316.1822, 
    317.0639, 317.953, 318.8494, 319.7529, 320.6637, 321.5815, 322.5063, 
    323.438, 324.3765, 325.3216, 326.2733, 327.2313, 328.1956, 329.1659, 
    330.1421, 331.1239, 332.1112, 333.1038, 334.1013, 335.1037, 336.1105, 
    337.1217, 338.1368, 339.1556, 340.1779, 341.2033, 342.2315, 343.2621, 
    344.295, 345.3297, 346.366, 347.4034, 348.4417, 349.4805, 350.5195, 
    351.5583, 352.5966, 353.634, 354.6703, 355.705, 356.7379, 357.7685, 
    358.7967, 359.8221, 0.8443567, 1.863194, 2.878321, 3.889457, 4.89633, 
    5.898679, 6.89625, 7.888804, 8.876112, 9.857955, 10.83413, 11.80443, 
    12.76869, 13.72673, 14.67839, 15.62353, 16.56201, 17.49371, 18.41851, 
    19.33633, 20.24706, 21.15064, 22.04699, 22.93606, 23.81781, 24.6922, 
    25.55919, 26.41879, 27.27096, 28.11573, 28.95308, 29.78305, 30.60565, 
    31.42092, 32.22888, 33.02958, 33.82308, 34.60942,
  305.3906, 306.1769, 306.9704, 307.7711, 308.579, 309.3943, 310.2169, 
    311.0469, 311.8842, 312.729, 313.5812, 314.4408, 315.3078, 316.1822, 
    317.0639, 317.953, 318.8493, 319.7529, 320.6636, 321.5815, 322.5063, 
    323.438, 324.3764, 325.3216, 326.2733, 327.2313, 328.1956, 329.1659, 
    330.142, 331.1239, 332.1112, 333.1037, 334.1013, 335.1037, 336.1105, 
    337.1217, 338.1368, 339.1556, 340.1779, 341.2033, 342.2314, 343.2621, 
    344.295, 345.3297, 346.366, 347.4034, 348.4417, 349.4805, 350.5195, 
    351.5583, 352.5966, 353.634, 354.6703, 355.705, 356.7379, 357.7686, 
    358.7967, 359.8221, 0.8443687, 1.863207, 2.878335, 3.889472, 4.896347, 
    5.898695, 6.896268, 7.888824, 8.876132, 9.857976, 10.83415, 11.80446, 
    12.76871, 13.72675, 14.67842, 15.62356, 16.56204, 17.49373, 18.41854, 
    19.33636, 20.24709, 21.15067, 22.04702, 22.93609, 23.81784, 24.69223, 
    25.55922, 26.41882, 27.27099, 28.11576, 28.95312, 29.78308, 30.60568, 
    31.42095, 32.22891, 33.02961, 33.82311, 34.60945,
  305.3905, 306.1768, 306.9704, 307.7711, 308.579, 309.3943, 310.2169, 
    311.0468, 311.8842, 312.729, 313.5811, 314.4407, 315.3077, 316.1821, 
    317.0639, 317.9529, 318.8493, 319.7529, 320.6636, 321.5814, 322.5062, 
    323.4379, 324.3764, 325.3216, 326.2732, 327.2313, 328.1955, 329.1658, 
    330.142, 331.1238, 332.1111, 333.1037, 334.1013, 335.1036, 336.1105, 
    337.1216, 338.1368, 339.1556, 340.1779, 341.2032, 342.2314, 343.2621, 
    344.295, 345.3297, 346.366, 347.4034, 348.4417, 349.4805, 350.5195, 
    351.5583, 352.5966, 353.634, 354.6703, 355.705, 356.7379, 357.7686, 
    358.7968, 359.8221, 0.8443806, 1.86322, 2.878349, 3.889488, 4.896363, 
    5.898713, 6.896286, 7.888842, 8.876152, 9.857996, 10.83417, 11.80448, 
    12.76874, 13.72678, 14.67844, 15.62358, 16.56206, 17.49376, 18.41857, 
    19.33638, 20.24712, 21.1507, 22.04705, 22.93612, 23.81787, 24.69226, 
    25.55925, 26.41885, 27.27102, 28.11579, 28.95315, 29.78312, 30.60571, 
    31.42098, 32.22894, 33.02964, 33.82314, 34.60948 ;

 grid_latt =
  -35.07925, -35.43988, -35.79544, -36.14578, -36.4908, -36.83038, -37.1644, 
    -37.49273, -37.81525, -38.13184, -38.44237, -38.74672, -39.04476, 
    -39.33637, -39.62142, -39.89979, -40.17135, -40.43598, -40.69355, 
    -40.94394, -41.18702, -41.42268, -41.65079, -41.87124, -42.08391, 
    -42.28868, -42.48545, -42.67411, -42.85454, -43.02665, -43.19033, 
    -43.34549, -43.49203, -43.62987, -43.75893, -43.87911, -43.99035, 
    -44.09258, -44.18572, -44.26973, -44.34454, -44.41011, -44.46639, 
    -44.51335, -44.55096, -44.57919, -44.59801, -44.60743, -44.60743, 
    -44.59801, -44.57919, -44.55096, -44.51335, -44.46639, -44.41011, 
    -44.34454, -44.26973, -44.18572, -44.09258, -43.99035, -43.87911, 
    -43.75893, -43.62987, -43.49203, -43.34549, -43.19033, -43.02665, 
    -42.85454, -42.67411, -42.48545, -42.28868, -42.08391, -41.87124, 
    -41.65079, -41.42268, -41.18702, -40.94394, -40.69355, -40.43598, 
    -40.17135, -39.89979, -39.62142, -39.33637, -39.04476, -38.74672, 
    -38.44237, -38.13184, -37.81525, -37.49273, -37.1644, -36.83038, 
    -36.4908, -36.14578, -35.79544, -35.43988, -35.07925,
  -34.34282, -34.70005, -35.05236, -35.39962, -35.7417, -36.0785, -36.40988, 
    -36.73572, -37.05589, -37.37026, -37.67871, -37.9811, -38.27731, 
    -38.56721, -38.85067, -39.12755, -39.39772, -39.66107, -39.91746, 
    -40.16676, -40.40884, -40.64358, -40.87085, -41.09053, -41.30251, 
    -41.50666, -41.70287, -41.89101, -42.07099, -42.24269, -42.40602, 
    -42.56086, -42.70713, -42.84472, -42.97356, -43.09357, -43.20465, 
    -43.30674, -43.39978, -43.48369, -43.55843, -43.62393, -43.68016, 
    -43.72708, -43.76466, -43.79286, -43.81168, -43.82109, -43.82109, 
    -43.81168, -43.79286, -43.76466, -43.72708, -43.68016, -43.62393, 
    -43.55843, -43.48369, -43.39978, -43.30674, -43.20465, -43.09357, 
    -42.97356, -42.84472, -42.70713, -42.56086, -42.40602, -42.24269, 
    -42.07099, -41.89101, -41.70287, -41.50666, -41.30251, -41.09053, 
    -40.87085, -40.64358, -40.40884, -40.16676, -39.91746, -39.66107, 
    -39.39772, -39.12755, -38.85067, -38.56721, -38.27731, -37.9811, 
    -37.67871, -37.37026, -37.05589, -36.73572, -36.40988, -36.0785, 
    -35.7417, -35.39962, -35.05236, -34.70005, -34.34282,
  -33.60628, -33.95987, -34.30869, -34.65261, -34.99154, -35.32531, 
    -35.65382, -35.97694, -36.29453, -36.60646, -36.91259, -37.21281, 
    -37.50697, -37.79493, -38.07658, -38.35176, -38.62035, -38.88222, 
    -39.13723, -39.38524, -39.62614, -39.85978, -40.08604, -40.30479, 
    -40.51591, -40.71927, -40.91476, -41.10225, -41.28164, -41.4528, 
    -41.61564, -41.77005, -41.91592, -42.05317, -42.18171, -42.30143, 
    -42.41228, -42.51416, -42.60701, -42.69076, -42.76536, -42.83075, 
    -42.88689, -42.93373, -42.97124, -42.9994, -43.01819, -43.02758, 
    -43.02758, -43.01819, -42.9994, -42.97124, -42.93373, -42.88689, 
    -42.83075, -42.76536, -42.69076, -42.60701, -42.51416, -42.41228, 
    -42.30143, -42.18171, -42.05317, -41.91592, -41.77005, -41.61564, 
    -41.4528, -41.28164, -41.10225, -40.91476, -40.71927, -40.51591, 
    -40.30479, -40.08604, -39.85978, -39.62614, -39.38524, -39.13723, 
    -38.88222, -38.62035, -38.35176, -38.07658, -37.79493, -37.50697, 
    -37.21281, -36.91259, -36.60646, -36.29453, -35.97694, -35.65382, 
    -35.32531, -34.99154, -34.65261, -34.30869, -33.95987, -33.60628,
  -32.86962, -33.21932, -33.56442, -33.90479, -34.2403, -34.57083, -34.89624, 
    -35.2164, -35.53117, -35.84042, -36.14403, -36.44184, -36.73372, 
    -37.01954, -37.29916, -37.57244, -37.83924, -38.09942, -38.35286, 
    -38.5994, -38.83891, -39.07127, -39.29634, -39.51399, -39.72409, 
    -39.9265, -40.12112, -40.30781, -40.48646, -40.65696, -40.81918, 
    -40.97303, -41.1184, -41.25519, -41.38331, -41.50267, -41.61318, 
    -41.71477, -41.80736, -41.89089, -41.96529, -42.03052, -42.08652, 
    -42.13324, -42.17067, -42.19876, -42.2175, -42.22688, -42.22688, 
    -42.2175, -42.19876, -42.17067, -42.13324, -42.08652, -42.03052, 
    -41.96529, -41.89089, -41.80736, -41.71477, -41.61318, -41.50267, 
    -41.38331, -41.25519, -41.1184, -40.97303, -40.81918, -40.65696, 
    -40.48646, -40.30781, -40.12112, -39.9265, -39.72409, -39.51399, 
    -39.29634, -39.07127, -38.83891, -38.5994, -38.35286, -38.09942, 
    -37.83924, -37.57244, -37.29916, -37.01954, -36.73372, -36.44184, 
    -36.14403, -35.84042, -35.53117, -35.2164, -34.89624, -34.57083, 
    -34.2403, -33.90479, -33.56442, -33.21932, -32.86962,
  -32.13284, -32.47842, -32.81957, -33.15614, -33.48802, -33.81506, 
    -34.13713, -34.4541, -34.76583, -35.07218, -35.37302, -35.66821, 
    -35.9576, -36.24105, -36.51843, -36.78959, -37.05439, -37.31269, 
    -37.56434, -37.80922, -38.04717, -38.27806, -38.50176, -38.71813, 
    -38.92703, -39.12834, -39.32193, -39.50767, -39.68544, -39.85512, 
    -40.0166, -40.16977, -40.31451, -40.45074, -40.57834, -40.69724, 
    -40.80733, -40.90854, -41.0008, -41.08404, -41.15818, -41.22319, -41.279, 
    -41.32558, -41.36288, -41.39089, -41.40957, -41.41891, -41.41891, 
    -41.40957, -41.39089, -41.36288, -41.32558, -41.279, -41.22319, 
    -41.15818, -41.08404, -41.0008, -40.90854, -40.80733, -40.69724, 
    -40.57834, -40.45074, -40.31451, -40.16977, -40.0166, -39.85512, 
    -39.68544, -39.50767, -39.32193, -39.12834, -38.92703, -38.71813, 
    -38.50176, -38.27806, -38.04717, -37.80922, -37.56434, -37.31269, 
    -37.05439, -36.78959, -36.51843, -36.24105, -35.9576, -35.66821, 
    -35.37302, -35.07218, -34.76583, -34.4541, -34.13713, -33.81506, 
    -33.48802, -33.15614, -32.81957, -32.47842, -32.13284,
  -31.39594, -31.73718, -32.07414, -32.40669, -32.73469, -33.05801, 
    -33.37651, -33.69006, -33.99852, -34.30174, -34.59959, -34.89193, 
    -35.1786, -35.45947, -35.73439, -36.00322, -36.26581, -36.52202, 
    -36.7717, -37.01471, -37.2509, -37.48015, -37.70229, -37.9172, -38.12474, 
    -38.32478, -38.51718, -38.70182, -38.87856, -39.04729, -39.20789, 
    -39.36025, -39.50425, -39.63979, -39.76678, -39.88511, -39.99469, 
    -40.09544, -40.18729, -40.27016, -40.34399, -40.40873, -40.46431, 
    -40.51069, -40.54784, -40.57574, -40.59435, -40.60365, -40.60365, 
    -40.59435, -40.57574, -40.54784, -40.51069, -40.46431, -40.40873, 
    -40.34399, -40.27016, -40.18729, -40.09544, -39.99469, -39.88511, 
    -39.76678, -39.63979, -39.50425, -39.36025, -39.20789, -39.04729, 
    -38.87856, -38.70182, -38.51718, -38.32478, -38.12474, -37.9172, 
    -37.70229, -37.48015, -37.2509, -37.01471, -36.7717, -36.52202, 
    -36.26581, -36.00322, -35.73439, -35.45947, -35.1786, -34.89193, 
    -34.59959, -34.30174, -33.99852, -33.69006, -33.37651, -33.05801, 
    -32.73469, -32.40669, -32.07414, -31.73718, -31.39594,
  -30.65893, -30.9956, -31.32814, -31.65643, -31.98032, -32.29969, -32.6144, 
    -32.9243, -33.22925, -33.52912, -33.82376, -34.11302, -34.39675, 
    -34.67482, -34.94707, -35.21335, -35.47353, -35.72744, -35.97494, 
    -36.21589, -36.45013, -36.67753, -36.89794, -37.11122, -37.31722, 
    -37.51582, -37.70687, -37.89024, -38.06581, -38.23346, -38.39304, 
    -38.54446, -38.6876, -38.82234, -38.94859, -39.06625, -39.17523, 
    -39.27544, -39.3668, -39.44924, -39.52269, -39.58709, -39.6424, 
    -39.68855, -39.72552, -39.75327, -39.77179, -39.78105, -39.78105, 
    -39.77179, -39.75327, -39.72552, -39.68855, -39.6424, -39.58709, 
    -39.52269, -39.44924, -39.3668, -39.27544, -39.17523, -39.06625, 
    -38.94859, -38.82234, -38.6876, -38.54446, -38.39304, -38.23346, 
    -38.06581, -37.89024, -37.70687, -37.51582, -37.31722, -37.11122, 
    -36.89794, -36.67753, -36.45013, -36.21589, -35.97494, -35.72744, 
    -35.47353, -35.21335, -34.94707, -34.67482, -34.39675, -34.11302, 
    -33.82376, -33.52912, -33.22925, -32.9243, -32.6144, -32.29969, 
    -31.98032, -31.65643, -31.32814, -30.9956, -30.65893,
  -29.92181, -30.25368, -30.58158, -30.90537, -31.22494, -31.54013, -31.8508, 
    -32.15683, -32.45805, -32.75434, -33.04553, -33.33149, -33.61207, 
    -33.88711, -34.15647, -34.42, -34.67754, -34.92895, -35.17407, -35.41275, 
    -35.64485, -35.87022, -36.08871, -36.30017, -36.50447, -36.70145, 
    -36.891, -37.07295, -37.2472, -37.4136, -37.57203, -37.72238, -37.86452, 
    -37.99836, -38.12377, -38.24066, -38.34894, -38.44851, -38.53931, 
    -38.62124, -38.69425, -38.75827, -38.81324, -38.85912, -38.89588, 
    -38.92347, -38.94188, -38.95109, -38.95109, -38.94188, -38.92347, 
    -38.89588, -38.85912, -38.81324, -38.75827, -38.69425, -38.62124, 
    -38.53931, -38.44851, -38.34894, -38.24066, -38.12377, -37.99836, 
    -37.86452, -37.72238, -37.57203, -37.4136, -37.2472, -37.07295, -36.891, 
    -36.70145, -36.50447, -36.30017, -36.08871, -35.87022, -35.64485, 
    -35.41275, -35.17407, -34.92895, -34.67754, -34.42, -34.15647, -33.88711, 
    -33.61207, -33.33149, -33.04553, -32.75434, -32.45805, -32.15683, 
    -31.8508, -31.54013, -31.22494, -30.90537, -30.58158, -30.25368, -29.92181,
  -29.18457, -29.51142, -29.83445, -30.15354, -30.46854, -30.77932, 
    -31.08575, -31.38766, -31.68493, -31.97741, -32.26494, -32.54737, 
    -32.82457, -33.09637, -33.36263, -33.62318, -33.87788, -34.12658, 
    -34.36911, -34.60533, -34.83509, -35.05824, -35.27462, -35.48409, 
    -35.68649, -35.8817, -36.06956, -36.24994, -36.42271, -36.58773, 
    -36.74487, -36.89401, -37.03504, -37.16784, -37.2923, -37.40832, 
    -37.5158, -37.61465, -37.7048, -37.78615, -37.85865, -37.92222, 
    -37.97682, -38.02239, -38.0589, -38.0863, -38.10459, -38.11374, 
    -38.11374, -38.10459, -38.0863, -38.0589, -38.02239, -37.97682, 
    -37.92222, -37.85865, -37.78615, -37.7048, -37.61465, -37.5158, 
    -37.40832, -37.2923, -37.16784, -37.03504, -36.89401, -36.74487, 
    -36.58773, -36.42271, -36.24994, -36.06956, -35.8817, -35.68649, 
    -35.48409, -35.27462, -35.05824, -34.83509, -34.60533, -34.36911, 
    -34.12658, -33.87788, -33.62318, -33.36263, -33.09637, -32.82457, 
    -32.54737, -32.26494, -31.97741, -31.68493, -31.38766, -31.08575, 
    -30.77932, -30.46854, -30.15354, -29.83445, -29.51142, -29.18457,
  -28.44723, -28.76883, -29.08677, -29.40093, -29.71115, -30.0173, -30.31924, 
    -30.61683, -30.90992, -31.19835, -31.482, -31.76069, -32.03428, 
    -32.30262, -32.56555, -32.82292, -33.07457, -33.32034, -33.56009, 
    -33.79364, -34.02087, -34.2416, -34.45568, -34.66297, -34.86331, 
    -35.05656, -35.24258, -35.42123, -35.59236, -35.75585, -35.91155, 
    -36.05936, -36.19914, -36.33079, -36.45418, -36.56922, -36.67581, 
    -36.77385, -36.86326, -36.94396, -37.01588, -37.07895, -37.13312, 
    -37.17834, -37.21456, -37.24176, -37.2599, -37.26898, -37.26898, 
    -37.2599, -37.24176, -37.21456, -37.17834, -37.13312, -37.07895, 
    -37.01588, -36.94396, -36.86326, -36.77385, -36.67581, -36.56922, 
    -36.45418, -36.33079, -36.19914, -36.05936, -35.91155, -35.75585, 
    -35.59236, -35.42123, -35.24258, -35.05656, -34.86331, -34.66297, 
    -34.45568, -34.2416, -34.02087, -33.79364, -33.56009, -33.32034, 
    -33.07457, -32.82292, -32.56555, -32.30262, -32.03428, -31.76069, 
    -31.482, -31.19835, -30.90992, -30.61683, -30.31924, -30.0173, -29.71115, 
    -29.40093, -29.08677, -28.76883, -28.44723,
  -27.70978, -28.02592, -28.33856, -28.64755, -28.95277, -29.25407, 
    -29.55131, -29.84434, -30.13302, -30.4172, -30.69673, -30.97146, 
    -31.24123, -31.50589, -31.76528, -32.01924, -32.26763, -32.51027, 
    -32.74702, -32.97771, -33.2022, -33.42032, -33.63192, -33.83684, 
    -34.03494, -34.22607, -34.41008, -34.58682, -34.75616, -34.91797, 
    -35.0721, -35.21843, -35.35684, -35.48721, -35.60942, -35.72337, 
    -35.82896, -35.9261, -36.01469, -36.09467, -36.16594, -36.22845, 
    -36.28214, -36.32696, -36.36287, -36.38982, -36.40781, -36.41681, 
    -36.41681, -36.40781, -36.38982, -36.36287, -36.32696, -36.28214, 
    -36.22845, -36.16594, -36.09467, -36.01469, -35.9261, -35.82896, 
    -35.72337, -35.60942, -35.48721, -35.35684, -35.21843, -35.0721, 
    -34.91797, -34.75616, -34.58682, -34.41008, -34.22607, -34.03494, 
    -33.83684, -33.63192, -33.42032, -33.2022, -32.97771, -32.74702, 
    -32.51027, -32.26763, -32.01924, -31.76528, -31.50589, -31.24123, 
    -30.97146, -30.69673, -30.4172, -30.13302, -29.84434, -29.55131, 
    -29.25407, -28.95277, -28.64755, -28.33856, -28.02592, -27.70978,
  -26.97222, -27.28269, -27.58981, -27.89343, -28.19342, -28.48965, 
    -28.78197, -29.07022, -29.35428, -29.63398, -29.90917, -30.17971, 
    -30.44544, -30.7062, -30.96183, -31.21218, -31.45709, -31.6964, 
    -31.92994, -32.15757, -32.37912, -32.59444, -32.80336, -33.00574, 
    -33.20141, -33.39024, -33.57207, -33.74675, -33.91414, -34.07411, 
    -34.22652, -34.37123, -34.50814, -34.6371, -34.75802, -34.87078, 
    -34.97528, -35.07141, -35.15911, -35.23827, -35.30883, -35.37072, 
    -35.42388, -35.46826, -35.50381, -35.53051, -35.54832, -35.55723, 
    -35.55723, -35.54832, -35.53051, -35.50381, -35.46826, -35.42388, 
    -35.37072, -35.30883, -35.23827, -35.15911, -35.07141, -34.97528, 
    -34.87078, -34.75802, -34.6371, -34.50814, -34.37123, -34.22652, 
    -34.07411, -33.91414, -33.74675, -33.57207, -33.39024, -33.20141, 
    -33.00574, -32.80336, -32.59444, -32.37912, -32.15757, -31.92994, 
    -31.6964, -31.45709, -31.21218, -30.96183, -30.7062, -30.44544, 
    -30.17971, -29.90917, -29.63398, -29.35428, -29.07022, -28.78197, 
    -28.48965, -28.19342, -27.89343, -27.58981, -27.28269, -26.97222,
  -26.23456, -26.53915, -26.84053, -27.13857, -27.43312, -27.72406, 
    -28.01123, -28.29449, -28.5737, -28.84871, -29.11935, -29.38548, 
    -29.64695, -29.90359, -30.15525, -30.40177, -30.643, -30.87876, 
    -31.10889, -31.33325, -31.55167, -31.76398, -31.97004, -32.16968, 
    -32.36275, -32.5491, -32.72858, -32.90103, -33.06631, -33.2243, 
    -33.37484, -33.5178, -33.65307, -33.78051, -33.90001, -34.01146, 
    -34.11476, -34.20981, -34.29651, -34.37479, -34.44456, -34.50577, 
    -34.55835, -34.60224, -34.63741, -34.66381, -34.68143, -34.69025, 
    -34.69025, -34.68143, -34.66381, -34.63741, -34.60224, -34.55835, 
    -34.50577, -34.44456, -34.37479, -34.29651, -34.20981, -34.11476, 
    -34.01146, -33.90001, -33.78051, -33.65307, -33.5178, -33.37484, 
    -33.2243, -33.06631, -32.90103, -32.72858, -32.5491, -32.36275, 
    -32.16968, -31.97004, -31.76398, -31.55167, -31.33325, -31.10889, 
    -30.87876, -30.643, -30.40177, -30.15525, -29.90359, -29.64695, 
    -29.38548, -29.11935, -28.84871, -28.5737, -28.29449, -28.01123, 
    -27.72406, -27.43312, -27.13857, -26.84053, -26.53915, -26.23456,
  -25.4968, -25.7953, -26.09074, -26.38298, -26.67189, -26.95732, -27.23913, 
    -27.51719, -27.79133, -28.06141, -28.32729, -28.5888, -28.84579, 
    -29.0981, -29.34557, -29.58805, -29.82537, -30.05738, -30.28391, 
    -30.50479, -30.71988, -30.929, -31.132, -31.32872, -31.519, -31.70269, 
    -31.87964, -32.0497, -32.21272, -32.36856, -32.51709, -32.65816, 
    -32.79165, -32.91744, -33.03541, -33.14545, -33.24744, -33.3413, 
    -33.42693, -33.50424, -33.57316, -33.63363, -33.68556, -33.72892, 
    -33.76367, -33.78976, -33.80717, -33.81588, -33.81588, -33.80717, 
    -33.78976, -33.76367, -33.72892, -33.68556, -33.63363, -33.57316, 
    -33.50424, -33.42693, -33.3413, -33.24744, -33.14545, -33.03541, 
    -32.91744, -32.79165, -32.65816, -32.51709, -32.36856, -32.21272, 
    -32.0497, -31.87964, -31.70269, -31.519, -31.32872, -31.132, -30.929, 
    -30.71988, -30.50479, -30.28391, -30.05738, -29.82537, -29.58805, 
    -29.34557, -29.0981, -28.84579, -28.5888, -28.32729, -28.06141, 
    -27.79133, -27.51719, -27.23913, -26.95732, -26.67189, -26.38298, 
    -26.09074, -25.7953, -25.4968,
  -24.75893, -25.05115, -25.34044, -25.62668, -25.90973, -26.18944, 
    -26.46569, -26.73832, -27.00718, -27.27213, -27.53302, -27.78969, 
    -28.04199, -28.28975, -28.53283, -28.77106, -29.00427, -29.23232, 
    -29.45502, -29.67224, -29.88379, -30.08952, -30.28927, -30.48288, 
    -30.6702, -30.85106, -31.02531, -31.19281, -31.3534, -31.50695, 
    -31.65331, -31.79235, -31.92393, -32.04794, -32.16426, -32.27277, 
    -32.37335, -32.46593, -32.55039, -32.62666, -32.69466, -32.75431, 
    -32.80555, -32.84834, -32.88263, -32.90837, -32.92555, -32.93415, 
    -32.93415, -32.92555, -32.90837, -32.88263, -32.84834, -32.80555, 
    -32.75431, -32.69466, -32.62666, -32.55039, -32.46593, -32.37335, 
    -32.27277, -32.16426, -32.04794, -31.92393, -31.79235, -31.65331, 
    -31.50695, -31.3534, -31.19281, -31.02531, -30.85106, -30.6702, 
    -30.48288, -30.28927, -30.08952, -29.88379, -29.67224, -29.45502, 
    -29.23232, -29.00427, -28.77106, -28.53283, -28.28975, -28.04199, 
    -27.78969, -27.53302, -27.27213, -27.00718, -26.73832, -26.46569, 
    -26.18944, -25.90973, -25.62668, -25.34044, -25.05115, -24.75893,
  -24.02097, -24.3067, -24.58965, -24.86968, -25.14667, -25.42046, -25.69092, 
    -25.95792, -26.22129, -26.4809, -26.73659, -26.98821, -27.2356, 
    -27.47861, -27.71707, -27.95084, -28.17974, -28.40361, -28.6223, 
    -28.83563, -29.04346, -29.2456, -29.44192, -29.63223, -29.81639, 
    -29.99424, -30.16563, -30.3304, -30.4884, -30.6395, -30.78355, -30.92041, 
    -31.04995, -31.17205, -31.28659, -31.39346, -31.49253, -31.58372, 
    -31.66694, -31.74208, -31.80908, -31.86786, -31.91836, -31.96053, 
    -31.99432, -32.01969, -32.03662, -32.04509, -32.04509, -32.03662, 
    -32.01969, -31.99432, -31.96053, -31.91836, -31.86786, -31.80908, 
    -31.74208, -31.66694, -31.58372, -31.49253, -31.39346, -31.28659, 
    -31.17205, -31.04995, -30.92041, -30.78355, -30.6395, -30.4884, -30.3304, 
    -30.16563, -29.99424, -29.81639, -29.63223, -29.44192, -29.2456, 
    -29.04346, -28.83563, -28.6223, -28.40361, -28.17974, -27.95084, 
    -27.71707, -27.47861, -27.2356, -26.98821, -26.73659, -26.4809, 
    -26.22129, -25.95792, -25.69092, -25.42046, -25.14667, -24.86968, 
    -24.58965, -24.3067, -24.02097,
  -23.28291, -23.56197, -23.83837, -24.112, -24.38272, -24.65038, -24.91487, 
    -25.17602, -25.43369, -25.68774, -25.93803, -26.18438, -26.42666, 
    -26.6647, -26.89834, -27.12744, -27.35181, -27.57131, -27.78577, 
    -27.99503, -28.19893, -28.3973, -28.58998, -28.77681, -28.95764, 
    -29.1323, -29.30065, -29.46252, -29.61777, -29.76627, -29.90785, 
    -30.04239, -30.16976, -30.28983, -30.40247, -30.50758, -30.60504, 
    -30.69475, -30.77662, -30.85055, -30.91648, -30.97433, -31.02403, 
    -31.06553, -31.09879, -31.12376, -31.14043, -31.14876, -31.14876, 
    -31.14043, -31.12376, -31.09879, -31.06553, -31.02403, -30.97433, 
    -30.91648, -30.85055, -30.77662, -30.69475, -30.60504, -30.50758, 
    -30.40247, -30.28983, -30.16976, -30.04239, -29.90785, -29.76627, 
    -29.61777, -29.46252, -29.30065, -29.1323, -28.95764, -28.77681, 
    -28.58998, -28.3973, -28.19893, -27.99503, -27.78577, -27.57131, 
    -27.35181, -27.12744, -26.89834, -26.6647, -26.42666, -26.18438, 
    -25.93803, -25.68774, -25.43369, -25.17602, -24.91487, -24.65038, 
    -24.38272, -24.112, -23.83837, -23.56197, -23.28291,
  -22.54476, -22.81695, -23.08662, -23.35365, -23.6179, -23.87924, -24.13754, 
    -24.39264, -24.64441, -24.89271, -25.13737, -25.37826, -25.61521, 
    -25.84807, -26.07669, -26.30091, -26.52055, -26.73548, -26.94551, 
    -27.1505, -27.35027, -27.54466, -27.73353, -27.91669, -28.094, -28.2653, 
    -28.43043, -28.58924, -28.74158, -28.88731, -29.02629, -29.15837, 
    -29.28342, -29.40132, -29.51195, -29.61518, -29.71092, -29.79905, 
    -29.87949, -29.95214, -30.01692, -30.07377, -30.12261, -30.1634, 
    -30.19609, -30.22064, -30.23702, -30.24521, -30.24521, -30.23702, 
    -30.22064, -30.19609, -30.1634, -30.12261, -30.07377, -30.01692, 
    -29.95214, -29.87949, -29.79905, -29.71092, -29.61518, -29.51195, 
    -29.40132, -29.28342, -29.15837, -29.02629, -28.88731, -28.74158, 
    -28.58924, -28.43043, -28.2653, -28.094, -27.91669, -27.73353, -27.54466, 
    -27.35027, -27.1505, -26.94551, -26.73548, -26.52055, -26.30091, 
    -26.07669, -25.84807, -25.61521, -25.37826, -25.13737, -24.89271, 
    -24.64441, -24.39264, -24.13754, -23.87924, -23.6179, -23.35365, 
    -23.08662, -22.81695, -22.54476,
  -21.80651, -22.07165, -22.33441, -22.59464, -22.85224, -23.10706, 
    -23.35897, -23.60783, -23.85349, -24.09582, -24.33467, -24.56988, 
    -24.8013, -25.02878, -25.25217, -25.4713, -25.68602, -25.89616, 
    -26.10157, -26.30208, -26.49753, -26.68777, -26.87262, -27.05193, 
    -27.22555, -27.3933, -27.55505, -27.71063, -27.8599, -28.00271, 
    -28.13892, -28.2684, -28.391, -28.50661, -28.6151, -28.71634, -28.81025, 
    -28.89671, -28.97562, -29.0469, -29.11047, -29.16625, -29.21418, 
    -29.25421, -29.28629, -29.31038, -29.32646, -29.33451, -29.33451, 
    -29.32646, -29.31038, -29.28629, -29.25421, -29.21418, -29.16625, 
    -29.11047, -29.0469, -28.97562, -28.89671, -28.81025, -28.71634, 
    -28.6151, -28.50661, -28.391, -28.2684, -28.13892, -28.00271, -27.8599, 
    -27.71063, -27.55505, -27.3933, -27.22555, -27.05193, -26.87262, 
    -26.68777, -26.49753, -26.30208, -26.10157, -25.89616, -25.68602, 
    -25.4713, -25.25217, -25.02878, -24.8013, -24.56988, -24.33467, 
    -24.09582, -23.85349, -23.60783, -23.35897, -23.10706, -22.85224, 
    -22.59464, -22.33441, -22.07165, -21.80651,
  -21.06818, -21.32609, -21.58174, -21.835, -22.08575, -22.33386, -22.57919, 
    -22.8216, -23.06096, -23.29713, -23.52995, -23.75929, -23.98498, 
    -24.20688, -24.42483, -24.63868, -24.84826, -25.05343, -25.25401, 
    -25.44986, -25.6408, -25.82668, -26.00734, -26.18261, -26.35234, 
    -26.51638, -26.67457, -26.82676, -26.9728, -27.11254, -27.24584, 
    -27.37256, -27.49258, -27.60576, -27.71199, -27.81114, -27.90311, 
    -27.98779, -28.06509, -28.13491, -28.19719, -28.25185, -28.29881, 
    -28.33804, -28.36947, -28.39308, -28.40884, -28.41672, -28.41672, 
    -28.40884, -28.39308, -28.36947, -28.33804, -28.29881, -28.25185, 
    -28.19719, -28.13491, -28.06509, -27.98779, -27.90311, -27.81114, 
    -27.71199, -27.60576, -27.49258, -27.37256, -27.24584, -27.11254, 
    -26.9728, -26.82676, -26.67457, -26.51638, -26.35234, -26.18261, 
    -26.00734, -25.82668, -25.6408, -25.44986, -25.25401, -25.05343, 
    -24.84826, -24.63868, -24.42483, -24.20688, -23.98498, -23.75929, 
    -23.52995, -23.29713, -23.06096, -22.8216, -22.57919, -22.33386, 
    -22.08575, -21.835, -21.58174, -21.32609, -21.06818,
  -20.32976, -20.58027, -20.82863, -21.07474, -21.31846, -21.55966, 
    -21.79822, -22.034, -22.26687, -22.49667, -22.72328, -22.94654, -23.1663, 
    -23.38242, -23.59474, -23.8031, -24.00736, -24.20735, -24.40292, 
    -24.5939, -24.78014, -24.96147, -25.13775, -25.3088, -25.47448, 
    -25.63463, -25.78909, -25.93772, -26.08036, -26.21687, -26.34712, 
    -26.47095, -26.58825, -26.69888, -26.80272, -26.89966, -26.98958, 
    -27.07239, -27.14798, -27.21628, -27.27719, -27.33065, -27.3766, 
    -27.41497, -27.44572, -27.46882, -27.48424, -27.49195, -27.49195, 
    -27.48424, -27.46882, -27.44572, -27.41497, -27.3766, -27.33065, 
    -27.27719, -27.21628, -27.14798, -27.07239, -26.98958, -26.89966, 
    -26.80272, -26.69888, -26.58825, -26.47095, -26.34712, -26.21687, 
    -26.08036, -25.93772, -25.78909, -25.63463, -25.47448, -25.3088, 
    -25.13775, -24.96147, -24.78014, -24.5939, -24.40292, -24.20735, 
    -24.00736, -23.8031, -23.59474, -23.38242, -23.1663, -22.94654, 
    -22.72328, -22.49667, -22.26687, -22.034, -21.79822, -21.55966, 
    -21.31846, -21.07474, -20.82863, -20.58027, -20.32976,
  -19.59126, -19.83419, -20.0751, -20.31387, -20.55038, -20.7845, -21.01611, 
    -21.24507, -21.47124, -21.6945, -21.91469, -22.13168, -22.34532, 
    -22.55546, -22.76195, -22.96464, -23.16337, -23.35799, -23.54835, 
    -23.73428, -23.91562, -24.09223, -24.26394, -24.43059, -24.59204, 
    -24.74813, -24.89869, -25.04359, -25.18268, -25.31582, -25.44285, 
    -25.56366, -25.6781, -25.78605, -25.88738, -25.98199, -26.06977, 
    -26.1506, -26.2244, -26.29108, -26.35056, -26.40276, -26.44763, -26.4851, 
    -26.51514, -26.5377, -26.55275, -26.56029, -26.56029, -26.55275, 
    -26.5377, -26.51514, -26.4851, -26.44763, -26.40276, -26.35056, 
    -26.29108, -26.2244, -26.1506, -26.06977, -25.98199, -25.88738, 
    -25.78605, -25.6781, -25.56366, -25.44285, -25.31582, -25.18268, 
    -25.04359, -24.89869, -24.74813, -24.59204, -24.43059, -24.26394, 
    -24.09223, -23.91562, -23.73428, -23.54835, -23.35799, -23.16337, 
    -22.96464, -22.76195, -22.55546, -22.34532, -22.13168, -21.91469, 
    -21.6945, -21.47124, -21.24507, -21.01611, -20.7845, -20.55038, 
    -20.31387, -20.0751, -19.83419, -19.59126,
  -18.85267, -19.08786, -19.32115, -19.55242, -19.78154, -20.0084, -20.23287, 
    -20.45482, -20.67413, -20.89065, -21.10424, -21.31477, -21.52209, 
    -21.72607, -21.92654, -22.12335, -22.31637, -22.50543, -22.69039, 
    -22.87107, -23.04734, -23.21904, -23.386, -23.54808, -23.70512, 
    -23.85697, -24.00347, -24.14449, -24.27987, -24.40947, -24.53315, 
    -24.65079, -24.76223, -24.86737, -24.96609, -25.05826, -25.14377, 
    -25.22254, -25.29446, -25.35944, -25.41741, -25.46829, -25.51202, 
    -25.54855, -25.57783, -25.59982, -25.6145, -25.62184, -25.62184, 
    -25.6145, -25.59982, -25.57783, -25.54855, -25.51202, -25.46829, 
    -25.41741, -25.35944, -25.29446, -25.22254, -25.14377, -25.05826, 
    -24.96609, -24.86737, -24.76223, -24.65079, -24.53315, -24.40947, 
    -24.27987, -24.14449, -24.00347, -23.85697, -23.70512, -23.54808, 
    -23.386, -23.21904, -23.04734, -22.87107, -22.69039, -22.50543, 
    -22.31637, -22.12335, -21.92654, -21.72607, -21.52209, -21.31477, 
    -21.10424, -20.89065, -20.67413, -20.45482, -20.23287, -20.0084, 
    -19.78154, -19.55242, -19.32115, -19.08786, -18.85267,
  -18.114, -18.3413, -18.5668, -18.79039, -19.01196, -19.23139, -19.44855, 
    -19.66332, -19.87557, -20.08517, -20.29198, -20.49586, -20.69669, 
    -20.8943, -21.08856, -21.27932, -21.46644, -21.64975, -21.82912, 
    -22.00438, -22.17539, -22.34199, -22.50403, -22.66135, -22.81381, 
    -22.96125, -23.10353, -23.2405, -23.37202, -23.49794, -23.61813, 
    -23.73245, -23.84077, -23.94298, -24.03895, -24.12856, -24.21172, 
    -24.28832, -24.35827, -24.42147, -24.47786, -24.52736, -24.5699, 
    -24.60544, -24.63392, -24.65532, -24.6696, -24.67674, -24.67674, 
    -24.6696, -24.65532, -24.63392, -24.60544, -24.5699, -24.52736, 
    -24.47786, -24.42147, -24.35827, -24.28832, -24.21172, -24.12856, 
    -24.03895, -23.94298, -23.84077, -23.73245, -23.61813, -23.49794, 
    -23.37202, -23.2405, -23.10353, -22.96125, -22.81381, -22.66135, 
    -22.50403, -22.34199, -22.17539, -22.00438, -21.82912, -21.64975, 
    -21.46644, -21.27932, -21.08856, -20.8943, -20.69669, -20.49586, 
    -20.29198, -20.08517, -19.87557, -19.66332, -19.44855, -19.23139, 
    -19.01196, -18.79039, -18.5668, -18.3413, -18.114,
  -17.37526, -17.59451, -17.81206, -18.02782, -18.24167, -18.45349, 
    -18.66317, -18.87058, -19.07561, -19.2781, -19.47795, -19.67501, 
    -19.86915, -20.06023, -20.2481, -20.43262, -20.61365, -20.79103, 
    -20.96463, -21.13428, -21.29985, -21.46118, -21.61812, -21.77052, 
    -21.91823, -22.0611, -22.19899, -22.33176, -22.45926, -22.58134, 
    -22.69789, -22.80877, -22.91384, -23.01299, -23.10609, -23.19304, 
    -23.27374, -23.34808, -23.41596, -23.47731, -23.53204, -23.58009, 
    -23.62139, -23.6559, -23.68355, -23.70432, -23.71819, -23.72513, 
    -23.72513, -23.71819, -23.70432, -23.68355, -23.6559, -23.62139, 
    -23.58009, -23.53204, -23.47731, -23.41596, -23.34808, -23.27374, 
    -23.19304, -23.10609, -23.01299, -22.91384, -22.80877, -22.69789, 
    -22.58134, -22.45926, -22.33176, -22.19899, -22.0611, -21.91823, 
    -21.77052, -21.61812, -21.46118, -21.29985, -21.13428, -20.96463, 
    -20.79103, -20.61365, -20.43262, -20.2481, -20.06023, -19.86915, 
    -19.67501, -19.47795, -19.2781, -19.07561, -18.87058, -18.66317, 
    -18.45349, -18.24167, -18.02782, -17.81206, -17.59451, -17.37526,
  -16.63645, -16.84749, -17.05695, -17.26471, -17.47068, -17.67474, 
    -17.87678, -18.07666, -18.27429, -18.46952, -18.66223, -18.85229, 
    -19.03956, -19.22392, -19.40522, -19.58332, -19.75808, -19.92936, 
    -20.09701, -20.26088, -20.42083, -20.57672, -20.72838, -20.87569, 
    -21.01848, -21.15662, -21.28997, -21.41838, -21.5417, -21.65982, 
    -21.77258, -21.87987, -21.98156, -22.07753, -22.16766, -22.25184, 
    -22.32997, -22.40195, -22.46768, -22.52709, -22.5801, -22.62664, 
    -22.66665, -22.70007, -22.72686, -22.74698, -22.76041, -22.76713, 
    -22.76713, -22.76041, -22.74698, -22.72686, -22.70007, -22.66665, 
    -22.62664, -22.5801, -22.52709, -22.46768, -22.40195, -22.32997, 
    -22.25184, -22.16766, -22.07753, -21.98156, -21.87987, -21.77258, 
    -21.65982, -21.5417, -21.41838, -21.28997, -21.15662, -21.01848, 
    -20.87569, -20.72838, -20.57672, -20.42083, -20.26088, -20.09701, 
    -19.92936, -19.75808, -19.58332, -19.40522, -19.22392, -19.03956, 
    -18.85229, -18.66223, -18.46952, -18.27429, -18.07666, -17.87678, 
    -17.67474, -17.47068, -17.26471, -17.05695, -16.84749, -16.63645,
  -15.89756, -16.10026, -16.30147, -16.50109, -16.69903, -16.89517, -17.0894, 
    -17.2816, -17.47165, -17.65945, -17.84485, -18.02774, -18.20799, 
    -18.38545, -18.56001, -18.73152, -18.89984, -19.06483, -19.22636, 
    -19.38427, -19.53844, -19.68871, -19.83493, -19.97698, -20.11469, 
    -20.24794, -20.37659, -20.50048, -20.61949, -20.73348, -20.84233, 
    -20.94591, -21.04409, -21.13675, -21.22379, -21.30509, -21.38055, 
    -21.45008, -21.51358, -21.57098, -21.6222, -21.66716, -21.70582, 
    -21.73811, -21.764, -21.78345, -21.79643, -21.80292, -21.80292, 
    -21.79643, -21.78345, -21.764, -21.73811, -21.70582, -21.66716, -21.6222, 
    -21.57098, -21.51358, -21.45008, -21.38055, -21.30509, -21.22379, 
    -21.13675, -21.04409, -20.94591, -20.84233, -20.73348, -20.61949, 
    -20.50048, -20.37659, -20.24794, -20.11469, -19.97698, -19.83493, 
    -19.68871, -19.53844, -19.38427, -19.22636, -19.06483, -18.89984, 
    -18.73152, -18.56001, -18.38545, -18.20799, -18.02774, -17.84485, 
    -17.65945, -17.47165, -17.2816, -17.0894, -16.89517, -16.69903, 
    -16.50109, -16.30147, -16.10026, -15.89756,
  -15.15861, -15.35282, -15.54564, -15.73699, -15.92674, -16.11481, 
    -16.30107, -16.48543, -16.66776, -16.84796, -17.02589, -17.20144, 
    -17.37449, -17.5449, -17.71254, -17.87728, -18.03899, -18.19754, 
    -18.35277, -18.50457, -18.65277, -18.79726, -18.93789, -19.07451, 
    -19.20699, -19.33519, -19.45897, -19.57821, -19.69276, -19.8025, 
    -19.90729, -20.00702, -20.10156, -20.19081, -20.27464, -20.35295, 
    -20.42565, -20.49264, -20.55383, -20.60913, -20.65849, -20.70182, 
    -20.73908, -20.7702, -20.79515, -20.81389, -20.8264, -20.83266, 
    -20.83266, -20.8264, -20.81389, -20.79515, -20.7702, -20.73908, 
    -20.70182, -20.65849, -20.60913, -20.55383, -20.49264, -20.42565, 
    -20.35295, -20.27464, -20.19081, -20.10156, -20.00702, -19.90729, 
    -19.8025, -19.69276, -19.57821, -19.45897, -19.33519, -19.20699, 
    -19.07451, -18.93789, -18.79726, -18.65277, -18.50457, -18.35277, 
    -18.19754, -18.03899, -17.87728, -17.71254, -17.5449, -17.37449, 
    -17.20144, -17.02589, -16.84796, -16.66776, -16.48543, -16.30107, 
    -16.11481, -15.92674, -15.73699, -15.54564, -15.35282, -15.15861,
  -14.41959, -14.60518, -14.78949, -14.9724, -15.15383, -15.33368, -15.51184, 
    -15.6882, -15.86266, -16.0351, -16.20541, -16.37346, -16.53915, 
    -16.70233, -16.8629, -17.02072, -17.17565, -17.32758, -17.47636, 
    -17.62187, -17.76396, -17.9025, -18.03736, -18.16841, -18.2955, -18.4185, 
    -18.53728, -18.65171, -18.76166, -18.867, -18.96761, -19.06337, 
    -19.15416, -19.23986, -19.32038, -19.39561, -19.46544, -19.5298, 
    -19.58859, -19.64173, -19.68916, -19.7308, -19.7666, -19.79651, 
    -19.82049, -19.8385, -19.85053, -19.85655, -19.85655, -19.85053, 
    -19.8385, -19.82049, -19.79651, -19.7666, -19.7308, -19.68916, -19.64173, 
    -19.58859, -19.5298, -19.46544, -19.39561, -19.32038, -19.23986, 
    -19.15416, -19.06337, -18.96761, -18.867, -18.76166, -18.65171, 
    -18.53728, -18.4185, -18.2955, -18.16841, -18.03736, -17.9025, -17.76396, 
    -17.62187, -17.47636, -17.32758, -17.17565, -17.02072, -16.8629, 
    -16.70233, -16.53915, -16.37346, -16.20541, -16.0351, -15.86266, 
    -15.6882, -15.51184, -15.33368, -15.15383, -14.9724, -14.78949, 
    -14.60518, -14.41959,
  -13.6805, -13.85736, -14.03301, -14.20737, -14.38034, -14.55183, -14.72173, 
    -14.88996, -15.05639, -15.22093, -15.38346, -15.54386, -15.70203, 
    -15.85784, -16.01117, -16.1619, -16.30991, -16.45506, -16.59723, 
    -16.73629, -16.87211, -17.00456, -17.1335, -17.25882, -17.38036, 
    -17.49802, -17.61165, -17.72114, -17.82635, -17.92716, -18.02345, 
    -18.11512, -18.20203, -18.28409, -18.36119, -18.43323, -18.50011, 
    -18.56174, -18.61805, -18.66896, -18.71439, -18.75428, -18.78858, 
    -18.81724, -18.84021, -18.85747, -18.86899, -18.87476, -18.87476, 
    -18.86899, -18.85747, -18.84021, -18.81724, -18.78858, -18.75428, 
    -18.71439, -18.66896, -18.61805, -18.56174, -18.50011, -18.43323, 
    -18.36119, -18.28409, -18.20203, -18.11512, -18.02345, -17.92716, 
    -17.82635, -17.72114, -17.61165, -17.49802, -17.38036, -17.25882, 
    -17.1335, -17.00456, -16.87211, -16.73629, -16.59723, -16.45506, 
    -16.30991, -16.1619, -16.01117, -15.85784, -15.70203, -15.54386, 
    -15.38346, -15.22093, -15.05639, -14.88996, -14.72173, -14.55183, 
    -14.38034, -14.20737, -14.03301, -13.85736, -13.6805,
  -12.94136, -13.10935, -13.27623, -13.4419, -13.60628, -13.76928, -13.9308, 
    -14.09074, -14.24901, -14.4055, -14.56011, -14.71272, -14.86322, 
    -15.0115, -15.15745, -15.30094, -15.44186, -15.58009, -15.71549, 
    -15.84795, -15.97735, -16.10355, -16.22643, -16.34587, -16.46173, 
    -16.57389, -16.68224, -16.78664, -16.88698, -16.98314, -17.075, 
    -17.16244, -17.24537, -17.32367, -17.39725, -17.466, -17.52983, 
    -17.58866, -17.64242, -17.69101, -17.73438, -17.77247, -17.80522, 
    -17.83258, -17.85452, -17.871, -17.882, -17.88751, -17.88751, -17.882, 
    -17.871, -17.85452, -17.83258, -17.80522, -17.77247, -17.73438, 
    -17.69101, -17.64242, -17.58866, -17.52983, -17.466, -17.39725, 
    -17.32367, -17.24537, -17.16244, -17.075, -16.98314, -16.88698, 
    -16.78664, -16.68224, -16.57389, -16.46173, -16.34587, -16.22643, 
    -16.10355, -15.97735, -15.84795, -15.71549, -15.58009, -15.44186, 
    -15.30094, -15.15745, -15.0115, -14.86322, -14.71272, -14.56011, 
    -14.4055, -14.24901, -14.09074, -13.9308, -13.76928, -13.60628, -13.4419, 
    -13.27623, -13.10935, -12.94136,
  -12.20216, -12.36118, -12.51916, -12.67602, -12.83169, -12.98607, 
    -13.13908, -13.29061, -13.44058, -13.58888, -13.73542, -13.88009, 
    -14.02279, -14.1634, -14.30182, -14.43793, -14.57162, -14.70277, 
    -14.83126, -14.95698, -15.07981, -15.19962, -15.31629, -15.42971, 
    -15.53974, -15.64629, -15.74921, -15.8484, -15.94374, -16.03511, 
    -16.12242, -16.20553, -16.28436, -16.3588, -16.42875, -16.49412, 
    -16.55482, -16.61077, -16.66188, -16.7081, -16.74936, -16.78558, 
    -16.81673, -16.84276, -16.86363, -16.87931, -16.88978, -16.89501, 
    -16.89501, -16.88978, -16.87931, -16.86363, -16.84276, -16.81673, 
    -16.78558, -16.74936, -16.7081, -16.66188, -16.61077, -16.55482, 
    -16.49412, -16.42875, -16.3588, -16.28436, -16.20553, -16.12242, 
    -16.03511, -15.94374, -15.8484, -15.74921, -15.64629, -15.53974, 
    -15.42971, -15.31629, -15.19962, -15.07981, -14.95698, -14.83126, 
    -14.70277, -14.57162, -14.43793, -14.30182, -14.1634, -14.02279, 
    -13.88009, -13.73542, -13.58888, -13.44058, -13.29061, -13.13908, 
    -12.98607, -12.83169, -12.67602, -12.51916, -12.36118, -12.20216,
  -11.46291, -11.61284, -11.76182, -11.90976, -12.05659, -12.20224, -12.3466, 
    -12.4896, -12.63114, -12.77113, -12.90947, -13.04607, -13.18083, 
    -13.31363, -13.44438, -13.57297, -13.69929, -13.82323, -13.94467, 
    -14.0635, -14.17962, -14.2929, -14.40323, -14.51049, -14.61457, 
    -14.71535, -14.81272, -14.90658, -14.99679, -15.08327, -15.1659, 
    -15.24457, -15.3192, -15.38967, -15.4559, -15.5178, -15.57528, -15.62826, 
    -15.67667, -15.72045, -15.75952, -15.79384, -15.82335, -15.84801, 
    -15.86777, -15.88263, -15.89254, -15.8975, -15.8975, -15.89254, 
    -15.88263, -15.86777, -15.84801, -15.82335, -15.79384, -15.75952, 
    -15.72045, -15.67667, -15.62826, -15.57528, -15.5178, -15.4559, 
    -15.38967, -15.3192, -15.24457, -15.1659, -15.08327, -14.99679, 
    -14.90658, -14.81272, -14.71535, -14.61457, -14.51049, -14.40323, 
    -14.2929, -14.17962, -14.0635, -13.94467, -13.82323, -13.69929, 
    -13.57297, -13.44438, -13.31363, -13.18083, -13.04607, -12.90947, 
    -12.77113, -12.63114, -12.4896, -12.3466, -12.20224, -12.05659, 
    -11.90976, -11.76182, -11.61284, -11.46291,
  -10.72361, -10.86435, -11.00421, -11.14313, -11.28102, -11.41781, 
    -11.55342, -11.68776, -11.82075, -11.9523, -12.08233, -12.21073, 
    -12.33741, -12.46228, -12.58523, -12.70616, -12.82498, -12.94157, 
    -13.05583, -13.16765, -13.27692, -13.38354, -13.48739, -13.58837, 
    -13.68636, -13.78126, -13.87296, -13.96135, -14.04633, -14.1278, 
    -14.20564, -14.27977, -14.35008, -14.4165, -14.47891, -14.53725, 
    -14.59143, -14.64138, -14.68701, -14.72828, -14.76512, -14.79747, 
    -14.8253, -14.84855, -14.86719, -14.88119, -14.89054, -14.89522, 
    -14.89522, -14.89054, -14.88119, -14.86719, -14.84855, -14.8253, 
    -14.79747, -14.76512, -14.72828, -14.68701, -14.64138, -14.59143, 
    -14.53725, -14.47891, -14.4165, -14.35008, -14.27977, -14.20564, 
    -14.1278, -14.04633, -13.96135, -13.87296, -13.78126, -13.68636, 
    -13.58837, -13.48739, -13.38354, -13.27692, -13.16765, -13.05583, 
    -12.94157, -12.82498, -12.70616, -12.58523, -12.46228, -12.33741, 
    -12.21073, -12.08233, -11.9523, -11.82075, -11.68776, -11.55342, 
    -11.41781, -11.28102, -11.14313, -11.00421, -10.86435, -10.72361,
  -9.984256, -10.11571, -10.24637, -10.37615, -10.505, -10.63283, -10.75957, 
    -10.88514, -11.00947, -11.13247, -11.25405, -11.37413, -11.49262, 
    -11.60943, -11.72446, -11.83762, -11.9488, -12.05792, -12.16487, 
    -12.26954, -12.37185, -12.47168, -12.56893, -12.66351, -12.75529, 
    -12.84419, -12.9301, -13.01292, -13.09255, -13.16889, -13.24185, 
    -13.31133, -13.37724, -13.43949, -13.49801, -13.55271, -13.60351, 
    -13.65034, -13.69314, -13.73184, -13.76639, -13.79673, -13.82283, 
    -13.84463, -13.86212, -13.87526, -13.88403, -13.88841, -13.88841, 
    -13.88403, -13.87526, -13.86212, -13.84463, -13.82283, -13.79673, 
    -13.76639, -13.73184, -13.69314, -13.65034, -13.60351, -13.55271, 
    -13.49801, -13.43949, -13.37724, -13.31133, -13.24185, -13.16889, 
    -13.09255, -13.01292, -12.9301, -12.84419, -12.75529, -12.66351, 
    -12.56893, -12.47168, -12.37185, -12.26954, -12.16487, -12.05792, 
    -11.9488, -11.83762, -11.72446, -11.60943, -11.49262, -11.37413, 
    -11.25405, -11.13247, -11.00947, -10.88514, -10.75957, -10.63283, 
    -10.505, -10.37615, -10.24637, -10.11571, -9.984256,
  -9.244861, -9.366945, -9.488298, -9.608856, -9.728554, -9.847324, 
    -9.965097, -10.0818, -10.19736, -10.31169, -10.42472, -10.53637, 
    -10.64656, -10.75519, -10.86218, -10.96744, -11.07087, -11.1724, 
    -11.27192, -11.36934, -11.46456, -11.55748, -11.64802, -11.73607, 
    -11.82154, -11.90432, -11.98433, -12.06147, -12.13564, -12.20676, 
    -12.27472, -12.33946, -12.40088, -12.45889, -12.51342, -12.5644, 
    -12.61175, -12.6554, -12.6953, -12.73137, -12.76358, -12.79187, -12.8162, 
    -12.83653, -12.85283, -12.86508, -12.87325, -12.87735, -12.87735, 
    -12.87325, -12.86508, -12.85283, -12.83653, -12.8162, -12.79187, 
    -12.76358, -12.73137, -12.6953, -12.6554, -12.61175, -12.5644, -12.51342, 
    -12.45889, -12.40088, -12.33946, -12.27472, -12.20676, -12.13564, 
    -12.06147, -11.98433, -11.90432, -11.82154, -11.73607, -11.64802, 
    -11.55748, -11.46456, -11.36934, -11.27192, -11.1724, -11.07087, 
    -10.96744, -10.86218, -10.75519, -10.64656, -10.53637, -10.42472, 
    -10.31169, -10.19736, -10.0818, -9.965097, -9.847324, -9.728554, 
    -9.608856, -9.488298, -9.366945, -9.244861,
  -8.505425, -8.618052, -8.730017, -8.84126, -8.951721, -9.061338, -9.170046, 
    -9.277779, -9.384465, -9.490034, -9.594414, -9.697527, -9.799295, 
    -9.899641, -9.998483, -10.09574, -10.19132, -10.28514, -10.37712, 
    -10.46716, -10.55519, -10.6411, -10.72481, -10.80623, -10.88527, 
    -10.96183, -11.03584, -11.10719, -11.17581, -11.2416, -11.30449, 
    -11.3644, -11.42123, -11.47492, -11.52539, -11.57257, -11.6164, 
    -11.65681, -11.69374, -11.72714, -11.75696, -11.78315, -11.80567, 
    -11.8245, -11.83959, -11.85093, -11.8585, -11.86229, -11.86229, -11.8585, 
    -11.85093, -11.83959, -11.8245, -11.80567, -11.78315, -11.75696, 
    -11.72714, -11.69374, -11.65681, -11.6164, -11.57257, -11.52539, 
    -11.47492, -11.42123, -11.3644, -11.30449, -11.2416, -11.17581, 
    -11.10719, -11.03584, -10.96183, -10.88527, -10.80623, -10.72481, 
    -10.6411, -10.55519, -10.46716, -10.37712, -10.28514, -10.19132, 
    -10.09574, -9.998483, -9.899641, -9.799295, -9.697527, -9.594414, 
    -9.490034, -9.384465, -9.277779, -9.170046, -9.061338, -8.951721, 
    -8.84126, -8.730017, -8.618052, -8.505425,
  -7.765951, -7.869044, -7.971541, -8.073387, -8.174527, -8.274905, -8.37446, 
    -8.473132, -8.570855, -8.667565, -8.763195, -8.857674, -8.95093, 
    -9.042892, -9.133484, -9.222629, -9.31025, -9.396269, -9.480604, 
    -9.563174, -9.643898, -9.722692, -9.799476, -9.874163, -9.946671, 
    -10.01692, -10.08482, -10.1503, -10.21327, -10.27365, -10.33138, 
    -10.38636, -10.43853, -10.48782, -10.53416, -10.57748, -10.61772, 
    -10.65482, -10.68873, -10.7194, -10.74679, -10.77084, -10.79152, 
    -10.80881, -10.82268, -10.83309, -10.84004, -10.84352, -10.84352, 
    -10.84004, -10.83309, -10.82268, -10.80881, -10.79152, -10.77084, 
    -10.74679, -10.7194, -10.68873, -10.65482, -10.61772, -10.57748, 
    -10.53416, -10.48782, -10.43853, -10.38636, -10.33138, -10.27365, 
    -10.21327, -10.1503, -10.08482, -10.01692, -9.946671, -9.874163, 
    -9.799476, -9.722692, -9.643898, -9.563174, -9.480604, -9.396269, 
    -9.31025, -9.222629, -9.133484, -9.042892, -8.95093, -8.857674, 
    -8.763195, -8.667565, -8.570855, -8.473132, -8.37446, -8.274905, 
    -8.174527, -8.073387, -7.971541, -7.869044, -7.765951,
  -7.026442, -7.119931, -7.212887, -7.305261, -7.397004, -7.488063, 
    -7.578384, -7.667912, -7.756588, -7.844352, -7.931143, -8.016898, 
    -8.101551, -8.185037, -8.267286, -8.34823, -8.427797, -8.505915, 
    -8.582511, -8.657512, -8.730841, -8.802423, -8.872184, -8.940046, 
    -9.005934, -9.069772, -9.131484, -9.190996, -9.248235, -9.303126, 
    -9.355601, -9.40559, -9.453025, -9.49784, -9.539974, -9.579368, 
    -9.615962, -9.649706, -9.680549, -9.708443, -9.733348, -9.755226, 
    -9.774042, -9.789767, -9.802377, -9.811852, -9.818177, -9.821342, 
    -9.821342, -9.818177, -9.811852, -9.802377, -9.789767, -9.774042, 
    -9.755226, -9.733348, -9.708443, -9.680549, -9.649706, -9.615962, 
    -9.579368, -9.539974, -9.49784, -9.453025, -9.40559, -9.355601, 
    -9.303126, -9.248235, -9.190996, -9.131484, -9.069772, -9.005934, 
    -8.940046, -8.872184, -8.802423, -8.730841, -8.657512, -8.582511, 
    -8.505915, -8.427797, -8.34823, -8.267286, -8.185037, -8.101551, 
    -8.016898, -7.931143, -7.844352, -7.756588, -7.667912, -7.578384, 
    -7.488063, -7.397004, -7.305261, -7.212887, -7.119931, -7.026442,
  -6.286901, -6.370722, -6.454072, -6.536906, -6.619181, -6.70085, -6.781863, 
    -6.862171, -6.941722, -7.020462, -7.098334, -7.175284, -7.251252, 
    -7.326178, -7.4, -7.472656, -7.544083, -7.614214, -7.682984, -7.750327, 
    -7.816175, -7.880459, -7.943112, -8.004064, -8.063247, -8.120593, 
    -8.176033, -8.229501, -8.280929, -8.330251, -8.377405, -8.422327, 
    -8.464956, -8.505234, -8.543103, -8.578511, -8.611405, -8.641738, 
    -8.669463, -8.69454, -8.716929, -8.736598, -8.753514, -8.767653, 
    -8.77899, -8.787509, -8.793196, -8.796041, -8.796041, -8.793196, 
    -8.787509, -8.77899, -8.767653, -8.753514, -8.736598, -8.716929, 
    -8.69454, -8.669463, -8.641738, -8.611405, -8.578511, -8.543103, 
    -8.505234, -8.464956, -8.422327, -8.377405, -8.330251, -8.280929, 
    -8.229501, -8.176033, -8.120593, -8.063247, -8.004064, -7.943112, 
    -7.880459, -7.816175, -7.750327, -7.682984, -7.614214, -7.544083, 
    -7.472656, -7.4, -7.326178, -7.251252, -7.175284, -7.098334, -7.020462, 
    -6.941722, -6.862171, -6.781863, -6.70085, -6.619181, -6.536906, 
    -6.454072, -6.370722, -6.286901,
  -5.547333, -5.621428, -5.695111, -5.768345, -5.84109, -5.913303, -5.984942, 
    -6.055964, -6.12632, -6.195964, -6.264847, -6.332918, -6.400125, 
    -6.466415, -6.531734, -6.596026, -6.659235, -6.721301, -6.782168, 
    -6.841775, -6.900063, -6.956971, -7.012438, -7.066403, -7.118805, 
    -7.169584, -7.218679, -7.266029, -7.311576, -7.355261, -7.397027, 
    -7.436818, -7.47458, -7.510261, -7.54381, -7.57518, -7.604323, -7.631198, 
    -7.655765, -7.677984, -7.697824, -7.715252, -7.730243, -7.742771, 
    -7.752818, -7.760367, -7.765407, -7.767929, -7.767929, -7.765407, 
    -7.760367, -7.752818, -7.742771, -7.730243, -7.715252, -7.697824, 
    -7.677984, -7.655765, -7.631198, -7.604323, -7.57518, -7.54381, 
    -7.510261, -7.47458, -7.436818, -7.397027, -7.355261, -7.311576, 
    -7.266029, -7.218679, -7.169584, -7.118805, -7.066403, -7.012438, 
    -6.956971, -6.900063, -6.841775, -6.782168, -6.721301, -6.659235, 
    -6.596026, -6.531734, -6.466415, -6.400125, -6.332918, -6.264847, 
    -6.195964, -6.12632, -6.055964, -5.984942, -5.913303, -5.84109, 
    -5.768345, -5.695111, -5.621428, -5.547333,
  -4.807739, -4.872057, -4.936023, -4.999602, -5.06276, -5.125462, -5.187668, 
    -5.249342, -5.310442, -5.370928, -5.430757, -5.489884, -5.548265, 
    -5.605854, -5.662601, -5.718461, -5.773382, -5.827315, -5.880208, 
    -5.93201, -5.982669, -6.032131, -6.080344, -6.127254, -6.172808, 
    -6.216953, -6.259636, -6.300805, -6.340407, -6.378393, -6.414712, 
    -6.449316, -6.482156, -6.513187, -6.542367, -6.56965, -6.594999, 
    -6.618376, -6.639744, -6.659072, -6.676331, -6.691492, -6.704533, 
    -6.715432, -6.724172, -6.73074, -6.735124, -6.737318, -6.737318, 
    -6.735124, -6.73074, -6.724172, -6.715432, -6.704533, -6.691492, 
    -6.676331, -6.659072, -6.639744, -6.618376, -6.594999, -6.56965, 
    -6.542367, -6.513187, -6.482156, -6.449316, -6.414712, -6.378393, 
    -6.340407, -6.300805, -6.259636, -6.216953, -6.172808, -6.127254, 
    -6.080344, -6.032131, -5.982669, -5.93201, -5.880208, -5.827315, 
    -5.773382, -5.718461, -5.662601, -5.605854, -5.548265, -5.489884, 
    -5.430757, -5.370928, -5.310442, -5.249342, -5.187668, -5.125462, 
    -5.06276, -4.999602, -4.936023, -4.872057, -4.807739,
  -4.068124, -4.122622, -4.176824, -4.230701, -4.284225, -4.337364, 
    -4.390087, -4.442361, -4.494153, -4.545426, -4.596145, -4.646272, 
    -4.695769, -4.744597, -4.792715, -4.840082, -4.886656, -4.932395, 
    -4.977254, -5.02119, -5.064158, -5.106114, -5.147013, -5.186808, 
    -5.225454, -5.262908, -5.299122, -5.334054, -5.367657, -5.399891, 
    -5.430711, -5.460076, -5.487947, -5.514283, -5.539048, -5.562205, 
    -5.58372, -5.603562, -5.6217, -5.638107, -5.652757, -5.665627, -5.676696, 
    -5.685948, -5.693368, -5.698944, -5.702665, -5.704528, -5.704528, 
    -5.702665, -5.698944, -5.693368, -5.685948, -5.676696, -5.665627, 
    -5.652757, -5.638107, -5.6217, -5.603562, -5.58372, -5.562205, -5.539048, 
    -5.514283, -5.487947, -5.460076, -5.430711, -5.399891, -5.367657, 
    -5.334054, -5.299122, -5.262908, -5.225454, -5.186808, -5.147013, 
    -5.106114, -5.064158, -5.02119, -4.977254, -4.932395, -4.886656, 
    -4.840082, -4.792715, -4.744597, -4.695769, -4.646272, -4.596145, 
    -4.545426, -4.494153, -4.442361, -4.390087, -4.337364, -4.284225, 
    -4.230701, -4.176824, -4.122622, -4.068124,
  -3.32849, -3.37313, -3.41753, -3.461666, -3.505514, -3.549049, -3.592245, 
    -3.635076, -3.677513, -3.719527, -3.761089, -3.802168, -3.842732, 
    -3.88275, -3.922188, -3.961012, -3.999188, -4.036681, -4.073455, 
    -4.109474, -4.144701, -4.179099, -4.212631, -4.245261, -4.27695, 
    -4.307662, -4.337358, -4.366004, -4.393563, -4.419998, -4.445276, 
    -4.46936, -4.49222, -4.513822, -4.534135, -4.55313, -4.570779, -4.587056, 
    -4.601935, -4.615394, -4.627412, -4.63797, -4.647052, -4.654643, 
    -4.660729, -4.665304, -4.668357, -4.669885, -4.669885, -4.668357, 
    -4.665304, -4.660729, -4.654643, -4.647052, -4.63797, -4.627412, 
    -4.615394, -4.601935, -4.587056, -4.570779, -4.55313, -4.534135, 
    -4.513822, -4.49222, -4.46936, -4.445276, -4.419998, -4.393563, 
    -4.366004, -4.337358, -4.307662, -4.27695, -4.245261, -4.212631, 
    -4.179099, -4.144701, -4.109474, -4.073455, -4.036681, -3.999188, 
    -3.961012, -3.922188, -3.88275, -3.842732, -3.802168, -3.761089, 
    -3.719527, -3.677513, -3.635076, -3.592245, -3.549049, -3.505514, 
    -3.461666, -3.41753, -3.37313, -3.32849,
  -2.588841, -2.623593, -2.658159, -2.692521, -2.72666, -2.760556, -2.79419, 
    -2.827541, -2.860586, -2.893303, -2.925669, -2.957661, -2.989253, 
    -3.02042, -3.051136, -3.081377, -3.111113, -3.140318, -3.168964, 
    -3.197022, -3.224465, -3.251263, -3.277388, -3.30281, -3.3275, -3.35143, 
    -3.374569, -3.39689, -3.418365, -3.438965, -3.458663, -3.477432, 
    -3.495247, -3.512082, -3.527913, -3.542717, -3.556473, -3.569159, 
    -3.580756, -3.591246, -3.600614, -3.608843, -3.615922, -3.621838, 
    -3.626583, -3.630148, -3.632529, -3.63372, -3.63372, -3.632529, 
    -3.630148, -3.626583, -3.621838, -3.615922, -3.608843, -3.600614, 
    -3.591246, -3.580756, -3.569159, -3.556473, -3.542717, -3.527913, 
    -3.512082, -3.495247, -3.477432, -3.458663, -3.438965, -3.418365, 
    -3.39689, -3.374569, -3.35143, -3.3275, -3.30281, -3.277388, -3.251263, 
    -3.224465, -3.197022, -3.168964, -3.140318, -3.111113, -3.081377, 
    -3.051136, -3.02042, -2.989253, -2.957661, -2.925669, -2.893303, 
    -2.860586, -2.827541, -2.79419, -2.760556, -2.72666, -2.692521, 
    -2.658159, -2.623593, -2.588841,
  -1.849181, -1.87402, -1.898728, -1.92329, -1.947694, -1.971925, -1.995969, 
    -2.019811, -2.043435, -2.066826, -2.089966, -2.112839, -2.135427, 
    -2.157712, -2.179676, -2.201299, -2.222563, -2.243447, -2.263932, 
    -2.283998, -2.303623, -2.322789, -2.341473, -2.359655, -2.377314, 
    -2.394429, -2.41098, -2.426945, -2.442306, -2.457041, -2.471131, 
    -2.484558, -2.497301, -2.509345, -2.52067, -2.53126, -2.541101, 
    -2.550177, -2.558473, -2.565979, -2.57268, -2.578568, -2.583632, 
    -2.587865, -2.59126, -2.593811, -2.595514, -2.596366, -2.596366, 
    -2.595514, -2.593811, -2.59126, -2.587865, -2.583632, -2.578568, 
    -2.57268, -2.565979, -2.558473, -2.550177, -2.541101, -2.53126, -2.52067, 
    -2.509345, -2.497301, -2.484558, -2.471131, -2.457041, -2.442306, 
    -2.426945, -2.41098, -2.394429, -2.377314, -2.359655, -2.341473, 
    -2.322789, -2.303623, -2.283998, -2.263932, -2.243447, -2.222563, 
    -2.201299, -2.179676, -2.157712, -2.135427, -2.112839, -2.089966, 
    -2.066826, -2.043435, -2.019811, -1.995969, -1.971925, -1.947694, 
    -1.92329, -1.898728, -1.87402, -1.849181,
  -1.109512, -1.124422, -1.139254, -1.153999, -1.168648, -1.183195, 
    -1.197629, -1.211942, -1.226125, -1.240168, -1.254061, -1.267794, 
    -1.281355, -1.294735, -1.307923, -1.320906, -1.333673, -1.346213, 
    -1.358514, -1.370563, -1.382348, -1.393856, -1.405076, -1.415995, 
    -1.4266, -1.436878, -1.446817, -1.456406, -1.46563, -1.47448, -1.482942, 
    -1.491006, -1.49866, -1.505893, -1.512695, -1.519056, -1.524966, 
    -1.530417, -1.535401, -1.539908, -1.543934, -1.54747, -1.550512, 
    -1.553055, -1.555094, -1.556626, -1.557649, -1.55816, -1.55816, 
    -1.557649, -1.556626, -1.555094, -1.553055, -1.550512, -1.54747, 
    -1.543934, -1.539908, -1.535401, -1.530417, -1.524966, -1.519056, 
    -1.512695, -1.505893, -1.49866, -1.491006, -1.482942, -1.47448, -1.46563, 
    -1.456406, -1.446817, -1.436878, -1.4266, -1.415995, -1.405076, 
    -1.393856, -1.382348, -1.370563, -1.358514, -1.346213, -1.333673, 
    -1.320906, -1.307923, -1.294735, -1.281355, -1.267794, -1.254061, 
    -1.240168, -1.226125, -1.211942, -1.197629, -1.183195, -1.168648, 
    -1.153999, -1.139254, -1.124422, -1.109512,
  -0.3698378, -0.3748092, -0.3797542, -0.3846703, -0.3895547, -0.3944048, 
    -0.3992176, -0.40399, -0.4087191, -0.4134014, -0.4180338, -0.4226128, 
    -0.4271349, -0.4315965, -0.4359938, -0.4403231, -0.4445804, -0.448762, 
    -0.4528638, -0.4568816, -0.4608116, -0.4646493, -0.4683909, -0.472032, 
    -0.4755684, -0.478996, -0.4823107, -0.4855082, -0.4885846, -0.4915359, 
    -0.494358, -0.4970472, -0.4995998, -0.502012, -0.5042805, -0.5064019, 
    -0.5083731, -0.510191, -0.511853, -0.5133564, -0.5146989, -0.5158784, 
    -0.5168929, -0.5177408, -0.5184209, -0.5189319, -0.519273, -0.5194437, 
    -0.5194437, -0.519273, -0.5189319, -0.5184209, -0.5177408, -0.5168929, 
    -0.5158784, -0.5146989, -0.5133564, -0.511853, -0.510191, -0.5083731, 
    -0.5064019, -0.5042805, -0.502012, -0.4995998, -0.4970472, -0.494358, 
    -0.4915359, -0.4885846, -0.4855082, -0.4823107, -0.478996, -0.4755684, 
    -0.472032, -0.4683909, -0.4646493, -0.4608116, -0.4568816, -0.4528638, 
    -0.448762, -0.4445804, -0.4403231, -0.4359938, -0.4315965, -0.4271349, 
    -0.4226128, -0.4180338, -0.4134014, -0.4087191, -0.40399, -0.3992176, 
    -0.3944048, -0.3895547, -0.3846703, -0.3797542, -0.3748092, -0.3698378,
  0.3698378, 0.3748092, 0.3797542, 0.3846703, 0.3895547, 0.3944048, 
    0.3992176, 0.40399, 0.4087191, 0.4134014, 0.4180338, 0.4226128, 
    0.4271349, 0.4315965, 0.4359938, 0.4403231, 0.4445804, 0.448762, 
    0.4528638, 0.4568816, 0.4608116, 0.4646493, 0.4683909, 0.472032, 
    0.4755684, 0.478996, 0.4823107, 0.4855082, 0.4885846, 0.4915359, 
    0.494358, 0.4970472, 0.4995998, 0.502012, 0.5042805, 0.5064019, 
    0.5083731, 0.510191, 0.511853, 0.5133564, 0.5146989, 0.5158784, 
    0.5168929, 0.5177408, 0.5184209, 0.5189319, 0.519273, 0.5194437, 
    0.5194437, 0.519273, 0.5189319, 0.5184209, 0.5177408, 0.5168929, 
    0.5158784, 0.5146989, 0.5133564, 0.511853, 0.510191, 0.5083731, 
    0.5064019, 0.5042805, 0.502012, 0.4995998, 0.4970472, 0.494358, 
    0.4915359, 0.4885846, 0.4855082, 0.4823107, 0.478996, 0.4755684, 
    0.472032, 0.4683909, 0.4646493, 0.4608116, 0.4568816, 0.4528638, 
    0.448762, 0.4445804, 0.4403231, 0.4359938, 0.4315965, 0.4271349, 
    0.4226128, 0.4180338, 0.4134014, 0.4087191, 0.40399, 0.3992176, 
    0.3944048, 0.3895547, 0.3846703, 0.3797542, 0.3748092, 0.3698378,
  1.109512, 1.124422, 1.139254, 1.153999, 1.168648, 1.183195, 1.197629, 
    1.211942, 1.226125, 1.240168, 1.254061, 1.267794, 1.281355, 1.294735, 
    1.307923, 1.320906, 1.333673, 1.346213, 1.358514, 1.370563, 1.382348, 
    1.393856, 1.405076, 1.415995, 1.4266, 1.436878, 1.446817, 1.456406, 
    1.46563, 1.47448, 1.482942, 1.491006, 1.49866, 1.505893, 1.512695, 
    1.519056, 1.524966, 1.530417, 1.535401, 1.539908, 1.543934, 1.54747, 
    1.550512, 1.553055, 1.555094, 1.556626, 1.557649, 1.55816, 1.55816, 
    1.557649, 1.556626, 1.555094, 1.553055, 1.550512, 1.54747, 1.543934, 
    1.539908, 1.535401, 1.530417, 1.524966, 1.519056, 1.512695, 1.505893, 
    1.49866, 1.491006, 1.482942, 1.47448, 1.46563, 1.456406, 1.446817, 
    1.436878, 1.4266, 1.415995, 1.405076, 1.393856, 1.382348, 1.370563, 
    1.358514, 1.346213, 1.333673, 1.320906, 1.307923, 1.294735, 1.281355, 
    1.267794, 1.254061, 1.240168, 1.226125, 1.211942, 1.197629, 1.183195, 
    1.168648, 1.153999, 1.139254, 1.124422, 1.109512,
  1.849181, 1.87402, 1.898728, 1.92329, 1.947694, 1.971925, 1.995969, 
    2.019811, 2.043435, 2.066826, 2.089966, 2.112839, 2.135427, 2.157712, 
    2.179676, 2.201299, 2.222563, 2.243447, 2.263932, 2.283998, 2.303623, 
    2.322789, 2.341473, 2.359655, 2.377314, 2.394429, 2.41098, 2.426945, 
    2.442306, 2.457041, 2.471131, 2.484558, 2.497301, 2.509345, 2.52067, 
    2.53126, 2.541101, 2.550177, 2.558473, 2.565979, 2.57268, 2.578568, 
    2.583632, 2.587865, 2.59126, 2.593811, 2.595514, 2.596366, 2.596366, 
    2.595514, 2.593811, 2.59126, 2.587865, 2.583632, 2.578568, 2.57268, 
    2.565979, 2.558473, 2.550177, 2.541101, 2.53126, 2.52067, 2.509345, 
    2.497301, 2.484558, 2.471131, 2.457041, 2.442306, 2.426945, 2.41098, 
    2.394429, 2.377314, 2.359655, 2.341473, 2.322789, 2.303623, 2.283998, 
    2.263932, 2.243447, 2.222563, 2.201299, 2.179676, 2.157712, 2.135427, 
    2.112839, 2.089966, 2.066826, 2.043435, 2.019811, 1.995969, 1.971925, 
    1.947694, 1.92329, 1.898728, 1.87402, 1.849181,
  2.588841, 2.623593, 2.658159, 2.692521, 2.72666, 2.760556, 2.79419, 
    2.827541, 2.860586, 2.893303, 2.925669, 2.957661, 2.989253, 3.02042, 
    3.051136, 3.081377, 3.111113, 3.140318, 3.168964, 3.197022, 3.224465, 
    3.251263, 3.277388, 3.30281, 3.3275, 3.35143, 3.374569, 3.39689, 
    3.418365, 3.438965, 3.458663, 3.477432, 3.495247, 3.512082, 3.527913, 
    3.542717, 3.556473, 3.569159, 3.580756, 3.591246, 3.600614, 3.608843, 
    3.615922, 3.621838, 3.626583, 3.630148, 3.632529, 3.63372, 3.63372, 
    3.632529, 3.630148, 3.626583, 3.621838, 3.615922, 3.608843, 3.600614, 
    3.591246, 3.580756, 3.569159, 3.556473, 3.542717, 3.527913, 3.512082, 
    3.495247, 3.477432, 3.458663, 3.438965, 3.418365, 3.39689, 3.374569, 
    3.35143, 3.3275, 3.30281, 3.277388, 3.251263, 3.224465, 3.197022, 
    3.168964, 3.140318, 3.111113, 3.081377, 3.051136, 3.02042, 2.989253, 
    2.957661, 2.925669, 2.893303, 2.860586, 2.827541, 2.79419, 2.760556, 
    2.72666, 2.692521, 2.658159, 2.623593, 2.588841,
  3.32849, 3.37313, 3.41753, 3.461666, 3.505514, 3.549049, 3.592245, 
    3.635076, 3.677513, 3.719527, 3.761089, 3.802168, 3.842732, 3.88275, 
    3.922188, 3.961012, 3.999188, 4.036681, 4.073455, 4.109474, 4.144701, 
    4.179099, 4.212631, 4.245261, 4.27695, 4.307662, 4.337358, 4.366004, 
    4.393563, 4.419998, 4.445276, 4.46936, 4.49222, 4.513822, 4.534135, 
    4.55313, 4.570779, 4.587056, 4.601935, 4.615394, 4.627412, 4.63797, 
    4.647052, 4.654643, 4.660729, 4.665304, 4.668357, 4.669885, 4.669885, 
    4.668357, 4.665304, 4.660729, 4.654643, 4.647052, 4.63797, 4.627412, 
    4.615394, 4.601935, 4.587056, 4.570779, 4.55313, 4.534135, 4.513822, 
    4.49222, 4.46936, 4.445276, 4.419998, 4.393563, 4.366004, 4.337358, 
    4.307662, 4.27695, 4.245261, 4.212631, 4.179099, 4.144701, 4.109474, 
    4.073455, 4.036681, 3.999188, 3.961012, 3.922188, 3.88275, 3.842732, 
    3.802168, 3.761089, 3.719527, 3.677513, 3.635076, 3.592245, 3.549049, 
    3.505514, 3.461666, 3.41753, 3.37313, 3.32849,
  4.068124, 4.122622, 4.176824, 4.230701, 4.284225, 4.337364, 4.390087, 
    4.442361, 4.494153, 4.545426, 4.596145, 4.646272, 4.695769, 4.744597, 
    4.792715, 4.840082, 4.886656, 4.932395, 4.977254, 5.02119, 5.064158, 
    5.106114, 5.147013, 5.186808, 5.225454, 5.262908, 5.299122, 5.334054, 
    5.367657, 5.399891, 5.430711, 5.460076, 5.487947, 5.514283, 5.539048, 
    5.562205, 5.58372, 5.603562, 5.6217, 5.638107, 5.652757, 5.665627, 
    5.676696, 5.685948, 5.693368, 5.698944, 5.702665, 5.704528, 5.704528, 
    5.702665, 5.698944, 5.693368, 5.685948, 5.676696, 5.665627, 5.652757, 
    5.638107, 5.6217, 5.603562, 5.58372, 5.562205, 5.539048, 5.514283, 
    5.487947, 5.460076, 5.430711, 5.399891, 5.367657, 5.334054, 5.299122, 
    5.262908, 5.225454, 5.186808, 5.147013, 5.106114, 5.064158, 5.02119, 
    4.977254, 4.932395, 4.886656, 4.840082, 4.792715, 4.744597, 4.695769, 
    4.646272, 4.596145, 4.545426, 4.494153, 4.442361, 4.390087, 4.337364, 
    4.284225, 4.230701, 4.176824, 4.122622, 4.068124,
  4.807739, 4.872057, 4.936023, 4.999602, 5.06276, 5.125462, 5.187668, 
    5.249342, 5.310442, 5.370928, 5.430757, 5.489884, 5.548265, 5.605854, 
    5.662601, 5.718461, 5.773382, 5.827315, 5.880208, 5.93201, 5.982669, 
    6.032131, 6.080344, 6.127254, 6.172808, 6.216953, 6.259636, 6.300805, 
    6.340407, 6.378393, 6.414712, 6.449316, 6.482156, 6.513187, 6.542367, 
    6.56965, 6.594999, 6.618376, 6.639744, 6.659072, 6.676331, 6.691492, 
    6.704533, 6.715432, 6.724172, 6.73074, 6.735124, 6.737318, 6.737318, 
    6.735124, 6.73074, 6.724172, 6.715432, 6.704533, 6.691492, 6.676331, 
    6.659072, 6.639744, 6.618376, 6.594999, 6.56965, 6.542367, 6.513187, 
    6.482156, 6.449316, 6.414712, 6.378393, 6.340407, 6.300805, 6.259636, 
    6.216953, 6.172808, 6.127254, 6.080344, 6.032131, 5.982669, 5.93201, 
    5.880208, 5.827315, 5.773382, 5.718461, 5.662601, 5.605854, 5.548265, 
    5.489884, 5.430757, 5.370928, 5.310442, 5.249342, 5.187668, 5.125462, 
    5.06276, 4.999602, 4.936023, 4.872057, 4.807739,
  5.547333, 5.621428, 5.695111, 5.768345, 5.84109, 5.913303, 5.984942, 
    6.055964, 6.12632, 6.195964, 6.264847, 6.332918, 6.400125, 6.466415, 
    6.531734, 6.596026, 6.659235, 6.721301, 6.782168, 6.841775, 6.900063, 
    6.956971, 7.012438, 7.066403, 7.118805, 7.169584, 7.218679, 7.266029, 
    7.311576, 7.355261, 7.397027, 7.436818, 7.47458, 7.510261, 7.54381, 
    7.57518, 7.604323, 7.631198, 7.655765, 7.677984, 7.697824, 7.715252, 
    7.730243, 7.742771, 7.752818, 7.760367, 7.765407, 7.767929, 7.767929, 
    7.765407, 7.760367, 7.752818, 7.742771, 7.730243, 7.715252, 7.697824, 
    7.677984, 7.655765, 7.631198, 7.604323, 7.57518, 7.54381, 7.510261, 
    7.47458, 7.436818, 7.397027, 7.355261, 7.311576, 7.266029, 7.218679, 
    7.169584, 7.118805, 7.066403, 7.012438, 6.956971, 6.900063, 6.841775, 
    6.782168, 6.721301, 6.659235, 6.596026, 6.531734, 6.466415, 6.400125, 
    6.332918, 6.264847, 6.195964, 6.12632, 6.055964, 5.984942, 5.913303, 
    5.84109, 5.768345, 5.695111, 5.621428, 5.547333,
  6.286901, 6.370722, 6.454072, 6.536906, 6.619181, 6.70085, 6.781863, 
    6.862171, 6.941722, 7.020462, 7.098334, 7.175284, 7.251252, 7.326178, 
    7.4, 7.472656, 7.544083, 7.614214, 7.682984, 7.750327, 7.816175, 
    7.880459, 7.943112, 8.004064, 8.063247, 8.120593, 8.176033, 8.229501, 
    8.280929, 8.330251, 8.377405, 8.422327, 8.464956, 8.505234, 8.543103, 
    8.578511, 8.611405, 8.641738, 8.669463, 8.69454, 8.716929, 8.736598, 
    8.753514, 8.767653, 8.77899, 8.787509, 8.793196, 8.796041, 8.796041, 
    8.793196, 8.787509, 8.77899, 8.767653, 8.753514, 8.736598, 8.716929, 
    8.69454, 8.669463, 8.641738, 8.611405, 8.578511, 8.543103, 8.505234, 
    8.464956, 8.422327, 8.377405, 8.330251, 8.280929, 8.229501, 8.176033, 
    8.120593, 8.063247, 8.004064, 7.943112, 7.880459, 7.816175, 7.750327, 
    7.682984, 7.614214, 7.544083, 7.472656, 7.4, 7.326178, 7.251252, 
    7.175284, 7.098334, 7.020462, 6.941722, 6.862171, 6.781863, 6.70085, 
    6.619181, 6.536906, 6.454072, 6.370722, 6.286901,
  7.026442, 7.119931, 7.212887, 7.305261, 7.397004, 7.488063, 7.578384, 
    7.667912, 7.756588, 7.844352, 7.931143, 8.016898, 8.101551, 8.185037, 
    8.267286, 8.34823, 8.427797, 8.505915, 8.582511, 8.657512, 8.730841, 
    8.802423, 8.872184, 8.940046, 9.005934, 9.069772, 9.131484, 9.190996, 
    9.248235, 9.303126, 9.355601, 9.40559, 9.453025, 9.49784, 9.539974, 
    9.579368, 9.615962, 9.649706, 9.680549, 9.708443, 9.733348, 9.755226, 
    9.774042, 9.789767, 9.802377, 9.811852, 9.818177, 9.821342, 9.821342, 
    9.818177, 9.811852, 9.802377, 9.789767, 9.774042, 9.755226, 9.733348, 
    9.708443, 9.680549, 9.649706, 9.615962, 9.579368, 9.539974, 9.49784, 
    9.453025, 9.40559, 9.355601, 9.303126, 9.248235, 9.190996, 9.131484, 
    9.069772, 9.005934, 8.940046, 8.872184, 8.802423, 8.730841, 8.657512, 
    8.582511, 8.505915, 8.427797, 8.34823, 8.267286, 8.185037, 8.101551, 
    8.016898, 7.931143, 7.844352, 7.756588, 7.667912, 7.578384, 7.488063, 
    7.397004, 7.305261, 7.212887, 7.119931, 7.026442,
  7.765951, 7.869044, 7.971541, 8.073387, 8.174527, 8.274905, 8.37446, 
    8.473132, 8.570855, 8.667565, 8.763195, 8.857674, 8.95093, 9.042892, 
    9.133484, 9.222629, 9.31025, 9.396269, 9.480604, 9.563174, 9.643898, 
    9.722692, 9.799476, 9.874163, 9.946671, 10.01692, 10.08482, 10.1503, 
    10.21327, 10.27365, 10.33138, 10.38636, 10.43853, 10.48782, 10.53416, 
    10.57748, 10.61772, 10.65482, 10.68873, 10.7194, 10.74679, 10.77084, 
    10.79152, 10.80881, 10.82268, 10.83309, 10.84004, 10.84352, 10.84352, 
    10.84004, 10.83309, 10.82268, 10.80881, 10.79152, 10.77084, 10.74679, 
    10.7194, 10.68873, 10.65482, 10.61772, 10.57748, 10.53416, 10.48782, 
    10.43853, 10.38636, 10.33138, 10.27365, 10.21327, 10.1503, 10.08482, 
    10.01692, 9.946671, 9.874163, 9.799476, 9.722692, 9.643898, 9.563174, 
    9.480604, 9.396269, 9.31025, 9.222629, 9.133484, 9.042892, 8.95093, 
    8.857674, 8.763195, 8.667565, 8.570855, 8.473132, 8.37446, 8.274905, 
    8.174527, 8.073387, 7.971541, 7.869044, 7.765951,
  8.505425, 8.618052, 8.730017, 8.84126, 8.951721, 9.061338, 9.170046, 
    9.277779, 9.384465, 9.490034, 9.594414, 9.697527, 9.799295, 9.899641, 
    9.998483, 10.09574, 10.19132, 10.28514, 10.37712, 10.46716, 10.55519, 
    10.6411, 10.72481, 10.80623, 10.88527, 10.96183, 11.03584, 11.10719, 
    11.17581, 11.2416, 11.30449, 11.3644, 11.42123, 11.47492, 11.52539, 
    11.57257, 11.6164, 11.65681, 11.69374, 11.72714, 11.75696, 11.78315, 
    11.80567, 11.8245, 11.83959, 11.85093, 11.8585, 11.86229, 11.86229, 
    11.8585, 11.85093, 11.83959, 11.8245, 11.80567, 11.78315, 11.75696, 
    11.72714, 11.69374, 11.65681, 11.6164, 11.57257, 11.52539, 11.47492, 
    11.42123, 11.3644, 11.30449, 11.2416, 11.17581, 11.10719, 11.03584, 
    10.96183, 10.88527, 10.80623, 10.72481, 10.6411, 10.55519, 10.46716, 
    10.37712, 10.28514, 10.19132, 10.09574, 9.998483, 9.899641, 9.799295, 
    9.697527, 9.594414, 9.490034, 9.384465, 9.277779, 9.170046, 9.061338, 
    8.951721, 8.84126, 8.730017, 8.618052, 8.505425,
  9.244861, 9.366945, 9.488298, 9.608856, 9.728554, 9.847324, 9.965097, 
    10.0818, 10.19736, 10.31169, 10.42472, 10.53637, 10.64656, 10.75519, 
    10.86218, 10.96744, 11.07087, 11.1724, 11.27192, 11.36934, 11.46456, 
    11.55748, 11.64802, 11.73607, 11.82154, 11.90432, 11.98433, 12.06147, 
    12.13564, 12.20676, 12.27472, 12.33946, 12.40088, 12.45889, 12.51342, 
    12.5644, 12.61175, 12.6554, 12.6953, 12.73137, 12.76358, 12.79187, 
    12.8162, 12.83653, 12.85283, 12.86508, 12.87325, 12.87735, 12.87735, 
    12.87325, 12.86508, 12.85283, 12.83653, 12.8162, 12.79187, 12.76358, 
    12.73137, 12.6953, 12.6554, 12.61175, 12.5644, 12.51342, 12.45889, 
    12.40088, 12.33946, 12.27472, 12.20676, 12.13564, 12.06147, 11.98433, 
    11.90432, 11.82154, 11.73607, 11.64802, 11.55748, 11.46456, 11.36934, 
    11.27192, 11.1724, 11.07087, 10.96744, 10.86218, 10.75519, 10.64656, 
    10.53637, 10.42472, 10.31169, 10.19736, 10.0818, 9.965097, 9.847324, 
    9.728554, 9.608856, 9.488298, 9.366945, 9.244861,
  9.984256, 10.11571, 10.24637, 10.37615, 10.505, 10.63283, 10.75957, 
    10.88514, 11.00947, 11.13247, 11.25405, 11.37413, 11.49262, 11.60943, 
    11.72446, 11.83762, 11.9488, 12.05792, 12.16487, 12.26954, 12.37185, 
    12.47168, 12.56893, 12.66351, 12.75529, 12.84419, 12.9301, 13.01292, 
    13.09255, 13.16889, 13.24185, 13.31133, 13.37724, 13.43949, 13.49801, 
    13.55271, 13.60351, 13.65034, 13.69314, 13.73184, 13.76639, 13.79673, 
    13.82283, 13.84463, 13.86212, 13.87526, 13.88403, 13.88841, 13.88841, 
    13.88403, 13.87526, 13.86212, 13.84463, 13.82283, 13.79673, 13.76639, 
    13.73184, 13.69314, 13.65034, 13.60351, 13.55271, 13.49801, 13.43949, 
    13.37724, 13.31133, 13.24185, 13.16889, 13.09255, 13.01292, 12.9301, 
    12.84419, 12.75529, 12.66351, 12.56893, 12.47168, 12.37185, 12.26954, 
    12.16487, 12.05792, 11.9488, 11.83762, 11.72446, 11.60943, 11.49262, 
    11.37413, 11.25405, 11.13247, 11.00947, 10.88514, 10.75957, 10.63283, 
    10.505, 10.37615, 10.24637, 10.11571, 9.984256,
  10.72361, 10.86435, 11.00421, 11.14313, 11.28102, 11.41781, 11.55342, 
    11.68776, 11.82075, 11.9523, 12.08233, 12.21073, 12.33741, 12.46228, 
    12.58523, 12.70616, 12.82498, 12.94157, 13.05583, 13.16765, 13.27692, 
    13.38354, 13.48739, 13.58837, 13.68636, 13.78126, 13.87296, 13.96135, 
    14.04633, 14.1278, 14.20564, 14.27977, 14.35008, 14.4165, 14.47891, 
    14.53725, 14.59143, 14.64138, 14.68701, 14.72828, 14.76512, 14.79747, 
    14.8253, 14.84855, 14.86719, 14.88119, 14.89054, 14.89522, 14.89522, 
    14.89054, 14.88119, 14.86719, 14.84855, 14.8253, 14.79747, 14.76512, 
    14.72828, 14.68701, 14.64138, 14.59143, 14.53725, 14.47891, 14.4165, 
    14.35008, 14.27977, 14.20564, 14.1278, 14.04633, 13.96135, 13.87296, 
    13.78126, 13.68636, 13.58837, 13.48739, 13.38354, 13.27692, 13.16765, 
    13.05583, 12.94157, 12.82498, 12.70616, 12.58523, 12.46228, 12.33741, 
    12.21073, 12.08233, 11.9523, 11.82075, 11.68776, 11.55342, 11.41781, 
    11.28102, 11.14313, 11.00421, 10.86435, 10.72361,
  11.46291, 11.61284, 11.76182, 11.90976, 12.05659, 12.20224, 12.3466, 
    12.4896, 12.63114, 12.77113, 12.90947, 13.04607, 13.18083, 13.31363, 
    13.44438, 13.57297, 13.69929, 13.82323, 13.94467, 14.0635, 14.17962, 
    14.2929, 14.40323, 14.51049, 14.61457, 14.71535, 14.81272, 14.90658, 
    14.99679, 15.08327, 15.1659, 15.24457, 15.3192, 15.38967, 15.4559, 
    15.5178, 15.57528, 15.62826, 15.67667, 15.72045, 15.75952, 15.79384, 
    15.82335, 15.84801, 15.86777, 15.88263, 15.89254, 15.8975, 15.8975, 
    15.89254, 15.88263, 15.86777, 15.84801, 15.82335, 15.79384, 15.75952, 
    15.72045, 15.67667, 15.62826, 15.57528, 15.5178, 15.4559, 15.38967, 
    15.3192, 15.24457, 15.1659, 15.08327, 14.99679, 14.90658, 14.81272, 
    14.71535, 14.61457, 14.51049, 14.40323, 14.2929, 14.17962, 14.0635, 
    13.94467, 13.82323, 13.69929, 13.57297, 13.44438, 13.31363, 13.18083, 
    13.04607, 12.90947, 12.77113, 12.63114, 12.4896, 12.3466, 12.20224, 
    12.05659, 11.90976, 11.76182, 11.61284, 11.46291,
  12.20216, 12.36118, 12.51916, 12.67602, 12.83169, 12.98607, 13.13908, 
    13.29061, 13.44058, 13.58888, 13.73542, 13.88009, 14.02279, 14.1634, 
    14.30182, 14.43793, 14.57162, 14.70277, 14.83126, 14.95698, 15.07981, 
    15.19962, 15.31629, 15.42971, 15.53974, 15.64629, 15.74921, 15.8484, 
    15.94374, 16.03511, 16.12242, 16.20553, 16.28436, 16.3588, 16.42875, 
    16.49412, 16.55482, 16.61077, 16.66188, 16.7081, 16.74936, 16.78558, 
    16.81673, 16.84276, 16.86363, 16.87931, 16.88978, 16.89501, 16.89501, 
    16.88978, 16.87931, 16.86363, 16.84276, 16.81673, 16.78558, 16.74936, 
    16.7081, 16.66188, 16.61077, 16.55482, 16.49412, 16.42875, 16.3588, 
    16.28436, 16.20553, 16.12242, 16.03511, 15.94374, 15.8484, 15.74921, 
    15.64629, 15.53974, 15.42971, 15.31629, 15.19962, 15.07981, 14.95698, 
    14.83126, 14.70277, 14.57162, 14.43793, 14.30182, 14.1634, 14.02279, 
    13.88009, 13.73542, 13.58888, 13.44058, 13.29061, 13.13908, 12.98607, 
    12.83169, 12.67602, 12.51916, 12.36118, 12.20216,
  12.94136, 13.10935, 13.27623, 13.4419, 13.60628, 13.76928, 13.9308, 
    14.09074, 14.24901, 14.4055, 14.56011, 14.71272, 14.86322, 15.0115, 
    15.15745, 15.30094, 15.44186, 15.58009, 15.71549, 15.84795, 15.97735, 
    16.10355, 16.22643, 16.34587, 16.46173, 16.57389, 16.68224, 16.78664, 
    16.88698, 16.98314, 17.075, 17.16244, 17.24537, 17.32367, 17.39725, 
    17.466, 17.52983, 17.58866, 17.64242, 17.69101, 17.73438, 17.77247, 
    17.80522, 17.83258, 17.85452, 17.871, 17.882, 17.88751, 17.88751, 17.882, 
    17.871, 17.85452, 17.83258, 17.80522, 17.77247, 17.73438, 17.69101, 
    17.64242, 17.58866, 17.52983, 17.466, 17.39725, 17.32367, 17.24537, 
    17.16244, 17.075, 16.98314, 16.88698, 16.78664, 16.68224, 16.57389, 
    16.46173, 16.34587, 16.22643, 16.10355, 15.97735, 15.84795, 15.71549, 
    15.58009, 15.44186, 15.30094, 15.15745, 15.0115, 14.86322, 14.71272, 
    14.56011, 14.4055, 14.24901, 14.09074, 13.9308, 13.76928, 13.60628, 
    13.4419, 13.27623, 13.10935, 12.94136,
  13.6805, 13.85736, 14.03301, 14.20737, 14.38034, 14.55183, 14.72173, 
    14.88996, 15.05639, 15.22093, 15.38346, 15.54386, 15.70203, 15.85784, 
    16.01117, 16.1619, 16.30991, 16.45506, 16.59723, 16.73629, 16.87211, 
    17.00456, 17.1335, 17.25882, 17.38036, 17.49802, 17.61165, 17.72114, 
    17.82635, 17.92716, 18.02345, 18.11512, 18.20203, 18.28409, 18.36119, 
    18.43323, 18.50011, 18.56174, 18.61805, 18.66896, 18.71439, 18.75428, 
    18.78858, 18.81724, 18.84021, 18.85747, 18.86899, 18.87476, 18.87476, 
    18.86899, 18.85747, 18.84021, 18.81724, 18.78858, 18.75428, 18.71439, 
    18.66896, 18.61805, 18.56174, 18.50011, 18.43323, 18.36119, 18.28409, 
    18.20203, 18.11512, 18.02345, 17.92716, 17.82635, 17.72114, 17.61165, 
    17.49802, 17.38036, 17.25882, 17.1335, 17.00456, 16.87211, 16.73629, 
    16.59723, 16.45506, 16.30991, 16.1619, 16.01117, 15.85784, 15.70203, 
    15.54386, 15.38346, 15.22093, 15.05639, 14.88996, 14.72173, 14.55183, 
    14.38034, 14.20737, 14.03301, 13.85736, 13.6805,
  14.41959, 14.60518, 14.78949, 14.9724, 15.15383, 15.33368, 15.51184, 
    15.6882, 15.86266, 16.0351, 16.20541, 16.37346, 16.53915, 16.70233, 
    16.8629, 17.02072, 17.17565, 17.32758, 17.47636, 17.62187, 17.76396, 
    17.9025, 18.03736, 18.16841, 18.2955, 18.4185, 18.53728, 18.65171, 
    18.76166, 18.867, 18.96761, 19.06337, 19.15416, 19.23986, 19.32038, 
    19.39561, 19.46544, 19.5298, 19.58859, 19.64173, 19.68916, 19.7308, 
    19.7666, 19.79651, 19.82049, 19.8385, 19.85053, 19.85655, 19.85655, 
    19.85053, 19.8385, 19.82049, 19.79651, 19.7666, 19.7308, 19.68916, 
    19.64173, 19.58859, 19.5298, 19.46544, 19.39561, 19.32038, 19.23986, 
    19.15416, 19.06337, 18.96761, 18.867, 18.76166, 18.65171, 18.53728, 
    18.4185, 18.2955, 18.16841, 18.03736, 17.9025, 17.76396, 17.62187, 
    17.47636, 17.32758, 17.17565, 17.02072, 16.8629, 16.70233, 16.53915, 
    16.37346, 16.20541, 16.0351, 15.86266, 15.6882, 15.51184, 15.33368, 
    15.15383, 14.9724, 14.78949, 14.60518, 14.41959,
  15.15861, 15.35282, 15.54564, 15.73699, 15.92674, 16.11481, 16.30107, 
    16.48543, 16.66776, 16.84796, 17.02589, 17.20144, 17.37449, 17.5449, 
    17.71254, 17.87728, 18.03899, 18.19754, 18.35277, 18.50457, 18.65277, 
    18.79726, 18.93789, 19.07451, 19.20699, 19.33519, 19.45897, 19.57821, 
    19.69276, 19.8025, 19.90729, 20.00702, 20.10156, 20.19081, 20.27464, 
    20.35295, 20.42565, 20.49264, 20.55383, 20.60913, 20.65849, 20.70182, 
    20.73908, 20.7702, 20.79515, 20.81389, 20.8264, 20.83266, 20.83266, 
    20.8264, 20.81389, 20.79515, 20.7702, 20.73908, 20.70182, 20.65849, 
    20.60913, 20.55383, 20.49264, 20.42565, 20.35295, 20.27464, 20.19081, 
    20.10156, 20.00702, 19.90729, 19.8025, 19.69276, 19.57821, 19.45897, 
    19.33519, 19.20699, 19.07451, 18.93789, 18.79726, 18.65277, 18.50457, 
    18.35277, 18.19754, 18.03899, 17.87728, 17.71254, 17.5449, 17.37449, 
    17.20144, 17.02589, 16.84796, 16.66776, 16.48543, 16.30107, 16.11481, 
    15.92674, 15.73699, 15.54564, 15.35282, 15.15861,
  15.89756, 16.10026, 16.30147, 16.50109, 16.69903, 16.89517, 17.0894, 
    17.2816, 17.47165, 17.65945, 17.84485, 18.02774, 18.20799, 18.38545, 
    18.56001, 18.73152, 18.89984, 19.06483, 19.22636, 19.38427, 19.53844, 
    19.68871, 19.83493, 19.97698, 20.11469, 20.24794, 20.37659, 20.50048, 
    20.61949, 20.73348, 20.84233, 20.94591, 21.04409, 21.13675, 21.22379, 
    21.30509, 21.38055, 21.45008, 21.51358, 21.57098, 21.6222, 21.66716, 
    21.70582, 21.73811, 21.764, 21.78345, 21.79643, 21.80292, 21.80292, 
    21.79643, 21.78345, 21.764, 21.73811, 21.70582, 21.66716, 21.6222, 
    21.57098, 21.51358, 21.45008, 21.38055, 21.30509, 21.22379, 21.13675, 
    21.04409, 20.94591, 20.84233, 20.73348, 20.61949, 20.50048, 20.37659, 
    20.24794, 20.11469, 19.97698, 19.83493, 19.68871, 19.53844, 19.38427, 
    19.22636, 19.06483, 18.89984, 18.73152, 18.56001, 18.38545, 18.20799, 
    18.02774, 17.84485, 17.65945, 17.47165, 17.2816, 17.0894, 16.89517, 
    16.69903, 16.50109, 16.30147, 16.10026, 15.89756,
  16.63645, 16.84749, 17.05695, 17.26471, 17.47068, 17.67474, 17.87678, 
    18.07666, 18.27429, 18.46952, 18.66223, 18.85229, 19.03956, 19.22392, 
    19.40522, 19.58332, 19.75808, 19.92936, 20.09701, 20.26088, 20.42083, 
    20.57672, 20.72838, 20.87569, 21.01848, 21.15662, 21.28997, 21.41838, 
    21.5417, 21.65982, 21.77258, 21.87987, 21.98156, 22.07753, 22.16766, 
    22.25184, 22.32997, 22.40195, 22.46768, 22.52709, 22.5801, 22.62664, 
    22.66665, 22.70007, 22.72686, 22.74698, 22.76041, 22.76713, 22.76713, 
    22.76041, 22.74698, 22.72686, 22.70007, 22.66665, 22.62664, 22.5801, 
    22.52709, 22.46768, 22.40195, 22.32997, 22.25184, 22.16766, 22.07753, 
    21.98156, 21.87987, 21.77258, 21.65982, 21.5417, 21.41838, 21.28997, 
    21.15662, 21.01848, 20.87569, 20.72838, 20.57672, 20.42083, 20.26088, 
    20.09701, 19.92936, 19.75808, 19.58332, 19.40522, 19.22392, 19.03956, 
    18.85229, 18.66223, 18.46952, 18.27429, 18.07666, 17.87678, 17.67474, 
    17.47068, 17.26471, 17.05695, 16.84749, 16.63645,
  17.37526, 17.59451, 17.81206, 18.02782, 18.24167, 18.45349, 18.66317, 
    18.87058, 19.07561, 19.2781, 19.47795, 19.67501, 19.86915, 20.06023, 
    20.2481, 20.43262, 20.61365, 20.79103, 20.96463, 21.13428, 21.29985, 
    21.46118, 21.61812, 21.77052, 21.91823, 22.0611, 22.19899, 22.33176, 
    22.45926, 22.58134, 22.69789, 22.80877, 22.91384, 23.01299, 23.10609, 
    23.19304, 23.27374, 23.34808, 23.41596, 23.47731, 23.53204, 23.58009, 
    23.62139, 23.6559, 23.68355, 23.70432, 23.71819, 23.72513, 23.72513, 
    23.71819, 23.70432, 23.68355, 23.6559, 23.62139, 23.58009, 23.53204, 
    23.47731, 23.41596, 23.34808, 23.27374, 23.19304, 23.10609, 23.01299, 
    22.91384, 22.80877, 22.69789, 22.58134, 22.45926, 22.33176, 22.19899, 
    22.0611, 21.91823, 21.77052, 21.61812, 21.46118, 21.29985, 21.13428, 
    20.96463, 20.79103, 20.61365, 20.43262, 20.2481, 20.06023, 19.86915, 
    19.67501, 19.47795, 19.2781, 19.07561, 18.87058, 18.66317, 18.45349, 
    18.24167, 18.02782, 17.81206, 17.59451, 17.37526,
  18.114, 18.3413, 18.5668, 18.79039, 19.01196, 19.23139, 19.44855, 19.66332, 
    19.87557, 20.08517, 20.29198, 20.49586, 20.69669, 20.8943, 21.08856, 
    21.27932, 21.46644, 21.64975, 21.82912, 22.00438, 22.17539, 22.34199, 
    22.50403, 22.66135, 22.81381, 22.96125, 23.10353, 23.2405, 23.37202, 
    23.49794, 23.61813, 23.73245, 23.84077, 23.94298, 24.03895, 24.12856, 
    24.21172, 24.28832, 24.35827, 24.42147, 24.47786, 24.52736, 24.5699, 
    24.60544, 24.63392, 24.65532, 24.6696, 24.67674, 24.67674, 24.6696, 
    24.65532, 24.63392, 24.60544, 24.5699, 24.52736, 24.47786, 24.42147, 
    24.35827, 24.28832, 24.21172, 24.12856, 24.03895, 23.94298, 23.84077, 
    23.73245, 23.61813, 23.49794, 23.37202, 23.2405, 23.10353, 22.96125, 
    22.81381, 22.66135, 22.50403, 22.34199, 22.17539, 22.00438, 21.82912, 
    21.64975, 21.46644, 21.27932, 21.08856, 20.8943, 20.69669, 20.49586, 
    20.29198, 20.08517, 19.87557, 19.66332, 19.44855, 19.23139, 19.01196, 
    18.79039, 18.5668, 18.3413, 18.114,
  18.85267, 19.08786, 19.32115, 19.55242, 19.78154, 20.0084, 20.23287, 
    20.45482, 20.67413, 20.89065, 21.10424, 21.31477, 21.52209, 21.72607, 
    21.92654, 22.12335, 22.31637, 22.50543, 22.69039, 22.87107, 23.04734, 
    23.21904, 23.386, 23.54808, 23.70512, 23.85697, 24.00347, 24.14449, 
    24.27987, 24.40947, 24.53315, 24.65079, 24.76223, 24.86737, 24.96609, 
    25.05826, 25.14377, 25.22254, 25.29446, 25.35944, 25.41741, 25.46829, 
    25.51202, 25.54855, 25.57783, 25.59982, 25.6145, 25.62184, 25.62184, 
    25.6145, 25.59982, 25.57783, 25.54855, 25.51202, 25.46829, 25.41741, 
    25.35944, 25.29446, 25.22254, 25.14377, 25.05826, 24.96609, 24.86737, 
    24.76223, 24.65079, 24.53315, 24.40947, 24.27987, 24.14449, 24.00347, 
    23.85697, 23.70512, 23.54808, 23.386, 23.21904, 23.04734, 22.87107, 
    22.69039, 22.50543, 22.31637, 22.12335, 21.92654, 21.72607, 21.52209, 
    21.31477, 21.10424, 20.89065, 20.67413, 20.45482, 20.23287, 20.0084, 
    19.78154, 19.55242, 19.32115, 19.08786, 18.85267,
  19.59126, 19.83419, 20.0751, 20.31387, 20.55038, 20.7845, 21.01611, 
    21.24507, 21.47124, 21.6945, 21.91469, 22.13168, 22.34532, 22.55546, 
    22.76195, 22.96464, 23.16337, 23.35799, 23.54835, 23.73428, 23.91562, 
    24.09223, 24.26394, 24.43059, 24.59204, 24.74813, 24.89869, 25.04359, 
    25.18268, 25.31582, 25.44285, 25.56366, 25.6781, 25.78605, 25.88738, 
    25.98199, 26.06977, 26.1506, 26.2244, 26.29108, 26.35056, 26.40276, 
    26.44763, 26.4851, 26.51514, 26.5377, 26.55275, 26.56029, 26.56029, 
    26.55275, 26.5377, 26.51514, 26.4851, 26.44763, 26.40276, 26.35056, 
    26.29108, 26.2244, 26.1506, 26.06977, 25.98199, 25.88738, 25.78605, 
    25.6781, 25.56366, 25.44285, 25.31582, 25.18268, 25.04359, 24.89869, 
    24.74813, 24.59204, 24.43059, 24.26394, 24.09223, 23.91562, 23.73428, 
    23.54835, 23.35799, 23.16337, 22.96464, 22.76195, 22.55546, 22.34532, 
    22.13168, 21.91469, 21.6945, 21.47124, 21.24507, 21.01611, 20.7845, 
    20.55038, 20.31387, 20.0751, 19.83419, 19.59126,
  20.32976, 20.58027, 20.82863, 21.07474, 21.31846, 21.55966, 21.79822, 
    22.034, 22.26687, 22.49667, 22.72328, 22.94654, 23.1663, 23.38242, 
    23.59474, 23.8031, 24.00736, 24.20735, 24.40292, 24.5939, 24.78014, 
    24.96147, 25.13775, 25.3088, 25.47448, 25.63463, 25.78909, 25.93772, 
    26.08036, 26.21687, 26.34712, 26.47095, 26.58825, 26.69888, 26.80272, 
    26.89966, 26.98958, 27.07239, 27.14798, 27.21628, 27.27719, 27.33065, 
    27.3766, 27.41497, 27.44572, 27.46882, 27.48424, 27.49195, 27.49195, 
    27.48424, 27.46882, 27.44572, 27.41497, 27.3766, 27.33065, 27.27719, 
    27.21628, 27.14798, 27.07239, 26.98958, 26.89966, 26.80272, 26.69888, 
    26.58825, 26.47095, 26.34712, 26.21687, 26.08036, 25.93772, 25.78909, 
    25.63463, 25.47448, 25.3088, 25.13775, 24.96147, 24.78014, 24.5939, 
    24.40292, 24.20735, 24.00736, 23.8031, 23.59474, 23.38242, 23.1663, 
    22.94654, 22.72328, 22.49667, 22.26687, 22.034, 21.79822, 21.55966, 
    21.31846, 21.07474, 20.82863, 20.58027, 20.32976,
  21.06818, 21.32609, 21.58174, 21.835, 22.08575, 22.33386, 22.57919, 
    22.8216, 23.06096, 23.29713, 23.52995, 23.75929, 23.98498, 24.20688, 
    24.42483, 24.63868, 24.84826, 25.05343, 25.25401, 25.44986, 25.6408, 
    25.82668, 26.00734, 26.18261, 26.35234, 26.51638, 26.67457, 26.82676, 
    26.9728, 27.11254, 27.24584, 27.37256, 27.49258, 27.60576, 27.71199, 
    27.81114, 27.90311, 27.98779, 28.06509, 28.13491, 28.19719, 28.25185, 
    28.29881, 28.33804, 28.36947, 28.39308, 28.40884, 28.41672, 28.41672, 
    28.40884, 28.39308, 28.36947, 28.33804, 28.29881, 28.25185, 28.19719, 
    28.13491, 28.06509, 27.98779, 27.90311, 27.81114, 27.71199, 27.60576, 
    27.49258, 27.37256, 27.24584, 27.11254, 26.9728, 26.82676, 26.67457, 
    26.51638, 26.35234, 26.18261, 26.00734, 25.82668, 25.6408, 25.44986, 
    25.25401, 25.05343, 24.84826, 24.63868, 24.42483, 24.20688, 23.98498, 
    23.75929, 23.52995, 23.29713, 23.06096, 22.8216, 22.57919, 22.33386, 
    22.08575, 21.835, 21.58174, 21.32609, 21.06818,
  21.80651, 22.07165, 22.33441, 22.59464, 22.85224, 23.10706, 23.35897, 
    23.60783, 23.85349, 24.09582, 24.33467, 24.56988, 24.8013, 25.02878, 
    25.25217, 25.4713, 25.68602, 25.89616, 26.10157, 26.30208, 26.49753, 
    26.68777, 26.87262, 27.05193, 27.22555, 27.3933, 27.55505, 27.71063, 
    27.8599, 28.00271, 28.13892, 28.2684, 28.391, 28.50661, 28.6151, 
    28.71634, 28.81025, 28.89671, 28.97562, 29.0469, 29.11047, 29.16625, 
    29.21418, 29.25421, 29.28629, 29.31038, 29.32646, 29.33451, 29.33451, 
    29.32646, 29.31038, 29.28629, 29.25421, 29.21418, 29.16625, 29.11047, 
    29.0469, 28.97562, 28.89671, 28.81025, 28.71634, 28.6151, 28.50661, 
    28.391, 28.2684, 28.13892, 28.00271, 27.8599, 27.71063, 27.55505, 
    27.3933, 27.22555, 27.05193, 26.87262, 26.68777, 26.49753, 26.30208, 
    26.10157, 25.89616, 25.68602, 25.4713, 25.25217, 25.02878, 24.8013, 
    24.56988, 24.33467, 24.09582, 23.85349, 23.60783, 23.35897, 23.10706, 
    22.85224, 22.59464, 22.33441, 22.07165, 21.80651,
  22.54476, 22.81695, 23.08662, 23.35365, 23.6179, 23.87924, 24.13754, 
    24.39264, 24.64441, 24.89271, 25.13737, 25.37826, 25.61521, 25.84807, 
    26.07669, 26.30091, 26.52055, 26.73548, 26.94551, 27.1505, 27.35027, 
    27.54466, 27.73353, 27.91669, 28.094, 28.2653, 28.43043, 28.58924, 
    28.74158, 28.88731, 29.02629, 29.15837, 29.28342, 29.40132, 29.51195, 
    29.61518, 29.71092, 29.79905, 29.87949, 29.95214, 30.01692, 30.07377, 
    30.12261, 30.1634, 30.19609, 30.22064, 30.23702, 30.24521, 30.24521, 
    30.23702, 30.22064, 30.19609, 30.1634, 30.12261, 30.07377, 30.01692, 
    29.95214, 29.87949, 29.79905, 29.71092, 29.61518, 29.51195, 29.40132, 
    29.28342, 29.15837, 29.02629, 28.88731, 28.74158, 28.58924, 28.43043, 
    28.2653, 28.094, 27.91669, 27.73353, 27.54466, 27.35027, 27.1505, 
    26.94551, 26.73548, 26.52055, 26.30091, 26.07669, 25.84807, 25.61521, 
    25.37826, 25.13737, 24.89271, 24.64441, 24.39264, 24.13754, 23.87924, 
    23.6179, 23.35365, 23.08662, 22.81695, 22.54476,
  23.28291, 23.56197, 23.83837, 24.112, 24.38272, 24.65038, 24.91487, 
    25.17602, 25.43369, 25.68774, 25.93803, 26.18438, 26.42666, 26.6647, 
    26.89834, 27.12744, 27.35181, 27.57131, 27.78577, 27.99503, 28.19893, 
    28.3973, 28.58998, 28.77681, 28.95764, 29.1323, 29.30065, 29.46252, 
    29.61777, 29.76627, 29.90785, 30.04239, 30.16976, 30.28983, 30.40247, 
    30.50758, 30.60504, 30.69475, 30.77662, 30.85055, 30.91648, 30.97433, 
    31.02403, 31.06553, 31.09879, 31.12376, 31.14043, 31.14876, 31.14876, 
    31.14043, 31.12376, 31.09879, 31.06553, 31.02403, 30.97433, 30.91648, 
    30.85055, 30.77662, 30.69475, 30.60504, 30.50758, 30.40247, 30.28983, 
    30.16976, 30.04239, 29.90785, 29.76627, 29.61777, 29.46252, 29.30065, 
    29.1323, 28.95764, 28.77681, 28.58998, 28.3973, 28.19893, 27.99503, 
    27.78577, 27.57131, 27.35181, 27.12744, 26.89834, 26.6647, 26.42666, 
    26.18438, 25.93803, 25.68774, 25.43369, 25.17602, 24.91487, 24.65038, 
    24.38272, 24.112, 23.83837, 23.56197, 23.28291,
  24.02097, 24.3067, 24.58965, 24.86968, 25.14667, 25.42046, 25.69092, 
    25.95792, 26.22129, 26.4809, 26.73659, 26.98821, 27.2356, 27.47861, 
    27.71707, 27.95084, 28.17974, 28.40361, 28.6223, 28.83563, 29.04346, 
    29.2456, 29.44192, 29.63223, 29.81639, 29.99424, 30.16563, 30.3304, 
    30.4884, 30.6395, 30.78355, 30.92041, 31.04995, 31.17205, 31.28659, 
    31.39346, 31.49253, 31.58372, 31.66694, 31.74208, 31.80908, 31.86786, 
    31.91836, 31.96053, 31.99432, 32.01969, 32.03662, 32.04509, 32.04509, 
    32.03662, 32.01969, 31.99432, 31.96053, 31.91836, 31.86786, 31.80908, 
    31.74208, 31.66694, 31.58372, 31.49253, 31.39346, 31.28659, 31.17205, 
    31.04995, 30.92041, 30.78355, 30.6395, 30.4884, 30.3304, 30.16563, 
    29.99424, 29.81639, 29.63223, 29.44192, 29.2456, 29.04346, 28.83563, 
    28.6223, 28.40361, 28.17974, 27.95084, 27.71707, 27.47861, 27.2356, 
    26.98821, 26.73659, 26.4809, 26.22129, 25.95792, 25.69092, 25.42046, 
    25.14667, 24.86968, 24.58965, 24.3067, 24.02097,
  24.75893, 25.05115, 25.34044, 25.62668, 25.90973, 26.18944, 26.46569, 
    26.73832, 27.00718, 27.27213, 27.53302, 27.78969, 28.04199, 28.28975, 
    28.53283, 28.77106, 29.00427, 29.23232, 29.45502, 29.67224, 29.88379, 
    30.08952, 30.28927, 30.48288, 30.6702, 30.85106, 31.02531, 31.19281, 
    31.3534, 31.50695, 31.65331, 31.79235, 31.92393, 32.04794, 32.16426, 
    32.27277, 32.37335, 32.46593, 32.55039, 32.62666, 32.69466, 32.75431, 
    32.80555, 32.84834, 32.88263, 32.90837, 32.92555, 32.93415, 32.93415, 
    32.92555, 32.90837, 32.88263, 32.84834, 32.80555, 32.75431, 32.69466, 
    32.62666, 32.55039, 32.46593, 32.37335, 32.27277, 32.16426, 32.04794, 
    31.92393, 31.79235, 31.65331, 31.50695, 31.3534, 31.19281, 31.02531, 
    30.85106, 30.6702, 30.48288, 30.28927, 30.08952, 29.88379, 29.67224, 
    29.45502, 29.23232, 29.00427, 28.77106, 28.53283, 28.28975, 28.04199, 
    27.78969, 27.53302, 27.27213, 27.00718, 26.73832, 26.46569, 26.18944, 
    25.90973, 25.62668, 25.34044, 25.05115, 24.75893,
  25.4968, 25.7953, 26.09074, 26.38298, 26.67189, 26.95732, 27.23913, 
    27.51719, 27.79133, 28.06141, 28.32729, 28.5888, 28.84579, 29.0981, 
    29.34557, 29.58805, 29.82537, 30.05738, 30.28391, 30.50479, 30.71988, 
    30.929, 31.132, 31.32872, 31.519, 31.70269, 31.87964, 32.0497, 32.21272, 
    32.36856, 32.51709, 32.65816, 32.79165, 32.91744, 33.03541, 33.14545, 
    33.24744, 33.3413, 33.42693, 33.50424, 33.57316, 33.63363, 33.68556, 
    33.72892, 33.76367, 33.78976, 33.80717, 33.81588, 33.81588, 33.80717, 
    33.78976, 33.76367, 33.72892, 33.68556, 33.63363, 33.57316, 33.50424, 
    33.42693, 33.3413, 33.24744, 33.14545, 33.03541, 32.91744, 32.79165, 
    32.65816, 32.51709, 32.36856, 32.21272, 32.0497, 31.87964, 31.70269, 
    31.519, 31.32872, 31.132, 30.929, 30.71988, 30.50479, 30.28391, 30.05738, 
    29.82537, 29.58805, 29.34557, 29.0981, 28.84579, 28.5888, 28.32729, 
    28.06141, 27.79133, 27.51719, 27.23913, 26.95732, 26.67189, 26.38298, 
    26.09074, 25.7953, 25.4968,
  26.23456, 26.53915, 26.84053, 27.13857, 27.43312, 27.72406, 28.01123, 
    28.29449, 28.5737, 28.84871, 29.11935, 29.38548, 29.64695, 29.90359, 
    30.15525, 30.40177, 30.643, 30.87876, 31.10889, 31.33325, 31.55167, 
    31.76398, 31.97004, 32.16968, 32.36275, 32.5491, 32.72858, 32.90103, 
    33.06631, 33.2243, 33.37484, 33.5178, 33.65307, 33.78051, 33.90001, 
    34.01146, 34.11476, 34.20981, 34.29651, 34.37479, 34.44456, 34.50577, 
    34.55835, 34.60224, 34.63741, 34.66381, 34.68143, 34.69025, 34.69025, 
    34.68143, 34.66381, 34.63741, 34.60224, 34.55835, 34.50577, 34.44456, 
    34.37479, 34.29651, 34.20981, 34.11476, 34.01146, 33.90001, 33.78051, 
    33.65307, 33.5178, 33.37484, 33.2243, 33.06631, 32.90103, 32.72858, 
    32.5491, 32.36275, 32.16968, 31.97004, 31.76398, 31.55167, 31.33325, 
    31.10889, 30.87876, 30.643, 30.40177, 30.15525, 29.90359, 29.64695, 
    29.38548, 29.11935, 28.84871, 28.5737, 28.29449, 28.01123, 27.72406, 
    27.43312, 27.13857, 26.84053, 26.53915, 26.23456,
  26.97222, 27.28269, 27.58981, 27.89343, 28.19342, 28.48965, 28.78197, 
    29.07022, 29.35428, 29.63398, 29.90917, 30.17971, 30.44544, 30.7062, 
    30.96183, 31.21218, 31.45709, 31.6964, 31.92994, 32.15757, 32.37912, 
    32.59444, 32.80336, 33.00574, 33.20141, 33.39024, 33.57207, 33.74675, 
    33.91414, 34.07411, 34.22652, 34.37123, 34.50814, 34.6371, 34.75802, 
    34.87078, 34.97528, 35.07141, 35.15911, 35.23827, 35.30883, 35.37072, 
    35.42388, 35.46826, 35.50381, 35.53051, 35.54832, 35.55723, 35.55723, 
    35.54832, 35.53051, 35.50381, 35.46826, 35.42388, 35.37072, 35.30883, 
    35.23827, 35.15911, 35.07141, 34.97528, 34.87078, 34.75802, 34.6371, 
    34.50814, 34.37123, 34.22652, 34.07411, 33.91414, 33.74675, 33.57207, 
    33.39024, 33.20141, 33.00574, 32.80336, 32.59444, 32.37912, 32.15757, 
    31.92994, 31.6964, 31.45709, 31.21218, 30.96183, 30.7062, 30.44544, 
    30.17971, 29.90917, 29.63398, 29.35428, 29.07022, 28.78197, 28.48965, 
    28.19342, 27.89343, 27.58981, 27.28269, 26.97222,
  27.70978, 28.02592, 28.33856, 28.64755, 28.95277, 29.25407, 29.55131, 
    29.84434, 30.13302, 30.4172, 30.69673, 30.97146, 31.24123, 31.50589, 
    31.76528, 32.01924, 32.26763, 32.51027, 32.74702, 32.97771, 33.2022, 
    33.42032, 33.63192, 33.83684, 34.03494, 34.22607, 34.41008, 34.58682, 
    34.75616, 34.91797, 35.0721, 35.21843, 35.35684, 35.48721, 35.60942, 
    35.72337, 35.82896, 35.9261, 36.01469, 36.09467, 36.16594, 36.22845, 
    36.28214, 36.32696, 36.36287, 36.38982, 36.40781, 36.41681, 36.41681, 
    36.40781, 36.38982, 36.36287, 36.32696, 36.28214, 36.22845, 36.16594, 
    36.09467, 36.01469, 35.9261, 35.82896, 35.72337, 35.60942, 35.48721, 
    35.35684, 35.21843, 35.0721, 34.91797, 34.75616, 34.58682, 34.41008, 
    34.22607, 34.03494, 33.83684, 33.63192, 33.42032, 33.2022, 32.97771, 
    32.74702, 32.51027, 32.26763, 32.01924, 31.76528, 31.50589, 31.24123, 
    30.97146, 30.69673, 30.4172, 30.13302, 29.84434, 29.55131, 29.25407, 
    28.95277, 28.64755, 28.33856, 28.02592, 27.70978,
  28.44723, 28.76883, 29.08677, 29.40093, 29.71115, 30.0173, 30.31924, 
    30.61683, 30.90992, 31.19835, 31.482, 31.76069, 32.03428, 32.30262, 
    32.56555, 32.82292, 33.07457, 33.32034, 33.56009, 33.79364, 34.02087, 
    34.2416, 34.45568, 34.66297, 34.86331, 35.05656, 35.24258, 35.42123, 
    35.59236, 35.75585, 35.91155, 36.05936, 36.19914, 36.33079, 36.45418, 
    36.56922, 36.67581, 36.77385, 36.86326, 36.94396, 37.01588, 37.07895, 
    37.13312, 37.17834, 37.21456, 37.24176, 37.2599, 37.26898, 37.26898, 
    37.2599, 37.24176, 37.21456, 37.17834, 37.13312, 37.07895, 37.01588, 
    36.94396, 36.86326, 36.77385, 36.67581, 36.56922, 36.45418, 36.33079, 
    36.19914, 36.05936, 35.91155, 35.75585, 35.59236, 35.42123, 35.24258, 
    35.05656, 34.86331, 34.66297, 34.45568, 34.2416, 34.02087, 33.79364, 
    33.56009, 33.32034, 33.07457, 32.82292, 32.56555, 32.30262, 32.03428, 
    31.76069, 31.482, 31.19835, 30.90992, 30.61683, 30.31924, 30.0173, 
    29.71115, 29.40093, 29.08677, 28.76883, 28.44723,
  29.18457, 29.51142, 29.83445, 30.15354, 30.46854, 30.77932, 31.08575, 
    31.38766, 31.68493, 31.97741, 32.26494, 32.54737, 32.82457, 33.09637, 
    33.36263, 33.62318, 33.87788, 34.12658, 34.36911, 34.60533, 34.83509, 
    35.05824, 35.27462, 35.48409, 35.68649, 35.8817, 36.06956, 36.24994, 
    36.42271, 36.58773, 36.74487, 36.89401, 37.03504, 37.16784, 37.2923, 
    37.40832, 37.5158, 37.61465, 37.7048, 37.78615, 37.85865, 37.92222, 
    37.97682, 38.02239, 38.0589, 38.0863, 38.10459, 38.11374, 38.11374, 
    38.10459, 38.0863, 38.0589, 38.02239, 37.97682, 37.92222, 37.85865, 
    37.78615, 37.7048, 37.61465, 37.5158, 37.40832, 37.2923, 37.16784, 
    37.03504, 36.89401, 36.74487, 36.58773, 36.42271, 36.24994, 36.06956, 
    35.8817, 35.68649, 35.48409, 35.27462, 35.05824, 34.83509, 34.60533, 
    34.36911, 34.12658, 33.87788, 33.62318, 33.36263, 33.09637, 32.82457, 
    32.54737, 32.26494, 31.97741, 31.68493, 31.38766, 31.08575, 30.77932, 
    30.46854, 30.15354, 29.83445, 29.51142, 29.18457,
  29.92181, 30.25368, 30.58158, 30.90537, 31.22494, 31.54013, 31.8508, 
    32.15683, 32.45805, 32.75434, 33.04553, 33.33149, 33.61207, 33.88711, 
    34.15647, 34.42, 34.67754, 34.92895, 35.17407, 35.41275, 35.64485, 
    35.87022, 36.08871, 36.30017, 36.50447, 36.70145, 36.891, 37.07295, 
    37.2472, 37.4136, 37.57203, 37.72238, 37.86452, 37.99836, 38.12377, 
    38.24066, 38.34894, 38.44851, 38.53931, 38.62124, 38.69425, 38.75827, 
    38.81324, 38.85912, 38.89588, 38.92347, 38.94188, 38.95109, 38.95109, 
    38.94188, 38.92347, 38.89588, 38.85912, 38.81324, 38.75827, 38.69425, 
    38.62124, 38.53931, 38.44851, 38.34894, 38.24066, 38.12377, 37.99836, 
    37.86452, 37.72238, 37.57203, 37.4136, 37.2472, 37.07295, 36.891, 
    36.70145, 36.50447, 36.30017, 36.08871, 35.87022, 35.64485, 35.41275, 
    35.17407, 34.92895, 34.67754, 34.42, 34.15647, 33.88711, 33.61207, 
    33.33149, 33.04553, 32.75434, 32.45805, 32.15683, 31.8508, 31.54013, 
    31.22494, 30.90537, 30.58158, 30.25368, 29.92181,
  30.65893, 30.9956, 31.32814, 31.65643, 31.98032, 32.29969, 32.6144, 
    32.9243, 33.22925, 33.52912, 33.82376, 34.11302, 34.39675, 34.67482, 
    34.94707, 35.21335, 35.47353, 35.72744, 35.97494, 36.21589, 36.45013, 
    36.67753, 36.89794, 37.11122, 37.31722, 37.51582, 37.70687, 37.89024, 
    38.06581, 38.23346, 38.39304, 38.54446, 38.6876, 38.82234, 38.94859, 
    39.06625, 39.17523, 39.27544, 39.3668, 39.44924, 39.52269, 39.58709, 
    39.6424, 39.68855, 39.72552, 39.75327, 39.77179, 39.78105, 39.78105, 
    39.77179, 39.75327, 39.72552, 39.68855, 39.6424, 39.58709, 39.52269, 
    39.44924, 39.3668, 39.27544, 39.17523, 39.06625, 38.94859, 38.82234, 
    38.6876, 38.54446, 38.39304, 38.23346, 38.06581, 37.89024, 37.70687, 
    37.51582, 37.31722, 37.11122, 36.89794, 36.67753, 36.45013, 36.21589, 
    35.97494, 35.72744, 35.47353, 35.21335, 34.94707, 34.67482, 34.39675, 
    34.11302, 33.82376, 33.52912, 33.22925, 32.9243, 32.6144, 32.29969, 
    31.98032, 31.65643, 31.32814, 30.9956, 30.65893,
  31.39594, 31.73718, 32.07414, 32.40669, 32.73469, 33.05801, 33.37651, 
    33.69006, 33.99852, 34.30174, 34.59959, 34.89193, 35.1786, 35.45947, 
    35.73439, 36.00322, 36.26581, 36.52202, 36.7717, 37.01471, 37.2509, 
    37.48015, 37.70229, 37.9172, 38.12474, 38.32478, 38.51718, 38.70182, 
    38.87856, 39.04729, 39.20789, 39.36025, 39.50425, 39.63979, 39.76678, 
    39.88511, 39.99469, 40.09544, 40.18729, 40.27016, 40.34399, 40.40873, 
    40.46431, 40.51069, 40.54784, 40.57574, 40.59435, 40.60365, 40.60365, 
    40.59435, 40.57574, 40.54784, 40.51069, 40.46431, 40.40873, 40.34399, 
    40.27016, 40.18729, 40.09544, 39.99469, 39.88511, 39.76678, 39.63979, 
    39.50425, 39.36025, 39.20789, 39.04729, 38.87856, 38.70182, 38.51718, 
    38.32478, 38.12474, 37.9172, 37.70229, 37.48015, 37.2509, 37.01471, 
    36.7717, 36.52202, 36.26581, 36.00322, 35.73439, 35.45947, 35.1786, 
    34.89193, 34.59959, 34.30174, 33.99852, 33.69006, 33.37651, 33.05801, 
    32.73469, 32.40669, 32.07414, 31.73718, 31.39594,
  32.13284, 32.47842, 32.81957, 33.15614, 33.48802, 33.81506, 34.13713, 
    34.4541, 34.76583, 35.07218, 35.37302, 35.66821, 35.9576, 36.24105, 
    36.51843, 36.78959, 37.05439, 37.31269, 37.56434, 37.80922, 38.04717, 
    38.27806, 38.50176, 38.71813, 38.92703, 39.12834, 39.32193, 39.50767, 
    39.68544, 39.85512, 40.0166, 40.16977, 40.31451, 40.45074, 40.57834, 
    40.69724, 40.80733, 40.90854, 41.0008, 41.08404, 41.15818, 41.22319, 
    41.279, 41.32558, 41.36288, 41.39089, 41.40957, 41.41891, 41.41891, 
    41.40957, 41.39089, 41.36288, 41.32558, 41.279, 41.22319, 41.15818, 
    41.08404, 41.0008, 40.90854, 40.80733, 40.69724, 40.57834, 40.45074, 
    40.31451, 40.16977, 40.0166, 39.85512, 39.68544, 39.50767, 39.32193, 
    39.12834, 38.92703, 38.71813, 38.50176, 38.27806, 38.04717, 37.80922, 
    37.56434, 37.31269, 37.05439, 36.78959, 36.51843, 36.24105, 35.9576, 
    35.66821, 35.37302, 35.07218, 34.76583, 34.4541, 34.13713, 33.81506, 
    33.48802, 33.15614, 32.81957, 32.47842, 32.13284,
  32.86962, 33.21932, 33.56442, 33.90479, 34.2403, 34.57083, 34.89624, 
    35.2164, 35.53117, 35.84042, 36.14403, 36.44184, 36.73372, 37.01954, 
    37.29916, 37.57244, 37.83924, 38.09942, 38.35286, 38.5994, 38.83891, 
    39.07127, 39.29634, 39.51399, 39.72409, 39.9265, 40.12112, 40.30781, 
    40.48646, 40.65696, 40.81918, 40.97303, 41.1184, 41.25519, 41.38331, 
    41.50267, 41.61318, 41.71477, 41.80736, 41.89089, 41.96529, 42.03052, 
    42.08652, 42.13324, 42.17067, 42.19876, 42.2175, 42.22688, 42.22688, 
    42.2175, 42.19876, 42.17067, 42.13324, 42.08652, 42.03052, 41.96529, 
    41.89089, 41.80736, 41.71477, 41.61318, 41.50267, 41.38331, 41.25519, 
    41.1184, 40.97303, 40.81918, 40.65696, 40.48646, 40.30781, 40.12112, 
    39.9265, 39.72409, 39.51399, 39.29634, 39.07127, 38.83891, 38.5994, 
    38.35286, 38.09942, 37.83924, 37.57244, 37.29916, 37.01954, 36.73372, 
    36.44184, 36.14403, 35.84042, 35.53117, 35.2164, 34.89624, 34.57083, 
    34.2403, 33.90479, 33.56442, 33.21932, 32.86962,
  33.60628, 33.95987, 34.30869, 34.65261, 34.99154, 35.32531, 35.65382, 
    35.97694, 36.29453, 36.60646, 36.91259, 37.21281, 37.50697, 37.79493, 
    38.07658, 38.35176, 38.62035, 38.88222, 39.13723, 39.38524, 39.62614, 
    39.85978, 40.08604, 40.30479, 40.51591, 40.71927, 40.91476, 41.10225, 
    41.28164, 41.4528, 41.61564, 41.77005, 41.91592, 42.05317, 42.18171, 
    42.30143, 42.41228, 42.51416, 42.60701, 42.69076, 42.76536, 42.83075, 
    42.88689, 42.93373, 42.97124, 42.9994, 43.01819, 43.02758, 43.02758, 
    43.01819, 42.9994, 42.97124, 42.93373, 42.88689, 42.83075, 42.76536, 
    42.69076, 42.60701, 42.51416, 42.41228, 42.30143, 42.18171, 42.05317, 
    41.91592, 41.77005, 41.61564, 41.4528, 41.28164, 41.10225, 40.91476, 
    40.71927, 40.51591, 40.30479, 40.08604, 39.85978, 39.62614, 39.38524, 
    39.13723, 38.88222, 38.62035, 38.35176, 38.07658, 37.79493, 37.50697, 
    37.21281, 36.91259, 36.60646, 36.29453, 35.97694, 35.65382, 35.32531, 
    34.99154, 34.65261, 34.30869, 33.95987, 33.60628,
  34.34282, 34.70005, 35.05236, 35.39962, 35.7417, 36.0785, 36.40988, 
    36.73572, 37.05589, 37.37026, 37.67871, 37.9811, 38.27731, 38.56721, 
    38.85067, 39.12755, 39.39772, 39.66107, 39.91746, 40.16676, 40.40884, 
    40.64358, 40.87085, 41.09053, 41.30251, 41.50666, 41.70287, 41.89101, 
    42.07099, 42.24269, 42.40602, 42.56086, 42.70713, 42.84472, 42.97356, 
    43.09357, 43.20465, 43.30674, 43.39978, 43.48369, 43.55843, 43.62393, 
    43.68016, 43.72708, 43.76466, 43.79286, 43.81168, 43.82109, 43.82109, 
    43.81168, 43.79286, 43.76466, 43.72708, 43.68016, 43.62393, 43.55843, 
    43.48369, 43.39978, 43.30674, 43.20465, 43.09357, 42.97356, 42.84472, 
    42.70713, 42.56086, 42.40602, 42.24269, 42.07099, 41.89101, 41.70287, 
    41.50666, 41.30251, 41.09053, 40.87085, 40.64358, 40.40884, 40.16676, 
    39.91746, 39.66107, 39.39772, 39.12755, 38.85067, 38.56721, 38.27731, 
    37.9811, 37.67871, 37.37026, 37.05589, 36.73572, 36.40988, 36.0785, 
    35.7417, 35.39962, 35.05236, 34.70005, 34.34282,
  35.07925, 35.43988, 35.79544, 36.14578, 36.4908, 36.83038, 37.1644, 
    37.49273, 37.81525, 38.13184, 38.44237, 38.74672, 39.04476, 39.33637, 
    39.62142, 39.89979, 40.17135, 40.43598, 40.69355, 40.94394, 41.18702, 
    41.42268, 41.65079, 41.87124, 42.08391, 42.28868, 42.48545, 42.67411, 
    42.85454, 43.02665, 43.19033, 43.34549, 43.49203, 43.62987, 43.75893, 
    43.87911, 43.99035, 44.09258, 44.18572, 44.26973, 44.34454, 44.41011, 
    44.46639, 44.51335, 44.55096, 44.57919, 44.59801, 44.60743, 44.60743, 
    44.59801, 44.57919, 44.55096, 44.51335, 44.46639, 44.41011, 44.34454, 
    44.26973, 44.18572, 44.09258, 43.99035, 43.87911, 43.75893, 43.62987, 
    43.49203, 43.34549, 43.19033, 43.02665, 42.85454, 42.67411, 42.48545, 
    42.28868, 42.08391, 41.87124, 41.65079, 41.42268, 41.18702, 40.94394, 
    40.69355, 40.43598, 40.17135, 39.89979, 39.62142, 39.33637, 39.04476, 
    38.74672, 38.44237, 38.13184, 37.81525, 37.49273, 37.1644, 36.83038, 
    36.4908, 36.14578, 35.79544, 35.43988, 35.07925 ;

 area =
  5.832426e+09, 5.885548e+09, 5.937712e+09, 5.988909e+09, 6.039129e+09, 
    6.088361e+09, 6.136596e+09, 6.183825e+09, 6.230037e+09, 6.275223e+09, 
    6.319373e+09, 6.362479e+09, 6.404531e+09, 6.445522e+09, 6.485442e+09, 
    6.524282e+09, 6.562035e+09, 6.598693e+09, 6.634248e+09, 6.668692e+09, 
    6.702019e+09, 6.734221e+09, 6.76529e+09, 6.795221e+09, 6.824007e+09, 
    6.851641e+09, 6.878117e+09, 6.903431e+09, 6.927576e+09, 6.950547e+09, 
    6.972339e+09, 6.992947e+09, 7.012366e+09, 7.030593e+09, 7.047623e+09, 
    7.063453e+09, 7.078078e+09, 7.091497e+09, 7.103705e+09, 7.1147e+09, 
    7.124479e+09, 7.133041e+09, 7.140384e+09, 7.146505e+09, 7.151404e+09, 
    7.155078e+09, 7.157529e+09, 7.158754e+09, 7.158754e+09, 7.157529e+09, 
    7.155078e+09, 7.151404e+09, 7.146505e+09, 7.140384e+09, 7.133041e+09, 
    7.124479e+09, 7.1147e+09, 7.103705e+09, 7.091497e+09, 7.078078e+09, 
    7.063453e+09, 7.047623e+09, 7.030593e+09, 7.012366e+09, 6.992947e+09, 
    6.972339e+09, 6.950547e+09, 6.927576e+09, 6.903431e+09, 6.878117e+09, 
    6.851641e+09, 6.824007e+09, 6.795221e+09, 6.76529e+09, 6.734221e+09, 
    6.702019e+09, 6.668692e+09, 6.634248e+09, 6.598693e+09, 6.562035e+09, 
    6.524282e+09, 6.485442e+09, 6.445522e+09, 6.404531e+09, 6.362479e+09, 
    6.319373e+09, 6.275223e+09, 6.230037e+09, 6.183825e+09, 6.136596e+09, 
    6.088361e+09, 6.039129e+09, 5.988909e+09, 5.937712e+09, 5.885548e+09, 
    5.832426e+09,
  5.885548e+09, 5.942029e+09, 5.99757e+09, 6.052155e+09, 6.105772e+09, 
    6.158404e+09, 6.210038e+09, 6.260659e+09, 6.310255e+09, 6.35881e+09, 
    6.406312e+09, 6.452746e+09, 6.4981e+09, 6.54236e+09, 6.585513e+09, 
    6.627547e+09, 6.668449e+09, 6.708208e+09, 6.74681e+09, 6.784244e+09, 
    6.8205e+09, 6.855565e+09, 6.889429e+09, 6.922081e+09, 6.953512e+09, 
    6.98371e+09, 7.012667e+09, 7.040374e+09, 7.066821e+09, 7.092e+09, 
    7.115902e+09, 7.138521e+09, 7.159848e+09, 7.179877e+09, 7.198601e+09, 
    7.216014e+09, 7.23211e+09, 7.246883e+09, 7.260329e+09, 7.272444e+09, 
    7.283223e+09, 7.292662e+09, 7.30076e+09, 7.307511e+09, 7.312915e+09, 
    7.316969e+09, 7.319673e+09, 7.321026e+09, 7.321026e+09, 7.319673e+09, 
    7.316969e+09, 7.312915e+09, 7.307511e+09, 7.30076e+09, 7.292662e+09, 
    7.283223e+09, 7.272444e+09, 7.260329e+09, 7.246883e+09, 7.23211e+09, 
    7.216014e+09, 7.198601e+09, 7.179877e+09, 7.159848e+09, 7.138521e+09, 
    7.115902e+09, 7.092e+09, 7.066821e+09, 7.040374e+09, 7.012667e+09, 
    6.98371e+09, 6.953512e+09, 6.922081e+09, 6.889429e+09, 6.855565e+09, 
    6.8205e+09, 6.784244e+09, 6.74681e+09, 6.708208e+09, 6.668449e+09, 
    6.627547e+09, 6.585513e+09, 6.54236e+09, 6.4981e+09, 6.452746e+09, 
    6.406312e+09, 6.35881e+09, 6.310255e+09, 6.260659e+09, 6.210038e+09, 
    6.158404e+09, 6.105772e+09, 6.052155e+09, 5.99757e+09, 5.942029e+09, 
    5.885548e+09,
  5.937712e+09, 5.99757e+09, 6.056508e+09, 6.114508e+09, 6.171552e+09, 
    6.227619e+09, 6.282692e+09, 6.336752e+09, 6.38978e+09, 6.441759e+09, 
    6.492669e+09, 6.542493e+09, 6.591213e+09, 6.638811e+09, 6.685269e+09, 
    6.730571e+09, 6.774699e+09, 6.817636e+09, 6.859367e+09, 6.899874e+09, 
    6.939143e+09, 6.977157e+09, 7.013901e+09, 7.049361e+09, 7.083523e+09, 
    7.116371e+09, 7.147894e+09, 7.178077e+09, 7.206909e+09, 7.234377e+09, 
    7.260469e+09, 7.285175e+09, 7.308484e+09, 7.330385e+09, 7.350871e+09, 
    7.36993e+09, 7.387556e+09, 7.403741e+09, 7.418477e+09, 7.431758e+09, 
    7.443579e+09, 7.453934e+09, 7.462817e+09, 7.470226e+09, 7.476158e+09, 
    7.480609e+09, 7.483577e+09, 7.485062e+09, 7.485062e+09, 7.483577e+09, 
    7.480609e+09, 7.476158e+09, 7.470226e+09, 7.462817e+09, 7.453934e+09, 
    7.443579e+09, 7.431758e+09, 7.418477e+09, 7.403741e+09, 7.387556e+09, 
    7.36993e+09, 7.350871e+09, 7.330385e+09, 7.308484e+09, 7.285175e+09, 
    7.260469e+09, 7.234377e+09, 7.206909e+09, 7.178077e+09, 7.147894e+09, 
    7.116371e+09, 7.083523e+09, 7.049361e+09, 7.013901e+09, 6.977157e+09, 
    6.939143e+09, 6.899874e+09, 6.859367e+09, 6.817636e+09, 6.774699e+09, 
    6.730571e+09, 6.685269e+09, 6.638811e+09, 6.591213e+09, 6.542493e+09, 
    6.492669e+09, 6.441759e+09, 6.38978e+09, 6.336752e+09, 6.282692e+09, 
    6.227619e+09, 6.171552e+09, 6.114508e+09, 6.056508e+09, 5.99757e+09, 
    5.937712e+09,
  5.988909e+09, 6.052155e+09, 6.114508e+09, 6.175945e+09, 6.236442e+09, 
    6.295976e+09, 6.354524e+09, 6.412062e+09, 6.468569e+09, 6.52402e+09, 
    6.578392e+09, 6.631664e+09, 6.683811e+09, 6.734811e+09, 6.784643e+09, 
    6.833284e+09, 6.880711e+09, 6.926904e+09, 6.971842e+09, 7.015503e+09, 
    7.057866e+09, 7.098912e+09, 7.13862e+09, 7.176973e+09, 7.21395e+09, 
    7.249533e+09, 7.283705e+09, 7.316448e+09, 7.347746e+09, 7.377583e+09, 
    7.405943e+09, 7.432813e+09, 7.458176e+09, 7.482021e+09, 7.504335e+09, 
    7.525106e+09, 7.544322e+09, 7.561974e+09, 7.578052e+09, 7.592547e+09, 
    7.605452e+09, 7.616759e+09, 7.626462e+09, 7.634556e+09, 7.641037e+09, 
    7.645901e+09, 7.649145e+09, 7.650767e+09, 7.650767e+09, 7.649145e+09, 
    7.645901e+09, 7.641037e+09, 7.634556e+09, 7.626462e+09, 7.616759e+09, 
    7.605452e+09, 7.592547e+09, 7.578052e+09, 7.561974e+09, 7.544322e+09, 
    7.525106e+09, 7.504335e+09, 7.482021e+09, 7.458176e+09, 7.432813e+09, 
    7.405943e+09, 7.377583e+09, 7.347746e+09, 7.316448e+09, 7.283705e+09, 
    7.249533e+09, 7.21395e+09, 7.176973e+09, 7.13862e+09, 7.098912e+09, 
    7.057866e+09, 7.015503e+09, 6.971842e+09, 6.926904e+09, 6.880711e+09, 
    6.833284e+09, 6.784643e+09, 6.734811e+09, 6.683811e+09, 6.631664e+09, 
    6.578392e+09, 6.52402e+09, 6.468569e+09, 6.412062e+09, 6.354524e+09, 
    6.295976e+09, 6.236442e+09, 6.175945e+09, 6.114508e+09, 6.052155e+09, 
    5.988909e+09,
  6.039129e+09, 6.105772e+09, 6.171552e+09, 6.236442e+09, 6.300414e+09, 
    6.363442e+09, 6.425497e+09, 6.486551e+09, 6.546576e+09, 6.605544e+09, 
    6.663429e+09, 6.720201e+09, 6.775833e+09, 6.830297e+09, 6.883567e+09, 
    6.935614e+09, 6.986412e+09, 7.035934e+09, 7.084154e+09, 7.131045e+09, 
    7.176583e+09, 7.220742e+09, 7.263496e+09, 7.304823e+09, 7.344698e+09, 
    7.383099e+09, 7.420003e+09, 7.455388e+09, 7.489233e+09, 7.521518e+09, 
    7.552224e+09, 7.581331e+09, 7.608822e+09, 7.634681e+09, 7.65889e+09, 
    7.681435e+09, 7.702302e+09, 7.721477e+09, 7.738948e+09, 7.754704e+09, 
    7.768736e+09, 7.781033e+09, 7.791588e+09, 7.800395e+09, 7.807448e+09, 
    7.812741e+09, 7.816271e+09, 7.818037e+09, 7.818037e+09, 7.816271e+09, 
    7.812741e+09, 7.807448e+09, 7.800395e+09, 7.791588e+09, 7.781033e+09, 
    7.768736e+09, 7.754704e+09, 7.738948e+09, 7.721477e+09, 7.702302e+09, 
    7.681435e+09, 7.65889e+09, 7.634681e+09, 7.608822e+09, 7.581331e+09, 
    7.552224e+09, 7.521518e+09, 7.489233e+09, 7.455388e+09, 7.420003e+09, 
    7.383099e+09, 7.344698e+09, 7.304823e+09, 7.263496e+09, 7.220742e+09, 
    7.176583e+09, 7.131045e+09, 7.084154e+09, 7.035934e+09, 6.986412e+09, 
    6.935614e+09, 6.883567e+09, 6.830297e+09, 6.775833e+09, 6.720201e+09, 
    6.663429e+09, 6.605544e+09, 6.546576e+09, 6.486551e+09, 6.425497e+09, 
    6.363442e+09, 6.300414e+09, 6.236442e+09, 6.171552e+09, 6.105772e+09, 
    6.039129e+09,
  6.088361e+09, 6.158404e+09, 6.227619e+09, 6.295976e+09, 6.363442e+09, 
    6.429985e+09, 6.495574e+09, 6.560175e+09, 6.623755e+09, 6.686283e+09, 
    6.747724e+09, 6.808046e+09, 6.867216e+09, 6.925201e+09, 6.981969e+09, 
    7.037487e+09, 7.091722e+09, 7.144643e+09, 7.196217e+09, 7.246414e+09, 
    7.295202e+09, 7.342552e+09, 7.388432e+09, 7.432814e+09, 7.475667e+09, 
    7.516966e+09, 7.556683e+09, 7.594789e+09, 7.631261e+09, 7.666072e+09, 
    7.699199e+09, 7.73062e+09, 7.760311e+09, 7.788252e+09, 7.814423e+09, 
    7.838806e+09, 7.861382e+09, 7.882135e+09, 7.901051e+09, 7.918115e+09, 
    7.933316e+09, 7.946641e+09, 7.958081e+09, 7.967627e+09, 7.975273e+09, 
    7.981012e+09, 7.984841e+09, 7.986756e+09, 7.986756e+09, 7.984841e+09, 
    7.981012e+09, 7.975273e+09, 7.967627e+09, 7.958081e+09, 7.946641e+09, 
    7.933316e+09, 7.918115e+09, 7.901051e+09, 7.882135e+09, 7.861382e+09, 
    7.838806e+09, 7.814423e+09, 7.788252e+09, 7.760311e+09, 7.73062e+09, 
    7.699199e+09, 7.666072e+09, 7.631261e+09, 7.594789e+09, 7.556683e+09, 
    7.516966e+09, 7.475667e+09, 7.432814e+09, 7.388432e+09, 7.342552e+09, 
    7.295202e+09, 7.246414e+09, 7.196217e+09, 7.144643e+09, 7.091722e+09, 
    7.037487e+09, 6.981969e+09, 6.925201e+09, 6.867216e+09, 6.808046e+09, 
    6.747724e+09, 6.686283e+09, 6.623755e+09, 6.560175e+09, 6.495574e+09, 
    6.429985e+09, 6.363442e+09, 6.295976e+09, 6.227619e+09, 6.158404e+09, 
    6.088361e+09,
  6.136596e+09, 6.210038e+09, 6.282692e+09, 6.354524e+09, 6.425497e+09, 
    6.495574e+09, 6.564719e+09, 6.632894e+09, 6.700061e+09, 6.766183e+09, 
    6.831222e+09, 6.895139e+09, 6.957896e+09, 7.019455e+09, 7.079777e+09, 
    7.138825e+09, 7.196561e+09, 7.252946e+09, 7.307944e+09, 7.361518e+09, 
    7.41363e+09, 7.464245e+09, 7.513327e+09, 7.56084e+09, 7.606751e+09, 
    7.651027e+09, 7.693634e+09, 7.734541e+09, 7.773715e+09, 7.811129e+09, 
    7.846753e+09, 7.880559e+09, 7.912521e+09, 7.942612e+09, 7.970811e+09, 
    7.997093e+09, 8.021437e+09, 8.043825e+09, 8.064236e+09, 8.082655e+09, 
    8.099066e+09, 8.113456e+09, 8.125813e+09, 8.136126e+09, 8.144387e+09, 
    8.150589e+09, 8.154726e+09, 8.156796e+09, 8.156796e+09, 8.154726e+09, 
    8.150589e+09, 8.144387e+09, 8.136126e+09, 8.125813e+09, 8.113456e+09, 
    8.099066e+09, 8.082655e+09, 8.064236e+09, 8.043825e+09, 8.021437e+09, 
    7.997093e+09, 7.970811e+09, 7.942612e+09, 7.912521e+09, 7.880559e+09, 
    7.846753e+09, 7.811129e+09, 7.773715e+09, 7.734541e+09, 7.693634e+09, 
    7.651027e+09, 7.606751e+09, 7.56084e+09, 7.513327e+09, 7.464245e+09, 
    7.41363e+09, 7.361518e+09, 7.307944e+09, 7.252946e+09, 7.196561e+09, 
    7.138825e+09, 7.079777e+09, 7.019455e+09, 6.957896e+09, 6.895139e+09, 
    6.831222e+09, 6.766183e+09, 6.700061e+09, 6.632894e+09, 6.564719e+09, 
    6.495574e+09, 6.425497e+09, 6.354524e+09, 6.282692e+09, 6.210038e+09, 
    6.136596e+09,
  6.183825e+09, 6.260659e+09, 6.336752e+09, 6.412062e+09, 6.486551e+09, 
    6.560175e+09, 6.632894e+09, 6.704666e+09, 6.775447e+09, 6.845195e+09, 
    6.913867e+09, 6.981418e+09, 7.047806e+09, 7.112987e+09, 7.176916e+09, 
    7.23955e+09, 7.300845e+09, 7.360757e+09, 7.419243e+09, 7.47626e+09, 
    7.531766e+09, 7.585717e+09, 7.638074e+09, 7.688794e+09, 7.737838e+09, 
    7.785166e+09, 7.830739e+09, 7.874522e+09, 7.916475e+09, 7.956566e+09, 
    7.994759e+09, 8.031022e+09, 8.065324e+09, 8.097633e+09, 8.127923e+09, 
    8.156166e+09, 8.182336e+09, 8.20641e+09, 8.228367e+09, 8.248187e+09, 
    8.26585e+09, 8.281342e+09, 8.294647e+09, 8.305754e+09, 8.314652e+09, 
    8.321333e+09, 8.32579e+09, 8.32802e+09, 8.32802e+09, 8.32579e+09, 
    8.321333e+09, 8.314652e+09, 8.305754e+09, 8.294647e+09, 8.281342e+09, 
    8.26585e+09, 8.248187e+09, 8.228367e+09, 8.20641e+09, 8.182336e+09, 
    8.156166e+09, 8.127923e+09, 8.097633e+09, 8.065324e+09, 8.031022e+09, 
    7.994759e+09, 7.956566e+09, 7.916475e+09, 7.874522e+09, 7.830739e+09, 
    7.785166e+09, 7.737838e+09, 7.688794e+09, 7.638074e+09, 7.585717e+09, 
    7.531766e+09, 7.47626e+09, 7.419243e+09, 7.360757e+09, 7.300845e+09, 
    7.23955e+09, 7.176916e+09, 7.112987e+09, 7.047806e+09, 6.981418e+09, 
    6.913867e+09, 6.845195e+09, 6.775447e+09, 6.704666e+09, 6.632894e+09, 
    6.560175e+09, 6.486551e+09, 6.412062e+09, 6.336752e+09, 6.260659e+09, 
    6.183825e+09,
  6.230037e+09, 6.310255e+09, 6.38978e+09, 6.468569e+09, 6.546576e+09, 
    6.623755e+09, 6.700061e+09, 6.775447e+09, 6.849864e+09, 6.923265e+09, 
    6.9956e+09, 7.066822e+09, 7.136881e+09, 7.205726e+09, 7.273309e+09, 
    7.339579e+09, 7.404488e+09, 7.467984e+09, 7.530018e+09, 7.590542e+09, 
    7.649507e+09, 7.706863e+09, 7.762563e+09, 7.816561e+09, 7.868808e+09, 
    7.919261e+09, 7.967875e+09, 8.014606e+09, 8.059411e+09, 8.10225e+09, 
    8.143084e+09, 8.181873e+09, 8.218582e+09, 8.253174e+09, 8.285618e+09, 
    8.31588e+09, 8.343933e+09, 8.369748e+09, 8.3933e+09, 8.414565e+09, 
    8.433522e+09, 8.450151e+09, 8.464436e+09, 8.476363e+09, 8.485919e+09, 
    8.493095e+09, 8.497883e+09, 8.500278e+09, 8.500278e+09, 8.497883e+09, 
    8.493095e+09, 8.485919e+09, 8.476363e+09, 8.464436e+09, 8.450151e+09, 
    8.433522e+09, 8.414565e+09, 8.3933e+09, 8.369748e+09, 8.343933e+09, 
    8.31588e+09, 8.285618e+09, 8.253174e+09, 8.218582e+09, 8.181873e+09, 
    8.143084e+09, 8.10225e+09, 8.059411e+09, 8.014606e+09, 7.967875e+09, 
    7.919261e+09, 7.868808e+09, 7.816561e+09, 7.762563e+09, 7.706863e+09, 
    7.649507e+09, 7.590542e+09, 7.530018e+09, 7.467984e+09, 7.404488e+09, 
    7.339579e+09, 7.273309e+09, 7.205726e+09, 7.136881e+09, 7.066822e+09, 
    6.9956e+09, 6.923265e+09, 6.849864e+09, 6.775447e+09, 6.700061e+09, 
    6.623755e+09, 6.546576e+09, 6.468569e+09, 6.38978e+09, 6.310255e+09, 
    6.230037e+09,
  6.275223e+09, 6.35881e+09, 6.441759e+09, 6.52402e+09, 6.605544e+09, 
    6.686283e+09, 6.766183e+09, 6.845195e+09, 6.923265e+09, 7.000339e+09, 
    7.076365e+09, 7.151286e+09, 7.225049e+09, 7.297597e+09, 7.368877e+09, 
    7.438829e+09, 7.5074e+09, 7.574533e+09, 7.640172e+09, 7.704261e+09, 
    7.766745e+09, 7.827569e+09, 7.886679e+09, 7.94402e+09, 7.99954e+09, 
    8.053188e+09, 8.10491e+09, 8.15466e+09, 8.202386e+09, 8.248043e+09, 
    8.291585e+09, 8.332967e+09, 8.372148e+09, 8.409087e+09, 8.443745e+09, 
    8.476086e+09, 8.506077e+09, 8.533684e+09, 8.558878e+09, 8.581632e+09, 
    8.601922e+09, 8.619724e+09, 8.63502e+09, 8.647793e+09, 8.658028e+09, 
    8.665715e+09, 8.670843e+09, 8.673409e+09, 8.673409e+09, 8.670843e+09, 
    8.665715e+09, 8.658028e+09, 8.647793e+09, 8.63502e+09, 8.619724e+09, 
    8.601922e+09, 8.581632e+09, 8.558878e+09, 8.533684e+09, 8.506077e+09, 
    8.476086e+09, 8.443745e+09, 8.409087e+09, 8.372148e+09, 8.332967e+09, 
    8.291585e+09, 8.248043e+09, 8.202386e+09, 8.15466e+09, 8.10491e+09, 
    8.053188e+09, 7.99954e+09, 7.94402e+09, 7.886679e+09, 7.827569e+09, 
    7.766745e+09, 7.704261e+09, 7.640172e+09, 7.574533e+09, 7.5074e+09, 
    7.438829e+09, 7.368877e+09, 7.297597e+09, 7.225049e+09, 7.151286e+09, 
    7.076365e+09, 7.000339e+09, 6.923265e+09, 6.845195e+09, 6.766183e+09, 
    6.686283e+09, 6.605544e+09, 6.52402e+09, 6.441759e+09, 6.35881e+09, 
    6.275223e+09,
  6.319373e+09, 6.406312e+09, 6.492669e+09, 6.578392e+09, 6.663429e+09, 
    6.747724e+09, 6.831222e+09, 6.913867e+09, 6.9956e+09, 7.076365e+09, 
    7.1561e+09, 7.234745e+09, 7.312241e+09, 7.388526e+09, 7.463537e+09, 
    7.537212e+09, 7.60949e+09, 7.680307e+09, 7.749601e+09, 7.817309e+09, 
    7.883369e+09, 7.94772e+09, 8.010299e+09, 8.071048e+09, 8.129904e+09, 
    8.186811e+09, 8.241709e+09, 8.294543e+09, 8.345257e+09, 8.393798e+09, 
    8.440113e+09, 8.484152e+09, 8.525868e+09, 8.565214e+09, 8.602145e+09, 
    8.636621e+09, 8.668601e+09, 8.698051e+09, 8.724934e+09, 8.749221e+09, 
    8.770882e+09, 8.789891e+09, 8.806228e+09, 8.819871e+09, 8.830806e+09, 
    8.839017e+09, 8.844498e+09, 8.84724e+09, 8.84724e+09, 8.844498e+09, 
    8.839017e+09, 8.830806e+09, 8.819871e+09, 8.806228e+09, 8.789891e+09, 
    8.770882e+09, 8.749221e+09, 8.724934e+09, 8.698051e+09, 8.668601e+09, 
    8.636621e+09, 8.602145e+09, 8.565214e+09, 8.525868e+09, 8.484152e+09, 
    8.440113e+09, 8.393798e+09, 8.345257e+09, 8.294543e+09, 8.241709e+09, 
    8.186811e+09, 8.129904e+09, 8.071048e+09, 8.010299e+09, 7.94772e+09, 
    7.883369e+09, 7.817309e+09, 7.749601e+09, 7.680307e+09, 7.60949e+09, 
    7.537212e+09, 7.463537e+09, 7.388526e+09, 7.312241e+09, 7.234745e+09, 
    7.1561e+09, 7.076365e+09, 6.9956e+09, 6.913867e+09, 6.831222e+09, 
    6.747724e+09, 6.663429e+09, 6.578392e+09, 6.492669e+09, 6.406312e+09, 
    6.319373e+09,
  6.362479e+09, 6.452746e+09, 6.542493e+09, 6.631664e+09, 6.720201e+09, 
    6.808046e+09, 6.895139e+09, 6.981418e+09, 7.066822e+09, 7.151286e+09, 
    7.234745e+09, 7.317134e+09, 7.398386e+09, 7.478433e+09, 7.557208e+09, 
    7.634641e+09, 7.710664e+09, 7.785207e+09, 7.858201e+09, 7.929576e+09, 
    7.999264e+09, 8.067195e+09, 8.133301e+09, 8.197513e+09, 8.259766e+09, 
    8.319992e+09, 8.378128e+09, 8.434108e+09, 8.487873e+09, 8.539359e+09, 
    8.58851e+09, 8.635267e+09, 8.679578e+09, 8.721389e+09, 8.760649e+09, 
    8.797313e+09, 8.831335e+09, 8.862674e+09, 8.891291e+09, 8.917151e+09, 
    8.940219e+09, 8.96047e+09, 8.977876e+09, 8.992415e+09, 9.004068e+09, 
    9.012821e+09, 9.018663e+09, 9.021585e+09, 9.021585e+09, 9.018663e+09, 
    9.012821e+09, 9.004068e+09, 8.992415e+09, 8.977876e+09, 8.96047e+09, 
    8.940219e+09, 8.917151e+09, 8.891291e+09, 8.862674e+09, 8.831335e+09, 
    8.797313e+09, 8.760649e+09, 8.721389e+09, 8.679578e+09, 8.635267e+09, 
    8.58851e+09, 8.539359e+09, 8.487873e+09, 8.434108e+09, 8.378128e+09, 
    8.319992e+09, 8.259766e+09, 8.197513e+09, 8.133301e+09, 8.067195e+09, 
    7.999264e+09, 7.929576e+09, 7.858201e+09, 7.785207e+09, 7.710664e+09, 
    7.634641e+09, 7.557208e+09, 7.478433e+09, 7.398386e+09, 7.317134e+09, 
    7.234745e+09, 7.151286e+09, 7.066822e+09, 6.981418e+09, 6.895139e+09, 
    6.808046e+09, 6.720201e+09, 6.631664e+09, 6.542493e+09, 6.452746e+09, 
    6.362479e+09,
  6.404531e+09, 6.4981e+09, 6.591213e+09, 6.683811e+09, 6.775833e+09, 
    6.867216e+09, 6.957896e+09, 7.047806e+09, 7.136881e+09, 7.225049e+09, 
    7.312241e+09, 7.398386e+09, 7.483411e+09, 7.567242e+09, 7.649805e+09, 
    7.731025e+09, 7.810825e+09, 7.889131e+09, 7.965864e+09, 8.04095e+09, 
    8.11431e+09, 8.18587e+09, 8.255552e+09, 8.323282e+09, 8.388985e+09, 
    8.452588e+09, 8.514017e+09, 8.573202e+09, 8.630074e+09, 8.684566e+09, 
    8.736609e+09, 8.786142e+09, 8.833104e+09, 8.877434e+09, 8.919077e+09, 
    8.95798e+09, 8.994092e+09, 9.027367e+09, 9.05776e+09, 9.085231e+09, 
    9.109745e+09, 9.131267e+09, 9.14977e+09, 9.165227e+09, 9.177618e+09, 
    9.186927e+09, 9.193139e+09, 9.196247e+09, 9.196247e+09, 9.193139e+09, 
    9.186927e+09, 9.177618e+09, 9.165227e+09, 9.14977e+09, 9.131267e+09, 
    9.109745e+09, 9.085231e+09, 9.05776e+09, 9.027367e+09, 8.994092e+09, 
    8.95798e+09, 8.919077e+09, 8.877434e+09, 8.833104e+09, 8.786142e+09, 
    8.736609e+09, 8.684566e+09, 8.630074e+09, 8.573202e+09, 8.514017e+09, 
    8.452588e+09, 8.388985e+09, 8.323282e+09, 8.255552e+09, 8.18587e+09, 
    8.11431e+09, 8.04095e+09, 7.965864e+09, 7.889131e+09, 7.810825e+09, 
    7.731025e+09, 7.649805e+09, 7.567242e+09, 7.483411e+09, 7.398386e+09, 
    7.312241e+09, 7.225049e+09, 7.136881e+09, 7.047806e+09, 6.957896e+09, 
    6.867216e+09, 6.775833e+09, 6.683811e+09, 6.591213e+09, 6.4981e+09, 
    6.404531e+09,
  6.445522e+09, 6.54236e+09, 6.638811e+09, 6.734811e+09, 6.830297e+09, 
    6.925201e+09, 7.019455e+09, 7.112987e+09, 7.205726e+09, 7.297597e+09, 
    7.388526e+09, 7.478433e+09, 7.567242e+09, 7.654872e+09, 7.741242e+09, 
    7.826271e+09, 7.909876e+09, 7.991974e+09, 8.072481e+09, 8.151313e+09, 
    8.228386e+09, 8.303616e+09, 8.37692e+09, 8.448214e+09, 8.517416e+09, 
    8.584445e+09, 8.649221e+09, 8.711665e+09, 8.771699e+09, 8.829247e+09, 
    8.884238e+09, 8.936601e+09, 8.986266e+09, 9.033167e+09, 9.077242e+09, 
    9.118431e+09, 9.156679e+09, 9.191932e+09, 9.224142e+09, 9.253263e+09, 
    9.279254e+09, 9.302078e+09, 9.321703e+09, 9.338102e+09, 9.351248e+09, 
    9.361125e+09, 9.367718e+09, 9.371016e+09, 9.371016e+09, 9.367718e+09, 
    9.361125e+09, 9.351248e+09, 9.338102e+09, 9.321703e+09, 9.302078e+09, 
    9.279254e+09, 9.253263e+09, 9.224142e+09, 9.191932e+09, 9.156679e+09, 
    9.118431e+09, 9.077242e+09, 9.033167e+09, 8.986266e+09, 8.936601e+09, 
    8.884238e+09, 8.829247e+09, 8.771699e+09, 8.711665e+09, 8.649221e+09, 
    8.584445e+09, 8.517416e+09, 8.448214e+09, 8.37692e+09, 8.303616e+09, 
    8.228386e+09, 8.151313e+09, 8.072481e+09, 7.991974e+09, 7.909876e+09, 
    7.826271e+09, 7.741242e+09, 7.654872e+09, 7.567242e+09, 7.478433e+09, 
    7.388526e+09, 7.297597e+09, 7.205726e+09, 7.112987e+09, 7.019455e+09, 
    6.925201e+09, 6.830297e+09, 6.734811e+09, 6.638811e+09, 6.54236e+09, 
    6.445522e+09,
  6.485442e+09, 6.585513e+09, 6.685269e+09, 6.784643e+09, 6.883567e+09, 
    6.981969e+09, 7.079777e+09, 7.176916e+09, 7.273309e+09, 7.368877e+09, 
    7.463537e+09, 7.557208e+09, 7.649805e+09, 7.741242e+09, 7.831433e+09, 
    7.920287e+09, 8.007716e+09, 8.093629e+09, 8.177936e+09, 8.260545e+09, 
    8.341364e+09, 8.420301e+09, 8.497266e+09, 8.572165e+09, 8.64491e+09, 
    8.715411e+09, 8.78358e+09, 8.849328e+09, 8.912572e+09, 8.973229e+09, 
    9.031216e+09, 9.086456e+09, 9.138871e+09, 9.188391e+09, 9.234944e+09, 
    9.278465e+09, 9.318892e+09, 9.356163e+09, 9.390226e+09, 9.421031e+09, 
    9.448532e+09, 9.472687e+09, 9.49346e+09, 9.510819e+09, 9.524738e+09, 
    9.535196e+09, 9.542177e+09, 9.54567e+09, 9.54567e+09, 9.542177e+09, 
    9.535196e+09, 9.524738e+09, 9.510819e+09, 9.49346e+09, 9.472687e+09, 
    9.448532e+09, 9.421031e+09, 9.390226e+09, 9.356163e+09, 9.318892e+09, 
    9.278465e+09, 9.234944e+09, 9.188391e+09, 9.138871e+09, 9.086456e+09, 
    9.031216e+09, 8.973229e+09, 8.912572e+09, 8.849328e+09, 8.78358e+09, 
    8.715411e+09, 8.64491e+09, 8.572165e+09, 8.497266e+09, 8.420301e+09, 
    8.341364e+09, 8.260545e+09, 8.177936e+09, 8.093629e+09, 8.007716e+09, 
    7.920287e+09, 7.831433e+09, 7.741242e+09, 7.649805e+09, 7.557208e+09, 
    7.463537e+09, 7.368877e+09, 7.273309e+09, 7.176916e+09, 7.079777e+09, 
    6.981969e+09, 6.883567e+09, 6.784643e+09, 6.685269e+09, 6.585513e+09, 
    6.485442e+09,
  6.524282e+09, 6.627547e+09, 6.730571e+09, 6.833284e+09, 6.935614e+09, 
    7.037487e+09, 7.138825e+09, 7.23955e+09, 7.339579e+09, 7.438829e+09, 
    7.537212e+09, 7.634641e+09, 7.731025e+09, 7.826271e+09, 7.920287e+09, 
    8.012976e+09, 8.104243e+09, 8.193989e+09, 8.282116e+09, 8.368525e+09, 
    8.453116e+09, 8.53579e+09, 8.616447e+09, 8.694987e+09, 8.771312e+09, 
    8.845323e+09, 8.916924e+09, 8.986021e+09, 9.052518e+09, 9.116325e+09, 
    9.177352e+09, 9.235513e+09, 9.290724e+09, 9.342905e+09, 9.391978e+09, 
    9.437871e+09, 9.480515e+09, 9.519842e+09, 9.555794e+09, 9.588315e+09, 
    9.617354e+09, 9.642865e+09, 9.664807e+09, 9.683147e+09, 9.697854e+09, 
    9.708905e+09, 9.716282e+09, 9.719975e+09, 9.719975e+09, 9.716282e+09, 
    9.708905e+09, 9.697854e+09, 9.683147e+09, 9.664807e+09, 9.642865e+09, 
    9.617354e+09, 9.588315e+09, 9.555794e+09, 9.519842e+09, 9.480515e+09, 
    9.437871e+09, 9.391978e+09, 9.342905e+09, 9.290724e+09, 9.235513e+09, 
    9.177352e+09, 9.116325e+09, 9.052518e+09, 8.986021e+09, 8.916924e+09, 
    8.845323e+09, 8.771312e+09, 8.694987e+09, 8.616447e+09, 8.53579e+09, 
    8.453116e+09, 8.368525e+09, 8.282116e+09, 8.193989e+09, 8.104243e+09, 
    8.012976e+09, 7.920287e+09, 7.826271e+09, 7.731025e+09, 7.634641e+09, 
    7.537212e+09, 7.438829e+09, 7.339579e+09, 7.23955e+09, 7.138825e+09, 
    7.037487e+09, 6.935614e+09, 6.833284e+09, 6.730571e+09, 6.627547e+09, 
    6.524282e+09,
  6.562035e+09, 6.668449e+09, 6.774699e+09, 6.880711e+09, 6.986412e+09, 
    7.091722e+09, 7.196561e+09, 7.300845e+09, 7.404488e+09, 7.5074e+09, 
    7.60949e+09, 7.710664e+09, 7.810825e+09, 7.909876e+09, 8.007716e+09, 
    8.104243e+09, 8.199353e+09, 8.292941e+09, 8.384902e+09, 8.475127e+09, 
    8.563511e+09, 8.649944e+09, 8.734319e+09, 8.816526e+09, 8.896461e+09, 
    8.974015e+09, 9.049084e+09, 9.121564e+09, 9.191351e+09, 9.258346e+09, 
    9.322452e+09, 9.383574e+09, 9.441618e+09, 9.496498e+09, 9.548129e+09, 
    9.596429e+09, 9.641325e+09, 9.68274e+09, 9.720613e+09, 9.754878e+09, 
    9.785482e+09, 9.812372e+09, 9.835507e+09, 9.854844e+09, 9.870353e+09, 
    9.882009e+09, 9.88979e+09, 9.893683e+09, 9.893683e+09, 9.88979e+09, 
    9.882009e+09, 9.870353e+09, 9.854844e+09, 9.835507e+09, 9.812372e+09, 
    9.785482e+09, 9.754878e+09, 9.720613e+09, 9.68274e+09, 9.641325e+09, 
    9.596429e+09, 9.548129e+09, 9.496498e+09, 9.441618e+09, 9.383574e+09, 
    9.322452e+09, 9.258346e+09, 9.191351e+09, 9.121564e+09, 9.049084e+09, 
    8.974015e+09, 8.896461e+09, 8.816526e+09, 8.734319e+09, 8.649944e+09, 
    8.563511e+09, 8.475127e+09, 8.384902e+09, 8.292941e+09, 8.199353e+09, 
    8.104243e+09, 8.007716e+09, 7.909876e+09, 7.810825e+09, 7.710664e+09, 
    7.60949e+09, 7.5074e+09, 7.404488e+09, 7.300845e+09, 7.196561e+09, 
    7.091722e+09, 6.986412e+09, 6.880711e+09, 6.774699e+09, 6.668449e+09, 
    6.562035e+09,
  6.598693e+09, 6.708208e+09, 6.817636e+09, 6.926904e+09, 7.035934e+09, 
    7.144643e+09, 7.252946e+09, 7.360757e+09, 7.467984e+09, 7.574533e+09, 
    7.680307e+09, 7.785207e+09, 7.889131e+09, 7.991974e+09, 8.093629e+09, 
    8.193989e+09, 8.292941e+09, 8.390374e+09, 8.486173e+09, 8.580225e+09, 
    8.672412e+09, 8.762619e+09, 8.85073e+09, 8.936627e+09, 9.020195e+09, 
    9.101317e+09, 9.17988e+09, 9.255772e+09, 9.32888e+09, 9.399095e+09, 
    9.466312e+09, 9.530426e+09, 9.591338e+09, 9.64895e+09, 9.703171e+09, 
    9.753911e+09, 9.801088e+09, 9.844622e+09, 9.884442e+09, 9.920478e+09, 
    9.95267e+09, 9.980962e+09, 1.00053e+10, 1.002566e+10, 1.004198e+10, 
    1.005425e+10, 1.006244e+10, 1.006654e+10, 1.006654e+10, 1.006244e+10, 
    1.005425e+10, 1.004198e+10, 1.002566e+10, 1.00053e+10, 9.980962e+09, 
    9.95267e+09, 9.920478e+09, 9.884442e+09, 9.844622e+09, 9.801088e+09, 
    9.753911e+09, 9.703171e+09, 9.64895e+09, 9.591338e+09, 9.530426e+09, 
    9.466312e+09, 9.399095e+09, 9.32888e+09, 9.255772e+09, 9.17988e+09, 
    9.101317e+09, 9.020195e+09, 8.936627e+09, 8.85073e+09, 8.762619e+09, 
    8.672412e+09, 8.580225e+09, 8.486173e+09, 8.390374e+09, 8.292941e+09, 
    8.193989e+09, 8.093629e+09, 7.991974e+09, 7.889131e+09, 7.785207e+09, 
    7.680307e+09, 7.574533e+09, 7.467984e+09, 7.360757e+09, 7.252946e+09, 
    7.144643e+09, 7.035934e+09, 6.926904e+09, 6.817636e+09, 6.708208e+09, 
    6.598693e+09,
  6.634248e+09, 6.74681e+09, 6.859367e+09, 6.971842e+09, 7.084154e+09, 
    7.196217e+09, 7.307944e+09, 7.419243e+09, 7.530018e+09, 7.640172e+09, 
    7.749601e+09, 7.858201e+09, 7.965864e+09, 8.072481e+09, 8.177936e+09, 
    8.282116e+09, 8.384902e+09, 8.486173e+09, 8.585809e+09, 8.683688e+09, 
    8.779684e+09, 8.873673e+09, 8.96553e+09, 9.055129e+09, 9.142345e+09, 
    9.227054e+09, 9.309132e+09, 9.388457e+09, 9.464909e+09, 9.53837e+09, 
    9.608722e+09, 9.675857e+09, 9.739662e+09, 9.800034e+09, 9.856871e+09, 
    9.910078e+09, 9.959563e+09, 1.000524e+10, 1.004703e+10, 1.008486e+10, 
    1.011866e+10, 1.014837e+10, 1.017394e+10, 1.019532e+10, 1.021247e+10, 
    1.022536e+10, 1.023397e+10, 1.023827e+10, 1.023827e+10, 1.023397e+10, 
    1.022536e+10, 1.021247e+10, 1.019532e+10, 1.017394e+10, 1.014837e+10, 
    1.011866e+10, 1.008486e+10, 1.004703e+10, 1.000524e+10, 9.959563e+09, 
    9.910078e+09, 9.856871e+09, 9.800034e+09, 9.739662e+09, 9.675857e+09, 
    9.608722e+09, 9.53837e+09, 9.464909e+09, 9.388457e+09, 9.309132e+09, 
    9.227054e+09, 9.142345e+09, 9.055129e+09, 8.96553e+09, 8.873673e+09, 
    8.779684e+09, 8.683688e+09, 8.585809e+09, 8.486173e+09, 8.384902e+09, 
    8.282116e+09, 8.177936e+09, 8.072481e+09, 7.965864e+09, 7.858201e+09, 
    7.749601e+09, 7.640172e+09, 7.530018e+09, 7.419243e+09, 7.307944e+09, 
    7.196217e+09, 7.084154e+09, 6.971842e+09, 6.859367e+09, 6.74681e+09, 
    6.634248e+09,
  6.668692e+09, 6.784244e+09, 6.899874e+09, 7.015503e+09, 7.131045e+09, 
    7.246414e+09, 7.361518e+09, 7.47626e+09, 7.590542e+09, 7.704261e+09, 
    7.817309e+09, 7.929576e+09, 8.04095e+09, 8.151313e+09, 8.260545e+09, 
    8.368525e+09, 8.475127e+09, 8.580225e+09, 8.683688e+09, 8.785385e+09, 
    8.885187e+09, 8.982957e+09, 9.078562e+09, 9.171869e+09, 9.262742e+09, 
    9.351046e+09, 9.436652e+09, 9.519426e+09, 9.599237e+09, 9.67596e+09, 
    9.749469e+09, 9.819643e+09, 9.886363e+09, 9.949515e+09, 1.000899e+10, 
    1.006469e+10, 1.01165e+10, 1.016434e+10, 1.020812e+10, 1.024776e+10, 
    1.028319e+10, 1.031433e+10, 1.034114e+10, 1.036355e+10, 1.038154e+10, 
    1.039506e+10, 1.040409e+10, 1.040861e+10, 1.040861e+10, 1.040409e+10, 
    1.039506e+10, 1.038154e+10, 1.036355e+10, 1.034114e+10, 1.031433e+10, 
    1.028319e+10, 1.024776e+10, 1.020812e+10, 1.016434e+10, 1.01165e+10, 
    1.006469e+10, 1.000899e+10, 9.949515e+09, 9.886363e+09, 9.819643e+09, 
    9.749469e+09, 9.67596e+09, 9.599237e+09, 9.519426e+09, 9.436652e+09, 
    9.351046e+09, 9.262742e+09, 9.171869e+09, 9.078562e+09, 8.982957e+09, 
    8.885187e+09, 8.785385e+09, 8.683688e+09, 8.580225e+09, 8.475127e+09, 
    8.368525e+09, 8.260545e+09, 8.151313e+09, 8.04095e+09, 7.929576e+09, 
    7.817309e+09, 7.704261e+09, 7.590542e+09, 7.47626e+09, 7.361518e+09, 
    7.246414e+09, 7.131045e+09, 7.015503e+09, 6.899874e+09, 6.784244e+09, 
    6.668692e+09,
  6.702019e+09, 6.8205e+09, 6.939143e+09, 7.057866e+09, 7.176583e+09, 
    7.295202e+09, 7.41363e+09, 7.531766e+09, 7.649507e+09, 7.766745e+09, 
    7.883369e+09, 7.999264e+09, 8.11431e+09, 8.228386e+09, 8.341364e+09, 
    8.453116e+09, 8.563511e+09, 8.672412e+09, 8.779684e+09, 8.885187e+09, 
    8.988781e+09, 9.090322e+09, 9.18967e+09, 9.286681e+09, 9.381209e+09, 
    9.473112e+09, 9.562249e+09, 9.648477e+09, 9.731658e+09, 9.811654e+09, 
    9.88833e+09, 9.961556e+09, 1.00312e+10, 1.009715e+10, 1.015928e+10, 
    1.021748e+10, 1.027164e+10, 1.032166e+10, 1.036744e+10, 1.040891e+10, 
    1.044597e+10, 1.047856e+10, 1.050662e+10, 1.053008e+10, 1.054891e+10, 
    1.056306e+10, 1.057252e+10, 1.057725e+10, 1.057725e+10, 1.057252e+10, 
    1.056306e+10, 1.054891e+10, 1.053008e+10, 1.050662e+10, 1.047856e+10, 
    1.044597e+10, 1.040891e+10, 1.036744e+10, 1.032166e+10, 1.027164e+10, 
    1.021748e+10, 1.015928e+10, 1.009715e+10, 1.00312e+10, 9.961556e+09, 
    9.88833e+09, 9.811654e+09, 9.731658e+09, 9.648477e+09, 9.562249e+09, 
    9.473112e+09, 9.381209e+09, 9.286681e+09, 9.18967e+09, 9.090322e+09, 
    8.988781e+09, 8.885187e+09, 8.779684e+09, 8.672412e+09, 8.563511e+09, 
    8.453116e+09, 8.341364e+09, 8.228386e+09, 8.11431e+09, 7.999264e+09, 
    7.883369e+09, 7.766745e+09, 7.649507e+09, 7.531766e+09, 7.41363e+09, 
    7.295202e+09, 7.176583e+09, 7.057866e+09, 6.939143e+09, 6.8205e+09, 
    6.702019e+09,
  6.734221e+09, 6.855565e+09, 6.977157e+09, 7.098912e+09, 7.220742e+09, 
    7.342552e+09, 7.464245e+09, 7.585717e+09, 7.706863e+09, 7.827569e+09, 
    7.94772e+09, 8.067195e+09, 8.18587e+09, 8.303616e+09, 8.420301e+09, 
    8.53579e+09, 8.649944e+09, 8.762619e+09, 8.873673e+09, 8.982957e+09, 
    9.090322e+09, 9.195619e+09, 9.298694e+09, 9.399396e+09, 9.497571e+09, 
    9.593066e+09, 9.68573e+09, 9.775411e+09, 9.861961e+09, 9.945231e+09, 
    1.002508e+10, 1.010136e+10, 1.017395e+10, 1.02427e+10, 1.030749e+10, 
    1.03682e+10, 1.042471e+10, 1.047692e+10, 1.052472e+10, 1.056802e+10, 
    1.060673e+10, 1.064077e+10, 1.067009e+10, 1.06946e+10, 1.071428e+10, 
    1.072907e+10, 1.073895e+10, 1.07439e+10, 1.07439e+10, 1.073895e+10, 
    1.072907e+10, 1.071428e+10, 1.06946e+10, 1.067009e+10, 1.064077e+10, 
    1.060673e+10, 1.056802e+10, 1.052472e+10, 1.047692e+10, 1.042471e+10, 
    1.03682e+10, 1.030749e+10, 1.02427e+10, 1.017395e+10, 1.010136e+10, 
    1.002508e+10, 9.945231e+09, 9.861961e+09, 9.775411e+09, 9.68573e+09, 
    9.593066e+09, 9.497571e+09, 9.399396e+09, 9.298694e+09, 9.195619e+09, 
    9.090322e+09, 8.982957e+09, 8.873673e+09, 8.762619e+09, 8.649944e+09, 
    8.53579e+09, 8.420301e+09, 8.303616e+09, 8.18587e+09, 8.067195e+09, 
    7.94772e+09, 7.827569e+09, 7.706863e+09, 7.585717e+09, 7.464245e+09, 
    7.342552e+09, 7.220742e+09, 7.098912e+09, 6.977157e+09, 6.855565e+09, 
    6.734221e+09,
  6.76529e+09, 6.889429e+09, 7.013901e+09, 7.13862e+09, 7.263496e+09, 
    7.388432e+09, 7.513327e+09, 7.638074e+09, 7.762563e+09, 7.886679e+09, 
    8.010299e+09, 8.133301e+09, 8.255552e+09, 8.37692e+09, 8.497266e+09, 
    8.616447e+09, 8.734319e+09, 8.85073e+09, 8.96553e+09, 9.078562e+09, 
    9.18967e+09, 9.298694e+09, 9.405474e+09, 9.509846e+09, 9.61165e+09, 
    9.710721e+09, 9.806899e+09, 9.900023e+09, 9.989933e+09, 1.007647e+10, 
    1.015949e+10, 1.023883e+10, 1.031435e+10, 1.03859e+10, 1.045336e+10, 
    1.051658e+10, 1.057545e+10, 1.062985e+10, 1.067967e+10, 1.07248e+10, 
    1.076517e+10, 1.080067e+10, 1.083124e+10, 1.085682e+10, 1.087735e+10, 
    1.089278e+10, 1.090309e+10, 1.090825e+10, 1.090825e+10, 1.090309e+10, 
    1.089278e+10, 1.087735e+10, 1.085682e+10, 1.083124e+10, 1.080067e+10, 
    1.076517e+10, 1.07248e+10, 1.067967e+10, 1.062985e+10, 1.057545e+10, 
    1.051658e+10, 1.045336e+10, 1.03859e+10, 1.031435e+10, 1.023883e+10, 
    1.015949e+10, 1.007647e+10, 9.989933e+09, 9.900023e+09, 9.806899e+09, 
    9.710721e+09, 9.61165e+09, 9.509846e+09, 9.405474e+09, 9.298694e+09, 
    9.18967e+09, 9.078562e+09, 8.96553e+09, 8.85073e+09, 8.734319e+09, 
    8.616447e+09, 8.497266e+09, 8.37692e+09, 8.255552e+09, 8.133301e+09, 
    8.010299e+09, 7.886679e+09, 7.762563e+09, 7.638074e+09, 7.513327e+09, 
    7.388432e+09, 7.263496e+09, 7.13862e+09, 7.013901e+09, 6.889429e+09, 
    6.76529e+09,
  6.795221e+09, 6.922081e+09, 7.049361e+09, 7.176973e+09, 7.304823e+09, 
    7.432814e+09, 7.56084e+09, 7.688794e+09, 7.816561e+09, 7.94402e+09, 
    8.071048e+09, 8.197513e+09, 8.323282e+09, 8.448214e+09, 8.572165e+09, 
    8.694987e+09, 8.816526e+09, 8.936627e+09, 9.055129e+09, 9.171869e+09, 
    9.286681e+09, 9.399396e+09, 9.509846e+09, 9.61786e+09, 9.723264e+09, 
    9.825887e+09, 9.925557e+09, 1.00221e+10, 1.011536e+10, 1.020515e+10, 
    1.029132e+10, 1.037371e+10, 1.045215e+10, 1.05265e+10, 1.059662e+10, 
    1.066235e+10, 1.072358e+10, 1.078017e+10, 1.0832e+10, 1.087898e+10, 
    1.092099e+10, 1.095795e+10, 1.098979e+10, 1.101642e+10, 1.10378e+10, 
    1.105388e+10, 1.106461e+10, 1.106999e+10, 1.106999e+10, 1.106461e+10, 
    1.105388e+10, 1.10378e+10, 1.101642e+10, 1.098979e+10, 1.095795e+10, 
    1.092099e+10, 1.087898e+10, 1.0832e+10, 1.078017e+10, 1.072358e+10, 
    1.066235e+10, 1.059662e+10, 1.05265e+10, 1.045215e+10, 1.037371e+10, 
    1.029132e+10, 1.020515e+10, 1.011536e+10, 1.00221e+10, 9.925557e+09, 
    9.825887e+09, 9.723264e+09, 9.61786e+09, 9.509846e+09, 9.399396e+09, 
    9.286681e+09, 9.171869e+09, 9.055129e+09, 8.936627e+09, 8.816526e+09, 
    8.694987e+09, 8.572165e+09, 8.448214e+09, 8.323282e+09, 8.197513e+09, 
    8.071048e+09, 7.94402e+09, 7.816561e+09, 7.688794e+09, 7.56084e+09, 
    7.432814e+09, 7.304823e+09, 7.176973e+09, 7.049361e+09, 6.922081e+09, 
    6.795221e+09,
  6.824007e+09, 6.953512e+09, 7.083523e+09, 7.21395e+09, 7.344698e+09, 
    7.475667e+09, 7.606751e+09, 7.737838e+09, 7.868808e+09, 7.99954e+09, 
    8.129904e+09, 8.259766e+09, 8.388985e+09, 8.517416e+09, 8.64491e+09, 
    8.771312e+09, 8.896461e+09, 9.020195e+09, 9.142345e+09, 9.262742e+09, 
    9.381209e+09, 9.497571e+09, 9.61165e+09, 9.723264e+09, 9.832232e+09, 
    9.938373e+09, 1.00415e+10, 1.014144e+10, 1.023802e+10, 1.033104e+10, 
    1.042034e+10, 1.050575e+10, 1.058711e+10, 1.066424e+10, 1.0737e+10, 
    1.080523e+10, 1.08688e+10, 1.092757e+10, 1.098142e+10, 1.103023e+10, 
    1.107389e+10, 1.111231e+10, 1.11454e+10, 1.117309e+10, 1.119532e+10, 
    1.121203e+10, 1.12232e+10, 1.122879e+10, 1.122879e+10, 1.12232e+10, 
    1.121203e+10, 1.119532e+10, 1.117309e+10, 1.11454e+10, 1.111231e+10, 
    1.107389e+10, 1.103023e+10, 1.098142e+10, 1.092757e+10, 1.08688e+10, 
    1.080523e+10, 1.0737e+10, 1.066424e+10, 1.058711e+10, 1.050575e+10, 
    1.042034e+10, 1.033104e+10, 1.023802e+10, 1.014144e+10, 1.00415e+10, 
    9.938373e+09, 9.832232e+09, 9.723264e+09, 9.61165e+09, 9.497571e+09, 
    9.381209e+09, 9.262742e+09, 9.142345e+09, 9.020195e+09, 8.896461e+09, 
    8.771312e+09, 8.64491e+09, 8.517416e+09, 8.388985e+09, 8.259766e+09, 
    8.129904e+09, 7.99954e+09, 7.868808e+09, 7.737838e+09, 7.606751e+09, 
    7.475667e+09, 7.344698e+09, 7.21395e+09, 7.083523e+09, 6.953512e+09, 
    6.824007e+09,
  6.851641e+09, 6.98371e+09, 7.116371e+09, 7.249533e+09, 7.383099e+09, 
    7.516966e+09, 7.651027e+09, 7.785166e+09, 7.919261e+09, 8.053188e+09, 
    8.186811e+09, 8.319992e+09, 8.452588e+09, 8.584445e+09, 8.715411e+09, 
    8.845323e+09, 8.974015e+09, 9.101317e+09, 9.227054e+09, 9.351046e+09, 
    9.473112e+09, 9.593066e+09, 9.710721e+09, 9.825887e+09, 9.938373e+09, 
    1.004799e+10, 1.015454e+10, 1.025783e+10, 1.035769e+10, 1.045391e+10, 
    1.054631e+10, 1.063472e+10, 1.071896e+10, 1.079885e+10, 1.087423e+10, 
    1.094495e+10, 1.101085e+10, 1.107179e+10, 1.112763e+10, 1.117826e+10, 
    1.122356e+10, 1.126342e+10, 1.129776e+10, 1.13265e+10, 1.134958e+10, 
    1.136693e+10, 1.137852e+10, 1.138432e+10, 1.138432e+10, 1.137852e+10, 
    1.136693e+10, 1.134958e+10, 1.13265e+10, 1.129776e+10, 1.126342e+10, 
    1.122356e+10, 1.117826e+10, 1.112763e+10, 1.107179e+10, 1.101085e+10, 
    1.094495e+10, 1.087423e+10, 1.079885e+10, 1.071896e+10, 1.063472e+10, 
    1.054631e+10, 1.045391e+10, 1.035769e+10, 1.025783e+10, 1.015454e+10, 
    1.004799e+10, 9.938373e+09, 9.825887e+09, 9.710721e+09, 9.593066e+09, 
    9.473112e+09, 9.351046e+09, 9.227054e+09, 9.101317e+09, 8.974015e+09, 
    8.845323e+09, 8.715411e+09, 8.584445e+09, 8.452588e+09, 8.319992e+09, 
    8.186811e+09, 8.053188e+09, 7.919261e+09, 7.785166e+09, 7.651027e+09, 
    7.516966e+09, 7.383099e+09, 7.249533e+09, 7.116371e+09, 6.98371e+09, 
    6.851641e+09,
  6.878117e+09, 7.012667e+09, 7.147894e+09, 7.283705e+09, 7.420003e+09, 
    7.556683e+09, 7.693634e+09, 7.830739e+09, 7.967875e+09, 8.10491e+09, 
    8.241709e+09, 8.378128e+09, 8.514017e+09, 8.649221e+09, 8.78358e+09, 
    8.916924e+09, 9.049084e+09, 9.17988e+09, 9.309132e+09, 9.436652e+09, 
    9.562249e+09, 9.68573e+09, 9.806899e+09, 9.925557e+09, 1.00415e+10, 
    1.015454e+10, 1.026446e+10, 1.037106e+10, 1.047415e+10, 1.057352e+10, 
    1.066899e+10, 1.076036e+10, 1.084745e+10, 1.093007e+10, 1.100805e+10, 
    1.108122e+10, 1.114942e+10, 1.12125e+10, 1.127033e+10, 1.132276e+10, 
    1.136968e+10, 1.141097e+10, 1.144656e+10, 1.147634e+10, 1.150025e+10, 
    1.151823e+10, 1.153025e+10, 1.153626e+10, 1.153626e+10, 1.153025e+10, 
    1.151823e+10, 1.150025e+10, 1.147634e+10, 1.144656e+10, 1.141097e+10, 
    1.136968e+10, 1.132276e+10, 1.127033e+10, 1.12125e+10, 1.114942e+10, 
    1.108122e+10, 1.100805e+10, 1.093007e+10, 1.084745e+10, 1.076036e+10, 
    1.066899e+10, 1.057352e+10, 1.047415e+10, 1.037106e+10, 1.026446e+10, 
    1.015454e+10, 1.00415e+10, 9.925557e+09, 9.806899e+09, 9.68573e+09, 
    9.562249e+09, 9.436652e+09, 9.309132e+09, 9.17988e+09, 9.049084e+09, 
    8.916924e+09, 8.78358e+09, 8.649221e+09, 8.514017e+09, 8.378128e+09, 
    8.241709e+09, 8.10491e+09, 7.967875e+09, 7.830739e+09, 7.693634e+09, 
    7.556683e+09, 7.420003e+09, 7.283705e+09, 7.147894e+09, 7.012667e+09, 
    6.878117e+09,
  6.903431e+09, 7.040374e+09, 7.178077e+09, 7.316448e+09, 7.455388e+09, 
    7.594789e+09, 7.734541e+09, 7.874522e+09, 8.014606e+09, 8.15466e+09, 
    8.294543e+09, 8.434108e+09, 8.573202e+09, 8.711665e+09, 8.849328e+09, 
    8.986021e+09, 9.121564e+09, 9.255772e+09, 9.388457e+09, 9.519426e+09, 
    9.648477e+09, 9.775411e+09, 9.900023e+09, 1.00221e+10, 1.014144e+10, 
    1.025783e+10, 1.037106e+10, 1.048091e+10, 1.058718e+10, 1.068966e+10, 
    1.078814e+10, 1.088243e+10, 1.097232e+10, 1.105763e+10, 1.113816e+10, 
    1.121375e+10, 1.128423e+10, 1.134943e+10, 1.14092e+10, 1.146341e+10, 
    1.151193e+10, 1.155465e+10, 1.159146e+10, 1.162227e+10, 1.164701e+10, 
    1.166561e+10, 1.167804e+10, 1.168427e+10, 1.168427e+10, 1.167804e+10, 
    1.166561e+10, 1.164701e+10, 1.162227e+10, 1.159146e+10, 1.155465e+10, 
    1.151193e+10, 1.146341e+10, 1.14092e+10, 1.134943e+10, 1.128423e+10, 
    1.121375e+10, 1.113816e+10, 1.105763e+10, 1.097232e+10, 1.088243e+10, 
    1.078814e+10, 1.068966e+10, 1.058718e+10, 1.048091e+10, 1.037106e+10, 
    1.025783e+10, 1.014144e+10, 1.00221e+10, 9.900023e+09, 9.775411e+09, 
    9.648477e+09, 9.519426e+09, 9.388457e+09, 9.255772e+09, 9.121564e+09, 
    8.986021e+09, 8.849328e+09, 8.711665e+09, 8.573202e+09, 8.434108e+09, 
    8.294543e+09, 8.15466e+09, 8.014606e+09, 7.874522e+09, 7.734541e+09, 
    7.594789e+09, 7.455388e+09, 7.316448e+09, 7.178077e+09, 7.040374e+09, 
    6.903431e+09,
  6.927576e+09, 7.066821e+09, 7.206909e+09, 7.347746e+09, 7.489233e+09, 
    7.631261e+09, 7.773715e+09, 7.916475e+09, 8.059411e+09, 8.202386e+09, 
    8.345257e+09, 8.487873e+09, 8.630074e+09, 8.771699e+09, 8.912572e+09, 
    9.052518e+09, 9.191351e+09, 9.32888e+09, 9.464909e+09, 9.599237e+09, 
    9.731658e+09, 9.861961e+09, 9.989933e+09, 1.011536e+10, 1.023802e+10, 
    1.035769e+10, 1.047415e+10, 1.058718e+10, 1.069657e+10, 1.080209e+10, 
    1.090352e+10, 1.100067e+10, 1.109331e+10, 1.118125e+10, 1.12643e+10, 
    1.134227e+10, 1.141498e+10, 1.148226e+10, 1.154395e+10, 1.159992e+10, 
    1.165001e+10, 1.169412e+10, 1.173213e+10, 1.176396e+10, 1.178951e+10, 
    1.180873e+10, 1.182158e+10, 1.1828e+10, 1.1828e+10, 1.182158e+10, 
    1.180873e+10, 1.178951e+10, 1.176396e+10, 1.173213e+10, 1.169412e+10, 
    1.165001e+10, 1.159992e+10, 1.154395e+10, 1.148226e+10, 1.141498e+10, 
    1.134227e+10, 1.12643e+10, 1.118125e+10, 1.109331e+10, 1.100067e+10, 
    1.090352e+10, 1.080209e+10, 1.069657e+10, 1.058718e+10, 1.047415e+10, 
    1.035769e+10, 1.023802e+10, 1.011536e+10, 9.989933e+09, 9.861961e+09, 
    9.731658e+09, 9.599237e+09, 9.464909e+09, 9.32888e+09, 9.191351e+09, 
    9.052518e+09, 8.912572e+09, 8.771699e+09, 8.630074e+09, 8.487873e+09, 
    8.345257e+09, 8.202386e+09, 8.059411e+09, 7.916475e+09, 7.773715e+09, 
    7.631261e+09, 7.489233e+09, 7.347746e+09, 7.206909e+09, 7.066821e+09, 
    6.927576e+09,
  6.950547e+09, 7.092e+09, 7.234377e+09, 7.377583e+09, 7.521518e+09, 
    7.666072e+09, 7.811129e+09, 7.956566e+09, 8.10225e+09, 8.248043e+09, 
    8.393798e+09, 8.539359e+09, 8.684566e+09, 8.829247e+09, 8.973229e+09, 
    9.116325e+09, 9.258346e+09, 9.399095e+09, 9.53837e+09, 9.67596e+09, 
    9.811654e+09, 9.945231e+09, 1.007647e+10, 1.020515e+10, 1.033104e+10, 
    1.045391e+10, 1.057352e+10, 1.068966e+10, 1.080209e+10, 1.091057e+10, 
    1.10149e+10, 1.111483e+10, 1.121017e+10, 1.130069e+10, 1.13862e+10, 
    1.146649e+10, 1.154138e+10, 1.16107e+10, 1.167428e+10, 1.173195e+10, 
    1.17836e+10, 1.182907e+10, 1.186826e+10, 1.190108e+10, 1.192743e+10, 
    1.194726e+10, 1.19605e+10, 1.196713e+10, 1.196713e+10, 1.19605e+10, 
    1.194726e+10, 1.192743e+10, 1.190108e+10, 1.186826e+10, 1.182907e+10, 
    1.17836e+10, 1.173195e+10, 1.167428e+10, 1.16107e+10, 1.154138e+10, 
    1.146649e+10, 1.13862e+10, 1.130069e+10, 1.121017e+10, 1.111483e+10, 
    1.10149e+10, 1.091057e+10, 1.080209e+10, 1.068966e+10, 1.057352e+10, 
    1.045391e+10, 1.033104e+10, 1.020515e+10, 1.007647e+10, 9.945231e+09, 
    9.811654e+09, 9.67596e+09, 9.53837e+09, 9.399095e+09, 9.258346e+09, 
    9.116325e+09, 8.973229e+09, 8.829247e+09, 8.684566e+09, 8.539359e+09, 
    8.393798e+09, 8.248043e+09, 8.10225e+09, 7.956566e+09, 7.811129e+09, 
    7.666072e+09, 7.521518e+09, 7.377583e+09, 7.234377e+09, 7.092e+09, 
    6.950547e+09,
  6.972339e+09, 7.115902e+09, 7.260469e+09, 7.405943e+09, 7.552224e+09, 
    7.699199e+09, 7.846753e+09, 7.994759e+09, 8.143084e+09, 8.291585e+09, 
    8.440113e+09, 8.58851e+09, 8.736609e+09, 8.884238e+09, 9.031216e+09, 
    9.177352e+09, 9.322452e+09, 9.466312e+09, 9.608722e+09, 9.749469e+09, 
    9.88833e+09, 1.002508e+10, 1.015949e+10, 1.029132e+10, 1.042034e+10, 
    1.054631e+10, 1.066899e+10, 1.078814e+10, 1.090352e+10, 1.10149e+10, 
    1.112203e+10, 1.122468e+10, 1.132264e+10, 1.141567e+10, 1.150357e+10, 
    1.158613e+10, 1.166315e+10, 1.173446e+10, 1.179987e+10, 1.185922e+10, 
    1.191237e+10, 1.195917e+10, 1.199952e+10, 1.203331e+10, 1.206044e+10, 
    1.208085e+10, 1.209449e+10, 1.210132e+10, 1.210132e+10, 1.209449e+10, 
    1.208085e+10, 1.206044e+10, 1.203331e+10, 1.199952e+10, 1.195917e+10, 
    1.191237e+10, 1.185922e+10, 1.179987e+10, 1.173446e+10, 1.166315e+10, 
    1.158613e+10, 1.150357e+10, 1.141567e+10, 1.132264e+10, 1.122468e+10, 
    1.112203e+10, 1.10149e+10, 1.090352e+10, 1.078814e+10, 1.066899e+10, 
    1.054631e+10, 1.042034e+10, 1.029132e+10, 1.015949e+10, 1.002508e+10, 
    9.88833e+09, 9.749469e+09, 9.608722e+09, 9.466312e+09, 9.322452e+09, 
    9.177352e+09, 9.031216e+09, 8.884238e+09, 8.736609e+09, 8.58851e+09, 
    8.440113e+09, 8.291585e+09, 8.143084e+09, 7.994759e+09, 7.846753e+09, 
    7.699199e+09, 7.552224e+09, 7.405943e+09, 7.260469e+09, 7.115902e+09, 
    6.972339e+09,
  6.992947e+09, 7.138521e+09, 7.285175e+09, 7.432813e+09, 7.581331e+09, 
    7.73062e+09, 7.880559e+09, 8.031022e+09, 8.181873e+09, 8.332967e+09, 
    8.484152e+09, 8.635267e+09, 8.786142e+09, 8.936601e+09, 9.086456e+09, 
    9.235513e+09, 9.383574e+09, 9.530426e+09, 9.675857e+09, 9.819643e+09, 
    9.961556e+09, 1.010136e+10, 1.023883e+10, 1.037371e+10, 1.050575e+10, 
    1.063472e+10, 1.076036e+10, 1.088243e+10, 1.100067e+10, 1.111483e+10, 
    1.122468e+10, 1.132997e+10, 1.143046e+10, 1.152593e+10, 1.161615e+10, 
    1.170091e+10, 1.178001e+10, 1.185324e+10, 1.192043e+10, 1.198141e+10, 
    1.203602e+10, 1.208412e+10, 1.212559e+10, 1.216031e+10, 1.218821e+10, 
    1.220919e+10, 1.222321e+10, 1.223023e+10, 1.223023e+10, 1.222321e+10, 
    1.220919e+10, 1.218821e+10, 1.216031e+10, 1.212559e+10, 1.208412e+10, 
    1.203602e+10, 1.198141e+10, 1.192043e+10, 1.185324e+10, 1.178001e+10, 
    1.170091e+10, 1.161615e+10, 1.152593e+10, 1.143046e+10, 1.132997e+10, 
    1.122468e+10, 1.111483e+10, 1.100067e+10, 1.088243e+10, 1.076036e+10, 
    1.063472e+10, 1.050575e+10, 1.037371e+10, 1.023883e+10, 1.010136e+10, 
    9.961556e+09, 9.819643e+09, 9.675857e+09, 9.530426e+09, 9.383574e+09, 
    9.235513e+09, 9.086456e+09, 8.936601e+09, 8.786142e+09, 8.635267e+09, 
    8.484152e+09, 8.332967e+09, 8.181873e+09, 8.031022e+09, 7.880559e+09, 
    7.73062e+09, 7.581331e+09, 7.432813e+09, 7.285175e+09, 7.138521e+09, 
    6.992947e+09,
  7.012366e+09, 7.159848e+09, 7.308484e+09, 7.458176e+09, 7.608822e+09, 
    7.760311e+09, 7.912521e+09, 8.065324e+09, 8.218582e+09, 8.372148e+09, 
    8.525868e+09, 8.679578e+09, 8.833104e+09, 8.986266e+09, 9.138871e+09, 
    9.290724e+09, 9.441618e+09, 9.591338e+09, 9.739662e+09, 9.886363e+09, 
    1.00312e+10, 1.017395e+10, 1.031435e+10, 1.045215e+10, 1.058711e+10, 
    1.071896e+10, 1.084745e+10, 1.097232e+10, 1.109331e+10, 1.121017e+10, 
    1.132264e+10, 1.143046e+10, 1.153341e+10, 1.163122e+10, 1.172369e+10, 
    1.181057e+10, 1.189166e+10, 1.196675e+10, 1.203567e+10, 1.209821e+10, 
    1.215424e+10, 1.220359e+10, 1.224615e+10, 1.228178e+10, 1.231041e+10, 
    1.233195e+10, 1.234634e+10, 1.235355e+10, 1.235355e+10, 1.234634e+10, 
    1.233195e+10, 1.231041e+10, 1.228178e+10, 1.224615e+10, 1.220359e+10, 
    1.215424e+10, 1.209821e+10, 1.203567e+10, 1.196675e+10, 1.189166e+10, 
    1.181057e+10, 1.172369e+10, 1.163122e+10, 1.153341e+10, 1.143046e+10, 
    1.132264e+10, 1.121017e+10, 1.109331e+10, 1.097232e+10, 1.084745e+10, 
    1.071896e+10, 1.058711e+10, 1.045215e+10, 1.031435e+10, 1.017395e+10, 
    1.00312e+10, 9.886363e+09, 9.739662e+09, 9.591338e+09, 9.441618e+09, 
    9.290724e+09, 9.138871e+09, 8.986266e+09, 8.833104e+09, 8.679578e+09, 
    8.525868e+09, 8.372148e+09, 8.218582e+09, 8.065324e+09, 7.912521e+09, 
    7.760311e+09, 7.608822e+09, 7.458176e+09, 7.308484e+09, 7.159848e+09, 
    7.012366e+09,
  7.030593e+09, 7.179877e+09, 7.330385e+09, 7.482021e+09, 7.634681e+09, 
    7.788252e+09, 7.942612e+09, 8.097633e+09, 8.253174e+09, 8.409087e+09, 
    8.565214e+09, 8.721389e+09, 8.877434e+09, 9.033167e+09, 9.188391e+09, 
    9.342905e+09, 9.496498e+09, 9.64895e+09, 9.800034e+09, 9.949515e+09, 
    1.009715e+10, 1.02427e+10, 1.03859e+10, 1.05265e+10, 1.066424e+10, 
    1.079885e+10, 1.093007e+10, 1.105763e+10, 1.118125e+10, 1.130069e+10, 
    1.141567e+10, 1.152593e+10, 1.163122e+10, 1.17313e+10, 1.182591e+10, 
    1.191483e+10, 1.199784e+10, 1.207473e+10, 1.214529e+10, 1.220935e+10, 
    1.226673e+10, 1.231729e+10, 1.236089e+10, 1.23974e+10, 1.242673e+10, 
    1.24488e+10, 1.246355e+10, 1.247093e+10, 1.247093e+10, 1.246355e+10, 
    1.24488e+10, 1.242673e+10, 1.23974e+10, 1.236089e+10, 1.231729e+10, 
    1.226673e+10, 1.220935e+10, 1.214529e+10, 1.207473e+10, 1.199784e+10, 
    1.191483e+10, 1.182591e+10, 1.17313e+10, 1.163122e+10, 1.152593e+10, 
    1.141567e+10, 1.130069e+10, 1.118125e+10, 1.105763e+10, 1.093007e+10, 
    1.079885e+10, 1.066424e+10, 1.05265e+10, 1.03859e+10, 1.02427e+10, 
    1.009715e+10, 9.949515e+09, 9.800034e+09, 9.64895e+09, 9.496498e+09, 
    9.342905e+09, 9.188391e+09, 9.033167e+09, 8.877434e+09, 8.721389e+09, 
    8.565214e+09, 8.409087e+09, 8.253174e+09, 8.097633e+09, 7.942612e+09, 
    7.788252e+09, 7.634681e+09, 7.482021e+09, 7.330385e+09, 7.179877e+09, 
    7.030593e+09,
  7.047623e+09, 7.198601e+09, 7.350871e+09, 7.504335e+09, 7.65889e+09, 
    7.814423e+09, 7.970811e+09, 8.127923e+09, 8.285618e+09, 8.443745e+09, 
    8.602145e+09, 8.760649e+09, 8.919077e+09, 9.077242e+09, 9.234944e+09, 
    9.391978e+09, 9.548129e+09, 9.703171e+09, 9.856871e+09, 1.000899e+10, 
    1.015928e+10, 1.030749e+10, 1.045336e+10, 1.059662e+10, 1.0737e+10, 
    1.087423e+10, 1.100805e+10, 1.113816e+10, 1.12643e+10, 1.13862e+10, 
    1.150357e+10, 1.161615e+10, 1.172369e+10, 1.182591e+10, 1.192258e+10, 
    1.201345e+10, 1.209829e+10, 1.217688e+10, 1.224902e+10, 1.231452e+10, 
    1.237321e+10, 1.242492e+10, 1.246951e+10, 1.250686e+10, 1.253687e+10, 
    1.255944e+10, 1.257453e+10, 1.258209e+10, 1.258209e+10, 1.257453e+10, 
    1.255944e+10, 1.253687e+10, 1.250686e+10, 1.246951e+10, 1.242492e+10, 
    1.237321e+10, 1.231452e+10, 1.224902e+10, 1.217688e+10, 1.209829e+10, 
    1.201345e+10, 1.192258e+10, 1.182591e+10, 1.172369e+10, 1.161615e+10, 
    1.150357e+10, 1.13862e+10, 1.12643e+10, 1.113816e+10, 1.100805e+10, 
    1.087423e+10, 1.0737e+10, 1.059662e+10, 1.045336e+10, 1.030749e+10, 
    1.015928e+10, 1.000899e+10, 9.856871e+09, 9.703171e+09, 9.548129e+09, 
    9.391978e+09, 9.234944e+09, 9.077242e+09, 8.919077e+09, 8.760649e+09, 
    8.602145e+09, 8.443745e+09, 8.285618e+09, 8.127923e+09, 7.970811e+09, 
    7.814423e+09, 7.65889e+09, 7.504335e+09, 7.350871e+09, 7.198601e+09, 
    7.047623e+09,
  7.063453e+09, 7.216014e+09, 7.36993e+09, 7.525106e+09, 7.681435e+09, 
    7.838806e+09, 7.997093e+09, 8.156166e+09, 8.31588e+09, 8.476086e+09, 
    8.636621e+09, 8.797313e+09, 8.95798e+09, 9.118431e+09, 9.278465e+09, 
    9.437871e+09, 9.596429e+09, 9.753911e+09, 9.910078e+09, 1.006469e+10, 
    1.021748e+10, 1.03682e+10, 1.051658e+10, 1.066235e+10, 1.080523e+10, 
    1.094495e+10, 1.108122e+10, 1.121375e+10, 1.134227e+10, 1.146649e+10, 
    1.158613e+10, 1.170091e+10, 1.181057e+10, 1.191483e+10, 1.201345e+10, 
    1.210616e+10, 1.219274e+10, 1.227295e+10, 1.234659e+10, 1.241347e+10, 
    1.247338e+10, 1.252618e+10, 1.257172e+10, 1.260987e+10, 1.264052e+10, 
    1.266358e+10, 1.267899e+10, 1.268671e+10, 1.268671e+10, 1.267899e+10, 
    1.266358e+10, 1.264052e+10, 1.260987e+10, 1.257172e+10, 1.252618e+10, 
    1.247338e+10, 1.241347e+10, 1.234659e+10, 1.227295e+10, 1.219274e+10, 
    1.210616e+10, 1.201345e+10, 1.191483e+10, 1.181057e+10, 1.170091e+10, 
    1.158613e+10, 1.146649e+10, 1.134227e+10, 1.121375e+10, 1.108122e+10, 
    1.094495e+10, 1.080523e+10, 1.066235e+10, 1.051658e+10, 1.03682e+10, 
    1.021748e+10, 1.006469e+10, 9.910078e+09, 9.753911e+09, 9.596429e+09, 
    9.437871e+09, 9.278465e+09, 9.118431e+09, 8.95798e+09, 8.797313e+09, 
    8.636621e+09, 8.476086e+09, 8.31588e+09, 8.156166e+09, 7.997093e+09, 
    7.838806e+09, 7.681435e+09, 7.525106e+09, 7.36993e+09, 7.216014e+09, 
    7.063453e+09,
  7.078078e+09, 7.23211e+09, 7.387556e+09, 7.544322e+09, 7.702302e+09, 
    7.861382e+09, 8.021437e+09, 8.182336e+09, 8.343933e+09, 8.506077e+09, 
    8.668601e+09, 8.831335e+09, 8.994092e+09, 9.156679e+09, 9.318892e+09, 
    9.480515e+09, 9.641325e+09, 9.801088e+09, 9.959563e+09, 1.01165e+10, 
    1.027164e+10, 1.042471e+10, 1.057545e+10, 1.072358e+10, 1.08688e+10, 
    1.101085e+10, 1.114942e+10, 1.128423e+10, 1.141498e+10, 1.154138e+10, 
    1.166315e+10, 1.178001e+10, 1.189166e+10, 1.199784e+10, 1.209829e+10, 
    1.219274e+10, 1.228095e+10, 1.236269e+10, 1.243775e+10, 1.250591e+10, 
    1.256699e+10, 1.262082e+10, 1.266725e+10, 1.270614e+10, 1.273739e+10, 
    1.276091e+10, 1.277663e+10, 1.27845e+10, 1.27845e+10, 1.277663e+10, 
    1.276091e+10, 1.273739e+10, 1.270614e+10, 1.266725e+10, 1.262082e+10, 
    1.256699e+10, 1.250591e+10, 1.243775e+10, 1.236269e+10, 1.228095e+10, 
    1.219274e+10, 1.209829e+10, 1.199784e+10, 1.189166e+10, 1.178001e+10, 
    1.166315e+10, 1.154138e+10, 1.141498e+10, 1.128423e+10, 1.114942e+10, 
    1.101085e+10, 1.08688e+10, 1.072358e+10, 1.057545e+10, 1.042471e+10, 
    1.027164e+10, 1.01165e+10, 9.959563e+09, 9.801088e+09, 9.641325e+09, 
    9.480515e+09, 9.318892e+09, 9.156679e+09, 8.994092e+09, 8.831335e+09, 
    8.668601e+09, 8.506077e+09, 8.343933e+09, 8.182336e+09, 8.021437e+09, 
    7.861382e+09, 7.702302e+09, 7.544322e+09, 7.387556e+09, 7.23211e+09, 
    7.078078e+09,
  7.091497e+09, 7.246883e+09, 7.403741e+09, 7.561974e+09, 7.721477e+09, 
    7.882135e+09, 8.043825e+09, 8.20641e+09, 8.369748e+09, 8.533684e+09, 
    8.698051e+09, 8.862674e+09, 9.027367e+09, 9.191932e+09, 9.356163e+09, 
    9.519842e+09, 9.68274e+09, 9.844622e+09, 1.000524e+10, 1.016434e+10, 
    1.032166e+10, 1.047692e+10, 1.062985e+10, 1.078017e+10, 1.092757e+10, 
    1.107179e+10, 1.12125e+10, 1.134943e+10, 1.148226e+10, 1.16107e+10, 
    1.173446e+10, 1.185324e+10, 1.196675e+10, 1.207473e+10, 1.217688e+10, 
    1.227295e+10, 1.236269e+10, 1.244586e+10, 1.252223e+10, 1.25916e+10, 
    1.265377e+10, 1.270856e+10, 1.275582e+10, 1.279542e+10, 1.282723e+10, 
    1.285118e+10, 1.286718e+10, 1.287519e+10, 1.287519e+10, 1.286718e+10, 
    1.285118e+10, 1.282723e+10, 1.279542e+10, 1.275582e+10, 1.270856e+10, 
    1.265377e+10, 1.25916e+10, 1.252223e+10, 1.244586e+10, 1.236269e+10, 
    1.227295e+10, 1.217688e+10, 1.207473e+10, 1.196675e+10, 1.185324e+10, 
    1.173446e+10, 1.16107e+10, 1.148226e+10, 1.134943e+10, 1.12125e+10, 
    1.107179e+10, 1.092757e+10, 1.078017e+10, 1.062985e+10, 1.047692e+10, 
    1.032166e+10, 1.016434e+10, 1.000524e+10, 9.844622e+09, 9.68274e+09, 
    9.519842e+09, 9.356163e+09, 9.191932e+09, 9.027367e+09, 8.862674e+09, 
    8.698051e+09, 8.533684e+09, 8.369748e+09, 8.20641e+09, 8.043825e+09, 
    7.882135e+09, 7.721477e+09, 7.561974e+09, 7.403741e+09, 7.246883e+09, 
    7.091497e+09,
  7.103705e+09, 7.260329e+09, 7.418477e+09, 7.578052e+09, 7.738948e+09, 
    7.901051e+09, 8.064236e+09, 8.228367e+09, 8.3933e+09, 8.558878e+09, 
    8.724934e+09, 8.891291e+09, 9.05776e+09, 9.224142e+09, 9.390226e+09, 
    9.555794e+09, 9.720613e+09, 9.884442e+09, 1.004703e+10, 1.020812e+10, 
    1.036744e+10, 1.052472e+10, 1.067967e+10, 1.0832e+10, 1.098142e+10, 
    1.112763e+10, 1.127033e+10, 1.14092e+10, 1.154395e+10, 1.167428e+10, 
    1.179987e+10, 1.192043e+10, 1.203567e+10, 1.214529e+10, 1.224902e+10, 
    1.234659e+10, 1.243775e+10, 1.252223e+10, 1.259983e+10, 1.267031e+10, 
    1.273348e+10, 1.278916e+10, 1.283719e+10, 1.287743e+10, 1.290977e+10, 
    1.293411e+10, 1.295038e+10, 1.295852e+10, 1.295852e+10, 1.295038e+10, 
    1.293411e+10, 1.290977e+10, 1.287743e+10, 1.283719e+10, 1.278916e+10, 
    1.273348e+10, 1.267031e+10, 1.259983e+10, 1.252223e+10, 1.243775e+10, 
    1.234659e+10, 1.224902e+10, 1.214529e+10, 1.203567e+10, 1.192043e+10, 
    1.179987e+10, 1.167428e+10, 1.154395e+10, 1.14092e+10, 1.127033e+10, 
    1.112763e+10, 1.098142e+10, 1.0832e+10, 1.067967e+10, 1.052472e+10, 
    1.036744e+10, 1.020812e+10, 1.004703e+10, 9.884442e+09, 9.720613e+09, 
    9.555794e+09, 9.390226e+09, 9.224142e+09, 9.05776e+09, 8.891291e+09, 
    8.724934e+09, 8.558878e+09, 8.3933e+09, 8.228367e+09, 8.064236e+09, 
    7.901051e+09, 7.738948e+09, 7.578052e+09, 7.418477e+09, 7.260329e+09, 
    7.103705e+09,
  7.1147e+09, 7.272444e+09, 7.431758e+09, 7.592547e+09, 7.754704e+09, 
    7.918115e+09, 8.082655e+09, 8.248187e+09, 8.414565e+09, 8.581632e+09, 
    8.749221e+09, 8.917151e+09, 9.085231e+09, 9.253263e+09, 9.421031e+09, 
    9.588315e+09, 9.754878e+09, 9.920478e+09, 1.008486e+10, 1.024776e+10, 
    1.040891e+10, 1.056802e+10, 1.07248e+10, 1.087898e+10, 1.103023e+10, 
    1.117826e+10, 1.132276e+10, 1.146341e+10, 1.159992e+10, 1.173195e+10, 
    1.185922e+10, 1.198141e+10, 1.209821e+10, 1.220935e+10, 1.231452e+10, 
    1.241347e+10, 1.250591e+10, 1.25916e+10, 1.267031e+10, 1.27418e+10, 
    1.280589e+10, 1.286239e+10, 1.291113e+10, 1.295196e+10, 1.298478e+10, 
    1.300948e+10, 1.302599e+10, 1.303425e+10, 1.303425e+10, 1.302599e+10, 
    1.300948e+10, 1.298478e+10, 1.295196e+10, 1.291113e+10, 1.286239e+10, 
    1.280589e+10, 1.27418e+10, 1.267031e+10, 1.25916e+10, 1.250591e+10, 
    1.241347e+10, 1.231452e+10, 1.220935e+10, 1.209821e+10, 1.198141e+10, 
    1.185922e+10, 1.173195e+10, 1.159992e+10, 1.146341e+10, 1.132276e+10, 
    1.117826e+10, 1.103023e+10, 1.087898e+10, 1.07248e+10, 1.056802e+10, 
    1.040891e+10, 1.024776e+10, 1.008486e+10, 9.920478e+09, 9.754878e+09, 
    9.588315e+09, 9.421031e+09, 9.253263e+09, 9.085231e+09, 8.917151e+09, 
    8.749221e+09, 8.581632e+09, 8.414565e+09, 8.248187e+09, 8.082655e+09, 
    7.918115e+09, 7.754704e+09, 7.592547e+09, 7.431758e+09, 7.272444e+09, 
    7.1147e+09,
  7.124479e+09, 7.283223e+09, 7.443579e+09, 7.605452e+09, 7.768736e+09, 
    7.933316e+09, 8.099066e+09, 8.26585e+09, 8.433522e+09, 8.601922e+09, 
    8.770882e+09, 8.940219e+09, 9.109745e+09, 9.279254e+09, 9.448532e+09, 
    9.617354e+09, 9.785482e+09, 9.95267e+09, 1.011866e+10, 1.028319e+10, 
    1.044597e+10, 1.060673e+10, 1.076517e+10, 1.092099e+10, 1.107389e+10, 
    1.122356e+10, 1.136968e+10, 1.151193e+10, 1.165001e+10, 1.17836e+10, 
    1.191237e+10, 1.203602e+10, 1.215424e+10, 1.226673e+10, 1.237321e+10, 
    1.247338e+10, 1.256699e+10, 1.265377e+10, 1.273348e+10, 1.280589e+10, 
    1.287081e+10, 1.292804e+10, 1.297741e+10, 1.301878e+10, 1.305203e+10, 
    1.307706e+10, 1.309378e+10, 1.310215e+10, 1.310215e+10, 1.309378e+10, 
    1.307706e+10, 1.305203e+10, 1.301878e+10, 1.297741e+10, 1.292804e+10, 
    1.287081e+10, 1.280589e+10, 1.273348e+10, 1.265377e+10, 1.256699e+10, 
    1.247338e+10, 1.237321e+10, 1.226673e+10, 1.215424e+10, 1.203602e+10, 
    1.191237e+10, 1.17836e+10, 1.165001e+10, 1.151193e+10, 1.136968e+10, 
    1.122356e+10, 1.107389e+10, 1.092099e+10, 1.076517e+10, 1.060673e+10, 
    1.044597e+10, 1.028319e+10, 1.011866e+10, 9.95267e+09, 9.785482e+09, 
    9.617354e+09, 9.448532e+09, 9.279254e+09, 9.109745e+09, 8.940219e+09, 
    8.770882e+09, 8.601922e+09, 8.433522e+09, 8.26585e+09, 8.099066e+09, 
    7.933316e+09, 7.768736e+09, 7.605452e+09, 7.443579e+09, 7.283223e+09, 
    7.124479e+09,
  7.133041e+09, 7.292662e+09, 7.453934e+09, 7.616759e+09, 7.781033e+09, 
    7.946641e+09, 8.113456e+09, 8.281342e+09, 8.450151e+09, 8.619724e+09, 
    8.789891e+09, 8.96047e+09, 9.131267e+09, 9.302078e+09, 9.472687e+09, 
    9.642865e+09, 9.812372e+09, 9.980962e+09, 1.014837e+10, 1.031433e+10, 
    1.047856e+10, 1.064077e+10, 1.080067e+10, 1.095795e+10, 1.111231e+10, 
    1.126342e+10, 1.141097e+10, 1.155465e+10, 1.169412e+10, 1.182907e+10, 
    1.195917e+10, 1.208412e+10, 1.220359e+10, 1.231729e+10, 1.242492e+10, 
    1.252618e+10, 1.262082e+10, 1.270856e+10, 1.278916e+10, 1.286239e+10, 
    1.292804e+10, 1.298592e+10, 1.303585e+10, 1.30777e+10, 1.311133e+10, 
    1.313664e+10, 1.315356e+10, 1.316203e+10, 1.316203e+10, 1.315356e+10, 
    1.313664e+10, 1.311133e+10, 1.30777e+10, 1.303585e+10, 1.298592e+10, 
    1.292804e+10, 1.286239e+10, 1.278916e+10, 1.270856e+10, 1.262082e+10, 
    1.252618e+10, 1.242492e+10, 1.231729e+10, 1.220359e+10, 1.208412e+10, 
    1.195917e+10, 1.182907e+10, 1.169412e+10, 1.155465e+10, 1.141097e+10, 
    1.126342e+10, 1.111231e+10, 1.095795e+10, 1.080067e+10, 1.064077e+10, 
    1.047856e+10, 1.031433e+10, 1.014837e+10, 9.980962e+09, 9.812372e+09, 
    9.642865e+09, 9.472687e+09, 9.302078e+09, 9.131267e+09, 8.96047e+09, 
    8.789891e+09, 8.619724e+09, 8.450151e+09, 8.281342e+09, 8.113456e+09, 
    7.946641e+09, 7.781033e+09, 7.616759e+09, 7.453934e+09, 7.292662e+09, 
    7.133041e+09,
  7.140384e+09, 7.30076e+09, 7.462817e+09, 7.626462e+09, 7.791588e+09, 
    7.958081e+09, 8.125813e+09, 8.294647e+09, 8.464436e+09, 8.63502e+09, 
    8.806228e+09, 8.977876e+09, 9.14977e+09, 9.321703e+09, 9.49346e+09, 
    9.664807e+09, 9.835507e+09, 1.00053e+10, 1.017394e+10, 1.034114e+10, 
    1.050662e+10, 1.067009e+10, 1.083124e+10, 1.098979e+10, 1.11454e+10, 
    1.129776e+10, 1.144656e+10, 1.159146e+10, 1.173213e+10, 1.186826e+10, 
    1.199952e+10, 1.212559e+10, 1.224615e+10, 1.236089e+10, 1.246951e+10, 
    1.257172e+10, 1.266725e+10, 1.275582e+10, 1.283719e+10, 1.291113e+10, 
    1.297741e+10, 1.303585e+10, 1.308628e+10, 1.312854e+10, 1.316249e+10, 
    1.318806e+10, 1.320514e+10, 1.32137e+10, 1.32137e+10, 1.320514e+10, 
    1.318806e+10, 1.316249e+10, 1.312854e+10, 1.308628e+10, 1.303585e+10, 
    1.297741e+10, 1.291113e+10, 1.283719e+10, 1.275582e+10, 1.266725e+10, 
    1.257172e+10, 1.246951e+10, 1.236089e+10, 1.224615e+10, 1.212559e+10, 
    1.199952e+10, 1.186826e+10, 1.173213e+10, 1.159146e+10, 1.144656e+10, 
    1.129776e+10, 1.11454e+10, 1.098979e+10, 1.083124e+10, 1.067009e+10, 
    1.050662e+10, 1.034114e+10, 1.017394e+10, 1.00053e+10, 9.835507e+09, 
    9.664807e+09, 9.49346e+09, 9.321703e+09, 9.14977e+09, 8.977876e+09, 
    8.806228e+09, 8.63502e+09, 8.464436e+09, 8.294647e+09, 8.125813e+09, 
    7.958081e+09, 7.791588e+09, 7.626462e+09, 7.462817e+09, 7.30076e+09, 
    7.140384e+09,
  7.146505e+09, 7.307511e+09, 7.470226e+09, 7.634556e+09, 7.800395e+09, 
    7.967627e+09, 8.136126e+09, 8.305754e+09, 8.476363e+09, 8.647793e+09, 
    8.819871e+09, 8.992415e+09, 9.165227e+09, 9.338102e+09, 9.510819e+09, 
    9.683147e+09, 9.854844e+09, 1.002566e+10, 1.019532e+10, 1.036355e+10, 
    1.053008e+10, 1.06946e+10, 1.085682e+10, 1.101642e+10, 1.117309e+10, 
    1.13265e+10, 1.147634e+10, 1.162227e+10, 1.176396e+10, 1.190108e+10, 
    1.203331e+10, 1.216031e+10, 1.228178e+10, 1.23974e+10, 1.250686e+10, 
    1.260987e+10, 1.270614e+10, 1.279542e+10, 1.287743e+10, 1.295196e+10, 
    1.301878e+10, 1.30777e+10, 1.312854e+10, 1.317114e+10, 1.320537e+10, 
    1.323115e+10, 1.324837e+10, 1.3257e+10, 1.3257e+10, 1.324837e+10, 
    1.323115e+10, 1.320537e+10, 1.317114e+10, 1.312854e+10, 1.30777e+10, 
    1.301878e+10, 1.295196e+10, 1.287743e+10, 1.279542e+10, 1.270614e+10, 
    1.260987e+10, 1.250686e+10, 1.23974e+10, 1.228178e+10, 1.216031e+10, 
    1.203331e+10, 1.190108e+10, 1.176396e+10, 1.162227e+10, 1.147634e+10, 
    1.13265e+10, 1.117309e+10, 1.101642e+10, 1.085682e+10, 1.06946e+10, 
    1.053008e+10, 1.036355e+10, 1.019532e+10, 1.002566e+10, 9.854844e+09, 
    9.683147e+09, 9.510819e+09, 9.338102e+09, 9.165227e+09, 8.992415e+09, 
    8.819871e+09, 8.647793e+09, 8.476363e+09, 8.305754e+09, 8.136126e+09, 
    7.967627e+09, 7.800395e+09, 7.634556e+09, 7.470226e+09, 7.307511e+09, 
    7.146505e+09,
  7.151404e+09, 7.312915e+09, 7.476158e+09, 7.641037e+09, 7.807448e+09, 
    7.975273e+09, 8.144387e+09, 8.314652e+09, 8.485919e+09, 8.658028e+09, 
    8.830806e+09, 9.004068e+09, 9.177618e+09, 9.351248e+09, 9.524738e+09, 
    9.697854e+09, 9.870353e+09, 1.004198e+10, 1.021247e+10, 1.038154e+10, 
    1.054891e+10, 1.071428e+10, 1.087735e+10, 1.10378e+10, 1.119532e+10, 
    1.134958e+10, 1.150025e+10, 1.164701e+10, 1.178951e+10, 1.192743e+10, 
    1.206044e+10, 1.218821e+10, 1.231041e+10, 1.242673e+10, 1.253687e+10, 
    1.264052e+10, 1.273739e+10, 1.282723e+10, 1.290977e+10, 1.298478e+10, 
    1.305203e+10, 1.311133e+10, 1.316249e+10, 1.320537e+10, 1.323984e+10, 
    1.326578e+10, 1.328312e+10, 1.32918e+10, 1.32918e+10, 1.328312e+10, 
    1.326578e+10, 1.323984e+10, 1.320537e+10, 1.316249e+10, 1.311133e+10, 
    1.305203e+10, 1.298478e+10, 1.290977e+10, 1.282723e+10, 1.273739e+10, 
    1.264052e+10, 1.253687e+10, 1.242673e+10, 1.231041e+10, 1.218821e+10, 
    1.206044e+10, 1.192743e+10, 1.178951e+10, 1.164701e+10, 1.150025e+10, 
    1.134958e+10, 1.119532e+10, 1.10378e+10, 1.087735e+10, 1.071428e+10, 
    1.054891e+10, 1.038154e+10, 1.021247e+10, 1.004198e+10, 9.870353e+09, 
    9.697854e+09, 9.524738e+09, 9.351248e+09, 9.177618e+09, 9.004068e+09, 
    8.830806e+09, 8.658028e+09, 8.485919e+09, 8.314652e+09, 8.144387e+09, 
    7.975273e+09, 7.807448e+09, 7.641037e+09, 7.476158e+09, 7.312915e+09, 
    7.151404e+09,
  7.155078e+09, 7.316969e+09, 7.480609e+09, 7.645901e+09, 7.812741e+09, 
    7.981012e+09, 8.150589e+09, 8.321333e+09, 8.493095e+09, 8.665715e+09, 
    8.839017e+09, 9.012821e+09, 9.186927e+09, 9.361125e+09, 9.535196e+09, 
    9.708905e+09, 9.882009e+09, 1.005425e+10, 1.022536e+10, 1.039506e+10, 
    1.056306e+10, 1.072907e+10, 1.089278e+10, 1.105388e+10, 1.121203e+10, 
    1.136693e+10, 1.151823e+10, 1.166561e+10, 1.180873e+10, 1.194726e+10, 
    1.208085e+10, 1.220919e+10, 1.233195e+10, 1.24488e+10, 1.255944e+10, 
    1.266358e+10, 1.276091e+10, 1.285118e+10, 1.293411e+10, 1.300948e+10, 
    1.307706e+10, 1.313664e+10, 1.318806e+10, 1.323115e+10, 1.326578e+10, 
    1.329185e+10, 1.330927e+10, 1.3318e+10, 1.3318e+10, 1.330927e+10, 
    1.329185e+10, 1.326578e+10, 1.323115e+10, 1.318806e+10, 1.313664e+10, 
    1.307706e+10, 1.300948e+10, 1.293411e+10, 1.285118e+10, 1.276091e+10, 
    1.266358e+10, 1.255944e+10, 1.24488e+10, 1.233195e+10, 1.220919e+10, 
    1.208085e+10, 1.194726e+10, 1.180873e+10, 1.166561e+10, 1.151823e+10, 
    1.136693e+10, 1.121203e+10, 1.105388e+10, 1.089278e+10, 1.072907e+10, 
    1.056306e+10, 1.039506e+10, 1.022536e+10, 1.005425e+10, 9.882009e+09, 
    9.708905e+09, 9.535196e+09, 9.361125e+09, 9.186927e+09, 9.012821e+09, 
    8.839017e+09, 8.665715e+09, 8.493095e+09, 8.321333e+09, 8.150589e+09, 
    7.981012e+09, 7.812741e+09, 7.645901e+09, 7.480609e+09, 7.316969e+09, 
    7.155078e+09,
  7.157529e+09, 7.319673e+09, 7.483577e+09, 7.649145e+09, 7.816271e+09, 
    7.984841e+09, 8.154726e+09, 8.32579e+09, 8.497883e+09, 8.670843e+09, 
    8.844498e+09, 9.018663e+09, 9.193139e+09, 9.367718e+09, 9.542177e+09, 
    9.716282e+09, 9.88979e+09, 1.006244e+10, 1.023397e+10, 1.040409e+10, 
    1.057252e+10, 1.073895e+10, 1.090309e+10, 1.106461e+10, 1.12232e+10, 
    1.137852e+10, 1.153025e+10, 1.167804e+10, 1.182158e+10, 1.19605e+10, 
    1.209449e+10, 1.222321e+10, 1.234634e+10, 1.246355e+10, 1.257453e+10, 
    1.267899e+10, 1.277663e+10, 1.286718e+10, 1.295038e+10, 1.302599e+10, 
    1.309378e+10, 1.315356e+10, 1.320514e+10, 1.324837e+10, 1.328312e+10, 
    1.330927e+10, 1.332675e+10, 1.333551e+10, 1.333551e+10, 1.332675e+10, 
    1.330927e+10, 1.328312e+10, 1.324837e+10, 1.320514e+10, 1.315356e+10, 
    1.309378e+10, 1.302599e+10, 1.295038e+10, 1.286718e+10, 1.277663e+10, 
    1.267899e+10, 1.257453e+10, 1.246355e+10, 1.234634e+10, 1.222321e+10, 
    1.209449e+10, 1.19605e+10, 1.182158e+10, 1.167804e+10, 1.153025e+10, 
    1.137852e+10, 1.12232e+10, 1.106461e+10, 1.090309e+10, 1.073895e+10, 
    1.057252e+10, 1.040409e+10, 1.023397e+10, 1.006244e+10, 9.88979e+09, 
    9.716282e+09, 9.542177e+09, 9.367718e+09, 9.193139e+09, 9.018663e+09, 
    8.844498e+09, 8.670843e+09, 8.497883e+09, 8.32579e+09, 8.154726e+09, 
    7.984841e+09, 7.816271e+09, 7.649145e+09, 7.483577e+09, 7.319673e+09, 
    7.157529e+09,
  7.158754e+09, 7.321026e+09, 7.485062e+09, 7.650767e+09, 7.818037e+09, 
    7.986756e+09, 8.156796e+09, 8.32802e+09, 8.500278e+09, 8.673409e+09, 
    8.84724e+09, 9.021585e+09, 9.196247e+09, 9.371016e+09, 9.54567e+09, 
    9.719975e+09, 9.893683e+09, 1.006654e+10, 1.023827e+10, 1.040861e+10, 
    1.057725e+10, 1.07439e+10, 1.090825e+10, 1.106999e+10, 1.122879e+10, 
    1.138432e+10, 1.153626e+10, 1.168427e+10, 1.1828e+10, 1.196713e+10, 
    1.210132e+10, 1.223023e+10, 1.235355e+10, 1.247093e+10, 1.258209e+10, 
    1.268671e+10, 1.27845e+10, 1.287519e+10, 1.295852e+10, 1.303425e+10, 
    1.310215e+10, 1.316203e+10, 1.32137e+10, 1.3257e+10, 1.32918e+10, 
    1.3318e+10, 1.333551e+10, 1.334428e+10, 1.334428e+10, 1.333551e+10, 
    1.3318e+10, 1.32918e+10, 1.3257e+10, 1.32137e+10, 1.316203e+10, 
    1.310215e+10, 1.303425e+10, 1.295852e+10, 1.287519e+10, 1.27845e+10, 
    1.268671e+10, 1.258209e+10, 1.247093e+10, 1.235355e+10, 1.223023e+10, 
    1.210132e+10, 1.196713e+10, 1.1828e+10, 1.168427e+10, 1.153626e+10, 
    1.138432e+10, 1.122879e+10, 1.106999e+10, 1.090825e+10, 1.07439e+10, 
    1.057725e+10, 1.040861e+10, 1.023827e+10, 1.006654e+10, 9.893683e+09, 
    9.719975e+09, 9.54567e+09, 9.371016e+09, 9.196247e+09, 9.021585e+09, 
    8.84724e+09, 8.673409e+09, 8.500278e+09, 8.32802e+09, 8.156796e+09, 
    7.986756e+09, 7.818037e+09, 7.650767e+09, 7.485062e+09, 7.321026e+09, 
    7.158754e+09,
  7.158754e+09, 7.321026e+09, 7.485062e+09, 7.650767e+09, 7.818037e+09, 
    7.986756e+09, 8.156796e+09, 8.32802e+09, 8.500278e+09, 8.673409e+09, 
    8.84724e+09, 9.021585e+09, 9.196247e+09, 9.371016e+09, 9.54567e+09, 
    9.719975e+09, 9.893683e+09, 1.006654e+10, 1.023827e+10, 1.040861e+10, 
    1.057725e+10, 1.07439e+10, 1.090825e+10, 1.106999e+10, 1.122879e+10, 
    1.138432e+10, 1.153626e+10, 1.168427e+10, 1.1828e+10, 1.196713e+10, 
    1.210132e+10, 1.223023e+10, 1.235355e+10, 1.247093e+10, 1.258209e+10, 
    1.268671e+10, 1.27845e+10, 1.287519e+10, 1.295852e+10, 1.303425e+10, 
    1.310215e+10, 1.316203e+10, 1.32137e+10, 1.3257e+10, 1.32918e+10, 
    1.3318e+10, 1.333551e+10, 1.334428e+10, 1.334428e+10, 1.333551e+10, 
    1.3318e+10, 1.32918e+10, 1.3257e+10, 1.32137e+10, 1.316203e+10, 
    1.310215e+10, 1.303425e+10, 1.295852e+10, 1.287519e+10, 1.27845e+10, 
    1.268671e+10, 1.258209e+10, 1.247093e+10, 1.235355e+10, 1.223023e+10, 
    1.210132e+10, 1.196713e+10, 1.1828e+10, 1.168427e+10, 1.153626e+10, 
    1.138432e+10, 1.122879e+10, 1.106999e+10, 1.090825e+10, 1.07439e+10, 
    1.057725e+10, 1.040861e+10, 1.023827e+10, 1.006654e+10, 9.893683e+09, 
    9.719975e+09, 9.54567e+09, 9.371016e+09, 9.196247e+09, 9.021585e+09, 
    8.84724e+09, 8.673409e+09, 8.500278e+09, 8.32802e+09, 8.156796e+09, 
    7.986756e+09, 7.818037e+09, 7.650767e+09, 7.485062e+09, 7.321026e+09, 
    7.158754e+09,
  7.157529e+09, 7.319673e+09, 7.483577e+09, 7.649145e+09, 7.816271e+09, 
    7.984841e+09, 8.154726e+09, 8.32579e+09, 8.497883e+09, 8.670843e+09, 
    8.844498e+09, 9.018663e+09, 9.193139e+09, 9.367718e+09, 9.542177e+09, 
    9.716282e+09, 9.88979e+09, 1.006244e+10, 1.023397e+10, 1.040409e+10, 
    1.057252e+10, 1.073895e+10, 1.090309e+10, 1.106461e+10, 1.12232e+10, 
    1.137852e+10, 1.153025e+10, 1.167804e+10, 1.182158e+10, 1.19605e+10, 
    1.209449e+10, 1.222321e+10, 1.234634e+10, 1.246355e+10, 1.257453e+10, 
    1.267899e+10, 1.277663e+10, 1.286718e+10, 1.295038e+10, 1.302599e+10, 
    1.309378e+10, 1.315356e+10, 1.320514e+10, 1.324837e+10, 1.328312e+10, 
    1.330927e+10, 1.332675e+10, 1.333551e+10, 1.333551e+10, 1.332675e+10, 
    1.330927e+10, 1.328312e+10, 1.324837e+10, 1.320514e+10, 1.315356e+10, 
    1.309378e+10, 1.302599e+10, 1.295038e+10, 1.286718e+10, 1.277663e+10, 
    1.267899e+10, 1.257453e+10, 1.246355e+10, 1.234634e+10, 1.222321e+10, 
    1.209449e+10, 1.19605e+10, 1.182158e+10, 1.167804e+10, 1.153025e+10, 
    1.137852e+10, 1.12232e+10, 1.106461e+10, 1.090309e+10, 1.073895e+10, 
    1.057252e+10, 1.040409e+10, 1.023397e+10, 1.006244e+10, 9.88979e+09, 
    9.716282e+09, 9.542177e+09, 9.367718e+09, 9.193139e+09, 9.018663e+09, 
    8.844498e+09, 8.670843e+09, 8.497883e+09, 8.32579e+09, 8.154726e+09, 
    7.984841e+09, 7.816271e+09, 7.649145e+09, 7.483577e+09, 7.319673e+09, 
    7.157529e+09,
  7.155078e+09, 7.316969e+09, 7.480609e+09, 7.645901e+09, 7.812741e+09, 
    7.981012e+09, 8.150589e+09, 8.321333e+09, 8.493095e+09, 8.665715e+09, 
    8.839017e+09, 9.012821e+09, 9.186927e+09, 9.361125e+09, 9.535196e+09, 
    9.708905e+09, 9.882009e+09, 1.005425e+10, 1.022536e+10, 1.039506e+10, 
    1.056306e+10, 1.072907e+10, 1.089278e+10, 1.105388e+10, 1.121203e+10, 
    1.136693e+10, 1.151823e+10, 1.166561e+10, 1.180873e+10, 1.194726e+10, 
    1.208085e+10, 1.220919e+10, 1.233195e+10, 1.24488e+10, 1.255944e+10, 
    1.266358e+10, 1.276091e+10, 1.285118e+10, 1.293411e+10, 1.300948e+10, 
    1.307706e+10, 1.313664e+10, 1.318806e+10, 1.323115e+10, 1.326578e+10, 
    1.329185e+10, 1.330927e+10, 1.3318e+10, 1.3318e+10, 1.330927e+10, 
    1.329185e+10, 1.326578e+10, 1.323115e+10, 1.318806e+10, 1.313664e+10, 
    1.307706e+10, 1.300948e+10, 1.293411e+10, 1.285118e+10, 1.276091e+10, 
    1.266358e+10, 1.255944e+10, 1.24488e+10, 1.233195e+10, 1.220919e+10, 
    1.208085e+10, 1.194726e+10, 1.180873e+10, 1.166561e+10, 1.151823e+10, 
    1.136693e+10, 1.121203e+10, 1.105388e+10, 1.089278e+10, 1.072907e+10, 
    1.056306e+10, 1.039506e+10, 1.022536e+10, 1.005425e+10, 9.882009e+09, 
    9.708905e+09, 9.535196e+09, 9.361125e+09, 9.186927e+09, 9.012821e+09, 
    8.839017e+09, 8.665715e+09, 8.493095e+09, 8.321333e+09, 8.150589e+09, 
    7.981012e+09, 7.812741e+09, 7.645901e+09, 7.480609e+09, 7.316969e+09, 
    7.155078e+09,
  7.151404e+09, 7.312915e+09, 7.476158e+09, 7.641037e+09, 7.807448e+09, 
    7.975273e+09, 8.144387e+09, 8.314652e+09, 8.485919e+09, 8.658028e+09, 
    8.830806e+09, 9.004068e+09, 9.177618e+09, 9.351248e+09, 9.524738e+09, 
    9.697854e+09, 9.870353e+09, 1.004198e+10, 1.021247e+10, 1.038154e+10, 
    1.054891e+10, 1.071428e+10, 1.087735e+10, 1.10378e+10, 1.119532e+10, 
    1.134958e+10, 1.150025e+10, 1.164701e+10, 1.178951e+10, 1.192743e+10, 
    1.206044e+10, 1.218821e+10, 1.231041e+10, 1.242673e+10, 1.253687e+10, 
    1.264052e+10, 1.273739e+10, 1.282723e+10, 1.290977e+10, 1.298478e+10, 
    1.305203e+10, 1.311133e+10, 1.316249e+10, 1.320537e+10, 1.323984e+10, 
    1.326578e+10, 1.328312e+10, 1.32918e+10, 1.32918e+10, 1.328312e+10, 
    1.326578e+10, 1.323984e+10, 1.320537e+10, 1.316249e+10, 1.311133e+10, 
    1.305203e+10, 1.298478e+10, 1.290977e+10, 1.282723e+10, 1.273739e+10, 
    1.264052e+10, 1.253687e+10, 1.242673e+10, 1.231041e+10, 1.218821e+10, 
    1.206044e+10, 1.192743e+10, 1.178951e+10, 1.164701e+10, 1.150025e+10, 
    1.134958e+10, 1.119532e+10, 1.10378e+10, 1.087735e+10, 1.071428e+10, 
    1.054891e+10, 1.038154e+10, 1.021247e+10, 1.004198e+10, 9.870353e+09, 
    9.697854e+09, 9.524738e+09, 9.351248e+09, 9.177618e+09, 9.004068e+09, 
    8.830806e+09, 8.658028e+09, 8.485919e+09, 8.314652e+09, 8.144387e+09, 
    7.975273e+09, 7.807448e+09, 7.641037e+09, 7.476158e+09, 7.312915e+09, 
    7.151404e+09,
  7.146505e+09, 7.307511e+09, 7.470226e+09, 7.634556e+09, 7.800395e+09, 
    7.967627e+09, 8.136126e+09, 8.305754e+09, 8.476363e+09, 8.647793e+09, 
    8.819871e+09, 8.992415e+09, 9.165227e+09, 9.338102e+09, 9.510819e+09, 
    9.683147e+09, 9.854844e+09, 1.002566e+10, 1.019532e+10, 1.036355e+10, 
    1.053008e+10, 1.06946e+10, 1.085682e+10, 1.101642e+10, 1.117309e+10, 
    1.13265e+10, 1.147634e+10, 1.162227e+10, 1.176396e+10, 1.190108e+10, 
    1.203331e+10, 1.216031e+10, 1.228178e+10, 1.23974e+10, 1.250686e+10, 
    1.260987e+10, 1.270614e+10, 1.279542e+10, 1.287743e+10, 1.295196e+10, 
    1.301878e+10, 1.30777e+10, 1.312854e+10, 1.317114e+10, 1.320537e+10, 
    1.323115e+10, 1.324837e+10, 1.3257e+10, 1.3257e+10, 1.324837e+10, 
    1.323115e+10, 1.320537e+10, 1.317114e+10, 1.312854e+10, 1.30777e+10, 
    1.301878e+10, 1.295196e+10, 1.287743e+10, 1.279542e+10, 1.270614e+10, 
    1.260987e+10, 1.250686e+10, 1.23974e+10, 1.228178e+10, 1.216031e+10, 
    1.203331e+10, 1.190108e+10, 1.176396e+10, 1.162227e+10, 1.147634e+10, 
    1.13265e+10, 1.117309e+10, 1.101642e+10, 1.085682e+10, 1.06946e+10, 
    1.053008e+10, 1.036355e+10, 1.019532e+10, 1.002566e+10, 9.854844e+09, 
    9.683147e+09, 9.510819e+09, 9.338102e+09, 9.165227e+09, 8.992415e+09, 
    8.819871e+09, 8.647793e+09, 8.476363e+09, 8.305754e+09, 8.136126e+09, 
    7.967627e+09, 7.800395e+09, 7.634556e+09, 7.470226e+09, 7.307511e+09, 
    7.146505e+09,
  7.140384e+09, 7.30076e+09, 7.462817e+09, 7.626462e+09, 7.791588e+09, 
    7.958081e+09, 8.125813e+09, 8.294647e+09, 8.464436e+09, 8.63502e+09, 
    8.806228e+09, 8.977876e+09, 9.14977e+09, 9.321703e+09, 9.49346e+09, 
    9.664807e+09, 9.835507e+09, 1.00053e+10, 1.017394e+10, 1.034114e+10, 
    1.050662e+10, 1.067009e+10, 1.083124e+10, 1.098979e+10, 1.11454e+10, 
    1.129776e+10, 1.144656e+10, 1.159146e+10, 1.173213e+10, 1.186826e+10, 
    1.199952e+10, 1.212559e+10, 1.224615e+10, 1.236089e+10, 1.246951e+10, 
    1.257172e+10, 1.266725e+10, 1.275582e+10, 1.283719e+10, 1.291113e+10, 
    1.297741e+10, 1.303585e+10, 1.308628e+10, 1.312854e+10, 1.316249e+10, 
    1.318806e+10, 1.320514e+10, 1.32137e+10, 1.32137e+10, 1.320514e+10, 
    1.318806e+10, 1.316249e+10, 1.312854e+10, 1.308628e+10, 1.303585e+10, 
    1.297741e+10, 1.291113e+10, 1.283719e+10, 1.275582e+10, 1.266725e+10, 
    1.257172e+10, 1.246951e+10, 1.236089e+10, 1.224615e+10, 1.212559e+10, 
    1.199952e+10, 1.186826e+10, 1.173213e+10, 1.159146e+10, 1.144656e+10, 
    1.129776e+10, 1.11454e+10, 1.098979e+10, 1.083124e+10, 1.067009e+10, 
    1.050662e+10, 1.034114e+10, 1.017394e+10, 1.00053e+10, 9.835507e+09, 
    9.664807e+09, 9.49346e+09, 9.321703e+09, 9.14977e+09, 8.977876e+09, 
    8.806228e+09, 8.63502e+09, 8.464436e+09, 8.294647e+09, 8.125813e+09, 
    7.958081e+09, 7.791588e+09, 7.626462e+09, 7.462817e+09, 7.30076e+09, 
    7.140384e+09,
  7.133041e+09, 7.292662e+09, 7.453934e+09, 7.616759e+09, 7.781033e+09, 
    7.946641e+09, 8.113456e+09, 8.281342e+09, 8.450151e+09, 8.619724e+09, 
    8.789891e+09, 8.96047e+09, 9.131267e+09, 9.302078e+09, 9.472687e+09, 
    9.642865e+09, 9.812372e+09, 9.980962e+09, 1.014837e+10, 1.031433e+10, 
    1.047856e+10, 1.064077e+10, 1.080067e+10, 1.095795e+10, 1.111231e+10, 
    1.126342e+10, 1.141097e+10, 1.155465e+10, 1.169412e+10, 1.182907e+10, 
    1.195917e+10, 1.208412e+10, 1.220359e+10, 1.231729e+10, 1.242492e+10, 
    1.252618e+10, 1.262082e+10, 1.270856e+10, 1.278916e+10, 1.286239e+10, 
    1.292804e+10, 1.298592e+10, 1.303585e+10, 1.30777e+10, 1.311133e+10, 
    1.313664e+10, 1.315356e+10, 1.316203e+10, 1.316203e+10, 1.315356e+10, 
    1.313664e+10, 1.311133e+10, 1.30777e+10, 1.303585e+10, 1.298592e+10, 
    1.292804e+10, 1.286239e+10, 1.278916e+10, 1.270856e+10, 1.262082e+10, 
    1.252618e+10, 1.242492e+10, 1.231729e+10, 1.220359e+10, 1.208412e+10, 
    1.195917e+10, 1.182907e+10, 1.169412e+10, 1.155465e+10, 1.141097e+10, 
    1.126342e+10, 1.111231e+10, 1.095795e+10, 1.080067e+10, 1.064077e+10, 
    1.047856e+10, 1.031433e+10, 1.014837e+10, 9.980962e+09, 9.812372e+09, 
    9.642865e+09, 9.472687e+09, 9.302078e+09, 9.131267e+09, 8.96047e+09, 
    8.789891e+09, 8.619724e+09, 8.450151e+09, 8.281342e+09, 8.113456e+09, 
    7.946641e+09, 7.781033e+09, 7.616759e+09, 7.453934e+09, 7.292662e+09, 
    7.133041e+09,
  7.124479e+09, 7.283223e+09, 7.443579e+09, 7.605452e+09, 7.768736e+09, 
    7.933316e+09, 8.099066e+09, 8.26585e+09, 8.433522e+09, 8.601922e+09, 
    8.770882e+09, 8.940219e+09, 9.109745e+09, 9.279254e+09, 9.448532e+09, 
    9.617354e+09, 9.785482e+09, 9.95267e+09, 1.011866e+10, 1.028319e+10, 
    1.044597e+10, 1.060673e+10, 1.076517e+10, 1.092099e+10, 1.107389e+10, 
    1.122356e+10, 1.136968e+10, 1.151193e+10, 1.165001e+10, 1.17836e+10, 
    1.191237e+10, 1.203602e+10, 1.215424e+10, 1.226673e+10, 1.237321e+10, 
    1.247338e+10, 1.256699e+10, 1.265377e+10, 1.273348e+10, 1.280589e+10, 
    1.287081e+10, 1.292804e+10, 1.297741e+10, 1.301878e+10, 1.305203e+10, 
    1.307706e+10, 1.309378e+10, 1.310215e+10, 1.310215e+10, 1.309378e+10, 
    1.307706e+10, 1.305203e+10, 1.301878e+10, 1.297741e+10, 1.292804e+10, 
    1.287081e+10, 1.280589e+10, 1.273348e+10, 1.265377e+10, 1.256699e+10, 
    1.247338e+10, 1.237321e+10, 1.226673e+10, 1.215424e+10, 1.203602e+10, 
    1.191237e+10, 1.17836e+10, 1.165001e+10, 1.151193e+10, 1.136968e+10, 
    1.122356e+10, 1.107389e+10, 1.092099e+10, 1.076517e+10, 1.060673e+10, 
    1.044597e+10, 1.028319e+10, 1.011866e+10, 9.95267e+09, 9.785482e+09, 
    9.617354e+09, 9.448532e+09, 9.279254e+09, 9.109745e+09, 8.940219e+09, 
    8.770882e+09, 8.601922e+09, 8.433522e+09, 8.26585e+09, 8.099066e+09, 
    7.933316e+09, 7.768736e+09, 7.605452e+09, 7.443579e+09, 7.283223e+09, 
    7.124479e+09,
  7.1147e+09, 7.272444e+09, 7.431758e+09, 7.592547e+09, 7.754704e+09, 
    7.918115e+09, 8.082655e+09, 8.248187e+09, 8.414565e+09, 8.581632e+09, 
    8.749221e+09, 8.917151e+09, 9.085231e+09, 9.253263e+09, 9.421031e+09, 
    9.588315e+09, 9.754878e+09, 9.920478e+09, 1.008486e+10, 1.024776e+10, 
    1.040891e+10, 1.056802e+10, 1.07248e+10, 1.087898e+10, 1.103023e+10, 
    1.117826e+10, 1.132276e+10, 1.146341e+10, 1.159992e+10, 1.173195e+10, 
    1.185922e+10, 1.198141e+10, 1.209821e+10, 1.220935e+10, 1.231452e+10, 
    1.241347e+10, 1.250591e+10, 1.25916e+10, 1.267031e+10, 1.27418e+10, 
    1.280589e+10, 1.286239e+10, 1.291113e+10, 1.295196e+10, 1.298478e+10, 
    1.300948e+10, 1.302599e+10, 1.303425e+10, 1.303425e+10, 1.302599e+10, 
    1.300948e+10, 1.298478e+10, 1.295196e+10, 1.291113e+10, 1.286239e+10, 
    1.280589e+10, 1.27418e+10, 1.267031e+10, 1.25916e+10, 1.250591e+10, 
    1.241347e+10, 1.231452e+10, 1.220935e+10, 1.209821e+10, 1.198141e+10, 
    1.185922e+10, 1.173195e+10, 1.159992e+10, 1.146341e+10, 1.132276e+10, 
    1.117826e+10, 1.103023e+10, 1.087898e+10, 1.07248e+10, 1.056802e+10, 
    1.040891e+10, 1.024776e+10, 1.008486e+10, 9.920478e+09, 9.754878e+09, 
    9.588315e+09, 9.421031e+09, 9.253263e+09, 9.085231e+09, 8.917151e+09, 
    8.749221e+09, 8.581632e+09, 8.414565e+09, 8.248187e+09, 8.082655e+09, 
    7.918115e+09, 7.754704e+09, 7.592547e+09, 7.431758e+09, 7.272444e+09, 
    7.1147e+09,
  7.103705e+09, 7.260329e+09, 7.418477e+09, 7.578052e+09, 7.738948e+09, 
    7.901051e+09, 8.064236e+09, 8.228367e+09, 8.3933e+09, 8.558878e+09, 
    8.724934e+09, 8.891291e+09, 9.05776e+09, 9.224142e+09, 9.390226e+09, 
    9.555794e+09, 9.720613e+09, 9.884442e+09, 1.004703e+10, 1.020812e+10, 
    1.036744e+10, 1.052472e+10, 1.067967e+10, 1.0832e+10, 1.098142e+10, 
    1.112763e+10, 1.127033e+10, 1.14092e+10, 1.154395e+10, 1.167428e+10, 
    1.179987e+10, 1.192043e+10, 1.203567e+10, 1.214529e+10, 1.224902e+10, 
    1.234659e+10, 1.243775e+10, 1.252223e+10, 1.259983e+10, 1.267031e+10, 
    1.273348e+10, 1.278916e+10, 1.283719e+10, 1.287743e+10, 1.290977e+10, 
    1.293411e+10, 1.295038e+10, 1.295852e+10, 1.295852e+10, 1.295038e+10, 
    1.293411e+10, 1.290977e+10, 1.287743e+10, 1.283719e+10, 1.278916e+10, 
    1.273348e+10, 1.267031e+10, 1.259983e+10, 1.252223e+10, 1.243775e+10, 
    1.234659e+10, 1.224902e+10, 1.214529e+10, 1.203567e+10, 1.192043e+10, 
    1.179987e+10, 1.167428e+10, 1.154395e+10, 1.14092e+10, 1.127033e+10, 
    1.112763e+10, 1.098142e+10, 1.0832e+10, 1.067967e+10, 1.052472e+10, 
    1.036744e+10, 1.020812e+10, 1.004703e+10, 9.884442e+09, 9.720613e+09, 
    9.555794e+09, 9.390226e+09, 9.224142e+09, 9.05776e+09, 8.891291e+09, 
    8.724934e+09, 8.558878e+09, 8.3933e+09, 8.228367e+09, 8.064236e+09, 
    7.901051e+09, 7.738948e+09, 7.578052e+09, 7.418477e+09, 7.260329e+09, 
    7.103705e+09,
  7.091497e+09, 7.246883e+09, 7.403741e+09, 7.561974e+09, 7.721477e+09, 
    7.882135e+09, 8.043825e+09, 8.20641e+09, 8.369748e+09, 8.533684e+09, 
    8.698051e+09, 8.862674e+09, 9.027367e+09, 9.191932e+09, 9.356163e+09, 
    9.519842e+09, 9.68274e+09, 9.844622e+09, 1.000524e+10, 1.016434e+10, 
    1.032166e+10, 1.047692e+10, 1.062985e+10, 1.078017e+10, 1.092757e+10, 
    1.107179e+10, 1.12125e+10, 1.134943e+10, 1.148226e+10, 1.16107e+10, 
    1.173446e+10, 1.185324e+10, 1.196675e+10, 1.207473e+10, 1.217688e+10, 
    1.227295e+10, 1.236269e+10, 1.244586e+10, 1.252223e+10, 1.25916e+10, 
    1.265377e+10, 1.270856e+10, 1.275582e+10, 1.279542e+10, 1.282723e+10, 
    1.285118e+10, 1.286718e+10, 1.287519e+10, 1.287519e+10, 1.286718e+10, 
    1.285118e+10, 1.282723e+10, 1.279542e+10, 1.275582e+10, 1.270856e+10, 
    1.265377e+10, 1.25916e+10, 1.252223e+10, 1.244586e+10, 1.236269e+10, 
    1.227295e+10, 1.217688e+10, 1.207473e+10, 1.196675e+10, 1.185324e+10, 
    1.173446e+10, 1.16107e+10, 1.148226e+10, 1.134943e+10, 1.12125e+10, 
    1.107179e+10, 1.092757e+10, 1.078017e+10, 1.062985e+10, 1.047692e+10, 
    1.032166e+10, 1.016434e+10, 1.000524e+10, 9.844622e+09, 9.68274e+09, 
    9.519842e+09, 9.356163e+09, 9.191932e+09, 9.027367e+09, 8.862674e+09, 
    8.698051e+09, 8.533684e+09, 8.369748e+09, 8.20641e+09, 8.043825e+09, 
    7.882135e+09, 7.721477e+09, 7.561974e+09, 7.403741e+09, 7.246883e+09, 
    7.091497e+09,
  7.078078e+09, 7.23211e+09, 7.387556e+09, 7.544322e+09, 7.702302e+09, 
    7.861382e+09, 8.021437e+09, 8.182336e+09, 8.343933e+09, 8.506077e+09, 
    8.668601e+09, 8.831335e+09, 8.994092e+09, 9.156679e+09, 9.318892e+09, 
    9.480515e+09, 9.641325e+09, 9.801088e+09, 9.959563e+09, 1.01165e+10, 
    1.027164e+10, 1.042471e+10, 1.057545e+10, 1.072358e+10, 1.08688e+10, 
    1.101085e+10, 1.114942e+10, 1.128423e+10, 1.141498e+10, 1.154138e+10, 
    1.166315e+10, 1.178001e+10, 1.189166e+10, 1.199784e+10, 1.209829e+10, 
    1.219274e+10, 1.228095e+10, 1.236269e+10, 1.243775e+10, 1.250591e+10, 
    1.256699e+10, 1.262082e+10, 1.266725e+10, 1.270614e+10, 1.273739e+10, 
    1.276091e+10, 1.277663e+10, 1.27845e+10, 1.27845e+10, 1.277663e+10, 
    1.276091e+10, 1.273739e+10, 1.270614e+10, 1.266725e+10, 1.262082e+10, 
    1.256699e+10, 1.250591e+10, 1.243775e+10, 1.236269e+10, 1.228095e+10, 
    1.219274e+10, 1.209829e+10, 1.199784e+10, 1.189166e+10, 1.178001e+10, 
    1.166315e+10, 1.154138e+10, 1.141498e+10, 1.128423e+10, 1.114942e+10, 
    1.101085e+10, 1.08688e+10, 1.072358e+10, 1.057545e+10, 1.042471e+10, 
    1.027164e+10, 1.01165e+10, 9.959563e+09, 9.801088e+09, 9.641325e+09, 
    9.480515e+09, 9.318892e+09, 9.156679e+09, 8.994092e+09, 8.831335e+09, 
    8.668601e+09, 8.506077e+09, 8.343933e+09, 8.182336e+09, 8.021437e+09, 
    7.861382e+09, 7.702302e+09, 7.544322e+09, 7.387556e+09, 7.23211e+09, 
    7.078078e+09,
  7.063453e+09, 7.216014e+09, 7.36993e+09, 7.525106e+09, 7.681435e+09, 
    7.838806e+09, 7.997093e+09, 8.156166e+09, 8.31588e+09, 8.476086e+09, 
    8.636621e+09, 8.797313e+09, 8.95798e+09, 9.118431e+09, 9.278465e+09, 
    9.437871e+09, 9.596429e+09, 9.753911e+09, 9.910078e+09, 1.006469e+10, 
    1.021748e+10, 1.03682e+10, 1.051658e+10, 1.066235e+10, 1.080523e+10, 
    1.094495e+10, 1.108122e+10, 1.121375e+10, 1.134227e+10, 1.146649e+10, 
    1.158613e+10, 1.170091e+10, 1.181057e+10, 1.191483e+10, 1.201345e+10, 
    1.210616e+10, 1.219274e+10, 1.227295e+10, 1.234659e+10, 1.241347e+10, 
    1.247338e+10, 1.252618e+10, 1.257172e+10, 1.260987e+10, 1.264052e+10, 
    1.266358e+10, 1.267899e+10, 1.268671e+10, 1.268671e+10, 1.267899e+10, 
    1.266358e+10, 1.264052e+10, 1.260987e+10, 1.257172e+10, 1.252618e+10, 
    1.247338e+10, 1.241347e+10, 1.234659e+10, 1.227295e+10, 1.219274e+10, 
    1.210616e+10, 1.201345e+10, 1.191483e+10, 1.181057e+10, 1.170091e+10, 
    1.158613e+10, 1.146649e+10, 1.134227e+10, 1.121375e+10, 1.108122e+10, 
    1.094495e+10, 1.080523e+10, 1.066235e+10, 1.051658e+10, 1.03682e+10, 
    1.021748e+10, 1.006469e+10, 9.910078e+09, 9.753911e+09, 9.596429e+09, 
    9.437871e+09, 9.278465e+09, 9.118431e+09, 8.95798e+09, 8.797313e+09, 
    8.636621e+09, 8.476086e+09, 8.31588e+09, 8.156166e+09, 7.997093e+09, 
    7.838806e+09, 7.681435e+09, 7.525106e+09, 7.36993e+09, 7.216014e+09, 
    7.063453e+09,
  7.047623e+09, 7.198601e+09, 7.350871e+09, 7.504335e+09, 7.65889e+09, 
    7.814423e+09, 7.970811e+09, 8.127923e+09, 8.285618e+09, 8.443745e+09, 
    8.602145e+09, 8.760649e+09, 8.919077e+09, 9.077242e+09, 9.234944e+09, 
    9.391978e+09, 9.548129e+09, 9.703171e+09, 9.856871e+09, 1.000899e+10, 
    1.015928e+10, 1.030749e+10, 1.045336e+10, 1.059662e+10, 1.0737e+10, 
    1.087423e+10, 1.100805e+10, 1.113816e+10, 1.12643e+10, 1.13862e+10, 
    1.150357e+10, 1.161615e+10, 1.172369e+10, 1.182591e+10, 1.192258e+10, 
    1.201345e+10, 1.209829e+10, 1.217688e+10, 1.224902e+10, 1.231452e+10, 
    1.237321e+10, 1.242492e+10, 1.246951e+10, 1.250686e+10, 1.253687e+10, 
    1.255944e+10, 1.257453e+10, 1.258209e+10, 1.258209e+10, 1.257453e+10, 
    1.255944e+10, 1.253687e+10, 1.250686e+10, 1.246951e+10, 1.242492e+10, 
    1.237321e+10, 1.231452e+10, 1.224902e+10, 1.217688e+10, 1.209829e+10, 
    1.201345e+10, 1.192258e+10, 1.182591e+10, 1.172369e+10, 1.161615e+10, 
    1.150357e+10, 1.13862e+10, 1.12643e+10, 1.113816e+10, 1.100805e+10, 
    1.087423e+10, 1.0737e+10, 1.059662e+10, 1.045336e+10, 1.030749e+10, 
    1.015928e+10, 1.000899e+10, 9.856871e+09, 9.703171e+09, 9.548129e+09, 
    9.391978e+09, 9.234944e+09, 9.077242e+09, 8.919077e+09, 8.760649e+09, 
    8.602145e+09, 8.443745e+09, 8.285618e+09, 8.127923e+09, 7.970811e+09, 
    7.814423e+09, 7.65889e+09, 7.504335e+09, 7.350871e+09, 7.198601e+09, 
    7.047623e+09,
  7.030593e+09, 7.179877e+09, 7.330385e+09, 7.482021e+09, 7.634681e+09, 
    7.788252e+09, 7.942612e+09, 8.097633e+09, 8.253174e+09, 8.409087e+09, 
    8.565214e+09, 8.721389e+09, 8.877434e+09, 9.033167e+09, 9.188391e+09, 
    9.342905e+09, 9.496498e+09, 9.64895e+09, 9.800034e+09, 9.949515e+09, 
    1.009715e+10, 1.02427e+10, 1.03859e+10, 1.05265e+10, 1.066424e+10, 
    1.079885e+10, 1.093007e+10, 1.105763e+10, 1.118125e+10, 1.130069e+10, 
    1.141567e+10, 1.152593e+10, 1.163122e+10, 1.17313e+10, 1.182591e+10, 
    1.191483e+10, 1.199784e+10, 1.207473e+10, 1.214529e+10, 1.220935e+10, 
    1.226673e+10, 1.231729e+10, 1.236089e+10, 1.23974e+10, 1.242673e+10, 
    1.24488e+10, 1.246355e+10, 1.247093e+10, 1.247093e+10, 1.246355e+10, 
    1.24488e+10, 1.242673e+10, 1.23974e+10, 1.236089e+10, 1.231729e+10, 
    1.226673e+10, 1.220935e+10, 1.214529e+10, 1.207473e+10, 1.199784e+10, 
    1.191483e+10, 1.182591e+10, 1.17313e+10, 1.163122e+10, 1.152593e+10, 
    1.141567e+10, 1.130069e+10, 1.118125e+10, 1.105763e+10, 1.093007e+10, 
    1.079885e+10, 1.066424e+10, 1.05265e+10, 1.03859e+10, 1.02427e+10, 
    1.009715e+10, 9.949515e+09, 9.800034e+09, 9.64895e+09, 9.496498e+09, 
    9.342905e+09, 9.188391e+09, 9.033167e+09, 8.877434e+09, 8.721389e+09, 
    8.565214e+09, 8.409087e+09, 8.253174e+09, 8.097633e+09, 7.942612e+09, 
    7.788252e+09, 7.634681e+09, 7.482021e+09, 7.330385e+09, 7.179877e+09, 
    7.030593e+09,
  7.012366e+09, 7.159848e+09, 7.308484e+09, 7.458176e+09, 7.608822e+09, 
    7.760311e+09, 7.912521e+09, 8.065324e+09, 8.218582e+09, 8.372148e+09, 
    8.525868e+09, 8.679578e+09, 8.833104e+09, 8.986266e+09, 9.138871e+09, 
    9.290724e+09, 9.441618e+09, 9.591338e+09, 9.739662e+09, 9.886363e+09, 
    1.00312e+10, 1.017395e+10, 1.031435e+10, 1.045215e+10, 1.058711e+10, 
    1.071896e+10, 1.084745e+10, 1.097232e+10, 1.109331e+10, 1.121017e+10, 
    1.132264e+10, 1.143046e+10, 1.153341e+10, 1.163122e+10, 1.172369e+10, 
    1.181057e+10, 1.189166e+10, 1.196675e+10, 1.203567e+10, 1.209821e+10, 
    1.215424e+10, 1.220359e+10, 1.224615e+10, 1.228178e+10, 1.231041e+10, 
    1.233195e+10, 1.234634e+10, 1.235355e+10, 1.235355e+10, 1.234634e+10, 
    1.233195e+10, 1.231041e+10, 1.228178e+10, 1.224615e+10, 1.220359e+10, 
    1.215424e+10, 1.209821e+10, 1.203567e+10, 1.196675e+10, 1.189166e+10, 
    1.181057e+10, 1.172369e+10, 1.163122e+10, 1.153341e+10, 1.143046e+10, 
    1.132264e+10, 1.121017e+10, 1.109331e+10, 1.097232e+10, 1.084745e+10, 
    1.071896e+10, 1.058711e+10, 1.045215e+10, 1.031435e+10, 1.017395e+10, 
    1.00312e+10, 9.886363e+09, 9.739662e+09, 9.591338e+09, 9.441618e+09, 
    9.290724e+09, 9.138871e+09, 8.986266e+09, 8.833104e+09, 8.679578e+09, 
    8.525868e+09, 8.372148e+09, 8.218582e+09, 8.065324e+09, 7.912521e+09, 
    7.760311e+09, 7.608822e+09, 7.458176e+09, 7.308484e+09, 7.159848e+09, 
    7.012366e+09,
  6.992947e+09, 7.138521e+09, 7.285175e+09, 7.432813e+09, 7.581331e+09, 
    7.73062e+09, 7.880559e+09, 8.031022e+09, 8.181873e+09, 8.332967e+09, 
    8.484152e+09, 8.635267e+09, 8.786142e+09, 8.936601e+09, 9.086456e+09, 
    9.235513e+09, 9.383574e+09, 9.530426e+09, 9.675857e+09, 9.819643e+09, 
    9.961556e+09, 1.010136e+10, 1.023883e+10, 1.037371e+10, 1.050575e+10, 
    1.063472e+10, 1.076036e+10, 1.088243e+10, 1.100067e+10, 1.111483e+10, 
    1.122468e+10, 1.132997e+10, 1.143046e+10, 1.152593e+10, 1.161615e+10, 
    1.170091e+10, 1.178001e+10, 1.185324e+10, 1.192043e+10, 1.198141e+10, 
    1.203602e+10, 1.208412e+10, 1.212559e+10, 1.216031e+10, 1.218821e+10, 
    1.220919e+10, 1.222321e+10, 1.223023e+10, 1.223023e+10, 1.222321e+10, 
    1.220919e+10, 1.218821e+10, 1.216031e+10, 1.212559e+10, 1.208412e+10, 
    1.203602e+10, 1.198141e+10, 1.192043e+10, 1.185324e+10, 1.178001e+10, 
    1.170091e+10, 1.161615e+10, 1.152593e+10, 1.143046e+10, 1.132997e+10, 
    1.122468e+10, 1.111483e+10, 1.100067e+10, 1.088243e+10, 1.076036e+10, 
    1.063472e+10, 1.050575e+10, 1.037371e+10, 1.023883e+10, 1.010136e+10, 
    9.961556e+09, 9.819643e+09, 9.675857e+09, 9.530426e+09, 9.383574e+09, 
    9.235513e+09, 9.086456e+09, 8.936601e+09, 8.786142e+09, 8.635267e+09, 
    8.484152e+09, 8.332967e+09, 8.181873e+09, 8.031022e+09, 7.880559e+09, 
    7.73062e+09, 7.581331e+09, 7.432813e+09, 7.285175e+09, 7.138521e+09, 
    6.992947e+09,
  6.972339e+09, 7.115902e+09, 7.260469e+09, 7.405943e+09, 7.552224e+09, 
    7.699199e+09, 7.846753e+09, 7.994759e+09, 8.143084e+09, 8.291585e+09, 
    8.440113e+09, 8.58851e+09, 8.736609e+09, 8.884238e+09, 9.031216e+09, 
    9.177352e+09, 9.322452e+09, 9.466312e+09, 9.608722e+09, 9.749469e+09, 
    9.88833e+09, 1.002508e+10, 1.015949e+10, 1.029132e+10, 1.042034e+10, 
    1.054631e+10, 1.066899e+10, 1.078814e+10, 1.090352e+10, 1.10149e+10, 
    1.112203e+10, 1.122468e+10, 1.132264e+10, 1.141567e+10, 1.150357e+10, 
    1.158613e+10, 1.166315e+10, 1.173446e+10, 1.179987e+10, 1.185922e+10, 
    1.191237e+10, 1.195917e+10, 1.199952e+10, 1.203331e+10, 1.206044e+10, 
    1.208085e+10, 1.209449e+10, 1.210132e+10, 1.210132e+10, 1.209449e+10, 
    1.208085e+10, 1.206044e+10, 1.203331e+10, 1.199952e+10, 1.195917e+10, 
    1.191237e+10, 1.185922e+10, 1.179987e+10, 1.173446e+10, 1.166315e+10, 
    1.158613e+10, 1.150357e+10, 1.141567e+10, 1.132264e+10, 1.122468e+10, 
    1.112203e+10, 1.10149e+10, 1.090352e+10, 1.078814e+10, 1.066899e+10, 
    1.054631e+10, 1.042034e+10, 1.029132e+10, 1.015949e+10, 1.002508e+10, 
    9.88833e+09, 9.749469e+09, 9.608722e+09, 9.466312e+09, 9.322452e+09, 
    9.177352e+09, 9.031216e+09, 8.884238e+09, 8.736609e+09, 8.58851e+09, 
    8.440113e+09, 8.291585e+09, 8.143084e+09, 7.994759e+09, 7.846753e+09, 
    7.699199e+09, 7.552224e+09, 7.405943e+09, 7.260469e+09, 7.115902e+09, 
    6.972339e+09,
  6.950547e+09, 7.092e+09, 7.234377e+09, 7.377583e+09, 7.521518e+09, 
    7.666072e+09, 7.811129e+09, 7.956566e+09, 8.10225e+09, 8.248043e+09, 
    8.393798e+09, 8.539359e+09, 8.684566e+09, 8.829247e+09, 8.973229e+09, 
    9.116325e+09, 9.258346e+09, 9.399095e+09, 9.53837e+09, 9.67596e+09, 
    9.811654e+09, 9.945231e+09, 1.007647e+10, 1.020515e+10, 1.033104e+10, 
    1.045391e+10, 1.057352e+10, 1.068966e+10, 1.080209e+10, 1.091057e+10, 
    1.10149e+10, 1.111483e+10, 1.121017e+10, 1.130069e+10, 1.13862e+10, 
    1.146649e+10, 1.154138e+10, 1.16107e+10, 1.167428e+10, 1.173195e+10, 
    1.17836e+10, 1.182907e+10, 1.186826e+10, 1.190108e+10, 1.192743e+10, 
    1.194726e+10, 1.19605e+10, 1.196713e+10, 1.196713e+10, 1.19605e+10, 
    1.194726e+10, 1.192743e+10, 1.190108e+10, 1.186826e+10, 1.182907e+10, 
    1.17836e+10, 1.173195e+10, 1.167428e+10, 1.16107e+10, 1.154138e+10, 
    1.146649e+10, 1.13862e+10, 1.130069e+10, 1.121017e+10, 1.111483e+10, 
    1.10149e+10, 1.091057e+10, 1.080209e+10, 1.068966e+10, 1.057352e+10, 
    1.045391e+10, 1.033104e+10, 1.020515e+10, 1.007647e+10, 9.945231e+09, 
    9.811654e+09, 9.67596e+09, 9.53837e+09, 9.399095e+09, 9.258346e+09, 
    9.116325e+09, 8.973229e+09, 8.829247e+09, 8.684566e+09, 8.539359e+09, 
    8.393798e+09, 8.248043e+09, 8.10225e+09, 7.956566e+09, 7.811129e+09, 
    7.666072e+09, 7.521518e+09, 7.377583e+09, 7.234377e+09, 7.092e+09, 
    6.950547e+09,
  6.927576e+09, 7.066821e+09, 7.206909e+09, 7.347746e+09, 7.489233e+09, 
    7.631261e+09, 7.773715e+09, 7.916475e+09, 8.059411e+09, 8.202386e+09, 
    8.345257e+09, 8.487873e+09, 8.630074e+09, 8.771699e+09, 8.912572e+09, 
    9.052518e+09, 9.191351e+09, 9.32888e+09, 9.464909e+09, 9.599237e+09, 
    9.731658e+09, 9.861961e+09, 9.989933e+09, 1.011536e+10, 1.023802e+10, 
    1.035769e+10, 1.047415e+10, 1.058718e+10, 1.069657e+10, 1.080209e+10, 
    1.090352e+10, 1.100067e+10, 1.109331e+10, 1.118125e+10, 1.12643e+10, 
    1.134227e+10, 1.141498e+10, 1.148226e+10, 1.154395e+10, 1.159992e+10, 
    1.165001e+10, 1.169412e+10, 1.173213e+10, 1.176396e+10, 1.178951e+10, 
    1.180873e+10, 1.182158e+10, 1.1828e+10, 1.1828e+10, 1.182158e+10, 
    1.180873e+10, 1.178951e+10, 1.176396e+10, 1.173213e+10, 1.169412e+10, 
    1.165001e+10, 1.159992e+10, 1.154395e+10, 1.148226e+10, 1.141498e+10, 
    1.134227e+10, 1.12643e+10, 1.118125e+10, 1.109331e+10, 1.100067e+10, 
    1.090352e+10, 1.080209e+10, 1.069657e+10, 1.058718e+10, 1.047415e+10, 
    1.035769e+10, 1.023802e+10, 1.011536e+10, 9.989933e+09, 9.861961e+09, 
    9.731658e+09, 9.599237e+09, 9.464909e+09, 9.32888e+09, 9.191351e+09, 
    9.052518e+09, 8.912572e+09, 8.771699e+09, 8.630074e+09, 8.487873e+09, 
    8.345257e+09, 8.202386e+09, 8.059411e+09, 7.916475e+09, 7.773715e+09, 
    7.631261e+09, 7.489233e+09, 7.347746e+09, 7.206909e+09, 7.066821e+09, 
    6.927576e+09,
  6.903431e+09, 7.040374e+09, 7.178077e+09, 7.316448e+09, 7.455388e+09, 
    7.594789e+09, 7.734541e+09, 7.874522e+09, 8.014606e+09, 8.15466e+09, 
    8.294543e+09, 8.434108e+09, 8.573202e+09, 8.711665e+09, 8.849328e+09, 
    8.986021e+09, 9.121564e+09, 9.255772e+09, 9.388457e+09, 9.519426e+09, 
    9.648477e+09, 9.775411e+09, 9.900023e+09, 1.00221e+10, 1.014144e+10, 
    1.025783e+10, 1.037106e+10, 1.048091e+10, 1.058718e+10, 1.068966e+10, 
    1.078814e+10, 1.088243e+10, 1.097232e+10, 1.105763e+10, 1.113816e+10, 
    1.121375e+10, 1.128423e+10, 1.134943e+10, 1.14092e+10, 1.146341e+10, 
    1.151193e+10, 1.155465e+10, 1.159146e+10, 1.162227e+10, 1.164701e+10, 
    1.166561e+10, 1.167804e+10, 1.168427e+10, 1.168427e+10, 1.167804e+10, 
    1.166561e+10, 1.164701e+10, 1.162227e+10, 1.159146e+10, 1.155465e+10, 
    1.151193e+10, 1.146341e+10, 1.14092e+10, 1.134943e+10, 1.128423e+10, 
    1.121375e+10, 1.113816e+10, 1.105763e+10, 1.097232e+10, 1.088243e+10, 
    1.078814e+10, 1.068966e+10, 1.058718e+10, 1.048091e+10, 1.037106e+10, 
    1.025783e+10, 1.014144e+10, 1.00221e+10, 9.900023e+09, 9.775411e+09, 
    9.648477e+09, 9.519426e+09, 9.388457e+09, 9.255772e+09, 9.121564e+09, 
    8.986021e+09, 8.849328e+09, 8.711665e+09, 8.573202e+09, 8.434108e+09, 
    8.294543e+09, 8.15466e+09, 8.014606e+09, 7.874522e+09, 7.734541e+09, 
    7.594789e+09, 7.455388e+09, 7.316448e+09, 7.178077e+09, 7.040374e+09, 
    6.903431e+09,
  6.878117e+09, 7.012667e+09, 7.147894e+09, 7.283705e+09, 7.420003e+09, 
    7.556683e+09, 7.693634e+09, 7.830739e+09, 7.967875e+09, 8.10491e+09, 
    8.241709e+09, 8.378128e+09, 8.514017e+09, 8.649221e+09, 8.78358e+09, 
    8.916924e+09, 9.049084e+09, 9.17988e+09, 9.309132e+09, 9.436652e+09, 
    9.562249e+09, 9.68573e+09, 9.806899e+09, 9.925557e+09, 1.00415e+10, 
    1.015454e+10, 1.026446e+10, 1.037106e+10, 1.047415e+10, 1.057352e+10, 
    1.066899e+10, 1.076036e+10, 1.084745e+10, 1.093007e+10, 1.100805e+10, 
    1.108122e+10, 1.114942e+10, 1.12125e+10, 1.127033e+10, 1.132276e+10, 
    1.136968e+10, 1.141097e+10, 1.144656e+10, 1.147634e+10, 1.150025e+10, 
    1.151823e+10, 1.153025e+10, 1.153626e+10, 1.153626e+10, 1.153025e+10, 
    1.151823e+10, 1.150025e+10, 1.147634e+10, 1.144656e+10, 1.141097e+10, 
    1.136968e+10, 1.132276e+10, 1.127033e+10, 1.12125e+10, 1.114942e+10, 
    1.108122e+10, 1.100805e+10, 1.093007e+10, 1.084745e+10, 1.076036e+10, 
    1.066899e+10, 1.057352e+10, 1.047415e+10, 1.037106e+10, 1.026446e+10, 
    1.015454e+10, 1.00415e+10, 9.925557e+09, 9.806899e+09, 9.68573e+09, 
    9.562249e+09, 9.436652e+09, 9.309132e+09, 9.17988e+09, 9.049084e+09, 
    8.916924e+09, 8.78358e+09, 8.649221e+09, 8.514017e+09, 8.378128e+09, 
    8.241709e+09, 8.10491e+09, 7.967875e+09, 7.830739e+09, 7.693634e+09, 
    7.556683e+09, 7.420003e+09, 7.283705e+09, 7.147894e+09, 7.012667e+09, 
    6.878117e+09,
  6.851641e+09, 6.98371e+09, 7.116371e+09, 7.249533e+09, 7.383099e+09, 
    7.516966e+09, 7.651027e+09, 7.785166e+09, 7.919261e+09, 8.053188e+09, 
    8.186811e+09, 8.319992e+09, 8.452588e+09, 8.584445e+09, 8.715411e+09, 
    8.845323e+09, 8.974015e+09, 9.101317e+09, 9.227054e+09, 9.351046e+09, 
    9.473112e+09, 9.593066e+09, 9.710721e+09, 9.825887e+09, 9.938373e+09, 
    1.004799e+10, 1.015454e+10, 1.025783e+10, 1.035769e+10, 1.045391e+10, 
    1.054631e+10, 1.063472e+10, 1.071896e+10, 1.079885e+10, 1.087423e+10, 
    1.094495e+10, 1.101085e+10, 1.107179e+10, 1.112763e+10, 1.117826e+10, 
    1.122356e+10, 1.126342e+10, 1.129776e+10, 1.13265e+10, 1.134958e+10, 
    1.136693e+10, 1.137852e+10, 1.138432e+10, 1.138432e+10, 1.137852e+10, 
    1.136693e+10, 1.134958e+10, 1.13265e+10, 1.129776e+10, 1.126342e+10, 
    1.122356e+10, 1.117826e+10, 1.112763e+10, 1.107179e+10, 1.101085e+10, 
    1.094495e+10, 1.087423e+10, 1.079885e+10, 1.071896e+10, 1.063472e+10, 
    1.054631e+10, 1.045391e+10, 1.035769e+10, 1.025783e+10, 1.015454e+10, 
    1.004799e+10, 9.938373e+09, 9.825887e+09, 9.710721e+09, 9.593066e+09, 
    9.473112e+09, 9.351046e+09, 9.227054e+09, 9.101317e+09, 8.974015e+09, 
    8.845323e+09, 8.715411e+09, 8.584445e+09, 8.452588e+09, 8.319992e+09, 
    8.186811e+09, 8.053188e+09, 7.919261e+09, 7.785166e+09, 7.651027e+09, 
    7.516966e+09, 7.383099e+09, 7.249533e+09, 7.116371e+09, 6.98371e+09, 
    6.851641e+09,
  6.824007e+09, 6.953512e+09, 7.083523e+09, 7.21395e+09, 7.344698e+09, 
    7.475667e+09, 7.606751e+09, 7.737838e+09, 7.868808e+09, 7.99954e+09, 
    8.129904e+09, 8.259766e+09, 8.388985e+09, 8.517416e+09, 8.64491e+09, 
    8.771312e+09, 8.896461e+09, 9.020195e+09, 9.142345e+09, 9.262742e+09, 
    9.381209e+09, 9.497571e+09, 9.61165e+09, 9.723264e+09, 9.832232e+09, 
    9.938373e+09, 1.00415e+10, 1.014144e+10, 1.023802e+10, 1.033104e+10, 
    1.042034e+10, 1.050575e+10, 1.058711e+10, 1.066424e+10, 1.0737e+10, 
    1.080523e+10, 1.08688e+10, 1.092757e+10, 1.098142e+10, 1.103023e+10, 
    1.107389e+10, 1.111231e+10, 1.11454e+10, 1.117309e+10, 1.119532e+10, 
    1.121203e+10, 1.12232e+10, 1.122879e+10, 1.122879e+10, 1.12232e+10, 
    1.121203e+10, 1.119532e+10, 1.117309e+10, 1.11454e+10, 1.111231e+10, 
    1.107389e+10, 1.103023e+10, 1.098142e+10, 1.092757e+10, 1.08688e+10, 
    1.080523e+10, 1.0737e+10, 1.066424e+10, 1.058711e+10, 1.050575e+10, 
    1.042034e+10, 1.033104e+10, 1.023802e+10, 1.014144e+10, 1.00415e+10, 
    9.938373e+09, 9.832232e+09, 9.723264e+09, 9.61165e+09, 9.497571e+09, 
    9.381209e+09, 9.262742e+09, 9.142345e+09, 9.020195e+09, 8.896461e+09, 
    8.771312e+09, 8.64491e+09, 8.517416e+09, 8.388985e+09, 8.259766e+09, 
    8.129904e+09, 7.99954e+09, 7.868808e+09, 7.737838e+09, 7.606751e+09, 
    7.475667e+09, 7.344698e+09, 7.21395e+09, 7.083523e+09, 6.953512e+09, 
    6.824007e+09,
  6.795221e+09, 6.922081e+09, 7.049361e+09, 7.176973e+09, 7.304823e+09, 
    7.432814e+09, 7.56084e+09, 7.688794e+09, 7.816561e+09, 7.94402e+09, 
    8.071048e+09, 8.197513e+09, 8.323282e+09, 8.448214e+09, 8.572165e+09, 
    8.694987e+09, 8.816526e+09, 8.936627e+09, 9.055129e+09, 9.171869e+09, 
    9.286681e+09, 9.399396e+09, 9.509846e+09, 9.61786e+09, 9.723264e+09, 
    9.825887e+09, 9.925557e+09, 1.00221e+10, 1.011536e+10, 1.020515e+10, 
    1.029132e+10, 1.037371e+10, 1.045215e+10, 1.05265e+10, 1.059662e+10, 
    1.066235e+10, 1.072358e+10, 1.078017e+10, 1.0832e+10, 1.087898e+10, 
    1.092099e+10, 1.095795e+10, 1.098979e+10, 1.101642e+10, 1.10378e+10, 
    1.105388e+10, 1.106461e+10, 1.106999e+10, 1.106999e+10, 1.106461e+10, 
    1.105388e+10, 1.10378e+10, 1.101642e+10, 1.098979e+10, 1.095795e+10, 
    1.092099e+10, 1.087898e+10, 1.0832e+10, 1.078017e+10, 1.072358e+10, 
    1.066235e+10, 1.059662e+10, 1.05265e+10, 1.045215e+10, 1.037371e+10, 
    1.029132e+10, 1.020515e+10, 1.011536e+10, 1.00221e+10, 9.925557e+09, 
    9.825887e+09, 9.723264e+09, 9.61786e+09, 9.509846e+09, 9.399396e+09, 
    9.286681e+09, 9.171869e+09, 9.055129e+09, 8.936627e+09, 8.816526e+09, 
    8.694987e+09, 8.572165e+09, 8.448214e+09, 8.323282e+09, 8.197513e+09, 
    8.071048e+09, 7.94402e+09, 7.816561e+09, 7.688794e+09, 7.56084e+09, 
    7.432814e+09, 7.304823e+09, 7.176973e+09, 7.049361e+09, 6.922081e+09, 
    6.795221e+09,
  6.76529e+09, 6.889429e+09, 7.013901e+09, 7.13862e+09, 7.263496e+09, 
    7.388432e+09, 7.513327e+09, 7.638074e+09, 7.762563e+09, 7.886679e+09, 
    8.010299e+09, 8.133301e+09, 8.255552e+09, 8.37692e+09, 8.497266e+09, 
    8.616447e+09, 8.734319e+09, 8.85073e+09, 8.96553e+09, 9.078562e+09, 
    9.18967e+09, 9.298694e+09, 9.405474e+09, 9.509846e+09, 9.61165e+09, 
    9.710721e+09, 9.806899e+09, 9.900023e+09, 9.989933e+09, 1.007647e+10, 
    1.015949e+10, 1.023883e+10, 1.031435e+10, 1.03859e+10, 1.045336e+10, 
    1.051658e+10, 1.057545e+10, 1.062985e+10, 1.067967e+10, 1.07248e+10, 
    1.076517e+10, 1.080067e+10, 1.083124e+10, 1.085682e+10, 1.087735e+10, 
    1.089278e+10, 1.090309e+10, 1.090825e+10, 1.090825e+10, 1.090309e+10, 
    1.089278e+10, 1.087735e+10, 1.085682e+10, 1.083124e+10, 1.080067e+10, 
    1.076517e+10, 1.07248e+10, 1.067967e+10, 1.062985e+10, 1.057545e+10, 
    1.051658e+10, 1.045336e+10, 1.03859e+10, 1.031435e+10, 1.023883e+10, 
    1.015949e+10, 1.007647e+10, 9.989933e+09, 9.900023e+09, 9.806899e+09, 
    9.710721e+09, 9.61165e+09, 9.509846e+09, 9.405474e+09, 9.298694e+09, 
    9.18967e+09, 9.078562e+09, 8.96553e+09, 8.85073e+09, 8.734319e+09, 
    8.616447e+09, 8.497266e+09, 8.37692e+09, 8.255552e+09, 8.133301e+09, 
    8.010299e+09, 7.886679e+09, 7.762563e+09, 7.638074e+09, 7.513327e+09, 
    7.388432e+09, 7.263496e+09, 7.13862e+09, 7.013901e+09, 6.889429e+09, 
    6.76529e+09,
  6.734221e+09, 6.855565e+09, 6.977157e+09, 7.098912e+09, 7.220742e+09, 
    7.342552e+09, 7.464245e+09, 7.585717e+09, 7.706863e+09, 7.827569e+09, 
    7.94772e+09, 8.067195e+09, 8.18587e+09, 8.303616e+09, 8.420301e+09, 
    8.53579e+09, 8.649944e+09, 8.762619e+09, 8.873673e+09, 8.982957e+09, 
    9.090322e+09, 9.195619e+09, 9.298694e+09, 9.399396e+09, 9.497571e+09, 
    9.593066e+09, 9.68573e+09, 9.775411e+09, 9.861961e+09, 9.945231e+09, 
    1.002508e+10, 1.010136e+10, 1.017395e+10, 1.02427e+10, 1.030749e+10, 
    1.03682e+10, 1.042471e+10, 1.047692e+10, 1.052472e+10, 1.056802e+10, 
    1.060673e+10, 1.064077e+10, 1.067009e+10, 1.06946e+10, 1.071428e+10, 
    1.072907e+10, 1.073895e+10, 1.07439e+10, 1.07439e+10, 1.073895e+10, 
    1.072907e+10, 1.071428e+10, 1.06946e+10, 1.067009e+10, 1.064077e+10, 
    1.060673e+10, 1.056802e+10, 1.052472e+10, 1.047692e+10, 1.042471e+10, 
    1.03682e+10, 1.030749e+10, 1.02427e+10, 1.017395e+10, 1.010136e+10, 
    1.002508e+10, 9.945231e+09, 9.861961e+09, 9.775411e+09, 9.68573e+09, 
    9.593066e+09, 9.497571e+09, 9.399396e+09, 9.298694e+09, 9.195619e+09, 
    9.090322e+09, 8.982957e+09, 8.873673e+09, 8.762619e+09, 8.649944e+09, 
    8.53579e+09, 8.420301e+09, 8.303616e+09, 8.18587e+09, 8.067195e+09, 
    7.94772e+09, 7.827569e+09, 7.706863e+09, 7.585717e+09, 7.464245e+09, 
    7.342552e+09, 7.220742e+09, 7.098912e+09, 6.977157e+09, 6.855565e+09, 
    6.734221e+09,
  6.702019e+09, 6.8205e+09, 6.939143e+09, 7.057866e+09, 7.176583e+09, 
    7.295202e+09, 7.41363e+09, 7.531766e+09, 7.649507e+09, 7.766745e+09, 
    7.883369e+09, 7.999264e+09, 8.11431e+09, 8.228386e+09, 8.341364e+09, 
    8.453116e+09, 8.563511e+09, 8.672412e+09, 8.779684e+09, 8.885187e+09, 
    8.988781e+09, 9.090322e+09, 9.18967e+09, 9.286681e+09, 9.381209e+09, 
    9.473112e+09, 9.562249e+09, 9.648477e+09, 9.731658e+09, 9.811654e+09, 
    9.88833e+09, 9.961556e+09, 1.00312e+10, 1.009715e+10, 1.015928e+10, 
    1.021748e+10, 1.027164e+10, 1.032166e+10, 1.036744e+10, 1.040891e+10, 
    1.044597e+10, 1.047856e+10, 1.050662e+10, 1.053008e+10, 1.054891e+10, 
    1.056306e+10, 1.057252e+10, 1.057725e+10, 1.057725e+10, 1.057252e+10, 
    1.056306e+10, 1.054891e+10, 1.053008e+10, 1.050662e+10, 1.047856e+10, 
    1.044597e+10, 1.040891e+10, 1.036744e+10, 1.032166e+10, 1.027164e+10, 
    1.021748e+10, 1.015928e+10, 1.009715e+10, 1.00312e+10, 9.961556e+09, 
    9.88833e+09, 9.811654e+09, 9.731658e+09, 9.648477e+09, 9.562249e+09, 
    9.473112e+09, 9.381209e+09, 9.286681e+09, 9.18967e+09, 9.090322e+09, 
    8.988781e+09, 8.885187e+09, 8.779684e+09, 8.672412e+09, 8.563511e+09, 
    8.453116e+09, 8.341364e+09, 8.228386e+09, 8.11431e+09, 7.999264e+09, 
    7.883369e+09, 7.766745e+09, 7.649507e+09, 7.531766e+09, 7.41363e+09, 
    7.295202e+09, 7.176583e+09, 7.057866e+09, 6.939143e+09, 6.8205e+09, 
    6.702019e+09,
  6.668692e+09, 6.784244e+09, 6.899874e+09, 7.015503e+09, 7.131045e+09, 
    7.246414e+09, 7.361518e+09, 7.47626e+09, 7.590542e+09, 7.704261e+09, 
    7.817309e+09, 7.929576e+09, 8.04095e+09, 8.151313e+09, 8.260545e+09, 
    8.368525e+09, 8.475127e+09, 8.580225e+09, 8.683688e+09, 8.785385e+09, 
    8.885187e+09, 8.982957e+09, 9.078562e+09, 9.171869e+09, 9.262742e+09, 
    9.351046e+09, 9.436652e+09, 9.519426e+09, 9.599237e+09, 9.67596e+09, 
    9.749469e+09, 9.819643e+09, 9.886363e+09, 9.949515e+09, 1.000899e+10, 
    1.006469e+10, 1.01165e+10, 1.016434e+10, 1.020812e+10, 1.024776e+10, 
    1.028319e+10, 1.031433e+10, 1.034114e+10, 1.036355e+10, 1.038154e+10, 
    1.039506e+10, 1.040409e+10, 1.040861e+10, 1.040861e+10, 1.040409e+10, 
    1.039506e+10, 1.038154e+10, 1.036355e+10, 1.034114e+10, 1.031433e+10, 
    1.028319e+10, 1.024776e+10, 1.020812e+10, 1.016434e+10, 1.01165e+10, 
    1.006469e+10, 1.000899e+10, 9.949515e+09, 9.886363e+09, 9.819643e+09, 
    9.749469e+09, 9.67596e+09, 9.599237e+09, 9.519426e+09, 9.436652e+09, 
    9.351046e+09, 9.262742e+09, 9.171869e+09, 9.078562e+09, 8.982957e+09, 
    8.885187e+09, 8.785385e+09, 8.683688e+09, 8.580225e+09, 8.475127e+09, 
    8.368525e+09, 8.260545e+09, 8.151313e+09, 8.04095e+09, 7.929576e+09, 
    7.817309e+09, 7.704261e+09, 7.590542e+09, 7.47626e+09, 7.361518e+09, 
    7.246414e+09, 7.131045e+09, 7.015503e+09, 6.899874e+09, 6.784244e+09, 
    6.668692e+09,
  6.634248e+09, 6.74681e+09, 6.859367e+09, 6.971842e+09, 7.084154e+09, 
    7.196217e+09, 7.307944e+09, 7.419243e+09, 7.530018e+09, 7.640172e+09, 
    7.749601e+09, 7.858201e+09, 7.965864e+09, 8.072481e+09, 8.177936e+09, 
    8.282116e+09, 8.384902e+09, 8.486173e+09, 8.585809e+09, 8.683688e+09, 
    8.779684e+09, 8.873673e+09, 8.96553e+09, 9.055129e+09, 9.142345e+09, 
    9.227054e+09, 9.309132e+09, 9.388457e+09, 9.464909e+09, 9.53837e+09, 
    9.608722e+09, 9.675857e+09, 9.739662e+09, 9.800034e+09, 9.856871e+09, 
    9.910078e+09, 9.959563e+09, 1.000524e+10, 1.004703e+10, 1.008486e+10, 
    1.011866e+10, 1.014837e+10, 1.017394e+10, 1.019532e+10, 1.021247e+10, 
    1.022536e+10, 1.023397e+10, 1.023827e+10, 1.023827e+10, 1.023397e+10, 
    1.022536e+10, 1.021247e+10, 1.019532e+10, 1.017394e+10, 1.014837e+10, 
    1.011866e+10, 1.008486e+10, 1.004703e+10, 1.000524e+10, 9.959563e+09, 
    9.910078e+09, 9.856871e+09, 9.800034e+09, 9.739662e+09, 9.675857e+09, 
    9.608722e+09, 9.53837e+09, 9.464909e+09, 9.388457e+09, 9.309132e+09, 
    9.227054e+09, 9.142345e+09, 9.055129e+09, 8.96553e+09, 8.873673e+09, 
    8.779684e+09, 8.683688e+09, 8.585809e+09, 8.486173e+09, 8.384902e+09, 
    8.282116e+09, 8.177936e+09, 8.072481e+09, 7.965864e+09, 7.858201e+09, 
    7.749601e+09, 7.640172e+09, 7.530018e+09, 7.419243e+09, 7.307944e+09, 
    7.196217e+09, 7.084154e+09, 6.971842e+09, 6.859367e+09, 6.74681e+09, 
    6.634248e+09,
  6.598693e+09, 6.708208e+09, 6.817636e+09, 6.926904e+09, 7.035934e+09, 
    7.144643e+09, 7.252946e+09, 7.360757e+09, 7.467984e+09, 7.574533e+09, 
    7.680307e+09, 7.785207e+09, 7.889131e+09, 7.991974e+09, 8.093629e+09, 
    8.193989e+09, 8.292941e+09, 8.390374e+09, 8.486173e+09, 8.580225e+09, 
    8.672412e+09, 8.762619e+09, 8.85073e+09, 8.936627e+09, 9.020195e+09, 
    9.101317e+09, 9.17988e+09, 9.255772e+09, 9.32888e+09, 9.399095e+09, 
    9.466312e+09, 9.530426e+09, 9.591338e+09, 9.64895e+09, 9.703171e+09, 
    9.753911e+09, 9.801088e+09, 9.844622e+09, 9.884442e+09, 9.920478e+09, 
    9.95267e+09, 9.980962e+09, 1.00053e+10, 1.002566e+10, 1.004198e+10, 
    1.005425e+10, 1.006244e+10, 1.006654e+10, 1.006654e+10, 1.006244e+10, 
    1.005425e+10, 1.004198e+10, 1.002566e+10, 1.00053e+10, 9.980962e+09, 
    9.95267e+09, 9.920478e+09, 9.884442e+09, 9.844622e+09, 9.801088e+09, 
    9.753911e+09, 9.703171e+09, 9.64895e+09, 9.591338e+09, 9.530426e+09, 
    9.466312e+09, 9.399095e+09, 9.32888e+09, 9.255772e+09, 9.17988e+09, 
    9.101317e+09, 9.020195e+09, 8.936627e+09, 8.85073e+09, 8.762619e+09, 
    8.672412e+09, 8.580225e+09, 8.486173e+09, 8.390374e+09, 8.292941e+09, 
    8.193989e+09, 8.093629e+09, 7.991974e+09, 7.889131e+09, 7.785207e+09, 
    7.680307e+09, 7.574533e+09, 7.467984e+09, 7.360757e+09, 7.252946e+09, 
    7.144643e+09, 7.035934e+09, 6.926904e+09, 6.817636e+09, 6.708208e+09, 
    6.598693e+09,
  6.562035e+09, 6.668449e+09, 6.774699e+09, 6.880711e+09, 6.986412e+09, 
    7.091722e+09, 7.196561e+09, 7.300845e+09, 7.404488e+09, 7.5074e+09, 
    7.60949e+09, 7.710664e+09, 7.810825e+09, 7.909876e+09, 8.007716e+09, 
    8.104243e+09, 8.199353e+09, 8.292941e+09, 8.384902e+09, 8.475127e+09, 
    8.563511e+09, 8.649944e+09, 8.734319e+09, 8.816526e+09, 8.896461e+09, 
    8.974015e+09, 9.049084e+09, 9.121564e+09, 9.191351e+09, 9.258346e+09, 
    9.322452e+09, 9.383574e+09, 9.441618e+09, 9.496498e+09, 9.548129e+09, 
    9.596429e+09, 9.641325e+09, 9.68274e+09, 9.720613e+09, 9.754878e+09, 
    9.785482e+09, 9.812372e+09, 9.835507e+09, 9.854844e+09, 9.870353e+09, 
    9.882009e+09, 9.88979e+09, 9.893683e+09, 9.893683e+09, 9.88979e+09, 
    9.882009e+09, 9.870353e+09, 9.854844e+09, 9.835507e+09, 9.812372e+09, 
    9.785482e+09, 9.754878e+09, 9.720613e+09, 9.68274e+09, 9.641325e+09, 
    9.596429e+09, 9.548129e+09, 9.496498e+09, 9.441618e+09, 9.383574e+09, 
    9.322452e+09, 9.258346e+09, 9.191351e+09, 9.121564e+09, 9.049084e+09, 
    8.974015e+09, 8.896461e+09, 8.816526e+09, 8.734319e+09, 8.649944e+09, 
    8.563511e+09, 8.475127e+09, 8.384902e+09, 8.292941e+09, 8.199353e+09, 
    8.104243e+09, 8.007716e+09, 7.909876e+09, 7.810825e+09, 7.710664e+09, 
    7.60949e+09, 7.5074e+09, 7.404488e+09, 7.300845e+09, 7.196561e+09, 
    7.091722e+09, 6.986412e+09, 6.880711e+09, 6.774699e+09, 6.668449e+09, 
    6.562035e+09,
  6.524282e+09, 6.627547e+09, 6.730571e+09, 6.833284e+09, 6.935614e+09, 
    7.037487e+09, 7.138825e+09, 7.23955e+09, 7.339579e+09, 7.438829e+09, 
    7.537212e+09, 7.634641e+09, 7.731025e+09, 7.826271e+09, 7.920287e+09, 
    8.012976e+09, 8.104243e+09, 8.193989e+09, 8.282116e+09, 8.368525e+09, 
    8.453116e+09, 8.53579e+09, 8.616447e+09, 8.694987e+09, 8.771312e+09, 
    8.845323e+09, 8.916924e+09, 8.986021e+09, 9.052518e+09, 9.116325e+09, 
    9.177352e+09, 9.235513e+09, 9.290724e+09, 9.342905e+09, 9.391978e+09, 
    9.437871e+09, 9.480515e+09, 9.519842e+09, 9.555794e+09, 9.588315e+09, 
    9.617354e+09, 9.642865e+09, 9.664807e+09, 9.683147e+09, 9.697854e+09, 
    9.708905e+09, 9.716282e+09, 9.719975e+09, 9.719975e+09, 9.716282e+09, 
    9.708905e+09, 9.697854e+09, 9.683147e+09, 9.664807e+09, 9.642865e+09, 
    9.617354e+09, 9.588315e+09, 9.555794e+09, 9.519842e+09, 9.480515e+09, 
    9.437871e+09, 9.391978e+09, 9.342905e+09, 9.290724e+09, 9.235513e+09, 
    9.177352e+09, 9.116325e+09, 9.052518e+09, 8.986021e+09, 8.916924e+09, 
    8.845323e+09, 8.771312e+09, 8.694987e+09, 8.616447e+09, 8.53579e+09, 
    8.453116e+09, 8.368525e+09, 8.282116e+09, 8.193989e+09, 8.104243e+09, 
    8.012976e+09, 7.920287e+09, 7.826271e+09, 7.731025e+09, 7.634641e+09, 
    7.537212e+09, 7.438829e+09, 7.339579e+09, 7.23955e+09, 7.138825e+09, 
    7.037487e+09, 6.935614e+09, 6.833284e+09, 6.730571e+09, 6.627547e+09, 
    6.524282e+09,
  6.485442e+09, 6.585513e+09, 6.685269e+09, 6.784643e+09, 6.883567e+09, 
    6.981969e+09, 7.079777e+09, 7.176916e+09, 7.273309e+09, 7.368877e+09, 
    7.463537e+09, 7.557208e+09, 7.649805e+09, 7.741242e+09, 7.831433e+09, 
    7.920287e+09, 8.007716e+09, 8.093629e+09, 8.177936e+09, 8.260545e+09, 
    8.341364e+09, 8.420301e+09, 8.497266e+09, 8.572165e+09, 8.64491e+09, 
    8.715411e+09, 8.78358e+09, 8.849328e+09, 8.912572e+09, 8.973229e+09, 
    9.031216e+09, 9.086456e+09, 9.138871e+09, 9.188391e+09, 9.234944e+09, 
    9.278465e+09, 9.318892e+09, 9.356163e+09, 9.390226e+09, 9.421031e+09, 
    9.448532e+09, 9.472687e+09, 9.49346e+09, 9.510819e+09, 9.524738e+09, 
    9.535196e+09, 9.542177e+09, 9.54567e+09, 9.54567e+09, 9.542177e+09, 
    9.535196e+09, 9.524738e+09, 9.510819e+09, 9.49346e+09, 9.472687e+09, 
    9.448532e+09, 9.421031e+09, 9.390226e+09, 9.356163e+09, 9.318892e+09, 
    9.278465e+09, 9.234944e+09, 9.188391e+09, 9.138871e+09, 9.086456e+09, 
    9.031216e+09, 8.973229e+09, 8.912572e+09, 8.849328e+09, 8.78358e+09, 
    8.715411e+09, 8.64491e+09, 8.572165e+09, 8.497266e+09, 8.420301e+09, 
    8.341364e+09, 8.260545e+09, 8.177936e+09, 8.093629e+09, 8.007716e+09, 
    7.920287e+09, 7.831433e+09, 7.741242e+09, 7.649805e+09, 7.557208e+09, 
    7.463537e+09, 7.368877e+09, 7.273309e+09, 7.176916e+09, 7.079777e+09, 
    6.981969e+09, 6.883567e+09, 6.784643e+09, 6.685269e+09, 6.585513e+09, 
    6.485442e+09,
  6.445522e+09, 6.54236e+09, 6.638811e+09, 6.734811e+09, 6.830297e+09, 
    6.925201e+09, 7.019455e+09, 7.112987e+09, 7.205726e+09, 7.297597e+09, 
    7.388526e+09, 7.478433e+09, 7.567242e+09, 7.654872e+09, 7.741242e+09, 
    7.826271e+09, 7.909876e+09, 7.991974e+09, 8.072481e+09, 8.151313e+09, 
    8.228386e+09, 8.303616e+09, 8.37692e+09, 8.448214e+09, 8.517416e+09, 
    8.584445e+09, 8.649221e+09, 8.711665e+09, 8.771699e+09, 8.829247e+09, 
    8.884238e+09, 8.936601e+09, 8.986266e+09, 9.033167e+09, 9.077242e+09, 
    9.118431e+09, 9.156679e+09, 9.191932e+09, 9.224142e+09, 9.253263e+09, 
    9.279254e+09, 9.302078e+09, 9.321703e+09, 9.338102e+09, 9.351248e+09, 
    9.361125e+09, 9.367718e+09, 9.371016e+09, 9.371016e+09, 9.367718e+09, 
    9.361125e+09, 9.351248e+09, 9.338102e+09, 9.321703e+09, 9.302078e+09, 
    9.279254e+09, 9.253263e+09, 9.224142e+09, 9.191932e+09, 9.156679e+09, 
    9.118431e+09, 9.077242e+09, 9.033167e+09, 8.986266e+09, 8.936601e+09, 
    8.884238e+09, 8.829247e+09, 8.771699e+09, 8.711665e+09, 8.649221e+09, 
    8.584445e+09, 8.517416e+09, 8.448214e+09, 8.37692e+09, 8.303616e+09, 
    8.228386e+09, 8.151313e+09, 8.072481e+09, 7.991974e+09, 7.909876e+09, 
    7.826271e+09, 7.741242e+09, 7.654872e+09, 7.567242e+09, 7.478433e+09, 
    7.388526e+09, 7.297597e+09, 7.205726e+09, 7.112987e+09, 7.019455e+09, 
    6.925201e+09, 6.830297e+09, 6.734811e+09, 6.638811e+09, 6.54236e+09, 
    6.445522e+09,
  6.404531e+09, 6.4981e+09, 6.591213e+09, 6.683811e+09, 6.775833e+09, 
    6.867216e+09, 6.957896e+09, 7.047806e+09, 7.136881e+09, 7.225049e+09, 
    7.312241e+09, 7.398386e+09, 7.483411e+09, 7.567242e+09, 7.649805e+09, 
    7.731025e+09, 7.810825e+09, 7.889131e+09, 7.965864e+09, 8.04095e+09, 
    8.11431e+09, 8.18587e+09, 8.255552e+09, 8.323282e+09, 8.388985e+09, 
    8.452588e+09, 8.514017e+09, 8.573202e+09, 8.630074e+09, 8.684566e+09, 
    8.736609e+09, 8.786142e+09, 8.833104e+09, 8.877434e+09, 8.919077e+09, 
    8.95798e+09, 8.994092e+09, 9.027367e+09, 9.05776e+09, 9.085231e+09, 
    9.109745e+09, 9.131267e+09, 9.14977e+09, 9.165227e+09, 9.177618e+09, 
    9.186927e+09, 9.193139e+09, 9.196247e+09, 9.196247e+09, 9.193139e+09, 
    9.186927e+09, 9.177618e+09, 9.165227e+09, 9.14977e+09, 9.131267e+09, 
    9.109745e+09, 9.085231e+09, 9.05776e+09, 9.027367e+09, 8.994092e+09, 
    8.95798e+09, 8.919077e+09, 8.877434e+09, 8.833104e+09, 8.786142e+09, 
    8.736609e+09, 8.684566e+09, 8.630074e+09, 8.573202e+09, 8.514017e+09, 
    8.452588e+09, 8.388985e+09, 8.323282e+09, 8.255552e+09, 8.18587e+09, 
    8.11431e+09, 8.04095e+09, 7.965864e+09, 7.889131e+09, 7.810825e+09, 
    7.731025e+09, 7.649805e+09, 7.567242e+09, 7.483411e+09, 7.398386e+09, 
    7.312241e+09, 7.225049e+09, 7.136881e+09, 7.047806e+09, 6.957896e+09, 
    6.867216e+09, 6.775833e+09, 6.683811e+09, 6.591213e+09, 6.4981e+09, 
    6.404531e+09,
  6.362479e+09, 6.452746e+09, 6.542493e+09, 6.631664e+09, 6.720201e+09, 
    6.808046e+09, 6.895139e+09, 6.981418e+09, 7.066822e+09, 7.151286e+09, 
    7.234745e+09, 7.317134e+09, 7.398386e+09, 7.478433e+09, 7.557208e+09, 
    7.634641e+09, 7.710664e+09, 7.785207e+09, 7.858201e+09, 7.929576e+09, 
    7.999264e+09, 8.067195e+09, 8.133301e+09, 8.197513e+09, 8.259766e+09, 
    8.319992e+09, 8.378128e+09, 8.434108e+09, 8.487873e+09, 8.539359e+09, 
    8.58851e+09, 8.635267e+09, 8.679578e+09, 8.721389e+09, 8.760649e+09, 
    8.797313e+09, 8.831335e+09, 8.862674e+09, 8.891291e+09, 8.917151e+09, 
    8.940219e+09, 8.96047e+09, 8.977876e+09, 8.992415e+09, 9.004068e+09, 
    9.012821e+09, 9.018663e+09, 9.021585e+09, 9.021585e+09, 9.018663e+09, 
    9.012821e+09, 9.004068e+09, 8.992415e+09, 8.977876e+09, 8.96047e+09, 
    8.940219e+09, 8.917151e+09, 8.891291e+09, 8.862674e+09, 8.831335e+09, 
    8.797313e+09, 8.760649e+09, 8.721389e+09, 8.679578e+09, 8.635267e+09, 
    8.58851e+09, 8.539359e+09, 8.487873e+09, 8.434108e+09, 8.378128e+09, 
    8.319992e+09, 8.259766e+09, 8.197513e+09, 8.133301e+09, 8.067195e+09, 
    7.999264e+09, 7.929576e+09, 7.858201e+09, 7.785207e+09, 7.710664e+09, 
    7.634641e+09, 7.557208e+09, 7.478433e+09, 7.398386e+09, 7.317134e+09, 
    7.234745e+09, 7.151286e+09, 7.066822e+09, 6.981418e+09, 6.895139e+09, 
    6.808046e+09, 6.720201e+09, 6.631664e+09, 6.542493e+09, 6.452746e+09, 
    6.362479e+09,
  6.319373e+09, 6.406312e+09, 6.492669e+09, 6.578392e+09, 6.663429e+09, 
    6.747724e+09, 6.831222e+09, 6.913867e+09, 6.9956e+09, 7.076365e+09, 
    7.1561e+09, 7.234745e+09, 7.312241e+09, 7.388526e+09, 7.463537e+09, 
    7.537212e+09, 7.60949e+09, 7.680307e+09, 7.749601e+09, 7.817309e+09, 
    7.883369e+09, 7.94772e+09, 8.010299e+09, 8.071048e+09, 8.129904e+09, 
    8.186811e+09, 8.241709e+09, 8.294543e+09, 8.345257e+09, 8.393798e+09, 
    8.440113e+09, 8.484152e+09, 8.525868e+09, 8.565214e+09, 8.602145e+09, 
    8.636621e+09, 8.668601e+09, 8.698051e+09, 8.724934e+09, 8.749221e+09, 
    8.770882e+09, 8.789891e+09, 8.806228e+09, 8.819871e+09, 8.830806e+09, 
    8.839017e+09, 8.844498e+09, 8.84724e+09, 8.84724e+09, 8.844498e+09, 
    8.839017e+09, 8.830806e+09, 8.819871e+09, 8.806228e+09, 8.789891e+09, 
    8.770882e+09, 8.749221e+09, 8.724934e+09, 8.698051e+09, 8.668601e+09, 
    8.636621e+09, 8.602145e+09, 8.565214e+09, 8.525868e+09, 8.484152e+09, 
    8.440113e+09, 8.393798e+09, 8.345257e+09, 8.294543e+09, 8.241709e+09, 
    8.186811e+09, 8.129904e+09, 8.071048e+09, 8.010299e+09, 7.94772e+09, 
    7.883369e+09, 7.817309e+09, 7.749601e+09, 7.680307e+09, 7.60949e+09, 
    7.537212e+09, 7.463537e+09, 7.388526e+09, 7.312241e+09, 7.234745e+09, 
    7.1561e+09, 7.076365e+09, 6.9956e+09, 6.913867e+09, 6.831222e+09, 
    6.747724e+09, 6.663429e+09, 6.578392e+09, 6.492669e+09, 6.406312e+09, 
    6.319373e+09,
  6.275223e+09, 6.35881e+09, 6.441759e+09, 6.52402e+09, 6.605544e+09, 
    6.686283e+09, 6.766183e+09, 6.845195e+09, 6.923265e+09, 7.000339e+09, 
    7.076365e+09, 7.151286e+09, 7.225049e+09, 7.297597e+09, 7.368877e+09, 
    7.438829e+09, 7.5074e+09, 7.574533e+09, 7.640172e+09, 7.704261e+09, 
    7.766745e+09, 7.827569e+09, 7.886679e+09, 7.94402e+09, 7.99954e+09, 
    8.053188e+09, 8.10491e+09, 8.15466e+09, 8.202386e+09, 8.248043e+09, 
    8.291585e+09, 8.332967e+09, 8.372148e+09, 8.409087e+09, 8.443745e+09, 
    8.476086e+09, 8.506077e+09, 8.533684e+09, 8.558878e+09, 8.581632e+09, 
    8.601922e+09, 8.619724e+09, 8.63502e+09, 8.647793e+09, 8.658028e+09, 
    8.665715e+09, 8.670843e+09, 8.673409e+09, 8.673409e+09, 8.670843e+09, 
    8.665715e+09, 8.658028e+09, 8.647793e+09, 8.63502e+09, 8.619724e+09, 
    8.601922e+09, 8.581632e+09, 8.558878e+09, 8.533684e+09, 8.506077e+09, 
    8.476086e+09, 8.443745e+09, 8.409087e+09, 8.372148e+09, 8.332967e+09, 
    8.291585e+09, 8.248043e+09, 8.202386e+09, 8.15466e+09, 8.10491e+09, 
    8.053188e+09, 7.99954e+09, 7.94402e+09, 7.886679e+09, 7.827569e+09, 
    7.766745e+09, 7.704261e+09, 7.640172e+09, 7.574533e+09, 7.5074e+09, 
    7.438829e+09, 7.368877e+09, 7.297597e+09, 7.225049e+09, 7.151286e+09, 
    7.076365e+09, 7.000339e+09, 6.923265e+09, 6.845195e+09, 6.766183e+09, 
    6.686283e+09, 6.605544e+09, 6.52402e+09, 6.441759e+09, 6.35881e+09, 
    6.275223e+09,
  6.230037e+09, 6.310255e+09, 6.38978e+09, 6.468569e+09, 6.546576e+09, 
    6.623755e+09, 6.700061e+09, 6.775447e+09, 6.849864e+09, 6.923265e+09, 
    6.9956e+09, 7.066822e+09, 7.136881e+09, 7.205726e+09, 7.273309e+09, 
    7.339579e+09, 7.404488e+09, 7.467984e+09, 7.530018e+09, 7.590542e+09, 
    7.649507e+09, 7.706863e+09, 7.762563e+09, 7.816561e+09, 7.868808e+09, 
    7.919261e+09, 7.967875e+09, 8.014606e+09, 8.059411e+09, 8.10225e+09, 
    8.143084e+09, 8.181873e+09, 8.218582e+09, 8.253174e+09, 8.285618e+09, 
    8.31588e+09, 8.343933e+09, 8.369748e+09, 8.3933e+09, 8.414565e+09, 
    8.433522e+09, 8.450151e+09, 8.464436e+09, 8.476363e+09, 8.485919e+09, 
    8.493095e+09, 8.497883e+09, 8.500278e+09, 8.500278e+09, 8.497883e+09, 
    8.493095e+09, 8.485919e+09, 8.476363e+09, 8.464436e+09, 8.450151e+09, 
    8.433522e+09, 8.414565e+09, 8.3933e+09, 8.369748e+09, 8.343933e+09, 
    8.31588e+09, 8.285618e+09, 8.253174e+09, 8.218582e+09, 8.181873e+09, 
    8.143084e+09, 8.10225e+09, 8.059411e+09, 8.014606e+09, 7.967875e+09, 
    7.919261e+09, 7.868808e+09, 7.816561e+09, 7.762563e+09, 7.706863e+09, 
    7.649507e+09, 7.590542e+09, 7.530018e+09, 7.467984e+09, 7.404488e+09, 
    7.339579e+09, 7.273309e+09, 7.205726e+09, 7.136881e+09, 7.066822e+09, 
    6.9956e+09, 6.923265e+09, 6.849864e+09, 6.775447e+09, 6.700061e+09, 
    6.623755e+09, 6.546576e+09, 6.468569e+09, 6.38978e+09, 6.310255e+09, 
    6.230037e+09,
  6.183825e+09, 6.260659e+09, 6.336752e+09, 6.412062e+09, 6.486551e+09, 
    6.560175e+09, 6.632894e+09, 6.704666e+09, 6.775447e+09, 6.845195e+09, 
    6.913867e+09, 6.981418e+09, 7.047806e+09, 7.112987e+09, 7.176916e+09, 
    7.23955e+09, 7.300845e+09, 7.360757e+09, 7.419243e+09, 7.47626e+09, 
    7.531766e+09, 7.585717e+09, 7.638074e+09, 7.688794e+09, 7.737838e+09, 
    7.785166e+09, 7.830739e+09, 7.874522e+09, 7.916475e+09, 7.956566e+09, 
    7.994759e+09, 8.031022e+09, 8.065324e+09, 8.097633e+09, 8.127923e+09, 
    8.156166e+09, 8.182336e+09, 8.20641e+09, 8.228367e+09, 8.248187e+09, 
    8.26585e+09, 8.281342e+09, 8.294647e+09, 8.305754e+09, 8.314652e+09, 
    8.321333e+09, 8.32579e+09, 8.32802e+09, 8.32802e+09, 8.32579e+09, 
    8.321333e+09, 8.314652e+09, 8.305754e+09, 8.294647e+09, 8.281342e+09, 
    8.26585e+09, 8.248187e+09, 8.228367e+09, 8.20641e+09, 8.182336e+09, 
    8.156166e+09, 8.127923e+09, 8.097633e+09, 8.065324e+09, 8.031022e+09, 
    7.994759e+09, 7.956566e+09, 7.916475e+09, 7.874522e+09, 7.830739e+09, 
    7.785166e+09, 7.737838e+09, 7.688794e+09, 7.638074e+09, 7.585717e+09, 
    7.531766e+09, 7.47626e+09, 7.419243e+09, 7.360757e+09, 7.300845e+09, 
    7.23955e+09, 7.176916e+09, 7.112987e+09, 7.047806e+09, 6.981418e+09, 
    6.913867e+09, 6.845195e+09, 6.775447e+09, 6.704666e+09, 6.632894e+09, 
    6.560175e+09, 6.486551e+09, 6.412062e+09, 6.336752e+09, 6.260659e+09, 
    6.183825e+09,
  6.136596e+09, 6.210038e+09, 6.282692e+09, 6.354524e+09, 6.425497e+09, 
    6.495574e+09, 6.564719e+09, 6.632894e+09, 6.700061e+09, 6.766183e+09, 
    6.831222e+09, 6.895139e+09, 6.957896e+09, 7.019455e+09, 7.079777e+09, 
    7.138825e+09, 7.196561e+09, 7.252946e+09, 7.307944e+09, 7.361518e+09, 
    7.41363e+09, 7.464245e+09, 7.513327e+09, 7.56084e+09, 7.606751e+09, 
    7.651027e+09, 7.693634e+09, 7.734541e+09, 7.773715e+09, 7.811129e+09, 
    7.846753e+09, 7.880559e+09, 7.912521e+09, 7.942612e+09, 7.970811e+09, 
    7.997093e+09, 8.021437e+09, 8.043825e+09, 8.064236e+09, 8.082655e+09, 
    8.099066e+09, 8.113456e+09, 8.125813e+09, 8.136126e+09, 8.144387e+09, 
    8.150589e+09, 8.154726e+09, 8.156796e+09, 8.156796e+09, 8.154726e+09, 
    8.150589e+09, 8.144387e+09, 8.136126e+09, 8.125813e+09, 8.113456e+09, 
    8.099066e+09, 8.082655e+09, 8.064236e+09, 8.043825e+09, 8.021437e+09, 
    7.997093e+09, 7.970811e+09, 7.942612e+09, 7.912521e+09, 7.880559e+09, 
    7.846753e+09, 7.811129e+09, 7.773715e+09, 7.734541e+09, 7.693634e+09, 
    7.651027e+09, 7.606751e+09, 7.56084e+09, 7.513327e+09, 7.464245e+09, 
    7.41363e+09, 7.361518e+09, 7.307944e+09, 7.252946e+09, 7.196561e+09, 
    7.138825e+09, 7.079777e+09, 7.019455e+09, 6.957896e+09, 6.895139e+09, 
    6.831222e+09, 6.766183e+09, 6.700061e+09, 6.632894e+09, 6.564719e+09, 
    6.495574e+09, 6.425497e+09, 6.354524e+09, 6.282692e+09, 6.210038e+09, 
    6.136596e+09,
  6.088361e+09, 6.158404e+09, 6.227619e+09, 6.295976e+09, 6.363442e+09, 
    6.429985e+09, 6.495574e+09, 6.560175e+09, 6.623755e+09, 6.686283e+09, 
    6.747724e+09, 6.808046e+09, 6.867216e+09, 6.925201e+09, 6.981969e+09, 
    7.037487e+09, 7.091722e+09, 7.144643e+09, 7.196217e+09, 7.246414e+09, 
    7.295202e+09, 7.342552e+09, 7.388432e+09, 7.432814e+09, 7.475667e+09, 
    7.516966e+09, 7.556683e+09, 7.594789e+09, 7.631261e+09, 7.666072e+09, 
    7.699199e+09, 7.73062e+09, 7.760311e+09, 7.788252e+09, 7.814423e+09, 
    7.838806e+09, 7.861382e+09, 7.882135e+09, 7.901051e+09, 7.918115e+09, 
    7.933316e+09, 7.946641e+09, 7.958081e+09, 7.967627e+09, 7.975273e+09, 
    7.981012e+09, 7.984841e+09, 7.986756e+09, 7.986756e+09, 7.984841e+09, 
    7.981012e+09, 7.975273e+09, 7.967627e+09, 7.958081e+09, 7.946641e+09, 
    7.933316e+09, 7.918115e+09, 7.901051e+09, 7.882135e+09, 7.861382e+09, 
    7.838806e+09, 7.814423e+09, 7.788252e+09, 7.760311e+09, 7.73062e+09, 
    7.699199e+09, 7.666072e+09, 7.631261e+09, 7.594789e+09, 7.556683e+09, 
    7.516966e+09, 7.475667e+09, 7.432814e+09, 7.388432e+09, 7.342552e+09, 
    7.295202e+09, 7.246414e+09, 7.196217e+09, 7.144643e+09, 7.091722e+09, 
    7.037487e+09, 6.981969e+09, 6.925201e+09, 6.867216e+09, 6.808046e+09, 
    6.747724e+09, 6.686283e+09, 6.623755e+09, 6.560175e+09, 6.495574e+09, 
    6.429985e+09, 6.363442e+09, 6.295976e+09, 6.227619e+09, 6.158404e+09, 
    6.088361e+09,
  6.039129e+09, 6.105772e+09, 6.171552e+09, 6.236442e+09, 6.300414e+09, 
    6.363442e+09, 6.425497e+09, 6.486551e+09, 6.546576e+09, 6.605544e+09, 
    6.663429e+09, 6.720201e+09, 6.775833e+09, 6.830297e+09, 6.883567e+09, 
    6.935614e+09, 6.986412e+09, 7.035934e+09, 7.084154e+09, 7.131045e+09, 
    7.176583e+09, 7.220742e+09, 7.263496e+09, 7.304823e+09, 7.344698e+09, 
    7.383099e+09, 7.420003e+09, 7.455388e+09, 7.489233e+09, 7.521518e+09, 
    7.552224e+09, 7.581331e+09, 7.608822e+09, 7.634681e+09, 7.65889e+09, 
    7.681435e+09, 7.702302e+09, 7.721477e+09, 7.738948e+09, 7.754704e+09, 
    7.768736e+09, 7.781033e+09, 7.791588e+09, 7.800395e+09, 7.807448e+09, 
    7.812741e+09, 7.816271e+09, 7.818037e+09, 7.818037e+09, 7.816271e+09, 
    7.812741e+09, 7.807448e+09, 7.800395e+09, 7.791588e+09, 7.781033e+09, 
    7.768736e+09, 7.754704e+09, 7.738948e+09, 7.721477e+09, 7.702302e+09, 
    7.681435e+09, 7.65889e+09, 7.634681e+09, 7.608822e+09, 7.581331e+09, 
    7.552224e+09, 7.521518e+09, 7.489233e+09, 7.455388e+09, 7.420003e+09, 
    7.383099e+09, 7.344698e+09, 7.304823e+09, 7.263496e+09, 7.220742e+09, 
    7.176583e+09, 7.131045e+09, 7.084154e+09, 7.035934e+09, 6.986412e+09, 
    6.935614e+09, 6.883567e+09, 6.830297e+09, 6.775833e+09, 6.720201e+09, 
    6.663429e+09, 6.605544e+09, 6.546576e+09, 6.486551e+09, 6.425497e+09, 
    6.363442e+09, 6.300414e+09, 6.236442e+09, 6.171552e+09, 6.105772e+09, 
    6.039129e+09,
  5.988909e+09, 6.052155e+09, 6.114508e+09, 6.175945e+09, 6.236442e+09, 
    6.295976e+09, 6.354524e+09, 6.412062e+09, 6.468569e+09, 6.52402e+09, 
    6.578392e+09, 6.631664e+09, 6.683811e+09, 6.734811e+09, 6.784643e+09, 
    6.833284e+09, 6.880711e+09, 6.926904e+09, 6.971842e+09, 7.015503e+09, 
    7.057866e+09, 7.098912e+09, 7.13862e+09, 7.176973e+09, 7.21395e+09, 
    7.249533e+09, 7.283705e+09, 7.316448e+09, 7.347746e+09, 7.377583e+09, 
    7.405943e+09, 7.432813e+09, 7.458176e+09, 7.482021e+09, 7.504335e+09, 
    7.525106e+09, 7.544322e+09, 7.561974e+09, 7.578052e+09, 7.592547e+09, 
    7.605452e+09, 7.616759e+09, 7.626462e+09, 7.634556e+09, 7.641037e+09, 
    7.645901e+09, 7.649145e+09, 7.650767e+09, 7.650767e+09, 7.649145e+09, 
    7.645901e+09, 7.641037e+09, 7.634556e+09, 7.626462e+09, 7.616759e+09, 
    7.605452e+09, 7.592547e+09, 7.578052e+09, 7.561974e+09, 7.544322e+09, 
    7.525106e+09, 7.504335e+09, 7.482021e+09, 7.458176e+09, 7.432813e+09, 
    7.405943e+09, 7.377583e+09, 7.347746e+09, 7.316448e+09, 7.283705e+09, 
    7.249533e+09, 7.21395e+09, 7.176973e+09, 7.13862e+09, 7.098912e+09, 
    7.057866e+09, 7.015503e+09, 6.971842e+09, 6.926904e+09, 6.880711e+09, 
    6.833284e+09, 6.784643e+09, 6.734811e+09, 6.683811e+09, 6.631664e+09, 
    6.578392e+09, 6.52402e+09, 6.468569e+09, 6.412062e+09, 6.354524e+09, 
    6.295976e+09, 6.236442e+09, 6.175945e+09, 6.114508e+09, 6.052155e+09, 
    5.988909e+09,
  5.937712e+09, 5.99757e+09, 6.056508e+09, 6.114508e+09, 6.171552e+09, 
    6.227619e+09, 6.282692e+09, 6.336752e+09, 6.38978e+09, 6.441759e+09, 
    6.492669e+09, 6.542493e+09, 6.591213e+09, 6.638811e+09, 6.685269e+09, 
    6.730571e+09, 6.774699e+09, 6.817636e+09, 6.859367e+09, 6.899874e+09, 
    6.939143e+09, 6.977157e+09, 7.013901e+09, 7.049361e+09, 7.083523e+09, 
    7.116371e+09, 7.147894e+09, 7.178077e+09, 7.206909e+09, 7.234377e+09, 
    7.260469e+09, 7.285175e+09, 7.308484e+09, 7.330385e+09, 7.350871e+09, 
    7.36993e+09, 7.387556e+09, 7.403741e+09, 7.418477e+09, 7.431758e+09, 
    7.443579e+09, 7.453934e+09, 7.462817e+09, 7.470226e+09, 7.476158e+09, 
    7.480609e+09, 7.483577e+09, 7.485062e+09, 7.485062e+09, 7.483577e+09, 
    7.480609e+09, 7.476158e+09, 7.470226e+09, 7.462817e+09, 7.453934e+09, 
    7.443579e+09, 7.431758e+09, 7.418477e+09, 7.403741e+09, 7.387556e+09, 
    7.36993e+09, 7.350871e+09, 7.330385e+09, 7.308484e+09, 7.285175e+09, 
    7.260469e+09, 7.234377e+09, 7.206909e+09, 7.178077e+09, 7.147894e+09, 
    7.116371e+09, 7.083523e+09, 7.049361e+09, 7.013901e+09, 6.977157e+09, 
    6.939143e+09, 6.899874e+09, 6.859367e+09, 6.817636e+09, 6.774699e+09, 
    6.730571e+09, 6.685269e+09, 6.638811e+09, 6.591213e+09, 6.542493e+09, 
    6.492669e+09, 6.441759e+09, 6.38978e+09, 6.336752e+09, 6.282692e+09, 
    6.227619e+09, 6.171552e+09, 6.114508e+09, 6.056508e+09, 5.99757e+09, 
    5.937712e+09,
  5.885548e+09, 5.942029e+09, 5.99757e+09, 6.052155e+09, 6.105772e+09, 
    6.158404e+09, 6.210038e+09, 6.260659e+09, 6.310255e+09, 6.35881e+09, 
    6.406312e+09, 6.452746e+09, 6.4981e+09, 6.54236e+09, 6.585513e+09, 
    6.627547e+09, 6.668449e+09, 6.708208e+09, 6.74681e+09, 6.784244e+09, 
    6.8205e+09, 6.855565e+09, 6.889429e+09, 6.922081e+09, 6.953512e+09, 
    6.98371e+09, 7.012667e+09, 7.040374e+09, 7.066821e+09, 7.092e+09, 
    7.115902e+09, 7.138521e+09, 7.159848e+09, 7.179877e+09, 7.198601e+09, 
    7.216014e+09, 7.23211e+09, 7.246883e+09, 7.260329e+09, 7.272444e+09, 
    7.283223e+09, 7.292662e+09, 7.30076e+09, 7.307511e+09, 7.312915e+09, 
    7.316969e+09, 7.319673e+09, 7.321026e+09, 7.321026e+09, 7.319673e+09, 
    7.316969e+09, 7.312915e+09, 7.307511e+09, 7.30076e+09, 7.292662e+09, 
    7.283223e+09, 7.272444e+09, 7.260329e+09, 7.246883e+09, 7.23211e+09, 
    7.216014e+09, 7.198601e+09, 7.179877e+09, 7.159848e+09, 7.138521e+09, 
    7.115902e+09, 7.092e+09, 7.066821e+09, 7.040374e+09, 7.012667e+09, 
    6.98371e+09, 6.953512e+09, 6.922081e+09, 6.889429e+09, 6.855565e+09, 
    6.8205e+09, 6.784244e+09, 6.74681e+09, 6.708208e+09, 6.668449e+09, 
    6.627547e+09, 6.585513e+09, 6.54236e+09, 6.4981e+09, 6.452746e+09, 
    6.406312e+09, 6.35881e+09, 6.310255e+09, 6.260659e+09, 6.210038e+09, 
    6.158404e+09, 6.105772e+09, 6.052155e+09, 5.99757e+09, 5.942029e+09, 
    5.885548e+09,
  5.832426e+09, 5.885548e+09, 5.937712e+09, 5.988909e+09, 6.039129e+09, 
    6.088361e+09, 6.136596e+09, 6.183825e+09, 6.230037e+09, 6.275223e+09, 
    6.319373e+09, 6.362479e+09, 6.404531e+09, 6.445522e+09, 6.485442e+09, 
    6.524282e+09, 6.562035e+09, 6.598693e+09, 6.634248e+09, 6.668692e+09, 
    6.702019e+09, 6.734221e+09, 6.76529e+09, 6.795221e+09, 6.824007e+09, 
    6.851641e+09, 6.878117e+09, 6.903431e+09, 6.927576e+09, 6.950547e+09, 
    6.972339e+09, 6.992947e+09, 7.012366e+09, 7.030593e+09, 7.047623e+09, 
    7.063453e+09, 7.078078e+09, 7.091497e+09, 7.103705e+09, 7.1147e+09, 
    7.124479e+09, 7.133041e+09, 7.140384e+09, 7.146505e+09, 7.151404e+09, 
    7.155078e+09, 7.157529e+09, 7.158754e+09, 7.158754e+09, 7.157529e+09, 
    7.155078e+09, 7.151404e+09, 7.146505e+09, 7.140384e+09, 7.133041e+09, 
    7.124479e+09, 7.1147e+09, 7.103705e+09, 7.091497e+09, 7.078078e+09, 
    7.063453e+09, 7.047623e+09, 7.030593e+09, 7.012366e+09, 6.992947e+09, 
    6.972339e+09, 6.950547e+09, 6.927576e+09, 6.903431e+09, 6.878117e+09, 
    6.851641e+09, 6.824007e+09, 6.795221e+09, 6.76529e+09, 6.734221e+09, 
    6.702019e+09, 6.668692e+09, 6.634248e+09, 6.598693e+09, 6.562035e+09, 
    6.524282e+09, 6.485442e+09, 6.445522e+09, 6.404531e+09, 6.362479e+09, 
    6.319373e+09, 6.275223e+09, 6.230037e+09, 6.183825e+09, 6.136596e+09, 
    6.088361e+09, 6.039129e+09, 5.988909e+09, 5.937712e+09, 5.885548e+09, 
    5.832426e+09 ;

 bk = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.01253, 0.04887, 0.10724, 0.18455, 0.27461, 0.36914, 
    0.46103, 0.54623, 0.62305, 0.69099, 0.75016, 0.8011, 0.84453, 0.88125, 
    0.9121, 0.93766, 0.95849, 0.97495, 0.98743, 0.9958, 1 ;

 pk = 1, 2.69722, 5.17136, 8.89455, 14.2479, 22.07157, 33.61283, 50.48096, 
    74.79993, 109.4006, 158.0046, 225.4411, 317.8956, 443.1935, 611.1156, 
    833.7439, 1125.834, 1505.208, 1993.158, 2614.863, 3399.784, 4382.062, 
    5600.87, 7100.731, 8931.782, 11149.97, 13817.17, 17001.21, 20775.82, 
    23967.34, 25527.65, 25671.22, 24609.3, 22640.51, 20147.13, 17477.63, 
    14859.86, 12414.93, 10201.44, 8241.503, 6534.432, 5066.179, 3815.607, 
    2758.603, 1880.646, 1169.339, 618.4799, 225, 10, 0 ;

 sftlf =
  0.3764576, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  0.9228161, 0.1739027, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  1, 0.8174675, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  1, 0.5504367, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  1, 0.9481694, 0.1901435, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  1, 1, 0.9983932, 0.2678785, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  1, 1, 1, 0.7833411, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.02900723, 0.3217153, 0.3830353, 
    0.5246126, 0.3472976, 0.1957928, 0.008647686, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 0.9731113, 0.3092794, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0006963735, 0.1754748, 0.4325673, 0.2951554, 
    0.6271494, 0.9393284, 1, 1, 1, 0.9934607, 0.9938456, 0.5638717, 
    0.02968918, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 0.9707108, 0.1046175, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0.06326846, 0.8031307, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 0.9995235, 0.7253351, 0.2813289, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 0.7709347, 0.06251514, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0.4201411, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 0.9849455, 0.1556062, 0.003983508, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 0.5608934, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.9381469, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.9549282, 0.5933414, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 0.8828677, 0.06657699, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0.6793007, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 0.8384063, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 0.669156, 0.0125583, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.1381188, 0.9697084, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 0.9104351, 0.2647975, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 0.04201834, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.00166111, 0.5541363, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 0.4645965, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 0.04201056, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.0307463, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 0.6972274, 0.5714607, 0.539219,
  1, 1, 1, 1, 1, 1, 1, 1, 0.04200291, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.2669835, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 0.5898379, 0.00854887, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.07485126, 0.9193581, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 0.4414221, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.0006397907, 0.4717199, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9447742, 0.2459255, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.1592281, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9522441, 0.693058, 0.077351, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.1598931, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.7353352, 0.09539028, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.6433973, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 0.6314353,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9975816, 0.8410712, 0.3690621, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.6869012, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9971337, 0.3079584, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.6868731, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.6658256, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.6868458, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9175764, 0.2185544, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.1822212, 0.9689022, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.7709059, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.651095, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9019616, 0.1664711, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.203948, 0.9547996, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.3274225, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.6748101, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.8615925, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.2362749, 0.9623896, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.8665756, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.7315421, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.8665628, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.7754121, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.8665506, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.2965498, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.8665391, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0509539, 0.8103296, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9383764, 0.2196166, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.7782937, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9603246, 
    0.0640404, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.2410026, 0.8761689, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.6294757, 
    0.007487927, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.7360525, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.266498, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.5350724, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9991729, 
    0.4061707, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.09449254, 0.8377889, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.9303989, 0.1264541, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.182272, 0.9179717, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.1799683, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.1560873, 0.8999666, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.3121897, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.4015228, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.159612, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.01152876, 0.7892212, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9283816, 
    0.6226964, 0.5535366, 0.06422334, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0.2964121, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.7704774, 
    0.05751295, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.03438287, 0.7932302, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9993793, 0.8113894, 0.6826136, 
    0.8702582, 0.5128348, 0.08204572, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.008766619, 0.6232422, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.7633693, 0.1774785, 0.2040459, 0, 0, 
    0.0009010995, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.6049436, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 0.9406916, 0.9853109, 0.9229649, 0.3723707, 
    0.03303384, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0.2605378, 0.9595606, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 0.9745548, 0.8413171, 0.115013, 0.1830149, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.3241267, 0.9822798, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 0.5268455, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.8645887, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 0.2353382, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.847726, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1,
  1, 1, 1, 1, 1, 0.7867104, 0.09881871, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.3535399, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 0.2738446, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1326434, 
    0.587546, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 0.01733101, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.01603992, 0.4454439, 0.6442813, 0.3830209, 0.05625193, 0, 
    0.03530673, 0.2579472, 0.08800853, 0, 0, 0, 0, 0, 0, 0.5546407, 
    0.6381541, 0.4571692, 0.7593831, 0.9919729, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 0.957557, 0.3666932, 0.001214215, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.06446161, 0.8062138, 1, 1, 1, 0.9404332, 0.9032256, 
    0.9204367, 1, 0.9587651, 0.5515207, 0.2075914, 0.002314975, 0, 0, 
    0.1886965, 0.9459232, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 0.9558364, 0.4539385, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.254573, 0.9151666, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.7619722, 
    0.6994123, 0.5289772, 0.9312455, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0.9320562, 0.7091275, 0.1623458, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.02540474, 0.619023, 0.9725087, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0.1557076, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.3710184, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.03056264, 
    0.5956897, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1148876, 0.5937533, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.07622165, 0.6823812, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.3449733, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.3805372, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.753692, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.3588129, 0.9958816, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.7856891, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.7856846, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01859863, 0.3884055, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.2158899, 0.9551845, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.3530129, 0.9508796, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.7544317, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.2654112, 0.9811226, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.6945245, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.07710309, 0.863272, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.6369579, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1824975, 
    0.7033954, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1683426, 
    0.8958945, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1531393, 
    0.5754542, 0.9937046, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.5226966, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.7708154, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.5950658, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.07487938, 0.8179564, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.03862339, 0.4152967, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 0.8500615, 0.946259, 0.884431, 0.7472318, 0.7092528, 
    0.9718166, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9999945, 
    0.4919434,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.004841657, 0.4270654, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 0.8776839, 0.7527315, 0.9694611, 0.8234424, 0.05545996, 0.01451342, 
    0.0766992, 0, 0, 0.7712654, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.740279, 0.0665665,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.1420659, 0.6810132, 0.2436509, 0.1621065, 0.2339793, 0.6901079, 
    0.9708213, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.8266005, 0.4517564, 0.04483075, 
    0.03248953, 0.1924889, 0.01307053, 0, 0, 0, 0, 0, 0.7712539, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9643438, 0.4936993, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.357605, 0.4481737, 0.01432, 0, 0, 0, 0.2996151, 0.8592404, 
    0.9996577, 1, 1, 1, 1, 1, 1, 1, 0.9999822, 0.3695327, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.1985431, 0.891767, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.4674213, 0.2888203, 0.163148,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.02609481, 0.6882609, 0.6668625, 0.8689135, 1, 0.997447, 0.9480262, 
    0.6412953, 0, 0, 0, 0.2262365, 0.6555864, 0.7921475, 0.9380791, 1, 1, 1, 
    1, 1, 0.6710668, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0618545, 0.7309781, 
    0.5937635, 0.3276973, 0.5878043, 0.4755114, 0.293394, 0.649609, 0.670538, 
    0.8472934, 1, 1, 1, 1, 0.942656, 0.977885, 0.3617498,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.03747177, 1, 1, 1, 1, 1, 1, 0.9728559, 0.7016522, 0.05877807, 0, 0, 0, 
    0, 0.0007180843, 0.2887189, 0.7476513, 0.6832384, 1, 1, 0.419323, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.009167003, 0, 0, 0, 0, 0, 0, 0.002281133, 
    0.2401035, 0.8190355, 1, 1, 1, 1, 0.6542072,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.4350484, 1, 1, 1, 1, 1, 1, 1, 1, 0.5818211, 0, 0, 0, 0, 0, 0, 0, 
    0.001013471, 0.1183226, 0.3208605, 0.3338135, 0, 0, 0, 0.006452882, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1757967, 0.6191416, 
    0.6542448, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.08844708, 1, 1, 1, 1, 1, 1, 1, 1, 0.4442382, 0, 0, 0.02307724, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.3639905, 0.6390771, 0.7038295, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.03658982, 0.4823922, 0.9029201, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.02019954, 0.7953823, 1, 1, 1, 1, 1, 1, 1, 0.8110214, 0.06406885, 0, 
    0.390024, 0.05420401, 0, 0, 0, 0, 0.4077412, 0.04842471, 0, 0, 0.1416207, 
    0.3410814, 0.6977392, 0.1285015, 0, 0, 0, 0, 0, 0, 0, 0, 0.1522885, 
    0.5140895, 0.258808, 0.0008218849, 0, 0, 0, 0, 0, 0, 0, 0, 0.02715651, 
    0.7257767,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.03747227, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.726593, 0.04869777, 0, 0, 0, 0, 
    0, 0, 0.8814211, 0.1349703, 0, 0, 0, 0, 0.01583155, 0.1170755, 0.247405, 
    0, 0, 0, 0, 0.0326486, 0.3860433, 0.1965477, 0, 0.00835224, 0.2670313, 
    0.005355601, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.4019571,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0374724, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.8357671, 0.2085238, 0, 0, 0, 
    0, 0, 0.809296, 0.1349555, 0, 0, 0, 0, 0, 0.09953156, 0.670812, 0, 0, 0, 
    0, 0.1109447, 1, 0.6344974, 0.005974696, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.2480379, 0.8815156, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.6203845, 0, 0, 0, 
    0, 0, 0.2954375, 0.07066895, 0, 0, 0, 0, 0.1317861, 0.6645802, 0.4592906, 
    0, 0.006340416, 0, 0.1393674, 0.7857525, 1, 1, 0.3672985, 0, 0, 0, 0, 
    0.000822613, 0.00348749, 0, 0, 0, 0.04631038, 0.06669453, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.14503, 0.4055507, 0.2551057, 0.3028015, 0.3623243, 0.4336107, 
    0.2924458, 0.9094968, 1, 1, 1, 0.7378889, 0.03122145, 0.001574896, 0, 0, 
    0, 0.7633188, 0.1349258, 0, 0.1208249, 0.5835989, 0.783038, 0.9167218, 1, 
    0.7098413, 0.4056285, 0.2833857, 0.1567454, 0.7330076, 1, 1, 0.9505261, 
    0.4874083, 0, 0, 0, 0.3619807, 0.7769179, 0.7792631, 0.6483424, 
    0.1295194, 0, 0.04274155, 0.6756219, 0.06986691, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.5567488, 1, 1, 1, 1, 0.7617028, 0.7580242, 
    0.8640846, 0.2590115, 0.01124508, 0.1238442, 0.05218257, 0.3791888, 
    0.9209204, 1, 1, 0.8919879, 0.9454092, 0.483057, 0.08077005, 0, 
    0.3203594, 1, 1, 1, 0.5728929, 0.0002312251, 0, 0, 0.5069734, 0.9029012, 
    1, 1, 1, 0.7427915, 0.221187, 0.2803968, 0.3342389, 0.03174093, 0 ;

 orog =
  8.54475, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  110.6839, 9.015973, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  118.8102, 18.13202, 0.007421071, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  130.705, 39.06387, 3.106806, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  141.0809, 84.24564, 11.19796, 0.4508977, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0,
  165.9822, 184.6116, 106.8482, 7.492514, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.08320683, 3.271346, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  180.4211, 249.8835, 220.8967, 76.21671, 1.021369, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    21.94272, 34.81591, 74.42256, 66.43814, 11.87937, 0, 0, 0, 0, 0, 0, 0, 0,
  149.0657, 196.1795, 177.1756, 126.4176, 11.39334, 0.5445582, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2.201014, 10.06274, 
    26.85098, 48.46229, 196.196, 446.1897, 398.605, 448.8601, 587.3398, 
    619.0617, 478.8845, 191.0291, 9.431361, 0, 0, 0, 0, 0, 0,
  247.4764, 260.0786, 196.9956, 132.1378, 48.361, 5.852092, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6.821061, 227.5061, 
    341.0564, 416.8428, 546.1491, 760.7002, 800.6117, 811.9203, 918.2296, 
    1199.078, 1194.457, 1065.196, 779.4019, 539.7784, 68.59048, 0, 0, 0, 0, 0,
  254.4188, 378.3603, 367.6226, 301.4343, 162.2049, 108.9995, 0.9085217, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8.392265, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    84.11958, 610.6379, 784.4166, 873.3272, 803.2366, 954.6566, 1133.667, 
    1193.683, 1333.627, 1518.089, 1657.062, 1719.367, 1548.189, 1097.09, 
    488.3766, 19.6729, 0, 0, 0, 0,
  282.803, 388.1694, 501.5489, 557.1978, 613.9719, 624.3671, 154.6011, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.850073, 136.7001, 
    621.1481, 1059.969, 1205.403, 1271.604, 1289.321, 1373.992, 1468.906, 
    1399.973, 1501.777, 1674.687, 2147.529, 2156.621, 1497.179, 907.9773, 
    341.0655, 33.16307, 0, 0, 0,
  281.039, 423.6907, 485.7559, 651.8676, 783.3052, 889.3768, 610.0162, 
    16.97377, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    129.3114, 660.4066, 997.0892, 1271.035, 1259.05, 1269.307, 1282.922, 
    1357.486, 1418.984, 1464.053, 1694.626, 2161.078, 2172.453, 1467.212, 
    1030.81, 612.332, 164.4304, 1.996331, 0, 0,
  322.6488, 427.8226, 549.0103, 681.7765, 829.639, 1022.879, 837.8648, 
    305.3638, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    9.138049, 280.6169, 659.5826, 1002.684, 1031.975, 1099.151, 1099.102, 
    1133.435, 1221.698, 1317.967, 1415.099, 1513.935, 1787.441, 1850.336, 
    1464.755, 1240.903, 696.9532, 172.8423, 13.54243, 0, 0,
  246.0376, 453.1236, 631.008, 871.3788, 1047.864, 932.1511, 816.0308, 
    317.9274, 6.631444, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    150.0291, 674.2753, 908.9203, 930.3144, 938.6702, 1006.137, 1124.25, 
    1170.841, 1154.932, 1264.449, 1330.767, 1451.47, 1585.219, 1689.979, 
    1656.847, 1377.684, 685.7067, 148.093, 7.893209, 0, 0,
  302.9081, 427.2077, 600.2842, 822.6921, 987.5324, 917.3104, 668.1157, 
    303.2888, 0.4759156, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.05529097, 404.3319, 849.9101, 942.0059, 899.2049, 892.3331, 1045.702, 
    1259.788, 1338.622, 1238.361, 1260.895, 1324.21, 1411.141, 1544.977, 
    1598.17, 1706.571, 1414.926, 652.4966, 175.4458, 20.1155, 25.00171, 
    36.41872,
  304.3976, 367.4553, 507.5162, 723.1177, 889.1189, 890.2856, 860.1849, 
    487.2796, 0.9306844, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    48.47385, 456.4773, 788.9446, 784.0788, 797.9801, 888.491, 1040.636, 
    1257.102, 1379.351, 1308.995, 1358.369, 1450.252, 1468.341, 1489.487, 
    1519.486, 1585.82, 1321.473, 545.1862, 138.8361, 40.63335, 49.9632, 
    84.77402,
  357.9227, 326.5664, 409.4615, 533.1976, 722.5844, 805.3265, 892.149, 
    651.6109, 85.95663, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6.497938, 272.2702, 615.2929, 908.9059, 917.061, 841.0509, 900.0991, 
    989.4551, 1097.285, 1229.295, 1245.714, 1381.851, 1374.066, 1291.548, 
    1248.401, 1166.31, 1273.148, 967.5308, 443.7959, 159.7697, 64.36124, 
    74.43269, 110.2169,
  374.3119, 313.8954, 345.6318, 445.4458, 583.0211, 721.8264, 795.6353, 
    683.6541, 309.0318, 22.92986, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 217.3822, 804.5779, 921.5053, 1073.372, 1032.455, 914.3887, 915.9861, 
    975.9174, 1025.77, 1091.464, 1183.756, 1203.829, 1146.519, 1118.986, 
    1206.85, 1186.365, 1061.127, 699.5498, 315.4096, 174.5182, 91.69196, 
    117.5326, 129.1317,
  384.2018, 316.835, 329.2943, 348.3972, 449.1535, 490.7008, 580.1392, 
    682.83, 561.0168, 450.0525, 74.4604, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 1.625334, 529.3156, 1179.003, 1083.251, 1046.369, 1010.433, 952.2749, 
    974.9957, 1008.044, 1025.375, 1088.216, 1136.371, 1137.306, 977.9841, 
    966.8591, 1095.862, 1080.748, 967.8829, 583.6017, 349.6461, 208.4064, 
    122.2884, 137.5921, 124.6154,
  425.9325, 402.693, 356.9512, 342.1429, 387.3358, 451.6554, 543.8193, 
    598.1646, 671.4254, 663.9327, 658.8842, 342.5872, 1.323529, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 55.75727, 723.3252, 1345.097, 1208.163, 1096.152, 
    1057.105, 1042.026, 1052.195, 1075.99, 1085.4, 1083.792, 1107.45, 
    1089.932, 1003.74, 908.7562, 881.2886, 806.4973, 725.7192, 521.3715, 
    374.6654, 268.3831, 172.0694, 131.0901, 57.53464,
  461.6035, 467.3536, 394.1595, 343.5833, 356.553, 412.9582, 456.8489, 
    546.8406, 586.7995, 714.7881, 969.0544, 855.0431, 500.8872, 32.52318, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 123.6441, 855.6476, 1413.006, 1269.892, 
    1172.559, 1156.56, 1149.75, 1151.305, 1144.381, 1103.469, 1061.514, 
    1045.96, 1102.312, 1112.108, 971.346, 808.2177, 695.4062, 630.5798, 
    525.356, 437.357, 384.1834, 350.2086, 123.1665, 31.22814,
  464.4684, 508.0797, 455.048, 373.7856, 366.4037, 387.9864, 443.3236, 
    495.3125, 589.3275, 739.6755, 988.6879, 1060.314, 904.9486, 528.0706, 
    225.8937, 27.69355, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 174.664, 879.7312, 1444.223, 
    1357.686, 1256.545, 1275.17, 1242.061, 1206.494, 1137.42, 1064.367, 
    1009.382, 1009.102, 1074.426, 1101.382, 1013.848, 935.0889, 872.3643, 
    823.5287, 742.5305, 702.767, 638.2717, 610.8529, 236.0903, 19.05215,
  377.5986, 476.2537, 554.4959, 498.4242, 421.1341, 410.7194, 460.7333, 
    508.1182, 604.0519, 780.8995, 940.6996, 912.0196, 1031.078, 860.0245, 
    593.0319, 288.8579, 12.86605, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 211.1246, 927.424, 
    1489.004, 1561.025, 1444.746, 1376.06, 1280.973, 1179.52, 1098.244, 
    1019.69, 975.9384, 963.2079, 978.0944, 1029.098, 1103.491, 1163.96, 
    1175.215, 1136.579, 1103.248, 1014.715, 943.465, 803.7495, 369.8148, 
    113.7734,
  332.751, 472.4073, 685.3926, 635.038, 517.4619, 464.7151, 489.6293, 
    589.0376, 704.1102, 888.3381, 946.3566, 843.2612, 937.7106, 952.2573, 
    593.1406, 408.6372, 87.12373, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 274.805, 948.42, 
    1506.014, 1601.052, 1578.846, 1456.921, 1284.965, 1163.84, 1079.576, 
    1015.096, 961.92, 924.3301, 919.1673, 969.1686, 1080.93, 1206.276, 
    1290.624, 1303.251, 1316.85, 1354.376, 1136.7, 970.1143, 487.621, 182.6047,
  386.6328, 599.5612, 743.3576, 737.4709, 670.9242, 536.273, 553.6517, 
    674.8468, 801.8613, 965.2466, 953.0202, 781.4857, 825.5333, 884.1866, 
    743.7918, 650.3617, 509.5243, 47.25615, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 34.19665, 536.6432, 
    1112.04, 1443.481, 1515.864, 1440.972, 1356.049, 1192.005, 1062.608, 
    976.4597, 953.9917, 942.6937, 942.3792, 969.4203, 966.9082, 1031.604, 
    1100.836, 1155.753, 1179.703, 1365.894, 1379.681, 1287.486, 922.5301, 
    544.6479, 214.8122,
  407.2789, 556.476, 691.2809, 737.9501, 749.3389, 662.7368, 563.8776, 
    667.7236, 775.2804, 860.3702, 857.4185, 735.3098, 719.4968, 858.9086, 
    655.9019, 560.5863, 441.2978, 138.1514, 0.004807308, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 245.0765, 
    740.5414, 1216.22, 1399.232, 1428.595, 1324.44, 1244.887, 1171.623, 
    1058.757, 978.5461, 948.2759, 945.5349, 979.3757, 1012.527, 980.8537, 
    912.5103, 983.9648, 1005.987, 1126.251, 1280.425, 1263.255, 944.915, 
    620.7706, 330.2798, 198.4007,
  485.9347, 536.7831, 520.842, 574.1156, 628.2961, 593.3192, 671.6805, 
    760.3802, 792.5333, 809.5409, 713.7068, 694.2451, 762.8157, 893.8396, 
    750.4239, 489.7271, 319.0528, 122.3887, 1.660121, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.1749505, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 36.20846, 
    639.6878, 1064.495, 1200.584, 1345.762, 1339.131, 1276.558, 1206.219, 
    1145.992, 1077.639, 997.5162, 966.3801, 956.3568, 970.2714, 1008.335, 
    951.059, 828.9758, 706.606, 863.0428, 1080.806, 1123.896, 920.291, 
    656.9827, 373.7796, 334.5416, 526.0103,
  571.2805, 576.3853, 467.4599, 411.0854, 392.3285, 505.7308, 722.9926, 
    869.4109, 931.8525, 811.3553, 662.9765, 604.0966, 688.219, 858.3245, 
    825.9299, 572.1747, 408.3769, 146.4941, 9.387668, 0.001074584, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    273.4626, 965.0869, 1142.758, 1166.024, 1121.857, 1187.254, 1166.343, 
    1151.341, 1121.571, 1066.005, 1020.396, 995.9119, 976.3922, 999.8099, 
    1080.855, 1153.143, 949.2833, 796.8798, 704.9807, 751.8674, 635.2756, 
    537.6038, 460.5406, 432.7109, 753.7834, 783.1511,
  541.8253, 527.6813, 442.9381, 349.75, 282.5704, 372.3629, 647.7617, 
    839.8668, 941.1125, 907.2533, 705.0693, 633.6419, 637.7145, 768.287, 
    809.7827, 674.5598, 493.8878, 279.3312, 44.60109, 0.003030813, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    59.35226, 753.0102, 1128.37, 1213.516, 1102.814, 1106.985, 1138.11, 
    1148.302, 1144.664, 1119.719, 1075.693, 1028.648, 1007.681, 1040.419, 
    1070.42, 1085.326, 1113.797, 1101.634, 964.3666, 826.3594, 688.6269, 
    581.0179, 749.9571, 747.4507, 813.9899, 1027.863, 909.4127,
  451.7546, 465.3449, 395.6716, 335.8462, 247.0956, 298.3383, 466.0626, 
    661.6984, 813.6958, 827.1074, 757.3602, 671.0699, 631.3232, 636.7422, 
    748.9434, 753.5067, 653.6973, 358.9735, 111.3765, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 237.6711, 881.6313, 
    1209.199, 1111.17, 1116.662, 1148.323, 1170.288, 1177.596, 1179.032, 
    1162.061, 1096.823, 1040.075, 1027.026, 1072.69, 1144.079, 1132.332, 
    1099.773, 1094.171, 1114.551, 970.8142, 812.7686, 713.1152, 878.1364, 
    977.2021, 1026.251, 1069.996, 736.0057,
  391.2837, 370.3196, 366.6443, 340.5762, 263.041, 234.9373, 359.7917, 
    485.6016, 684.4538, 736.9855, 740.4536, 781.7585, 658.1667, 565.2335, 
    713.5017, 808.0051, 692.545, 472.7854, 120.2969, 0.03788849, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 152.0637, 
    745.3533, 1129.647, 1190.232, 1165.257, 1217.449, 1233.613, 1242.039, 
    1225.1, 1190.186, 1129.522, 1051.2, 1039.217, 1088.383, 1158.137, 
    1160.562, 1157.639, 1146.778, 1176.388, 1196.262, 1103.755, 939.6448, 
    773.607, 786.1696, 1066.588, 999.4681, 658.9298,
  343.9839, 329.1209, 326.8227, 338.2211, 268.4422, 231.5902, 273.1661, 
    411.1793, 556.3333, 647.4001, 724.2601, 776.667, 679.067, 508.2994, 
    620.4402, 716.1536, 666.8013, 484.4005, 195.8266, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 49.35054, 549.8828, 
    1179.242, 1286.947, 1285.081, 1347.293, 1373.125, 1342.854, 1282.255, 
    1234.189, 1156.042, 1075.134, 1044.677, 1093.778, 1146.635, 1190.949, 
    1194.665, 1203.338, 1225.234, 1270.81, 1379.499, 1236.873, 994.0289, 
    744.1392, 1000.295, 1032.345, 591.7537,
  341.9223, 323.5297, 312.363, 327.7422, 256.121, 211.4899, 232.2774, 
    293.0904, 373.0227, 483.3326, 649.4127, 771.75, 673.2164, 571.9428, 
    626.7587, 791.145, 642.7789, 521.3182, 201.4202, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 3.703202, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10.91209, 
    566.6647, 1165.319, 1443.802, 1442.337, 1513.629, 1471.694, 1443.57, 
    1354.923, 1276.675, 1185.226, 1087.362, 1080.905, 1145.881, 1175.568, 
    1221.021, 1282.013, 1268.265, 1230.614, 1228.024, 1211.29, 1307.737, 
    1161.229, 873.0657, 933.2297, 1159.808, 670.6091,
  346.7993, 338.6057, 314.9171, 289.7007, 236.9087, 190.2888, 202.9013, 
    268.8091, 310.8858, 411.589, 656.1295, 740.801, 656.6727, 541.4875, 
    678.8455, 853.9406, 730.4851, 459.3751, 220.1203, 13.96118, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    413.7036, 981.3401, 1411.613, 1624.979, 1620.908, 1479.521, 1444.335, 
    1392.403, 1297.059, 1161.221, 1098.89, 1153.009, 1254.525, 1302.453, 
    1335.512, 1364.571, 1280.526, 1204.677, 1180.655, 1170.281, 1240.504, 
    1336.752, 1084.095, 1070.497, 1113.52, 930.3657,
  373.4141, 339.6274, 318.1039, 291.9559, 260.7186, 191.6193, 197.949, 
    276.8808, 356.4713, 444.8528, 671.9672, 707.4572, 541.8743, 515.196, 
    593.6595, 844.5728, 740.3514, 450.5794, 236.8895, 126.5775, 12.02609, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    74.79279, 582.2818, 1387.929, 1653.479, 1656.323, 1452.037, 1384.894, 
    1380.74, 1263.157, 1129.277, 1087.819, 1140.283, 1291.528, 1349.267, 
    1427.148, 1380.747, 1211.18, 1182.415, 1173.129, 1242.567, 1253.907, 
    1328.973, 1235.93, 1102.579, 1212.149, 1188.651,
  411.907, 359.5694, 312.9021, 316.0843, 319.7564, 228.2056, 193.8342, 
    296.6815, 321.6121, 390.0383, 586.1972, 616.8071, 522.6686, 497.1555, 
    514.1055, 625.6185, 709.9496, 500.6991, 322.1615, 233.313, 73.02024, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 251.8302, 1240.724, 1602.32, 1519.831, 1331.846, 1307.905, 1319.815, 
    1247.846, 1123.754, 1088.791, 1091.119, 1166.166, 1236.438, 1262.825, 
    1296.363, 1122.022, 1172.453, 1197.705, 1311.24, 1400.86, 1405.443, 
    1374.509, 1337.278, 1486.886, 1500.223,
  361.1769, 319.2283, 308.7516, 344.1496, 351.8325, 252.6501, 205.3004, 
    264.0542, 284.5062, 319.0981, 459.6907, 492.8576, 454.6547, 494.1764, 
    467.236, 499.1732, 633.0408, 550.3798, 449.2036, 364.1278, 174.6403, 
    28.89057, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 104.2696, 1010.841, 1362.054, 1315.101, 1130.426, 1149.357, 
    1245.088, 1169.575, 1095.747, 1041.157, 1027.792, 1023.939, 991.415, 
    1043.899, 1006.476, 1261.374, 1189.962, 1103.186, 1205.096, 1273.994, 
    1571.499, 1265.122, 1354.616, 1342.277, 1499.963,
  288.3837, 296.7624, 328.1481, 349.2853, 354.0044, 300.8336, 209.8271, 
    242.339, 257.6059, 315.6365, 438.6422, 454.057, 469.7331, 499.5292, 
    472.8086, 418.0537, 492.4049, 451.988, 414.6512, 387.9483, 298.7437, 
    224.9868, 30.84828, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.8451669, 71.35338, 642.9059, 1073.645, 1063.941, 
    943.9172, 1026.204, 1114.221, 1073.748, 1012.559, 1027.82, 1014.382, 
    1057.285, 1027.442, 823.2462, 941.8942, 1091.702, 1226.689, 1104.525, 
    1242.194, 1126.849, 1339.002, 1262.845, 1232.307, 1363.345, 1223.546,
  260.1389, 284.7289, 287.6657, 321.2379, 323.3841, 321.9951, 239.3829, 
    211.8097, 231.2988, 276.1485, 389.8618, 400.1599, 419.2465, 413.5182, 
    379.3967, 365.7533, 402.7262, 476.0164, 436.6118, 442.7455, 523.3729, 
    513.603, 263.7818, 2.99741, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 6.84726, 127.0682, 564.7839, 1027.651, 923.8217, 
    809.4365, 946.3239, 1098.568, 971.295, 901.8392, 924.174, 968.075, 
    986.755, 1009.199, 898.538, 673.96, 868.1624, 893.8102, 1322.028, 
    1317.703, 1118.277, 1254.662, 1102.685, 1225.965, 1365.095, 1100.581,
  256.0101, 258.5121, 265.4595, 271.6456, 281.9239, 339.2019, 239.4398, 
    201.6286, 231.9184, 272.3331, 346.6201, 365.2863, 335.9691, 301.0338, 
    258.306, 271.6318, 450.0833, 557.5646, 531.2784, 522.4316, 549.2473, 
    622.1465, 329.0093, 25.54767, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 6.427928, 262.789, 692.8567, 1032.231, 824.3097, 
    711.4518, 954.0336, 994.9745, 852.847, 765.702, 840.2001, 873.9611, 
    851.5475, 920.1156, 891.8646, 743.049, 630.5678, 807.291, 1051.364, 
    1174.423, 1034.36, 1105.102, 1130.744, 1221.451, 1312.698, 1236.457,
  244.8726, 235.7898, 238.6499, 250.9584, 264.177, 304.3681, 231.7038, 
    171.5492, 194.0964, 237.4297, 322.8626, 324.8877, 315.0707, 258.6005, 
    236.6363, 277.2534, 457.8071, 528.7694, 405.2236, 342.8656, 385.32, 
    442.8686, 295.1935, 24.17916, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 1.293201, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 52.95097, 347.3517, 720.2449, 929.5432, 
    735.391, 780.5626, 910.9541, 885.9318, 687.3369, 662.2593, 723.8735, 
    755.4806, 723.0743, 769.8126, 788.1163, 702.8589, 630.3057, 768.6213, 
    1059.849, 972.3868, 1188.259, 1177.481, 1121.192, 1184.726, 1279.616, 
    1302.242,
  235.042, 217.7554, 200.0201, 218.5201, 210.6107, 214.8637, 159.0711, 
    132.8887, 194.6062, 222.7486, 255.3079, 243.1668, 189.8971, 189.5496, 
    151.8132, 254.9043, 441.0879, 450.9707, 312.1183, 209.6811, 199.2862, 
    258.3366, 160.7645, 4.592148, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.1700515, 92.22056, 366.6779, 594.3502, 777.5218, 
    693.3395, 719.6742, 801.9887, 715.3484, 599.9813, 555.8511, 606.0909, 
    628.077, 622.9703, 659.368, 666.463, 613.6947, 660.4321, 819.1418, 
    1024.8, 1005.07, 1167.154, 1107.55, 1131.997, 1173.377, 1208.152, 1350.651,
  196.7365, 204.5998, 198.4898, 193.5049, 169.7109, 154.1599, 121.315, 
    140.5267, 197.9303, 241.7397, 228.9246, 149.1499, 105.5863, 101.0614, 
    123.9294, 166.2768, 433.4229, 365.3992, 271.7154, 133.414, 51.558, 
    55.21501, 35.0076, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 13.58836, 185.3467, 334.9186, 518.5123, 624.0504, 611.5664, 
    573.1268, 551.8474, 545.7886, 508.7069, 509.3336, 518.7409, 552.8677, 
    565.2957, 587.2665, 552.8708, 585.5536, 619.3701, 901.4293, 1212.324, 
    1221.37, 1192.156, 1120.597, 1169.473, 1176.514, 1126.01, 1376.636,
  146.6925, 179.7951, 169.8683, 144.5109, 115.9851, 100.912, 77.22723, 
    96.99864, 139.7948, 160.3108, 134.8792, 69.91695, 26.29307, 64.91444, 
    76.29048, 164.2859, 290.0237, 281.2162, 184.3736, 70.43913, 2.701435, 0, 
    0, 0, 0, 0.09234287, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 2.41791, 93.65132, 238.9857, 412.0441, 452.2166, 553.3406, 506.5167, 
    421.6122, 392.6665, 425.7772, 440.7444, 462.4359, 492.6555, 517.598, 
    531.2183, 527.7665, 529.114, 571.4398, 752.8386, 1117.882, 1654.942, 
    1618.519, 1398.75, 1202.588, 1191.508, 1195.801, 1221.172, 1415.927,
  69.31319, 104.212, 110.316, 83.84324, 63.33185, 52.58361, 41.60804, 
    45.76586, 76.87368, 101.9827, 93.67348, 33.04323, 20.12624, 46.1826, 
    54.88905, 34.84738, 115.9459, 49.21751, 40.83882, 0.5943004, 0, 0, 0, 0, 
    0, 0.0057942, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.398386, 
    119.9112, 199.3601, 411.994, 476.3767, 578.0508, 529.0004, 436.2539, 
    335.8598, 335.8933, 358.957, 401.7341, 439.7245, 481.3549, 499.7074, 
    519.8088, 515.3641, 502.7769, 560.4839, 723.5606, 1163.4, 1705.951, 
    1771.096, 1455.29, 1286.019, 1198.102, 1179.159, 1260.96, 1461.374,
  79.25274, 98.79363, 46.67113, 25.34361, 28.43618, 24.51583, 16.18622, 
    19.50146, 37.39209, 67.61229, 56.61288, 32.74178, 14.21986, 3.174914, 
    2.647948, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.01747818, 46.90157, 207.9118, 460.4455, 514.9199, 
    602.9887, 590.7431, 513.9005, 364.6547, 319.0529, 315.5271, 335.9451, 
    373.1736, 425.5178, 449.45, 464.8029, 490.2738, 503.6892, 494.0532, 
    586.5953, 751.3316, 1115.167, 1723.364, 1792.263, 1481.577, 1256.694, 
    1160.092, 1138.162, 1189.935, 1531.006,
  304.3052, 225.9071, 146.4976, 49.22798, 14.06787, 15.70426, 14.31254, 
    10.55259, 21.65571, 34.42345, 26.47721, 10.16362, 1.715719, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.3261773, 0, 0, 5.140869, 66.8336, 316.336, 486.2376, 557.2535, 
    481.0815, 482.611, 398.9484, 317.3685, 310.7681, 323.2128, 329.6191, 
    362.9882, 389.781, 416.3743, 421.8354, 456.8871, 480.976, 483.8488, 
    540.1299, 714.4539, 990.8341, 1670.664, 1620.258, 1494.627, 1232.962, 
    1134.55, 1134, 1203.068, 1431.174,
  377.3476, 300.3462, 179.3239, 123.5264, 29.18042, 8.49296, 10.41877, 
    2.594529, 2.675612, 3.391332, 0.1138654, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.007269558, 0, 
    7.853471, 62.3085, 274.8862, 413.5488, 423.2161, 435.7926, 444.4748, 
    361.6428, 308.9561, 319.7975, 321.1809, 340.5662, 354.3437, 378.4564, 
    404.6211, 438.1272, 444.1309, 457.4094, 472.3898, 582.7078, 713.5034, 
    965.1596, 1325.418, 1513.297, 1287.996, 1268.213, 1155.886, 1135.109, 
    1137.983, 1441.737,
  397.6618, 290.1455, 262.0854, 164.1737, 72.91979, 9.641136, 3.297817, 
    0.002408294, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24.52353, 0, 1.134986, 131.7988, 
    413.9996, 487.4259, 485.74, 514.1754, 483.7487, 398.7583, 334.6064, 
    318.3876, 329.1971, 343.4026, 364.3184, 386.8412, 433.8055, 462.0353, 
    443.1543, 453.2259, 475.2897, 560.871, 675.3644, 778.7476, 1195.336, 
    1219.456, 1293.797, 1255.619, 1167.165, 1128.763, 1127.737, 1605.608,
  359.7442, 322.1634, 256.7101, 190.8573, 99.29717, 20.20619, 2.261762, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 1.042433, 1.061284, 0.06026918, 221.4693, 588.1027, 
    609.5046, 567.6266, 539.7374, 519.683, 443.9848, 375.9164, 330.9009, 
    328.2888, 345.5885, 367.2719, 396.1122, 425.6252, 436.9988, 445.1413, 
    455.4268, 478.2379, 538.37, 618.6725, 704.752, 879.9337, 1044.206, 
    1143.218, 1000.543, 1114.351, 1055.759, 1244.916, 1644.584,
  339.5918, 283.2596, 244.217, 182.1556, 115.8238, 16.9204, 1.281723, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 118.1892, 542.7286, 664.8825, 616.7386, 
    595.4612, 551.9771, 495.2496, 416.2375, 373.1087, 345.3355, 352.5166, 
    377.2891, 390.3913, 413.6357, 444.6428, 442.3636, 488.6983, 526.4742, 
    581.7993, 665.6102, 783.5282, 909.798, 1160.341, 1189.347, 1036.943, 
    1004.612, 1053.218, 1059.908, 1416.363,
  279.6242, 227.4193, 199.1174, 149.1774, 83.37285, 3.592551, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 101.2812, 60.90662, 478.8484, 643.0255, 690.905, 
    652.9017, 619.0784, 549.6542, 517.7484, 445.3293, 372.7345, 391.3872, 
    396.3501, 434.3335, 453.7928, 469.5943, 484.0396, 513.5276, 579.3093, 
    651.2834, 708.0594, 776.8271, 870.302, 1036.794, 1245.989, 901.5364, 
    940.5923, 1070.94, 1195.01, 1146.841,
  196.4323, 187.7343, 179.3497, 120.5639, 39.21375, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2.005413, 45.81821, 62.24737, 21.02495, 
    3.207724, 0.02404907, 1.234567, 12.24459, 1.728072, 0, 0, 0, 0, 0, 0, 
    3.453561, 7.352701, 19.79626, 158.7443, 296.7885, 521.1622, 627.5361, 
    662.5475, 682.7275, 655.5103, 590.583, 580.2885, 526.9755, 427.6072, 
    407.3717, 430.1629, 446.7533, 474.6825, 500.0133, 519.8837, 559.5943, 
    617.9446, 655.3353, 686.9636, 713.472, 753.1322, 906.1678, 1018.012, 
    815.1847, 882.2279, 1056.679, 1259.787, 1045.098,
  141.7976, 159.4438, 144.7507, 76.36758, 7.418705, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5.733681, 94.68479, 175.18, 187.5313, 
    155.0462, 110.0206, 72.29835, 93.21919, 121.2557, 115.5466, 66.30669, 
    6.150113, 0, 0, 0, 3.670892, 28.15756, 46.06707, 79.14339, 305.7281, 
    712.5394, 940.3807, 751.7666, 698.2665, 746.433, 768.7173, 723.7104, 
    672.3049, 616.0403, 509.8206, 453.0623, 453.5248, 504.1813, 528.5236, 
    544.4155, 565.7984, 598.8699, 625.6595, 655.5828, 686.7064, 683.7915, 
    732.2036, 789.5637, 840.5327, 723.5177, 745.4189, 965.6844, 1038.274, 
    796.5178,
  95.12392, 103.6217, 82.47251, 13.03405, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.002540734, 15.74638, 122.9433, 222.9018, 302.6361, 
    279.6983, 224.5893, 190.8986, 149.559, 188.5142, 236.7475, 212.6731, 
    150.321, 153.6949, 48.69242, 25.20141, 29.67488, 91.25098, 132.1451, 
    112.2913, 103.7838, 263.8452, 764.3199, 1062.096, 1009.38, 884.1952, 
    931.0499, 977.1282, 882.8214, 713.9742, 616.5552, 536.9384, 509.7403, 
    500.2069, 555.3665, 585.5272, 600.3098, 607.6362, 615.286, 634.0374, 
    661.1276, 645.6732, 626.6214, 638.4325, 669.1021, 625.0273, 530.0295, 
    528.0609, 601.1044, 644.5855, 548.4876,
  30.5022, 27.99392, 7.313161, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.7658302, 12.3739, 142.0602, 300.8344, 465.4789, 498.4969, 
    391.7122, 316.7618, 249.2353, 219.1284, 259.9997, 244.4664, 174.3858, 
    179.9653, 249.7257, 193.2922, 150.1301, 234.5797, 302.7541, 285.0494, 
    207.801, 158.7262, 115.508, 347.3649, 690.9739, 928.4409, 982.3543, 
    1030.41, 1034.681, 877.8196, 652.1367, 503.6282, 493.2419, 491.9219, 
    520.8734, 593.4538, 643.876, 652.7304, 662.8006, 652.0361, 676.1411, 
    653.5867, 602.203, 551.5805, 537.899, 522.2339, 492.5406, 445.3781, 
    430.9313, 431.1991, 487.3873, 602.6268,
  0.766829, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7.8648, 
    83.18796, 276.2613, 500.1916, 600.5903, 597.6884, 475.5048, 352.7767, 
    314.1613, 281.9288, 287.8528, 237.377, 131.9863, 144.99, 306.4143, 
    294.3946, 305.1169, 332.2526, 310.4181, 229.8286, 185.2745, 224.0371, 
    255.049, 135.4041, 273.2138, 527.6912, 587.1231, 611.7789, 642.2618, 
    595.1403, 463.5603, 424.1609, 415.3838, 429.1796, 490.9037, 608.7256, 
    694.1671, 728.9787, 711.6575, 716.4285, 701.124, 642.769, 552.2159, 
    495.597, 465.6459, 440.4718, 429.3813, 424.0435, 422.3978, 418.5041, 
    446.8545, 718.7314,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.295444, 78.97375, 
    275.3757, 455.0948, 458.2011, 506.2027, 494.194, 412.8863, 375.2495, 
    355.046, 307.8675, 307.6067, 255.4145, 162.655, 174.7049, 269.6479, 
    362.2924, 358.3284, 318.2245, 211.9518, 198.9956, 327.952, 577.7234, 
    678.533, 449.4442, 258.9631, 309.9615, 318.2204, 354.7622, 372.4727, 
    407.3471, 409.3253, 394.0547, 388.1353, 397.6263, 455.2305, 588.9576, 
    706.325, 787.8987, 810.1958, 757.8834, 690.1829, 588.7928, 504.9205, 
    456.3733, 419.4193, 401.9965, 409.1686, 411.8871, 415.8695, 412.8529, 
    415.983, 653.3243,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.04495476, 1.543852, 
    40.60966, 249.5493, 570.8077, 624.9529, 503.8392, 404.5659, 388.5279, 
    371.8024, 372.5071, 373.0171, 344.5746, 314.8991, 279.2988, 232.3392, 
    204.3131, 251.619, 321.1378, 336.9094, 265.9687, 241.0423, 314.6817, 
    503.8398, 693.5359, 810.1852, 579.9879, 386.7859, 384.9114, 418.0108, 
    446.1444, 373.0016, 350.7278, 352.2296, 366.1898, 378.6504, 386.957, 
    403.5961, 448.4445, 545.6042, 676.7407, 741.8482, 705.261, 612.5644, 
    508.2358, 457.7974, 419.8724, 397.5679, 394.2395, 399.4266, 405.9669, 
    407.882, 402.7976, 410.4689, 789.8555,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.7914926, 10.71653, 
    37.00443, 201.4314, 448.087, 531.7697, 431.7727, 398.7067, 393.9764, 
    349.5272, 333.6953, 360.2705, 337.4265, 298.6373, 309.2917, 282.9134, 
    270.9925, 231.9091, 272.6257, 235.9534, 234.1443, 273.3409, 414.232, 
    561.9924, 633.738, 604.2332, 478.0908, 428.5763, 404.8661, 464.5562, 
    464.1216, 373.5608, 319.6164, 329.3439, 353.2355, 408.3477, 412.724, 
    410.5272, 419.3637, 448.9814, 538.6779, 576.0292, 562.1622, 501.3907, 
    457.8747, 424.4431, 405.648, 395.4491, 393.9858, 397.7108, 400.8848, 
    400.0156, 396.7203, 474.1039, 980.1252,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6.459178, 23.89642, 
    39.5673, 52.56926, 168.347, 227.195, 285.7491, 353.7228, 381.3757, 
    362.791, 311.1005, 312.541, 320.0593, 289.4526, 308.0459, 311.635, 
    295.6172, 265.5541, 242.1341, 228.7672, 222.6893, 264.653, 356.3772, 
    481.8984, 514.7236, 444.572, 376.3537, 375.8529, 367.9664, 341.9634, 
    351.7896, 291.5329, 307.0333, 322.6101, 365.6251, 444.1953, 465.1169, 
    441.8697, 452.7754, 478.7091, 527.0575, 540.0756, 491.8977, 461.4532, 
    433.0887, 417.837, 414.4355, 413.9627, 410.6415, 421.8182, 400.1716, 
    394.3721, 399.2646, 611.9307, 1308.194,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6.790205, 27.87427, 
    37.87522, 49.99376, 77.3848, 129.5688, 225.8023, 291.5181, 345.4376, 
    327.5065, 299.076, 285.3165, 292.4263, 320.6955, 306.0085, 310.2983, 
    291.4063, 262.9675, 246.8307, 238.5132, 249.1621, 271.4966, 326.77, 
    393.712, 450.9673, 416.2671, 374.2629, 344.2727, 333.5673, 305.9854, 
    280.9805, 285.871, 292.4921, 298.5072, 329.7079, 419.0633, 450.0066, 
    465.448, 502.8485, 574.8007, 637.0599, 703.0728, 587.3303, 483.8123, 
    452.7943, 442.7585, 455.8902, 478.3641, 513.434, 528.1032, 446.6922, 
    395.0017, 396.0436, 580.3947, 1096.152,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 7.539374, 13.82793, 0, 0, 0, 0, 0, 0.3629586, 
    22.22618, 38.05198, 50.36842, 51.9423, 55.76481, 123.9351, 200.9567, 
    248.0657, 288.369, 296.5797, 284.997, 272.4008, 306.0285, 313.191, 
    326.7126, 292.9926, 277.2778, 264.6691, 265.5726, 260.786, 272.6996, 
    322.4322, 380.3541, 402.2595, 439.8839, 455.1393, 427.6396, 381.3865, 
    336.1739, 308.6934, 286.1038, 296.1768, 298.6016, 292.2509, 297.8213, 
    348.2343, 392.0045, 441.4889, 561.517, 686.3062, 815.3308, 935.5671, 
    875.5865, 574.7263, 510.7076, 481.0591, 505.4455, 569.8447, 637.2155, 
    645.5725, 578.0183, 406.8309, 416.0845, 555.6661, 828.242,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 6.968982, 31.56356, 1.362759, 0, 0, 0, 0, 0, 
    9.483889, 33.60556, 38.53296, 50.37358, 74.38406, 139.3567, 205.6824, 
    215.1312, 223.8199, 264.2617, 295.2328, 280.9891, 269.5547, 301.0195, 
    283.1612, 300.8699, 290.1711, 288.1376, 298.2253, 296.4409, 301.7662, 
    372.0651, 450.2336, 467.1264, 467.0771, 487.0597, 462.8398, 408.4555, 
    374.192, 332.696, 321.5491, 328.5142, 322.4901, 299.8736, 293.3217, 
    324.0511, 366.8441, 447.5163, 626.8708, 836.7401, 890.7211, 1096.81, 
    1047.843, 760.592, 575.9907, 540.1681, 540.2332, 595.8331, 628.45, 
    649.7249, 568.4493, 455.0399, 431.6068, 517.0565, 601.8608,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 1.797053, 7.747849, 3.450143, 0, 0, 0, 0, 0, 
    0.9109401, 18.42504, 39.59516, 52.26551, 97.90691, 235.892, 219.3992, 
    208.2924, 216.5296, 262.5898, 292.2108, 286.3712, 274.5794, 269.5547, 
    279.5371, 287.6822, 293.7041, 308.5545, 345.3323, 335.1651, 328.9469, 
    369.3367, 444.4053, 470.777, 502.3892, 510.839, 472.6234, 420.1351, 
    393.2463, 375.5051, 344.6975, 341.879, 320.9992, 295.3217, 288.8875, 
    310.2828, 356.9085, 436.3004, 643.2478, 908.5942, 908.9702, 1001.605, 
    1072.39, 855.878, 706.8087, 615.7324, 594.7244, 607.8818, 589.8001, 
    519.1802, 495.0875, 398.2069, 416.0681, 481.5428, 468.7679,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 45.77684, 0, 0, 0, 0, 0, 0, 0, 0, 19.37672, 
    35.37803, 69.18604, 153.2726, 288.3199, 317.8352, 244.572, 258.4949, 
    287.7384, 311.5768, 297.4268, 289.1551, 278.5264, 276.3994, 304.6932, 
    323.0869, 346.2746, 396.4057, 380.4884, 341.7323, 349.6577, 376.4726, 
    426.947, 504.5984, 651.9197, 501.9165, 434.0541, 415.7284, 411.0024, 
    387.9035, 340.0662, 290.0233, 265.8179, 252.4831, 284.6985, 349.8331, 
    406.4402, 572.5109, 805.2451, 886.5491, 902.3984, 984.8835, 957.6617, 
    842.1849, 709.3141, 604.957, 577.4132, 542.0748, 476.5501, 421.5896, 
    398.5287, 416.1053, 436.3309, 444.6508,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.2233779, 7.883308, 
    46.45991, 63.79469, 184.3558, 336.8821, 374.0247, 374.8209, 335.6512, 
    339.178, 324.0201, 312.332, 293.5074, 275.675, 291.9893, 330.8283, 
    374.3214, 414.9174, 493.441, 464.5028, 388.4646, 358.354, 358.3539, 
    399.2584, 604.8146, 824.4387, 636.0546, 425.0211, 422.0507, 444.4562, 
    444.8008, 388.2694, 300.7451, 240.5886, 216.5688, 229.7297, 312.2461, 
    400.7599, 488.0696, 759.7354, 869.7776, 810.3863, 836.918, 927.7097, 
    906.3384, 778.0356, 610.2334, 542.7169, 508.4426, 490.6646, 424.6607, 
    396.6208, 405.9286, 424.3958, 467.8904,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.524688, 44.15213, 
    88.41959, 159.127, 276.4428, 370.4227, 392.6274, 382.1442, 366.4334, 
    336.8749, 317.2722, 299.4598, 286.5885, 283.6873, 292.2945, 335.28, 
    393.107, 469.711, 592.4265, 585.6436, 482.2569, 415.559, 389.8748, 
    408.3621, 619.8497, 895.7261, 639.1478, 447.5954, 410.7881, 450.1098, 
    465.333, 443.5472, 380.2547, 332.284, 295.5856, 256.3805, 299.0791, 
    379.3657, 547.1831, 780.5206, 955.9313, 825.8504, 679.0082, 745.6443, 
    771.3798, 700.3216, 547.1471, 488.1773, 493.5975, 534.8677, 465.9749, 
    408.6629, 406.9938, 428.9316, 486.2154,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8.648079, 90.31952, 
    139.5776, 213.0849, 372.9224, 415.0632, 410.2803, 377.4778, 360.1422, 
    341.8087, 303.7456, 280.1181, 284.2162, 290.7113, 310.3253, 325.1641, 
    379.646, 458.2865, 595.5748, 642.431, 599.8919, 527.5738, 473.18, 
    483.1668, 614.2881, 799.8925, 603.7574, 431.5247, 413.0665, 434.388, 
    454.1592, 461.4271, 468.4397, 452.5511, 440.9289, 400.6418, 349.5063, 
    404.0337, 485.1346, 668.6317, 844.2675, 779.2899, 658.3606, 603.169, 
    619.9202, 579.0063, 475.0612, 424.7502, 455.7198, 513.4985, 468.9218, 
    415.5838, 421.0052, 460.8036, 482.3849,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26.58741, 141.5162, 
    204.9548, 236.1427, 343.1058, 379.2624, 360.7214, 335.7108, 336.3476, 
    332.6995, 308.2321, 285.1463, 271.4974, 292.8643, 320.6105, 328.3786, 
    355.2569, 397.3354, 482.0117, 568.8033, 603.5388, 619.1583, 583.2557, 
    547.499, 603.738, 696.2391, 558.0874, 454.7069, 434.771, 488.2554, 
    465.5451, 480.1592, 528.2115, 662.0346, 767.2975, 774.6315, 505.6811, 
    453.9677, 500.7877, 584.0219, 721.4752, 757.2107, 622.8404, 564.5931, 
    553.7775, 544.0915, 438.6134, 401.1854, 402.1854, 448.803, 413.0183, 
    422.9466, 438.3102, 442.5483, 441.3457,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9.301848, 158.3098, 
    258.9337, 303.8173, 299.6194, 299.056, 279.9115, 262.4927, 294.193, 
    317.6132, 308.028, 282.2506, 265.0864, 268.781, 299.4977, 330.493, 
    349.1855, 376.8177, 421.5884, 502.247, 599.8027, 734.8414, 890.7762, 
    678.5621, 700.035, 677.1342, 600.2327, 509.2974, 559.8538, 608.821, 
    538.714, 488.7658, 668.5876, 1060.59, 1373.92, 1418.137, 819.2729, 
    541.28, 535.3813, 612.2632, 721.4976, 746.7157, 652.4662, 555.7067, 
    576.511, 582.4625, 469.2462, 383.6081, 342.5653, 332.923, 354.656, 
    407.8102, 443.4485, 401.7837, 378.6187,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 86.89892, 228.9686, 
    307.1906, 284.381, 247.07, 238.9294, 245.0831, 292.1502, 321.7906, 
    317.2473, 299.972, 288.464, 279.9789, 285.0193, 296.3184, 328.2048, 
    358.1512, 417.3985, 513.0966, 649.8973, 1018.273, 1282.382, 1139.754, 
    900.5889, 797.8112, 659.6571, 681.5824, 716.9097, 741.9376, 622.0638, 
    551.46, 815.8694, 1147.539, 1486.932, 1523.49, 1029.805, 601.8781, 
    552.1006, 578.9692, 660.6729, 721.0251, 691.4706, 615.808, 579.7531, 
    580.8895, 447.5938, 336.6733, 275.8545, 256.4472, 302.6965, 384.8403, 
    451.3116, 391.0798, 372.3258,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5.010157, 137.2761, 
    246.5296, 275.4832, 286.3332, 281.9478, 285.9474, 335.5515, 358.7326, 
    329.0612, 289.5595, 278.5055, 274.489, 270.4537, 278.7563, 306.5069, 
    345.374, 407.7699, 519.6101, 695.6252, 1020.536, 1431.428, 1296.497, 
    1159.715, 894.8511, 889.3289, 837.659, 898.1722, 824.8221, 688.373, 
    685.1447, 783.9781, 882.051, 899.179, 1132.87, 975.0953, 703.803, 
    579.3523, 556.1559, 602.6837, 672.3351, 701.9514, 668.7778, 612.2599, 
    538.6722, 430.2552, 334.1217, 260.4696, 247.4416, 300.6423, 367.5648, 
    419.1653, 385.3712, 385.5648,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 57.55773, 181.7126, 
    294.1019, 358.642, 376.2969, 381.9689, 378.035, 391.0516, 372.8776, 
    348.465, 324.6873, 307.1947, 273.0872, 273.6699, 274.8869, 275.7082, 
    315.3789, 463.814, 693.0596, 959.1632, 1143.813, 1204.84, 1186.019, 
    1113.179, 1009.146, 981.3286, 895.3462, 765.3611, 644.151, 603.1124, 
    711.8834, 624.4473, 590.9575, 727.5765, 872.574, 675.1846, 577.9081, 
    544.3901, 554.0104, 578.1396, 636.2142, 666.0281, 591.5745, 499.7725, 
    416.1812, 362.9875, 301.6709, 266.8849, 341.4141, 365.0664, 373.7022, 
    355.0049, 393.6327,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7.672453, 76.61076, 
    200.5678, 304.525, 397.0667, 442.379, 428.145, 388.1142, 388.5081, 
    408.9069, 422.5594, 380.0047, 325.1395, 271.7728, 229.48, 221.3898, 
    214.3802, 330.7382, 597.4027, 826.9779, 1010.901, 1106.384, 1267.898, 
    1164.386, 1014.269, 812.2874, 856.5626, 721.2389, 588.0623, 545.859, 
    605.4478, 543.02, 491.1708, 537.3549, 686.0102, 599.1124, 549.1641, 
    530.5813, 510.3197, 549.0093, 608.9304, 682.692, 603.2574, 419.0844, 
    360.2815, 332.0342, 312.2987, 297.1729, 354.3885, 423.995, 364.6626, 
    357.3581, 429.184,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4.492652, 0, 5.913332, 0, 
    9.827749, 122.8932, 239.9646, 413.3958, 469.7688, 442.4698, 411.2574, 
    384.8907, 404.1997, 419.0803, 395.6619, 331.3684, 275.5099, 249.502, 
    270.0858, 300.564, 302.8828, 432.2428, 627.8237, 685.1678, 758.2089, 
    829.3271, 816.4886, 691.1724, 675.4188, 734.3888, 674.1106, 540.9742, 
    509.9907, 540.2866, 512.6861, 438.8988, 428.1956, 510.8031, 492.1108, 
    477.0582, 467.651, 481.3288, 477.3205, 570.1652, 742.3004, 660.6039, 
    434.6603, 307.3639, 286.5654, 295.7912, 296.1364, 355.3662, 457.1753, 
    393.4307, 396.5924, 493.4605,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 38.18091, 177.9759, 
    78.61066, 5.231147, 20.97725, 4.670784, 80.24761, 276.9565, 515.89, 
    480.1449, 420.3515, 475.0774, 450.7651, 429.4347, 397.8179, 353.9267, 
    293.7534, 272.3435, 388.218, 463.1545, 491.6412, 475.5977, 481.5441, 
    496.2309, 455.1932, 510.3101, 537.7867, 541.0651, 539.1157, 607.288, 
    534.366, 475.9772, 458.8337, 508.1748, 500.2999, 470.7975, 373.0616, 
    372.9929, 372.6212, 339.7219, 379.8255, 402.0655, 426.9336, 542.4205, 
    772.5742, 775.2917, 518.3701, 319.2849, 250.5893, 235.3483, 234.3458, 
    282.5884, 389.9496, 389.2494, 430.362, 541.4569,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 42.64318, 0, 0, 0, 14.13362, 
    0, 0, 97.32533, 567.0143, 755.1489, 660.1171, 552.6977, 559.0915, 
    519.6163, 501.7351, 442.0413, 369.866, 317.342, 371.9945, 499.4051, 
    535.2877, 491.8406, 421.9243, 376.5453, 400.5975, 453.606, 510.7452, 
    552.5534, 541.176, 503.5962, 466.0743, 452.3511, 428.7473, 469.4224, 
    558.7114, 555.1274, 362.4989, 286.6256, 277.3649, 257.8876, 279.6031, 
    357.494, 406.6543, 470.3801, 647.2722, 685.0935, 537.283, 372.8993, 
    288.5817, 221.9755, 181.4825, 209.1741, 291.7701, 287.4789, 395.4302, 
    561.2106,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01953389, 0, 0, 0, 
    0, 0, 455.7978, 1051.609, 1211.341, 1040.144, 739.9411, 620.1765, 
    620.5828, 543.5131, 502.523, 425.7497, 412.7139, 442.9023, 449.829, 
    379.7539, 314.4379, 297.9188, 320.5314, 397.3131, 505.9446, 602.7551, 
    619.6101, 569.6279, 539.3142, 520.7625, 497.6906, 523.4991, 613.6224, 
    612.6038, 400.595, 262.5043, 224.5589, 204.1281, 205.329, 279.9945, 
    355.9917, 390.6264, 461.2118, 514.0649, 484.4973, 380.1658, 331.9442, 
    259.4583, 192.7791, 282.2837, 280.4692, 273.8584, 398.2701, 491.5527,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    524.9088, 1227.854, 1514.503, 1593.471, 1283.125, 835.2573, 726.7971, 
    681.4029, 629.7035, 589.2842, 510.3927, 473.1457, 430.4084, 306.1007, 
    237.6619, 228.5278, 244.4046, 284.5834, 374.7751, 497.4753, 605.6686, 
    636.1135, 616.2618, 595.865, 525.5728, 477.7885, 496.7985, 413.9014, 
    286.8343, 221.6673, 207.5997, 165.5916, 149.3675, 196.3652, 251.1849, 
    278.328, 301.5162, 361.5432, 350.5833, 304.2287, 281.5658, 276.7146, 
    189.8026, 362.6567, 363.6728, 247.8723, 372.7149, 441.053,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    109.9336, 398.2949, 940.3243, 1436.861, 1731.173, 1299.493, 1035.062, 
    902.295, 892.6244, 738.1326, 628.37, 557.6457, 490.0444, 346.9488, 
    207.4061, 175.4873, 181.6765, 210.3732, 258.1815, 368.8855, 533.0062, 
    620.7709, 626.9582, 508.8629, 400.888, 363.2095, 333.2734, 270.4286, 
    219.8917, 179.2967, 159.2247, 142.6616, 109.0908, 142.8433, 178.4309, 
    190.0326, 221.8169, 245.1929, 268.4247, 231.8128, 307.9815, 330.6054, 
    275.8257, 397.8697, 359.8254, 219.364, 334.6523, 463.7612,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.06423091, 57.11491, 0, 0, 
    0, 0, 0, 0, 7.836217, 136.0153, 314.1614, 994.2757, 1493.946, 1517.679, 
    1301.398, 1272.304, 1158.99, 1018.497, 845.142, 688.6971, 603.6498, 
    439.0118, 236.4267, 146.054, 144.4927, 163.0123, 225.2119, 349.3079, 
    489.0631, 592.2128, 608.7792, 410.0895, 244.743, 193.4141, 256.4616, 
    227.5397, 197.2503, 107.2875, 83.52959, 68.98138, 80.46129, 115.9747, 
    132.9302, 145.9669, 152.7381, 174.7173, 173.7455, 175.6978, 235.3297, 
    318.201, 276.576, 340.2295, 316.9229, 225.2303, 420.5147, 420.0156,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2.182514, 89.51676, 343.4627, 955.3691, 1260.624, 1151.738, 1138.569, 
    1236.952, 1157.061, 1085.779, 1005.899, 794.526, 562.4872, 299.4979, 
    123.4399, 98.68906, 119.4459, 185.4302, 329.3733, 361.4457, 432.3123, 
    502.7655, 379.1094, 146.3032, 62.53582, 92.53636, 99.53645, 60.84525, 
    11.73829, 14.53334, 21.45396, 50.65263, 84.13147, 89.0048, 93.22248, 
    110.0247, 112.9956, 145.8865, 186.0687, 228.4272, 220.4345, 204.2188, 
    252.7047, 291.9086, 311.514, 407.4745, 196.5356,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 37.47989, 422.1205, 709.343, 683.818, 813.1848, 1012.258, 1090.199, 
    1166.657, 1117.992, 963.0756, 744.8711, 327.3204, 67.59232, 51.20574, 
    51.10489, 136.7648, 215.8003, 145.3761, 67.80409, 186.2934, 218.4242, 
    88.11556, 0.4354767, 0, 0, 0, 0, 34.36349, 48.50853, 69.10825, 73.94706, 
    66.00063, 75.26979, 83.438, 52.38344, 29.00477, 151.119, 204.1204, 
    143.2567, 130.4681, 270.9427, 483.1219, 465.0688, 362.5184, 4.126702,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 17.66449, 261.7532, 151.233, 91.45276, 90.23305, 372.949, 595.9958, 
    811.2404, 1056.335, 1019.892, 820.1436, 449.4274, 159.2536, 109.9366, 
    231.9172, 190.1881, 121.1451, 13.04661, 0.002457884, 0.07684267, 
    1.469449, 0.02487941, 0, 0, 0, 0, 0, 69.92484, 163.3495, 125.5531, 
    119.3953, 127.3019, 150.9474, 169.9525, 115.3876, -54.83441, 78.6655, 
    169.3711, 172.5084, 110.4562, 298.2401, 618.7454, 450.6016, 111.6259, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 18.18774, 198.2974, 24.82351, 0.01659623, 0, 9.641451, 62.01321, 
    362.3916, 663.819, 745.0246, 764.4761, 729.5575, 860.1415, 989.5406, 
    901.2372, 633.0322, 214.5284, 22.94515, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    71.94882, 276.9225, 273.4788, 160.4362, 155.9303, 183.5391, 191.451, 
    188.135, 115.3398, 35.40816, 124.8625, 162.5711, 94.14777, 280.8703, 
    519.7524, 233.8496, 268.5618, 36.8153,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.1127852, 103.1683, 83.84983, 125.6781, 310.4157, 588.7912, 843.4153, 
    526.3326, 1.147217, 0, 31.65186, 188.915, 342.4284, 556.4823, 714.2188, 
    878.2565, 858.4985, 833.0258, 646.3763, 302.5152, 38.86568, 0, 
    0.01003916, 0, 0, 0, 0, 0, 0, 0, 0, 50.22194, 269.6366, 109.4844, 
    37.02338, 59.75043, 26.35164, 79.59688, 104.9516, 76.24226, 67.52459, 
    111.2902, 103.7956, 226.3943, 374.5558, 285.326, 834.7192, 451.0992,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 2.3265, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3.225108, 103.0244, 258.1696, 347.2978, 418.1593, 560.3155, 894.6843, 
    791.2195, 306.0076, 0.8998873, 0, 0, 0, 14.49841, 35.44591, 118.7575, 
    200.4224, 258.1529, 344.5415, 204.937, 28.87837, 0, 0.1383204, 0, 
    2.479101, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01911015, 
    8.849098, 12.94733, 55.8584, 180.516, 374.3842, 761.2708, 606.065,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 15.89997, 14.70358, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 37.67767, 140.6756, 246.9203, 375.567, 456.3772, 603.2179, 
    768.8178, 926.5468, 582.7935, 196.5176, 0, 0.4811277, 0, 0, 0, 0, 0, 0, 
    24.83666, 45.255, 12.15549, 2.415782, 0, 0.09825284, 1.407857, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.6392468, 2.363386, 28.96285, 
    234.0622, 386.0693, 563.9972,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 17.55955, 29.1074, 15.34933, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 10.62364, 190.7695, 391.3156, 404.325, 600.9966, 680.045, 
    704.8675, 862.8046, 749.6393, 130.0502, 3.100419, 5.116066, 6.17757, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.4328433, 76.46776, 242.6619, 291.0963, 5.134037, 
    0, 0, 0, 0, 0, 0, 0, 0, 0.8376673, 0, 0, 0, 0, 0, 0, 0, 0, 0.008186113, 
    0.07604827, 15.87589, 119.0556, 379.1627,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 1.163343, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 255.9357, 568.2272, 791.1302, 892.6254, 903.9981, 891.0063, 
    1059.328, 1098.428, 617.2275, 6.932829, 0.3629374, 65.03675, 7.93887, 0, 
    0, 0, 0.8275996, 112.0045, 17.52323, 0, 0, 57.19586, 246.4086, 451.7093, 
    100.6016, 0.06041526, 0, 0, 0, 0, 0, 0, 0.5732526, 182.9803, 198.6564, 
    161.3975, 11.53954, 0, 0, 0, 0, 0, 0, 0, 0, 0.992954, 173.7827,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 8.585627, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 257.8992, 621.7795, 752.3851, 846.557, 900.2053, 1019.242, 1113.99, 
    880.9015, 529.3146, 159.8383, 6.419941, 0, 0, 0, 0, 0, 0.03464887, 
    317.7343, 145.3232, 0, 0, 0.1035934, 0, 5.595896, 134.9415, 159.4373, 0, 
    0, 0, 0, 0.5597559, 213.3741, 71.13373, 0, 0, 10.51704, 18.63104, 
    3.763446, 0, 0, 0, 0, 0, 0, 0, 0, 34.35713,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1.43994, 381.3143, 748.3234, 941.8181, 893.6531, 933.1523, 1035.22, 
    860.355, 610.6863, 554.7979, 525.4812, 498.002, 75.12685, 0, 0, 0, 0, 
    11.73125, 325.2318, 124.1923, 0, 0, 0, 0, 0, 42.32673, 450.324, 9.972672, 
    0, 0, 34.3005, 62.80934, 603.7728, 328.5521, 8.121914, 9.169447, 
    6.230115, 1.321965, 11.59744, 3.048517, 0, 0, 0, 0, 0, 0, 0, 6.704556,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    30.85074, 297.304, 660.8721, 966.9948, 998.4858, 885.1306, 751.5646, 
    655.1858, 732.1314, 1084.44, 1349.639, 1119.806, 408.8793, 0, 0, 0, 0, 0, 
    140.0299, 7.918328, 0, 0, 0.1702392, 1.991248, 53.83979, 472.2008, 
    346.2012, 2.112901, 0.005206824, 0, 24.37175, 219.4124, 598.756, 
    329.5864, 98.26838, 18.94595, 28.95024, 2.492014, 22.5628, 50.42095, 0, 
    0, 0, 0, 22.81216, 24.65398, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    26.93062, 106.7775, 98.48605, 75.9237, 51.93491, 62.07972, 66.57274, 
    176.725, 422.3495, 479.3473, 519.7673, 215.12, 2.231832, 0.004072465, 
    1.405816, 0.08232938, 0, 495.7819, 40.24272, 0, 7.263184, 112.9553, 
    325.7667, 421.6084, 533.7393, 301.4734, 91.60561, 24.09392, 33.98492, 
    380.9341, 705.0402, 632.1104, 263.1127, 138.8074, 37.80578, 1.129739, 
    35.61073, 95.76726, 325.1597, 511.9413, 832.47, 77.51266, 0, 41.77975, 
    292.1154, 30.66951, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 23.8246, 73.93395, 126.2193, 321.1346, 494.5471, 
    282.6015, 106.8233, 331.644, 202.062, 0, 24.80076, 24.1915, 49.88836, 
    269.6974, 671.1443, 778.3289, 494.5531, 183.3987, 40.72751, 10.41955, 0, 
    92.49084, 767.71, 1000.381, 579.1232, 178.2135, 9.95975, 6.408473, 
    10.95331, 70.58002, 197.3521, 552.4769, 928.8527, 1256.867, 539.4283, 
    47.92098, 154.266, 98.49847, 27.90792, 1.357446 ;

 land_mask =
  0.3764576, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  0.9228161, 0.1739027, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  1, 0.8174675, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  1, 0.5504367, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  1, 0.9481694, 0.1901435, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  1, 1, 0.9983932, 0.2678785, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  1, 1, 1, 0.7833411, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.02900723, 0.3217153, 0.3830353, 
    0.5246126, 0.3472976, 0.1957928, 0.008647686, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 0.9731113, 0.3092794, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0006963735, 0.1754748, 0.4325673, 0.2951554, 
    0.6271494, 0.9393284, 1, 1, 1, 0.9934607, 0.9938456, 0.5638717, 
    0.02968918, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 0.9707108, 0.1046175, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0.06326846, 0.8031307, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 0.9995235, 0.7253351, 0.2813289, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 0.7709347, 0.06251514, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0.4201411, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 0.9849455, 0.1556062, 0.003983508, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 0.5608934, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.9381469, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.9549282, 0.5933414, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 0.8828677, 0.06657699, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0.6793007, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 0.8384063, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 0.669156, 0.0125583, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.1381188, 0.9697084, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 0.9104351, 0.2647975, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 0.04201834, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.00166111, 0.5541363, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 0.4645965, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 0.04201056, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.0307463, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 0.6972274, 0.5714607, 0.539219,
  1, 1, 1, 1, 1, 1, 1, 1, 0.04200291, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.2669835, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 0.5898379, 0.00854887, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.07485126, 0.9193581, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 0.4414221, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.0006397907, 0.4717199, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9447742, 0.2459255, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.1592281, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9522441, 0.693058, 0.077351, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.1598931, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.7353352, 0.09539028, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.6433973, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 0.6314353,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9975816, 0.8410712, 0.3690621, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.6869012, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9971337, 0.3079584, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.6868731, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.6658256, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.6868458, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9175764, 0.2185544, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.1822212, 0.9689022, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.7709059, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.651095, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9019616, 0.1664711, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.203948, 0.9547996, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.3274225, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.6748101, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.8615925, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.2362749, 0.9623896, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.8665756, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.7315421, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.8665628, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.7754121, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.8665506, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.2965498, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.8665391, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0509539, 0.8103296, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9383764, 0.2196166, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.7782937, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9603246, 
    0.0640404, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.2410026, 0.8761689, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.6294757, 
    0.007487927, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.7360525, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.266498, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.5350724, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9991729, 
    0.4061707, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.09449254, 0.8377889, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.9303989, 0.1264541, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.182272, 0.9179717, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.1799683, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.1560873, 0.8999666, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.3121897, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.4015228, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.159612, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.01152876, 0.7892212, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9283816, 
    0.6226964, 0.5535366, 0.06422334, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0.2964121, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.7704774, 
    0.05751295, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.03438287, 0.7932302, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9993793, 0.8113894, 0.6826136, 
    0.8702582, 0.5128348, 0.08204572, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.008766619, 0.6232422, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.7633693, 0.1774785, 0.2040459, 0, 0, 
    0.0009010995, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.6049436, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 0.9406916, 0.9853109, 0.9229649, 0.3723707, 
    0.03303384, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0.2605378, 0.9595606, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 0.9745548, 0.8413171, 0.115013, 0.1830149, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.3241267, 0.9822798, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 0.5268455, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.8645887, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 0.2353382, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.847726, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1,
  1, 1, 1, 1, 1, 0.7867104, 0.09881871, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.3535399, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 0.2738446, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1326434, 
    0.587546, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 0.01733101, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.01603992, 0.4454439, 0.6442813, 0.3830209, 0.05625193, 0, 
    0.03530673, 0.2579472, 0.08800853, 0, 0, 0, 0, 0, 0, 0.5546407, 
    0.6381541, 0.4571692, 0.7593831, 0.9919729, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 0.957557, 0.3666932, 0.001214215, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.06446161, 0.8062138, 1, 1, 1, 0.9404332, 0.9032256, 
    0.9204367, 1, 0.9587651, 0.5515207, 0.2075914, 0.002314975, 0, 0, 
    0.1886965, 0.9459232, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 0.9558364, 0.4539385, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.254573, 0.9151666, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.7619722, 
    0.6994123, 0.5289772, 0.9312455, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0.9320562, 0.7091275, 0.1623458, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.02540474, 0.619023, 0.9725087, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0.1557076, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.3710184, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.03056264, 
    0.5956897, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1148876, 0.5937533, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.07622165, 0.6823812, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.3449733, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.3805372, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.753692, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.3588129, 0.9958816, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.7856891, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.7856846, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01859863, 0.3884055, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.2158899, 0.9551845, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.3530129, 0.9508796, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.7544317, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.2654112, 0.9811226, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.6945245, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.07710309, 0.863272, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.6369579, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1824975, 
    0.7033954, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1683426, 
    0.8958945, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1531393, 
    0.5754542, 0.9937046, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.5226966, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.7708154, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.5950658, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.07487938, 0.8179564, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.03862339, 0.4152967, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 0.8500615, 0.946259, 0.884431, 0.7472318, 0.7092528, 
    0.9718166, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9999945, 
    0.4919434,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.004841657, 0.4270654, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 0.8776839, 0.7527315, 0.9694611, 0.8234424, 0.05545996, 0.01451342, 
    0.0766992, 0, 0, 0.7712654, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.740279, 0.0665665,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.1420659, 0.6810132, 0.2436509, 0.1621065, 0.2339793, 0.6901079, 
    0.9708213, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.8266005, 0.4517564, 0.04483075, 
    0.03248953, 0.1924889, 0.01307053, 0, 0, 0, 0, 0, 0.7712539, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9643438, 0.4936993, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.357605, 0.4481737, 0.01432, 0, 0, 0, 0.2996151, 0.8592404, 
    0.9996577, 1, 1, 1, 1, 1, 1, 1, 0.9999822, 0.3695327, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.1985431, 0.891767, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.4674213, 0.2888203, 0.163148,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.02609481, 0.6882609, 0.6668625, 0.8689135, 1, 0.997447, 0.9480262, 
    0.6412953, 0, 0, 0, 0.2262365, 0.6555864, 0.7921475, 0.9380791, 1, 1, 1, 
    1, 1, 0.6710668, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0618545, 0.7309781, 
    0.5937635, 0.3276973, 0.5878043, 0.4755114, 0.293394, 0.649609, 0.670538, 
    0.8472934, 1, 1, 1, 1, 0.942656, 0.977885, 0.3617498,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.03747177, 1, 1, 1, 1, 1, 1, 0.9728559, 0.7016522, 0.05877807, 0, 0, 0, 
    0, 0.0007180843, 0.2887189, 0.7476513, 0.6832384, 1, 1, 0.419323, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.009167003, 0, 0, 0, 0, 0, 0, 0.002281133, 
    0.2401035, 0.8190355, 1, 1, 1, 1, 0.6542072,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.4350484, 1, 1, 1, 1, 1, 1, 1, 1, 0.5818211, 0, 0, 0, 0, 0, 0, 0, 
    0.001013471, 0.1183226, 0.3208605, 0.3338135, 0, 0, 0, 0.006452882, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1757967, 0.6191416, 
    0.6542448, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.08844708, 1, 1, 1, 1, 1, 1, 1, 1, 0.4442382, 0, 0, 0.02307724, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.3639905, 0.6390771, 0.7038295, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.03658982, 0.4823922, 0.9029201, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.02019954, 0.7953823, 1, 1, 1, 1, 1, 1, 1, 0.8110214, 0.06406885, 0, 
    0.390024, 0.05420401, 0, 0, 0, 0, 0.4077412, 0.04842471, 0, 0, 0.1416207, 
    0.3410814, 0.6977392, 0.1285015, 0, 0, 0, 0, 0, 0, 0, 0, 0.1522885, 
    0.5140895, 0.258808, 0.0008218849, 0, 0, 0, 0, 0, 0, 0, 0, 0.02715651, 
    0.7257767,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.03747227, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.726593, 0.04869777, 0, 0, 0, 0, 
    0, 0, 0.8814211, 0.1349703, 0, 0, 0, 0, 0.01583155, 0.1170755, 0.247405, 
    0, 0, 0, 0, 0.0326486, 0.3860433, 0.1965477, 0, 0.00835224, 0.2670313, 
    0.005355601, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.4019571,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0374724, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.8357671, 0.2085238, 0, 0, 0, 
    0, 0, 0.809296, 0.1349555, 0, 0, 0, 0, 0, 0.09953156, 0.670812, 0, 0, 0, 
    0, 0.1109447, 1, 0.6344974, 0.005974696, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.2480379, 0.8815156, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.6203845, 0, 0, 0, 
    0, 0, 0.2954375, 0.07066895, 0, 0, 0, 0, 0.1317861, 0.6645802, 0.4592906, 
    0, 0.006340416, 0, 0.1393674, 0.7857525, 1, 1, 0.3672985, 0, 0, 0, 0, 
    0.000822613, 0.00348749, 0, 0, 0, 0.04631038, 0.06669453, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.14503, 0.4055507, 0.2551057, 0.3028015, 0.3623243, 0.4336107, 
    0.2924458, 0.9094968, 1, 1, 1, 0.7378889, 0.03122145, 0.001574896, 0, 0, 
    0, 0.7633188, 0.1349258, 0, 0.1208249, 0.5835989, 0.783038, 0.9167218, 1, 
    0.7098413, 0.4056285, 0.2833857, 0.1567454, 0.7330076, 1, 1, 0.9505261, 
    0.4874083, 0, 0, 0, 0.3619807, 0.7769179, 0.7792631, 0.6483424, 
    0.1295194, 0, 0.04274155, 0.6756219, 0.06986691, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.5567488, 1, 1, 1, 1, 0.7617028, 0.7580242, 
    0.8640846, 0.2590115, 0.01124508, 0.1238442, 0.05218257, 0.3791888, 
    0.9209204, 1, 1, 0.8919879, 0.9454092, 0.483057, 0.08077005, 0, 
    0.3203594, 1, 1, 1, 0.5728929, 0.0002312251, 0, 0, 0.5069734, 0.9029012, 
    1, 1, 1, 0.7427915, 0.221187, 0.2803968, 0.3342389, 0.03174093, 0 ;

 zsurf =
  8.54475, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  110.6839, 9.015973, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  118.8102, 18.13202, 0.007421071, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  130.705, 39.06387, 3.106806, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  141.0809, 84.24564, 11.19796, 0.4508977, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0,
  165.9822, 184.6116, 106.8482, 7.492514, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.08320683, 3.271346, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  180.4211, 249.8835, 220.8967, 76.21671, 1.021369, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    21.94272, 34.81591, 74.42256, 66.43814, 11.87937, 0, 0, 0, 0, 0, 0, 0, 0,
  149.0657, 196.1795, 177.1756, 126.4176, 11.39334, 0.5445582, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2.201014, 10.06274, 
    26.85098, 48.46229, 196.196, 446.1897, 398.605, 448.8601, 587.3398, 
    619.0617, 478.8845, 191.0291, 9.431361, 0, 0, 0, 0, 0, 0,
  247.4764, 260.0786, 196.9956, 132.1378, 48.361, 5.852092, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6.821061, 227.5061, 
    341.0564, 416.8428, 546.1491, 760.7002, 800.6117, 811.9203, 918.2296, 
    1199.078, 1194.457, 1065.196, 779.4019, 539.7784, 68.59048, 0, 0, 0, 0, 0,
  254.4188, 378.3603, 367.6226, 301.4343, 162.2049, 108.9995, 0.9085217, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8.392265, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    84.11958, 610.6379, 784.4166, 873.3272, 803.2366, 954.6566, 1133.667, 
    1193.683, 1333.627, 1518.089, 1657.062, 1719.367, 1548.189, 1097.09, 
    488.3766, 19.6729, 0, 0, 0, 0,
  282.803, 388.1694, 501.5489, 557.1978, 613.9719, 624.3671, 154.6011, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.850073, 136.7001, 
    621.1481, 1059.969, 1205.403, 1271.604, 1289.321, 1373.992, 1468.906, 
    1399.973, 1501.777, 1674.687, 2147.529, 2156.621, 1497.179, 907.9773, 
    341.0655, 33.16307, 0, 0, 0,
  281.039, 423.6907, 485.7559, 651.8676, 783.3052, 889.3768, 610.0162, 
    16.97377, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    129.3114, 660.4066, 997.0892, 1271.035, 1259.05, 1269.307, 1282.922, 
    1357.486, 1418.984, 1464.053, 1694.626, 2161.078, 2172.453, 1467.212, 
    1030.81, 612.332, 164.4304, 1.996331, 0, 0,
  322.6488, 427.8226, 549.0103, 681.7765, 829.639, 1022.879, 837.8648, 
    305.3638, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    9.138049, 280.6169, 659.5826, 1002.684, 1031.975, 1099.151, 1099.102, 
    1133.435, 1221.698, 1317.967, 1415.099, 1513.935, 1787.441, 1850.336, 
    1464.755, 1240.903, 696.9532, 172.8423, 13.54243, 0, 0,
  246.0376, 453.1236, 631.008, 871.3788, 1047.864, 932.1511, 816.0308, 
    317.9274, 6.631444, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    150.0291, 674.2753, 908.9203, 930.3144, 938.6702, 1006.137, 1124.25, 
    1170.841, 1154.932, 1264.449, 1330.767, 1451.47, 1585.219, 1689.979, 
    1656.847, 1377.684, 685.7067, 148.093, 7.893209, 0, 0,
  302.9081, 427.2077, 600.2842, 822.6921, 987.5324, 917.3104, 668.1157, 
    303.2888, 0.4759156, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.05529097, 404.3319, 849.9101, 942.0059, 899.2049, 892.3331, 1045.702, 
    1259.788, 1338.622, 1238.361, 1260.895, 1324.21, 1411.141, 1544.977, 
    1598.17, 1706.571, 1414.926, 652.4966, 175.4458, 20.1155, 25.00171, 
    36.41872,
  304.3976, 367.4553, 507.5162, 723.1177, 889.1189, 890.2856, 860.1849, 
    487.2796, 0.9306844, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    48.47385, 456.4773, 788.9446, 784.0788, 797.9801, 888.491, 1040.636, 
    1257.102, 1379.351, 1308.995, 1358.369, 1450.252, 1468.341, 1489.487, 
    1519.486, 1585.82, 1321.473, 545.1862, 138.8361, 40.63335, 49.9632, 
    84.77402,
  357.9227, 326.5664, 409.4615, 533.1976, 722.5844, 805.3265, 892.149, 
    651.6109, 85.95663, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6.497938, 272.2702, 615.2929, 908.9059, 917.061, 841.0509, 900.0991, 
    989.4551, 1097.285, 1229.295, 1245.714, 1381.851, 1374.066, 1291.548, 
    1248.401, 1166.31, 1273.148, 967.5308, 443.7959, 159.7697, 64.36124, 
    74.43269, 110.2169,
  374.3119, 313.8954, 345.6318, 445.4458, 583.0211, 721.8264, 795.6353, 
    683.6541, 309.0318, 22.92986, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 217.3822, 804.5779, 921.5053, 1073.372, 1032.455, 914.3887, 915.9861, 
    975.9174, 1025.77, 1091.464, 1183.756, 1203.829, 1146.519, 1118.986, 
    1206.85, 1186.365, 1061.127, 699.5498, 315.4096, 174.5182, 91.69196, 
    117.5326, 129.1317,
  384.2018, 316.835, 329.2943, 348.3972, 449.1535, 490.7008, 580.1392, 
    682.83, 561.0168, 450.0525, 74.4604, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 1.625334, 529.3156, 1179.003, 1083.251, 1046.369, 1010.433, 952.2749, 
    974.9957, 1008.044, 1025.375, 1088.216, 1136.371, 1137.306, 977.9841, 
    966.8591, 1095.862, 1080.748, 967.8829, 583.6017, 349.6461, 208.4064, 
    122.2884, 137.5921, 124.6154,
  425.9325, 402.693, 356.9512, 342.1429, 387.3358, 451.6554, 543.8193, 
    598.1646, 671.4254, 663.9327, 658.8842, 342.5872, 1.323529, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 55.75727, 723.3252, 1345.097, 1208.163, 1096.152, 
    1057.105, 1042.026, 1052.195, 1075.99, 1085.4, 1083.792, 1107.45, 
    1089.932, 1003.74, 908.7562, 881.2886, 806.4973, 725.7192, 521.3715, 
    374.6654, 268.3831, 172.0694, 131.0901, 57.53464,
  461.6035, 467.3536, 394.1595, 343.5833, 356.553, 412.9582, 456.8489, 
    546.8406, 586.7995, 714.7881, 969.0544, 855.0431, 500.8872, 32.52318, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 123.6441, 855.6476, 1413.006, 1269.892, 
    1172.559, 1156.56, 1149.75, 1151.305, 1144.381, 1103.469, 1061.514, 
    1045.96, 1102.312, 1112.108, 971.346, 808.2177, 695.4062, 630.5798, 
    525.356, 437.357, 384.1834, 350.2086, 123.1665, 31.22814,
  464.4684, 508.0797, 455.048, 373.7856, 366.4037, 387.9864, 443.3236, 
    495.3125, 589.3275, 739.6755, 988.6879, 1060.314, 904.9486, 528.0706, 
    225.8937, 27.69355, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 174.664, 879.7312, 1444.223, 
    1357.686, 1256.545, 1275.17, 1242.061, 1206.494, 1137.42, 1064.367, 
    1009.382, 1009.102, 1074.426, 1101.382, 1013.848, 935.0889, 872.3643, 
    823.5287, 742.5305, 702.767, 638.2717, 610.8529, 236.0903, 19.05215,
  377.5986, 476.2537, 554.4959, 498.4242, 421.1341, 410.7194, 460.7333, 
    508.1182, 604.0519, 780.8995, 940.6996, 912.0196, 1031.078, 860.0245, 
    593.0319, 288.8579, 12.86605, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 211.1246, 927.424, 
    1489.004, 1561.025, 1444.746, 1376.06, 1280.973, 1179.52, 1098.244, 
    1019.69, 975.9384, 963.2079, 978.0944, 1029.098, 1103.491, 1163.96, 
    1175.215, 1136.579, 1103.248, 1014.715, 943.465, 803.7495, 369.8148, 
    113.7734,
  332.751, 472.4073, 685.3926, 635.038, 517.4619, 464.7151, 489.6293, 
    589.0376, 704.1102, 888.3381, 946.3566, 843.2612, 937.7106, 952.2573, 
    593.1406, 408.6372, 87.12373, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 274.805, 948.42, 
    1506.014, 1601.052, 1578.846, 1456.921, 1284.965, 1163.84, 1079.576, 
    1015.096, 961.92, 924.3301, 919.1673, 969.1686, 1080.93, 1206.276, 
    1290.624, 1303.251, 1316.85, 1354.376, 1136.7, 970.1143, 487.621, 182.6047,
  386.6328, 599.5612, 743.3576, 737.4709, 670.9242, 536.273, 553.6517, 
    674.8468, 801.8613, 965.2466, 953.0202, 781.4857, 825.5333, 884.1866, 
    743.7918, 650.3617, 509.5243, 47.25615, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 34.19665, 536.6432, 
    1112.04, 1443.481, 1515.864, 1440.972, 1356.049, 1192.005, 1062.608, 
    976.4597, 953.9917, 942.6937, 942.3792, 969.4203, 966.9082, 1031.604, 
    1100.836, 1155.753, 1179.703, 1365.894, 1379.681, 1287.486, 922.5301, 
    544.6479, 214.8122,
  407.2789, 556.476, 691.2809, 737.9501, 749.3389, 662.7368, 563.8776, 
    667.7236, 775.2804, 860.3702, 857.4185, 735.3098, 719.4968, 858.9086, 
    655.9019, 560.5863, 441.2978, 138.1514, 0.004807308, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 245.0765, 
    740.5414, 1216.22, 1399.232, 1428.595, 1324.44, 1244.887, 1171.623, 
    1058.757, 978.5461, 948.2759, 945.5349, 979.3757, 1012.527, 980.8537, 
    912.5103, 983.9648, 1005.987, 1126.251, 1280.425, 1263.255, 944.915, 
    620.7706, 330.2798, 198.4007,
  485.9347, 536.7831, 520.842, 574.1156, 628.2961, 593.3192, 671.6805, 
    760.3802, 792.5333, 809.5409, 713.7068, 694.2451, 762.8157, 893.8396, 
    750.4239, 489.7271, 319.0528, 122.3887, 1.660121, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.1749505, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 36.20846, 
    639.6878, 1064.495, 1200.584, 1345.762, 1339.131, 1276.558, 1206.219, 
    1145.992, 1077.639, 997.5162, 966.3801, 956.3568, 970.2714, 1008.335, 
    951.059, 828.9758, 706.606, 863.0428, 1080.806, 1123.896, 920.291, 
    656.9827, 373.7796, 334.5416, 526.0103,
  571.2805, 576.3853, 467.4599, 411.0854, 392.3285, 505.7308, 722.9926, 
    869.4109, 931.8525, 811.3553, 662.9765, 604.0966, 688.219, 858.3245, 
    825.9299, 572.1747, 408.3769, 146.4941, 9.387668, 0.001074584, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    273.4626, 965.0869, 1142.758, 1166.024, 1121.857, 1187.254, 1166.343, 
    1151.341, 1121.571, 1066.005, 1020.396, 995.9119, 976.3922, 999.8099, 
    1080.855, 1153.143, 949.2833, 796.8798, 704.9807, 751.8674, 635.2756, 
    537.6038, 460.5406, 432.7109, 753.7834, 783.1511,
  541.8253, 527.6813, 442.9381, 349.75, 282.5704, 372.3629, 647.7617, 
    839.8668, 941.1125, 907.2533, 705.0693, 633.6419, 637.7145, 768.287, 
    809.7827, 674.5598, 493.8878, 279.3312, 44.60109, 0.003030813, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    59.35226, 753.0102, 1128.37, 1213.516, 1102.814, 1106.985, 1138.11, 
    1148.302, 1144.664, 1119.719, 1075.693, 1028.648, 1007.681, 1040.419, 
    1070.42, 1085.326, 1113.797, 1101.634, 964.3666, 826.3594, 688.6269, 
    581.0179, 749.9571, 747.4507, 813.9899, 1027.863, 909.4127,
  451.7546, 465.3449, 395.6716, 335.8462, 247.0956, 298.3383, 466.0626, 
    661.6984, 813.6958, 827.1074, 757.3602, 671.0699, 631.3232, 636.7422, 
    748.9434, 753.5067, 653.6973, 358.9735, 111.3765, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 237.6711, 881.6313, 
    1209.199, 1111.17, 1116.662, 1148.323, 1170.288, 1177.596, 1179.032, 
    1162.061, 1096.823, 1040.075, 1027.026, 1072.69, 1144.079, 1132.332, 
    1099.773, 1094.171, 1114.551, 970.8142, 812.7686, 713.1152, 878.1364, 
    977.2021, 1026.251, 1069.996, 736.0057,
  391.2837, 370.3196, 366.6443, 340.5762, 263.041, 234.9373, 359.7917, 
    485.6016, 684.4538, 736.9855, 740.4536, 781.7585, 658.1667, 565.2335, 
    713.5017, 808.0051, 692.545, 472.7854, 120.2969, 0.03788849, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 152.0637, 
    745.3533, 1129.647, 1190.232, 1165.257, 1217.449, 1233.613, 1242.039, 
    1225.1, 1190.186, 1129.522, 1051.2, 1039.217, 1088.383, 1158.137, 
    1160.562, 1157.639, 1146.778, 1176.388, 1196.262, 1103.755, 939.6448, 
    773.607, 786.1696, 1066.588, 999.4681, 658.9298,
  343.9839, 329.1209, 326.8227, 338.2211, 268.4422, 231.5902, 273.1661, 
    411.1793, 556.3333, 647.4001, 724.2601, 776.667, 679.067, 508.2994, 
    620.4402, 716.1536, 666.8013, 484.4005, 195.8266, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 49.35054, 549.8828, 
    1179.242, 1286.947, 1285.081, 1347.293, 1373.125, 1342.854, 1282.255, 
    1234.189, 1156.042, 1075.134, 1044.677, 1093.778, 1146.635, 1190.949, 
    1194.665, 1203.338, 1225.234, 1270.81, 1379.499, 1236.873, 994.0289, 
    744.1392, 1000.295, 1032.345, 591.7537,
  341.9223, 323.5297, 312.363, 327.7422, 256.121, 211.4899, 232.2774, 
    293.0904, 373.0227, 483.3326, 649.4127, 771.75, 673.2164, 571.9428, 
    626.7587, 791.145, 642.7789, 521.3182, 201.4202, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 3.703202, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10.91209, 
    566.6647, 1165.319, 1443.802, 1442.337, 1513.629, 1471.694, 1443.57, 
    1354.923, 1276.675, 1185.226, 1087.362, 1080.905, 1145.881, 1175.568, 
    1221.021, 1282.013, 1268.265, 1230.614, 1228.024, 1211.29, 1307.737, 
    1161.229, 873.0657, 933.2297, 1159.808, 670.6091,
  346.7993, 338.6057, 314.9171, 289.7007, 236.9087, 190.2888, 202.9013, 
    268.8091, 310.8858, 411.589, 656.1295, 740.801, 656.6727, 541.4875, 
    678.8455, 853.9406, 730.4851, 459.3751, 220.1203, 13.96118, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    413.7036, 981.3401, 1411.613, 1624.979, 1620.908, 1479.521, 1444.335, 
    1392.403, 1297.059, 1161.221, 1098.89, 1153.009, 1254.525, 1302.453, 
    1335.512, 1364.571, 1280.526, 1204.677, 1180.655, 1170.281, 1240.504, 
    1336.752, 1084.095, 1070.497, 1113.52, 930.3657,
  373.4141, 339.6274, 318.1039, 291.9559, 260.7186, 191.6193, 197.949, 
    276.8808, 356.4713, 444.8528, 671.9672, 707.4572, 541.8743, 515.196, 
    593.6595, 844.5728, 740.3514, 450.5794, 236.8895, 126.5775, 12.02609, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    74.79279, 582.2818, 1387.929, 1653.479, 1656.323, 1452.037, 1384.894, 
    1380.74, 1263.157, 1129.277, 1087.819, 1140.283, 1291.528, 1349.267, 
    1427.148, 1380.747, 1211.18, 1182.415, 1173.129, 1242.567, 1253.907, 
    1328.973, 1235.93, 1102.579, 1212.149, 1188.651,
  411.907, 359.5694, 312.9021, 316.0843, 319.7564, 228.2056, 193.8342, 
    296.6815, 321.6121, 390.0383, 586.1972, 616.8071, 522.6686, 497.1555, 
    514.1055, 625.6185, 709.9496, 500.6991, 322.1615, 233.313, 73.02024, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 251.8302, 1240.724, 1602.32, 1519.831, 1331.846, 1307.905, 1319.815, 
    1247.846, 1123.754, 1088.791, 1091.119, 1166.166, 1236.438, 1262.825, 
    1296.363, 1122.022, 1172.453, 1197.705, 1311.24, 1400.86, 1405.443, 
    1374.509, 1337.278, 1486.886, 1500.223,
  361.1769, 319.2283, 308.7516, 344.1496, 351.8325, 252.6501, 205.3004, 
    264.0542, 284.5062, 319.0981, 459.6907, 492.8576, 454.6547, 494.1764, 
    467.236, 499.1732, 633.0408, 550.3798, 449.2036, 364.1278, 174.6403, 
    28.89057, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 104.2696, 1010.841, 1362.054, 1315.101, 1130.426, 1149.357, 
    1245.088, 1169.575, 1095.747, 1041.157, 1027.792, 1023.939, 991.415, 
    1043.899, 1006.476, 1261.374, 1189.962, 1103.186, 1205.096, 1273.994, 
    1571.499, 1265.122, 1354.616, 1342.277, 1499.963,
  288.3837, 296.7624, 328.1481, 349.2853, 354.0044, 300.8336, 209.8271, 
    242.339, 257.6059, 315.6365, 438.6422, 454.057, 469.7331, 499.5292, 
    472.8086, 418.0537, 492.4049, 451.988, 414.6512, 387.9483, 298.7437, 
    224.9868, 30.84828, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.8451669, 71.35338, 642.9059, 1073.645, 1063.941, 
    943.9172, 1026.204, 1114.221, 1073.748, 1012.559, 1027.82, 1014.382, 
    1057.285, 1027.442, 823.2462, 941.8942, 1091.702, 1226.689, 1104.525, 
    1242.194, 1126.849, 1339.002, 1262.845, 1232.307, 1363.345, 1223.546,
  260.1389, 284.7289, 287.6657, 321.2379, 323.3841, 321.9951, 239.3829, 
    211.8097, 231.2988, 276.1485, 389.8618, 400.1599, 419.2465, 413.5182, 
    379.3967, 365.7533, 402.7262, 476.0164, 436.6118, 442.7455, 523.3729, 
    513.603, 263.7818, 2.99741, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 6.84726, 127.0682, 564.7839, 1027.651, 923.8217, 
    809.4365, 946.3239, 1098.568, 971.295, 901.8392, 924.174, 968.075, 
    986.755, 1009.199, 898.538, 673.96, 868.1624, 893.8102, 1322.028, 
    1317.703, 1118.277, 1254.662, 1102.685, 1225.965, 1365.095, 1100.581,
  256.0101, 258.5121, 265.4595, 271.6456, 281.9239, 339.2019, 239.4398, 
    201.6286, 231.9184, 272.3331, 346.6201, 365.2863, 335.9691, 301.0338, 
    258.306, 271.6318, 450.0833, 557.5646, 531.2784, 522.4316, 549.2473, 
    622.1465, 329.0093, 25.54767, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 6.427928, 262.789, 692.8567, 1032.231, 824.3097, 
    711.4518, 954.0336, 994.9745, 852.847, 765.702, 840.2001, 873.9611, 
    851.5475, 920.1156, 891.8646, 743.049, 630.5678, 807.291, 1051.364, 
    1174.423, 1034.36, 1105.102, 1130.744, 1221.451, 1312.698, 1236.457,
  244.8726, 235.7898, 238.6499, 250.9584, 264.177, 304.3681, 231.7038, 
    171.5492, 194.0964, 237.4297, 322.8626, 324.8877, 315.0707, 258.6005, 
    236.6363, 277.2534, 457.8071, 528.7694, 405.2236, 342.8656, 385.32, 
    442.8686, 295.1935, 24.17916, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 1.293201, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 52.95097, 347.3517, 720.2449, 929.5432, 
    735.391, 780.5626, 910.9541, 885.9318, 687.3369, 662.2593, 723.8735, 
    755.4806, 723.0743, 769.8126, 788.1163, 702.8589, 630.3057, 768.6213, 
    1059.849, 972.3868, 1188.259, 1177.481, 1121.192, 1184.726, 1279.616, 
    1302.242,
  235.042, 217.7554, 200.0201, 218.5201, 210.6107, 214.8637, 159.0711, 
    132.8887, 194.6062, 222.7486, 255.3079, 243.1668, 189.8971, 189.5496, 
    151.8132, 254.9043, 441.0879, 450.9707, 312.1183, 209.6811, 199.2862, 
    258.3366, 160.7645, 4.592148, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.1700515, 92.22056, 366.6779, 594.3502, 777.5218, 
    693.3395, 719.6742, 801.9887, 715.3484, 599.9813, 555.8511, 606.0909, 
    628.077, 622.9703, 659.368, 666.463, 613.6947, 660.4321, 819.1418, 
    1024.8, 1005.07, 1167.154, 1107.55, 1131.997, 1173.377, 1208.152, 1350.651,
  196.7365, 204.5998, 198.4898, 193.5049, 169.7109, 154.1599, 121.315, 
    140.5267, 197.9303, 241.7397, 228.9246, 149.1499, 105.5863, 101.0614, 
    123.9294, 166.2768, 433.4229, 365.3992, 271.7154, 133.414, 51.558, 
    55.21501, 35.0076, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 13.58836, 185.3467, 334.9186, 518.5123, 624.0504, 611.5664, 
    573.1268, 551.8474, 545.7886, 508.7069, 509.3336, 518.7409, 552.8677, 
    565.2957, 587.2665, 552.8708, 585.5536, 619.3701, 901.4293, 1212.324, 
    1221.37, 1192.156, 1120.597, 1169.473, 1176.514, 1126.01, 1376.636,
  146.6925, 179.7951, 169.8683, 144.5109, 115.9851, 100.912, 77.22723, 
    96.99864, 139.7948, 160.3108, 134.8792, 69.91695, 26.29307, 64.91444, 
    76.29048, 164.2859, 290.0237, 281.2162, 184.3736, 70.43913, 2.701435, 0, 
    0, 0, 0, 0.09234287, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 2.41791, 93.65132, 238.9857, 412.0441, 452.2166, 553.3406, 506.5167, 
    421.6122, 392.6665, 425.7772, 440.7444, 462.4359, 492.6555, 517.598, 
    531.2183, 527.7665, 529.114, 571.4398, 752.8386, 1117.882, 1654.942, 
    1618.519, 1398.75, 1202.588, 1191.508, 1195.801, 1221.172, 1415.927,
  69.31319, 104.212, 110.316, 83.84324, 63.33185, 52.58361, 41.60804, 
    45.76586, 76.87368, 101.9827, 93.67348, 33.04323, 20.12624, 46.1826, 
    54.88905, 34.84738, 115.9459, 49.21751, 40.83882, 0.5943004, 0, 0, 0, 0, 
    0, 0.0057942, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.398386, 
    119.9112, 199.3601, 411.994, 476.3767, 578.0508, 529.0004, 436.2539, 
    335.8598, 335.8933, 358.957, 401.7341, 439.7245, 481.3549, 499.7074, 
    519.8088, 515.3641, 502.7769, 560.4839, 723.5606, 1163.4, 1705.951, 
    1771.096, 1455.29, 1286.019, 1198.102, 1179.159, 1260.96, 1461.374,
  79.25274, 98.79363, 46.67113, 25.34361, 28.43618, 24.51583, 16.18622, 
    19.50146, 37.39209, 67.61229, 56.61288, 32.74178, 14.21986, 3.174914, 
    2.647948, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.01747818, 46.90157, 207.9118, 460.4455, 514.9199, 
    602.9887, 590.7431, 513.9005, 364.6547, 319.0529, 315.5271, 335.9451, 
    373.1736, 425.5178, 449.45, 464.8029, 490.2738, 503.6892, 494.0532, 
    586.5953, 751.3316, 1115.167, 1723.364, 1792.263, 1481.577, 1256.694, 
    1160.092, 1138.162, 1189.935, 1531.006,
  304.3052, 225.9071, 146.4976, 49.22798, 14.06787, 15.70426, 14.31254, 
    10.55259, 21.65571, 34.42345, 26.47721, 10.16362, 1.715719, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.3261773, 0, 0, 5.140869, 66.8336, 316.336, 486.2376, 557.2535, 
    481.0815, 482.611, 398.9484, 317.3685, 310.7681, 323.2128, 329.6191, 
    362.9882, 389.781, 416.3743, 421.8354, 456.8871, 480.976, 483.8488, 
    540.1299, 714.4539, 990.8341, 1670.664, 1620.258, 1494.627, 1232.962, 
    1134.55, 1134, 1203.068, 1431.174,
  377.3476, 300.3462, 179.3239, 123.5264, 29.18042, 8.49296, 10.41877, 
    2.594529, 2.675612, 3.391332, 0.1138654, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.007269558, 0, 
    7.853471, 62.3085, 274.8862, 413.5488, 423.2161, 435.7926, 444.4748, 
    361.6428, 308.9561, 319.7975, 321.1809, 340.5662, 354.3437, 378.4564, 
    404.6211, 438.1272, 444.1309, 457.4094, 472.3898, 582.7078, 713.5034, 
    965.1596, 1325.418, 1513.297, 1287.996, 1268.213, 1155.886, 1135.109, 
    1137.983, 1441.737,
  397.6618, 290.1455, 262.0854, 164.1737, 72.91979, 9.641136, 3.297817, 
    0.002408294, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24.52353, 0, 1.134986, 131.7988, 
    413.9996, 487.4259, 485.74, 514.1754, 483.7487, 398.7583, 334.6064, 
    318.3876, 329.1971, 343.4026, 364.3184, 386.8412, 433.8055, 462.0353, 
    443.1543, 453.2259, 475.2897, 560.871, 675.3644, 778.7476, 1195.336, 
    1219.456, 1293.797, 1255.619, 1167.165, 1128.763, 1127.737, 1605.608,
  359.7442, 322.1634, 256.7101, 190.8573, 99.29717, 20.20619, 2.261762, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 1.042433, 1.061284, 0.06026918, 221.4693, 588.1027, 
    609.5046, 567.6266, 539.7374, 519.683, 443.9848, 375.9164, 330.9009, 
    328.2888, 345.5885, 367.2719, 396.1122, 425.6252, 436.9988, 445.1413, 
    455.4268, 478.2379, 538.37, 618.6725, 704.752, 879.9337, 1044.206, 
    1143.218, 1000.543, 1114.351, 1055.759, 1244.916, 1644.584,
  339.5918, 283.2596, 244.217, 182.1556, 115.8238, 16.9204, 1.281723, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 118.1892, 542.7286, 664.8825, 616.7386, 
    595.4612, 551.9771, 495.2496, 416.2375, 373.1087, 345.3355, 352.5166, 
    377.2891, 390.3913, 413.6357, 444.6428, 442.3636, 488.6983, 526.4742, 
    581.7993, 665.6102, 783.5282, 909.798, 1160.341, 1189.347, 1036.943, 
    1004.612, 1053.218, 1059.908, 1416.363,
  279.6242, 227.4193, 199.1174, 149.1774, 83.37285, 3.592551, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 101.2812, 60.90662, 478.8484, 643.0255, 690.905, 
    652.9017, 619.0784, 549.6542, 517.7484, 445.3293, 372.7345, 391.3872, 
    396.3501, 434.3335, 453.7928, 469.5943, 484.0396, 513.5276, 579.3093, 
    651.2834, 708.0594, 776.8271, 870.302, 1036.794, 1245.989, 901.5364, 
    940.5923, 1070.94, 1195.01, 1146.841,
  196.4323, 187.7343, 179.3497, 120.5639, 39.21375, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2.005413, 45.81821, 62.24737, 21.02495, 
    3.207724, 0.02404907, 1.234567, 12.24459, 1.728072, 0, 0, 0, 0, 0, 0, 
    3.453561, 7.352701, 19.79626, 158.7443, 296.7885, 521.1622, 627.5361, 
    662.5475, 682.7275, 655.5103, 590.583, 580.2885, 526.9755, 427.6072, 
    407.3717, 430.1629, 446.7533, 474.6825, 500.0133, 519.8837, 559.5943, 
    617.9446, 655.3353, 686.9636, 713.472, 753.1322, 906.1678, 1018.012, 
    815.1847, 882.2279, 1056.679, 1259.787, 1045.098,
  141.7976, 159.4438, 144.7507, 76.36758, 7.418705, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5.733681, 94.68479, 175.18, 187.5313, 
    155.0462, 110.0206, 72.29835, 93.21919, 121.2557, 115.5466, 66.30669, 
    6.150113, 0, 0, 0, 3.670892, 28.15756, 46.06707, 79.14339, 305.7281, 
    712.5394, 940.3807, 751.7666, 698.2665, 746.433, 768.7173, 723.7104, 
    672.3049, 616.0403, 509.8206, 453.0623, 453.5248, 504.1813, 528.5236, 
    544.4155, 565.7984, 598.8699, 625.6595, 655.5828, 686.7064, 683.7915, 
    732.2036, 789.5637, 840.5327, 723.5177, 745.4189, 965.6844, 1038.274, 
    796.5178,
  95.12392, 103.6217, 82.47251, 13.03405, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.002540734, 15.74638, 122.9433, 222.9018, 302.6361, 
    279.6983, 224.5893, 190.8986, 149.559, 188.5142, 236.7475, 212.6731, 
    150.321, 153.6949, 48.69242, 25.20141, 29.67488, 91.25098, 132.1451, 
    112.2913, 103.7838, 263.8452, 764.3199, 1062.096, 1009.38, 884.1952, 
    931.0499, 977.1282, 882.8214, 713.9742, 616.5552, 536.9384, 509.7403, 
    500.2069, 555.3665, 585.5272, 600.3098, 607.6362, 615.286, 634.0374, 
    661.1276, 645.6732, 626.6214, 638.4325, 669.1021, 625.0273, 530.0295, 
    528.0609, 601.1044, 644.5855, 548.4876,
  30.5022, 27.99392, 7.313161, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.7658302, 12.3739, 142.0602, 300.8344, 465.4789, 498.4969, 
    391.7122, 316.7618, 249.2353, 219.1284, 259.9997, 244.4664, 174.3858, 
    179.9653, 249.7257, 193.2922, 150.1301, 234.5797, 302.7541, 285.0494, 
    207.801, 158.7262, 115.508, 347.3649, 690.9739, 928.4409, 982.3543, 
    1030.41, 1034.681, 877.8196, 652.1367, 503.6282, 493.2419, 491.9219, 
    520.8734, 593.4538, 643.876, 652.7304, 662.8006, 652.0361, 676.1411, 
    653.5867, 602.203, 551.5805, 537.899, 522.2339, 492.5406, 445.3781, 
    430.9313, 431.1991, 487.3873, 602.6268,
  0.766829, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7.8648, 
    83.18796, 276.2613, 500.1916, 600.5903, 597.6884, 475.5048, 352.7767, 
    314.1613, 281.9288, 287.8528, 237.377, 131.9863, 144.99, 306.4143, 
    294.3946, 305.1169, 332.2526, 310.4181, 229.8286, 185.2745, 224.0371, 
    255.049, 135.4041, 273.2138, 527.6912, 587.1231, 611.7789, 642.2618, 
    595.1403, 463.5603, 424.1609, 415.3838, 429.1796, 490.9037, 608.7256, 
    694.1671, 728.9787, 711.6575, 716.4285, 701.124, 642.769, 552.2159, 
    495.597, 465.6459, 440.4718, 429.3813, 424.0435, 422.3978, 418.5041, 
    446.8545, 718.7314,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.295444, 78.97375, 
    275.3757, 455.0948, 458.2011, 506.2027, 494.194, 412.8863, 375.2495, 
    355.046, 307.8675, 307.6067, 255.4145, 162.655, 174.7049, 269.6479, 
    362.2924, 358.3284, 318.2245, 211.9518, 198.9956, 327.952, 577.7234, 
    678.533, 449.4442, 258.9631, 309.9615, 318.2204, 354.7622, 372.4727, 
    407.3471, 409.3253, 394.0547, 388.1353, 397.6263, 455.2305, 588.9576, 
    706.325, 787.8987, 810.1958, 757.8834, 690.1829, 588.7928, 504.9205, 
    456.3733, 419.4193, 401.9965, 409.1686, 411.8871, 415.8695, 412.8529, 
    415.983, 653.3243,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.04495476, 1.543852, 
    40.60966, 249.5493, 570.8077, 624.9529, 503.8392, 404.5659, 388.5279, 
    371.8024, 372.5071, 373.0171, 344.5746, 314.8991, 279.2988, 232.3392, 
    204.3131, 251.619, 321.1378, 336.9094, 265.9687, 241.0423, 314.6817, 
    503.8398, 693.5359, 810.1852, 579.9879, 386.7859, 384.9114, 418.0108, 
    446.1444, 373.0016, 350.7278, 352.2296, 366.1898, 378.6504, 386.957, 
    403.5961, 448.4445, 545.6042, 676.7407, 741.8482, 705.261, 612.5644, 
    508.2358, 457.7974, 419.8724, 397.5679, 394.2395, 399.4266, 405.9669, 
    407.882, 402.7976, 410.4689, 789.8555,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.7914926, 10.71653, 
    37.00443, 201.4314, 448.087, 531.7697, 431.7727, 398.7067, 393.9764, 
    349.5272, 333.6953, 360.2705, 337.4265, 298.6373, 309.2917, 282.9134, 
    270.9925, 231.9091, 272.6257, 235.9534, 234.1443, 273.3409, 414.232, 
    561.9924, 633.738, 604.2332, 478.0908, 428.5763, 404.8661, 464.5562, 
    464.1216, 373.5608, 319.6164, 329.3439, 353.2355, 408.3477, 412.724, 
    410.5272, 419.3637, 448.9814, 538.6779, 576.0292, 562.1622, 501.3907, 
    457.8747, 424.4431, 405.648, 395.4491, 393.9858, 397.7108, 400.8848, 
    400.0156, 396.7203, 474.1039, 980.1252,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6.459178, 23.89642, 
    39.5673, 52.56926, 168.347, 227.195, 285.7491, 353.7228, 381.3757, 
    362.791, 311.1005, 312.541, 320.0593, 289.4526, 308.0459, 311.635, 
    295.6172, 265.5541, 242.1341, 228.7672, 222.6893, 264.653, 356.3772, 
    481.8984, 514.7236, 444.572, 376.3537, 375.8529, 367.9664, 341.9634, 
    351.7896, 291.5329, 307.0333, 322.6101, 365.6251, 444.1953, 465.1169, 
    441.8697, 452.7754, 478.7091, 527.0575, 540.0756, 491.8977, 461.4532, 
    433.0887, 417.837, 414.4355, 413.9627, 410.6415, 421.8182, 400.1716, 
    394.3721, 399.2646, 611.9307, 1308.194,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6.790205, 27.87427, 
    37.87522, 49.99376, 77.3848, 129.5688, 225.8023, 291.5181, 345.4376, 
    327.5065, 299.076, 285.3165, 292.4263, 320.6955, 306.0085, 310.2983, 
    291.4063, 262.9675, 246.8307, 238.5132, 249.1621, 271.4966, 326.77, 
    393.712, 450.9673, 416.2671, 374.2629, 344.2727, 333.5673, 305.9854, 
    280.9805, 285.871, 292.4921, 298.5072, 329.7079, 419.0633, 450.0066, 
    465.448, 502.8485, 574.8007, 637.0599, 703.0728, 587.3303, 483.8123, 
    452.7943, 442.7585, 455.8902, 478.3641, 513.434, 528.1032, 446.6922, 
    395.0017, 396.0436, 580.3947, 1096.152,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 7.539374, 13.82793, 0, 0, 0, 0, 0, 0.3629586, 
    22.22618, 38.05198, 50.36842, 51.9423, 55.76481, 123.9351, 200.9567, 
    248.0657, 288.369, 296.5797, 284.997, 272.4008, 306.0285, 313.191, 
    326.7126, 292.9926, 277.2778, 264.6691, 265.5726, 260.786, 272.6996, 
    322.4322, 380.3541, 402.2595, 439.8839, 455.1393, 427.6396, 381.3865, 
    336.1739, 308.6934, 286.1038, 296.1768, 298.6016, 292.2509, 297.8213, 
    348.2343, 392.0045, 441.4889, 561.517, 686.3062, 815.3308, 935.5671, 
    875.5865, 574.7263, 510.7076, 481.0591, 505.4455, 569.8447, 637.2155, 
    645.5725, 578.0183, 406.8309, 416.0845, 555.6661, 828.242,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 6.968982, 31.56356, 1.362759, 0, 0, 0, 0, 0, 
    9.483889, 33.60556, 38.53296, 50.37358, 74.38406, 139.3567, 205.6824, 
    215.1312, 223.8199, 264.2617, 295.2328, 280.9891, 269.5547, 301.0195, 
    283.1612, 300.8699, 290.1711, 288.1376, 298.2253, 296.4409, 301.7662, 
    372.0651, 450.2336, 467.1264, 467.0771, 487.0597, 462.8398, 408.4555, 
    374.192, 332.696, 321.5491, 328.5142, 322.4901, 299.8736, 293.3217, 
    324.0511, 366.8441, 447.5163, 626.8708, 836.7401, 890.7211, 1096.81, 
    1047.843, 760.592, 575.9907, 540.1681, 540.2332, 595.8331, 628.45, 
    649.7249, 568.4493, 455.0399, 431.6068, 517.0565, 601.8608,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 1.797053, 7.747849, 3.450143, 0, 0, 0, 0, 0, 
    0.9109401, 18.42504, 39.59516, 52.26551, 97.90691, 235.892, 219.3992, 
    208.2924, 216.5296, 262.5898, 292.2108, 286.3712, 274.5794, 269.5547, 
    279.5371, 287.6822, 293.7041, 308.5545, 345.3323, 335.1651, 328.9469, 
    369.3367, 444.4053, 470.777, 502.3892, 510.839, 472.6234, 420.1351, 
    393.2463, 375.5051, 344.6975, 341.879, 320.9992, 295.3217, 288.8875, 
    310.2828, 356.9085, 436.3004, 643.2478, 908.5942, 908.9702, 1001.605, 
    1072.39, 855.878, 706.8087, 615.7324, 594.7244, 607.8818, 589.8001, 
    519.1802, 495.0875, 398.2069, 416.0681, 481.5428, 468.7679,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 45.77684, 0, 0, 0, 0, 0, 0, 0, 0, 19.37672, 
    35.37803, 69.18604, 153.2726, 288.3199, 317.8352, 244.572, 258.4949, 
    287.7384, 311.5768, 297.4268, 289.1551, 278.5264, 276.3994, 304.6932, 
    323.0869, 346.2746, 396.4057, 380.4884, 341.7323, 349.6577, 376.4726, 
    426.947, 504.5984, 651.9197, 501.9165, 434.0541, 415.7284, 411.0024, 
    387.9035, 340.0662, 290.0233, 265.8179, 252.4831, 284.6985, 349.8331, 
    406.4402, 572.5109, 805.2451, 886.5491, 902.3984, 984.8835, 957.6617, 
    842.1849, 709.3141, 604.957, 577.4132, 542.0748, 476.5501, 421.5896, 
    398.5287, 416.1053, 436.3309, 444.6508,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.2233779, 7.883308, 
    46.45991, 63.79469, 184.3558, 336.8821, 374.0247, 374.8209, 335.6512, 
    339.178, 324.0201, 312.332, 293.5074, 275.675, 291.9893, 330.8283, 
    374.3214, 414.9174, 493.441, 464.5028, 388.4646, 358.354, 358.3539, 
    399.2584, 604.8146, 824.4387, 636.0546, 425.0211, 422.0507, 444.4562, 
    444.8008, 388.2694, 300.7451, 240.5886, 216.5688, 229.7297, 312.2461, 
    400.7599, 488.0696, 759.7354, 869.7776, 810.3863, 836.918, 927.7097, 
    906.3384, 778.0356, 610.2334, 542.7169, 508.4426, 490.6646, 424.6607, 
    396.6208, 405.9286, 424.3958, 467.8904,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.524688, 44.15213, 
    88.41959, 159.127, 276.4428, 370.4227, 392.6274, 382.1442, 366.4334, 
    336.8749, 317.2722, 299.4598, 286.5885, 283.6873, 292.2945, 335.28, 
    393.107, 469.711, 592.4265, 585.6436, 482.2569, 415.559, 389.8748, 
    408.3621, 619.8497, 895.7261, 639.1478, 447.5954, 410.7881, 450.1098, 
    465.333, 443.5472, 380.2547, 332.284, 295.5856, 256.3805, 299.0791, 
    379.3657, 547.1831, 780.5206, 955.9313, 825.8504, 679.0082, 745.6443, 
    771.3798, 700.3216, 547.1471, 488.1773, 493.5975, 534.8677, 465.9749, 
    408.6629, 406.9938, 428.9316, 486.2154,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8.648079, 90.31952, 
    139.5776, 213.0849, 372.9224, 415.0632, 410.2803, 377.4778, 360.1422, 
    341.8087, 303.7456, 280.1181, 284.2162, 290.7113, 310.3253, 325.1641, 
    379.646, 458.2865, 595.5748, 642.431, 599.8919, 527.5738, 473.18, 
    483.1668, 614.2881, 799.8925, 603.7574, 431.5247, 413.0665, 434.388, 
    454.1592, 461.4271, 468.4397, 452.5511, 440.9289, 400.6418, 349.5063, 
    404.0337, 485.1346, 668.6317, 844.2675, 779.2899, 658.3606, 603.169, 
    619.9202, 579.0063, 475.0612, 424.7502, 455.7198, 513.4985, 468.9218, 
    415.5838, 421.0052, 460.8036, 482.3849,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26.58741, 141.5162, 
    204.9548, 236.1427, 343.1058, 379.2624, 360.7214, 335.7108, 336.3476, 
    332.6995, 308.2321, 285.1463, 271.4974, 292.8643, 320.6105, 328.3786, 
    355.2569, 397.3354, 482.0117, 568.8033, 603.5388, 619.1583, 583.2557, 
    547.499, 603.738, 696.2391, 558.0874, 454.7069, 434.771, 488.2554, 
    465.5451, 480.1592, 528.2115, 662.0346, 767.2975, 774.6315, 505.6811, 
    453.9677, 500.7877, 584.0219, 721.4752, 757.2107, 622.8404, 564.5931, 
    553.7775, 544.0915, 438.6134, 401.1854, 402.1854, 448.803, 413.0183, 
    422.9466, 438.3102, 442.5483, 441.3457,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9.301848, 158.3098, 
    258.9337, 303.8173, 299.6194, 299.056, 279.9115, 262.4927, 294.193, 
    317.6132, 308.028, 282.2506, 265.0864, 268.781, 299.4977, 330.493, 
    349.1855, 376.8177, 421.5884, 502.247, 599.8027, 734.8414, 890.7762, 
    678.5621, 700.035, 677.1342, 600.2327, 509.2974, 559.8538, 608.821, 
    538.714, 488.7658, 668.5876, 1060.59, 1373.92, 1418.137, 819.2729, 
    541.28, 535.3813, 612.2632, 721.4976, 746.7157, 652.4662, 555.7067, 
    576.511, 582.4625, 469.2462, 383.6081, 342.5653, 332.923, 354.656, 
    407.8102, 443.4485, 401.7837, 378.6187,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 86.89892, 228.9686, 
    307.1906, 284.381, 247.07, 238.9294, 245.0831, 292.1502, 321.7906, 
    317.2473, 299.972, 288.464, 279.9789, 285.0193, 296.3184, 328.2048, 
    358.1512, 417.3985, 513.0966, 649.8973, 1018.273, 1282.382, 1139.754, 
    900.5889, 797.8112, 659.6571, 681.5824, 716.9097, 741.9376, 622.0638, 
    551.46, 815.8694, 1147.539, 1486.932, 1523.49, 1029.805, 601.8781, 
    552.1006, 578.9692, 660.6729, 721.0251, 691.4706, 615.808, 579.7531, 
    580.8895, 447.5938, 336.6733, 275.8545, 256.4472, 302.6965, 384.8403, 
    451.3116, 391.0798, 372.3258,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5.010157, 137.2761, 
    246.5296, 275.4832, 286.3332, 281.9478, 285.9474, 335.5515, 358.7326, 
    329.0612, 289.5595, 278.5055, 274.489, 270.4537, 278.7563, 306.5069, 
    345.374, 407.7699, 519.6101, 695.6252, 1020.536, 1431.428, 1296.497, 
    1159.715, 894.8511, 889.3289, 837.659, 898.1722, 824.8221, 688.373, 
    685.1447, 783.9781, 882.051, 899.179, 1132.87, 975.0953, 703.803, 
    579.3523, 556.1559, 602.6837, 672.3351, 701.9514, 668.7778, 612.2599, 
    538.6722, 430.2552, 334.1217, 260.4696, 247.4416, 300.6423, 367.5648, 
    419.1653, 385.3712, 385.5648,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 57.55773, 181.7126, 
    294.1019, 358.642, 376.2969, 381.9689, 378.035, 391.0516, 372.8776, 
    348.465, 324.6873, 307.1947, 273.0872, 273.6699, 274.8869, 275.7082, 
    315.3789, 463.814, 693.0596, 959.1632, 1143.813, 1204.84, 1186.019, 
    1113.179, 1009.146, 981.3286, 895.3462, 765.3611, 644.151, 603.1124, 
    711.8834, 624.4473, 590.9575, 727.5765, 872.574, 675.1846, 577.9081, 
    544.3901, 554.0104, 578.1396, 636.2142, 666.0281, 591.5745, 499.7725, 
    416.1812, 362.9875, 301.6709, 266.8849, 341.4141, 365.0664, 373.7022, 
    355.0049, 393.6327,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7.672453, 76.61076, 
    200.5678, 304.525, 397.0667, 442.379, 428.145, 388.1142, 388.5081, 
    408.9069, 422.5594, 380.0047, 325.1395, 271.7728, 229.48, 221.3898, 
    214.3802, 330.7382, 597.4027, 826.9779, 1010.901, 1106.384, 1267.898, 
    1164.386, 1014.269, 812.2874, 856.5626, 721.2389, 588.0623, 545.859, 
    605.4478, 543.02, 491.1708, 537.3549, 686.0102, 599.1124, 549.1641, 
    530.5813, 510.3197, 549.0093, 608.9304, 682.692, 603.2574, 419.0844, 
    360.2815, 332.0342, 312.2987, 297.1729, 354.3885, 423.995, 364.6626, 
    357.3581, 429.184,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4.492652, 0, 5.913332, 0, 
    9.827749, 122.8932, 239.9646, 413.3958, 469.7688, 442.4698, 411.2574, 
    384.8907, 404.1997, 419.0803, 395.6619, 331.3684, 275.5099, 249.502, 
    270.0858, 300.564, 302.8828, 432.2428, 627.8237, 685.1678, 758.2089, 
    829.3271, 816.4886, 691.1724, 675.4188, 734.3888, 674.1106, 540.9742, 
    509.9907, 540.2866, 512.6861, 438.8988, 428.1956, 510.8031, 492.1108, 
    477.0582, 467.651, 481.3288, 477.3205, 570.1652, 742.3004, 660.6039, 
    434.6603, 307.3639, 286.5654, 295.7912, 296.1364, 355.3662, 457.1753, 
    393.4307, 396.5924, 493.4605,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 38.18091, 177.9759, 
    78.61066, 5.231147, 20.97725, 4.670784, 80.24761, 276.9565, 515.89, 
    480.1449, 420.3515, 475.0774, 450.7651, 429.4347, 397.8179, 353.9267, 
    293.7534, 272.3435, 388.218, 463.1545, 491.6412, 475.5977, 481.5441, 
    496.2309, 455.1932, 510.3101, 537.7867, 541.0651, 539.1157, 607.288, 
    534.366, 475.9772, 458.8337, 508.1748, 500.2999, 470.7975, 373.0616, 
    372.9929, 372.6212, 339.7219, 379.8255, 402.0655, 426.9336, 542.4205, 
    772.5742, 775.2917, 518.3701, 319.2849, 250.5893, 235.3483, 234.3458, 
    282.5884, 389.9496, 389.2494, 430.362, 541.4569,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 42.64318, 0, 0, 0, 14.13362, 
    0, 0, 97.32533, 567.0143, 755.1489, 660.1171, 552.6977, 559.0915, 
    519.6163, 501.7351, 442.0413, 369.866, 317.342, 371.9945, 499.4051, 
    535.2877, 491.8406, 421.9243, 376.5453, 400.5975, 453.606, 510.7452, 
    552.5534, 541.176, 503.5962, 466.0743, 452.3511, 428.7473, 469.4224, 
    558.7114, 555.1274, 362.4989, 286.6256, 277.3649, 257.8876, 279.6031, 
    357.494, 406.6543, 470.3801, 647.2722, 685.0935, 537.283, 372.8993, 
    288.5817, 221.9755, 181.4825, 209.1741, 291.7701, 287.4789, 395.4302, 
    561.2106,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01953389, 0, 0, 0, 
    0, 0, 455.7978, 1051.609, 1211.341, 1040.144, 739.9411, 620.1765, 
    620.5828, 543.5131, 502.523, 425.7497, 412.7139, 442.9023, 449.829, 
    379.7539, 314.4379, 297.9188, 320.5314, 397.3131, 505.9446, 602.7551, 
    619.6101, 569.6279, 539.3142, 520.7625, 497.6906, 523.4991, 613.6224, 
    612.6038, 400.595, 262.5043, 224.5589, 204.1281, 205.329, 279.9945, 
    355.9917, 390.6264, 461.2118, 514.0649, 484.4973, 380.1658, 331.9442, 
    259.4583, 192.7791, 282.2837, 280.4692, 273.8584, 398.2701, 491.5527,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    524.9088, 1227.854, 1514.503, 1593.471, 1283.125, 835.2573, 726.7971, 
    681.4029, 629.7035, 589.2842, 510.3927, 473.1457, 430.4084, 306.1007, 
    237.6619, 228.5278, 244.4046, 284.5834, 374.7751, 497.4753, 605.6686, 
    636.1135, 616.2618, 595.865, 525.5728, 477.7885, 496.7985, 413.9014, 
    286.8343, 221.6673, 207.5997, 165.5916, 149.3675, 196.3652, 251.1849, 
    278.328, 301.5162, 361.5432, 350.5833, 304.2287, 281.5658, 276.7146, 
    189.8026, 362.6567, 363.6728, 247.8723, 372.7149, 441.053,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    109.9336, 398.2949, 940.3243, 1436.861, 1731.173, 1299.493, 1035.062, 
    902.295, 892.6244, 738.1326, 628.37, 557.6457, 490.0444, 346.9488, 
    207.4061, 175.4873, 181.6765, 210.3732, 258.1815, 368.8855, 533.0062, 
    620.7709, 626.9582, 508.8629, 400.888, 363.2095, 333.2734, 270.4286, 
    219.8917, 179.2967, 159.2247, 142.6616, 109.0908, 142.8433, 178.4309, 
    190.0326, 221.8169, 245.1929, 268.4247, 231.8128, 307.9815, 330.6054, 
    275.8257, 397.8697, 359.8254, 219.364, 334.6523, 463.7612,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.06423091, 57.11491, 0, 0, 
    0, 0, 0, 0, 7.836217, 136.0153, 314.1614, 994.2757, 1493.946, 1517.679, 
    1301.398, 1272.304, 1158.99, 1018.497, 845.142, 688.6971, 603.6498, 
    439.0118, 236.4267, 146.054, 144.4927, 163.0123, 225.2119, 349.3079, 
    489.0631, 592.2128, 608.7792, 410.0895, 244.743, 193.4141, 256.4616, 
    227.5397, 197.2503, 107.2875, 83.52959, 68.98138, 80.46129, 115.9747, 
    132.9302, 145.9669, 152.7381, 174.7173, 173.7455, 175.6978, 235.3297, 
    318.201, 276.576, 340.2295, 316.9229, 225.2303, 420.5147, 420.0156,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2.182514, 89.51676, 343.4627, 955.3691, 1260.624, 1151.738, 1138.569, 
    1236.952, 1157.061, 1085.779, 1005.899, 794.526, 562.4872, 299.4979, 
    123.4399, 98.68906, 119.4459, 185.4302, 329.3733, 361.4457, 432.3123, 
    502.7655, 379.1094, 146.3032, 62.53582, 92.53636, 99.53645, 60.84525, 
    11.73829, 14.53334, 21.45396, 50.65263, 84.13147, 89.0048, 93.22248, 
    110.0247, 112.9956, 145.8865, 186.0687, 228.4272, 220.4345, 204.2188, 
    252.7047, 291.9086, 311.514, 407.4745, 196.5356,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 37.47989, 422.1205, 709.343, 683.818, 813.1848, 1012.258, 1090.199, 
    1166.657, 1117.992, 963.0756, 744.8711, 327.3204, 67.59232, 51.20574, 
    51.10489, 136.7648, 215.8003, 145.3761, 67.80409, 186.2934, 218.4242, 
    88.11556, 0.4354767, 0, 0, 0, 0, 34.36349, 48.50853, 69.10825, 73.94706, 
    66.00063, 75.26979, 83.438, 52.38344, 29.00477, 151.119, 204.1204, 
    143.2567, 130.4681, 270.9427, 483.1219, 465.0688, 362.5184, 4.126702,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 17.66449, 261.7532, 151.233, 91.45276, 90.23305, 372.949, 595.9958, 
    811.2404, 1056.335, 1019.892, 820.1436, 449.4274, 159.2536, 109.9366, 
    231.9172, 190.1881, 121.1451, 13.04661, 0.002457884, 0.07684267, 
    1.469449, 0.02487941, 0, 0, 0, 0, 0, 69.92484, 163.3495, 125.5531, 
    119.3953, 127.3019, 150.9474, 169.9525, 115.3876, -54.83441, 78.6655, 
    169.3711, 172.5084, 110.4562, 298.2401, 618.7454, 450.6016, 111.6259, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 18.18774, 198.2974, 24.82351, 0.01659623, 0, 9.641451, 62.01321, 
    362.3916, 663.819, 745.0246, 764.4761, 729.5575, 860.1415, 989.5406, 
    901.2372, 633.0322, 214.5284, 22.94515, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    71.94882, 276.9225, 273.4788, 160.4362, 155.9303, 183.5391, 191.451, 
    188.135, 115.3398, 35.40816, 124.8625, 162.5711, 94.14777, 280.8703, 
    519.7524, 233.8496, 268.5618, 36.8153,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.1127852, 103.1683, 83.84983, 125.6781, 310.4157, 588.7912, 843.4153, 
    526.3326, 1.147217, 0, 31.65186, 188.915, 342.4284, 556.4823, 714.2188, 
    878.2565, 858.4985, 833.0258, 646.3763, 302.5152, 38.86568, 0, 
    0.01003916, 0, 0, 0, 0, 0, 0, 0, 0, 50.22194, 269.6366, 109.4844, 
    37.02338, 59.75043, 26.35164, 79.59688, 104.9516, 76.24226, 67.52459, 
    111.2902, 103.7956, 226.3943, 374.5558, 285.326, 834.7192, 451.0992,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 2.3265, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3.225108, 103.0244, 258.1696, 347.2978, 418.1593, 560.3155, 894.6843, 
    791.2195, 306.0076, 0.8998873, 0, 0, 0, 14.49841, 35.44591, 118.7575, 
    200.4224, 258.1529, 344.5415, 204.937, 28.87837, 0, 0.1383204, 0, 
    2.479101, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01911015, 
    8.849098, 12.94733, 55.8584, 180.516, 374.3842, 761.2708, 606.065,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 15.89997, 14.70358, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 37.67767, 140.6756, 246.9203, 375.567, 456.3772, 603.2179, 
    768.8178, 926.5468, 582.7935, 196.5176, 0, 0.4811277, 0, 0, 0, 0, 0, 0, 
    24.83666, 45.255, 12.15549, 2.415782, 0, 0.09825284, 1.407857, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.6392468, 2.363386, 28.96285, 
    234.0622, 386.0693, 563.9972,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 17.55955, 29.1074, 15.34933, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 10.62364, 190.7695, 391.3156, 404.325, 600.9966, 680.045, 
    704.8675, 862.8046, 749.6393, 130.0502, 3.100419, 5.116066, 6.17757, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.4328433, 76.46776, 242.6619, 291.0963, 5.134037, 
    0, 0, 0, 0, 0, 0, 0, 0, 0.8376673, 0, 0, 0, 0, 0, 0, 0, 0, 0.008186113, 
    0.07604827, 15.87589, 119.0556, 379.1627,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 1.163343, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 255.9357, 568.2272, 791.1302, 892.6254, 903.9981, 891.0063, 
    1059.328, 1098.428, 617.2275, 6.932829, 0.3629374, 65.03675, 7.93887, 0, 
    0, 0, 0.8275996, 112.0045, 17.52323, 0, 0, 57.19586, 246.4086, 451.7093, 
    100.6016, 0.06041526, 0, 0, 0, 0, 0, 0, 0.5732526, 182.9803, 198.6564, 
    161.3975, 11.53954, 0, 0, 0, 0, 0, 0, 0, 0, 0.992954, 173.7827,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 8.585627, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 257.8992, 621.7795, 752.3851, 846.557, 900.2053, 1019.242, 1113.99, 
    880.9015, 529.3146, 159.8383, 6.419941, 0, 0, 0, 0, 0, 0.03464887, 
    317.7343, 145.3232, 0, 0, 0.1035934, 0, 5.595896, 134.9415, 159.4373, 0, 
    0, 0, 0, 0.5597559, 213.3741, 71.13373, 0, 0, 10.51704, 18.63104, 
    3.763446, 0, 0, 0, 0, 0, 0, 0, 0, 34.35713,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1.43994, 381.3143, 748.3234, 941.8181, 893.6531, 933.1523, 1035.22, 
    860.355, 610.6863, 554.7979, 525.4812, 498.002, 75.12685, 0, 0, 0, 0, 
    11.73125, 325.2318, 124.1923, 0, 0, 0, 0, 0, 42.32673, 450.324, 9.972672, 
    0, 0, 34.3005, 62.80934, 603.7728, 328.5521, 8.121914, 9.169447, 
    6.230115, 1.321965, 11.59744, 3.048517, 0, 0, 0, 0, 0, 0, 0, 6.704556,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    30.85074, 297.304, 660.8721, 966.9948, 998.4858, 885.1306, 751.5646, 
    655.1858, 732.1314, 1084.44, 1349.639, 1119.806, 408.8793, 0, 0, 0, 0, 0, 
    140.0299, 7.918328, 0, 0, 0.1702392, 1.991248, 53.83979, 472.2008, 
    346.2012, 2.112901, 0.005206824, 0, 24.37175, 219.4124, 598.756, 
    329.5864, 98.26838, 18.94595, 28.95024, 2.492014, 22.5628, 50.42095, 0, 
    0, 0, 0, 22.81216, 24.65398, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    26.93062, 106.7775, 98.48605, 75.9237, 51.93491, 62.07972, 66.57274, 
    176.725, 422.3495, 479.3473, 519.7673, 215.12, 2.231832, 0.004072465, 
    1.405816, 0.08232938, 0, 495.7819, 40.24272, 0, 7.263184, 112.9553, 
    325.7667, 421.6084, 533.7393, 301.4734, 91.60561, 24.09392, 33.98492, 
    380.9341, 705.0402, 632.1104, 263.1127, 138.8074, 37.80578, 1.129739, 
    35.61073, 95.76726, 325.1597, 511.9413, 832.47, 77.51266, 0, 41.77975, 
    292.1154, 30.66951, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 23.8246, 73.93395, 126.2193, 321.1346, 494.5471, 
    282.6015, 106.8233, 331.644, 202.062, 0, 24.80076, 24.1915, 49.88836, 
    269.6974, 671.1443, 778.3289, 494.5531, 183.3987, 40.72751, 10.41955, 0, 
    92.49084, 767.71, 1000.381, 579.1232, 178.2135, 9.95975, 6.408473, 
    10.95331, 70.58002, 197.3521, 552.4769, 928.8527, 1256.867, 539.4283, 
    47.92098, 154.266, 98.49847, 27.90792, 1.357446 ;
}
