netcdf atmos_month.198001-198012.alb_sfc {
dimensions:
	time = UNLIMITED ; // (12 currently)
	lat = 18 ;
	lon = 29 ;
	bnds = 2 ;
variables:
	float alb_sfc(time, lat, lon) ;
		alb_sfc:long_name = "Surface Albedo for  Flux" ;
		alb_sfc:units = "percent" ;
		alb_sfc:_FillValue = 1.e+20f ;
		alb_sfc:missing_value = 1.e+20f ;
		alb_sfc:cell_methods = "time: mean" ;
		alb_sfc:cell_measures = "area: area" ;
		alb_sfc:interp_method = "conserve_order1" ;
	double lat(lat) ;
		lat:standard_name = "latitude" ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_N" ;
		lat:axis = "Y" ;
		lat:bounds = "lat_bnds" ;
	double lat_bnds(lat, bnds) ;
	double lon(lon) ;
		lon:standard_name = "longitude" ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_E" ;
		lon:axis = "X" ;
		lon:bounds = "lon_bnds" ;
	double lon_bnds(lon, bnds) ;
	double time(time) ;
		time:standard_name = "time" ;
		time:long_name = "time" ;
		time:bounds = "time_bnds" ;
		time:units = "days since 1979-01-01 00:00:00" ;
		time:calendar = "standard" ;
		time:axis = "T" ;
	double time_bnds(time, bnds) ;

// global attributes:
		:CDI = "Climate Data Interface version 2.4.4 (https://mpimet.mpg.de/cdi)" ;
		:Conventions = "CF-1.6" ;
		:title = "c96L65_am5f9d8r0_amip" ;
		:associated_files = "area: 19800101.grid_spec.nc" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
		:code_release_version = "2024.05" ;
		:git_hash = "5d306c05d9fe755cab04eedc8fd3de0d3c8355a0" ;
		:creationtime = "Mon Aug 11 19:59:10 2025" ;
		:hostname = "pp033" ;
		:history = "Mon Aug 11 16:13:43 2025: ncks -d lat,,,10 -d lon,,,10 atmos_month.198001-198012.alb_sfc.nc reduced/atmos_month.198001-198012.alb_sfc.nc\n",
			"Mon Aug 11 20:02:14 2025: cdo --history splitname 19800101.atmos_month.nc /home/Chris.Blanton/cylc-run/c96L65_am5f9d8r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run1/share/cycle/19800101T0000Z/split/regrid-xy/180_288.conserve_order2/19800101.atmos_month.\n",
			"fregrid --debug --standard_dimension --input_mosaic C96_mosaic.nc --input_dir /home/Chris.Blanton/cylc-run/c96L65_am5f9d8r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run1/share/cycle/19800101T0000Z/history/native --input_file 19800101.atmos_month --associated_file_dir /home/Chris.Blanton/cylc-run/c96L65_am5f9d8r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run1/share/cycle/19800101T0000Z/history/native --interp_method conserve_order2 --remap_file fregrid_remap_file_288_by_180.nc --nlon 288 --nlat 180 --scalar_field (**please see the field list in this file**) --output_file 19800101.atmos_month.nc" ;
		:CDO = "Climate Data Operators version 2.4.4 (https://mpimet.mpg.de/cdo)" ;
		:NCO = "netCDF Operators version 5.2.4 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco, Citation = 10.1016/j.envsoft.2008.03.004)" ;
data:

 alb_sfc =
  76.21249, 76.21249, 76.21249, 76.21249, 76.21249, 76.21249, 76.21249, 
    76.2067, 76.2067, 76.2067, 76.2067, 76.2067, 76.2067, 76.2067, 76.20618, 
    76.20618, 76.20618, 76.20618, 76.20618, 76.20618, 76.20618, 76.22049, 
    76.22049, 76.22049, 76.22049, 76.22049, 76.22049, 76.22049, 76.21249,
  76.5369, 76.35718, 76.23174, 76.10892, 76.10101, 76.08167, 76.05757, 
    76.01556, 76.03475, 76.10069, 76.13761, 76.25919, 76.36391, 74.80975, 
    76.22225, 70.45061, 72.72987, 70.20911, 67.06656, 73.40981, 74.84594, 
    75.86151, 74.76565, 65.86028, 72.43765, 67.02516, 71.26469, 68.82244, 
    76.55497,
  51.43897, 60.99732, 38.65466, 64.09626, 72.40456, 72.73711, 53.51461, 
    72.80325, 72.66396, 72.08009, 72.7183, 73.06756, 68.82347, 25.47618, 
    6.310994, 6.287273, 6.188186, 6.40295, 6.345472, 40.47618, 48.00944, 
    37.99785, 59.14075, 61.76669, 61.29424, 60.35058, 53.38457, 6.341237, 
    11.61759,
  4.584107, 4.622993, 4.815651, 4.85297, 4.736935, 4.608834, 4.689611, 
    4.663966, 4.732478, 4.913521, 4.805801, 4.686138, 4.733097, 4.791592, 
    4.823448, 4.757921, 4.587622, 4.728386, 4.739498, 4.89659, 5.09698, 
    4.924362, 5.034412, 4.946849, 4.902513, 4.661936, 18.9911, 4.721068, 
    4.634075,
  4.176626, 4.266893, 4.226772, 4.273165, 4.334706, 4.292007, 4.357611, 
    4.247204, 4.304564, 4.255612, 4.303858, 4.410933, 4.568583, 4.389814, 
    4.393828, 4.621373, 4.339199, 4.349639, 4.305265, 4.272543, 4.297712, 
    4.22269, 4.342278, 8.659232, 4.840526, 4.434886, 4.38345, 4.265073, 
    4.299405,
  4.356071, 4.202331, 4.264299, 4.122086, 3.973567, 4.03682, 4.108491, 
    4.330956, 3.958149, 4.225961, 3.932641, 4.286959, 4.098232, 4.146395, 
    10.42426, 4.088362, 4.222639, 4.029999, 4.073057, 3.914867, 4.115468, 
    4.028337, 4.180781, 9.999311, 4.54083, 4.18158, 3.942292, 3.930175, 
    4.129374,
  4.030599, 4.133832, 12.66912, 3.775947, 3.916299, 4.163543, 3.790476, 
    3.997024, 3.86202, 4.048335, 10.20615, 15.79773, 10.34978, 3.861449, 
    3.918101, 3.842443, 3.749597, 3.522948, 3.62639, 3.725332, 4.295681, 
    4.164379, 4.065354, 4.653529, 9.61346, 3.666675, 3.828869, 3.936225, 
    4.018545,
  3.636105, 10.12084, 12.41177, 3.730566, 3.601546, 3.604157, 3.871427, 
    3.829409, 3.693151, 3.459607, 12.14845, 11.25358, 3.504437, 3.392504, 
    3.66571, 3.742146, 3.362797, 3.645343, 3.544976, 3.935373, 3.878034, 
    3.97615, 3.364853, 3.286826, 9.228889, 9.311712, 3.946262, 3.849511, 
    4.032434,
  3.356254, 6.490816, 8.660058, 9.409101, 3.384045, 3.267991, 3.41915, 
    3.349215, 3.463663, 3.276826, 4.574463, 3.308344, 4.349068, 3.729162, 
    3.491187, 3.358585, 3.3162, 3.787813, 3.605729, 4.005332, 3.699137, 
    3.83112, 3.521028, 8.746784, 8.47916, 9.027272, 3.64309, 3.52108, 3.794034,
  3.272268, 8.928912, 8.70536, 9.986491, 3.425856, 3.524868, 3.158233, 
    3.343197, 8.665392, 8.234029, 3.602675, 3.570207, 3.30008, 3.484152, 
    3.392289, 3.49744, 3.607059, 3.873033, 3.731937, 3.863287, 3.631095, 
    3.429137, 3.364611, 8.588988, 8.381393, 3.253352, 3.324705, 3.47948, 
    3.261089,
  10.20084, 10.30241, 10.59198, 9.733245, 14.32778, 3.513367, 5.362089, 
    3.535958, 3.423971, 3.403905, 4.055064, 3.5247, 3.31671, 3.475969, 
    3.64768, 3.604045, 3.815579, 3.639285, 3.907879, 3.539376, 3.445787, 
    3.565281, 8.599044, 7.277642, 3.656084, 3.816393, 3.356907, 3.869777, 
    9.011524,
  16.08762, 18.65469, 20.70734, 3.771494, 20.81906, 4.048032, 10.02926, 
    3.971389, 8.982236, 3.38551, 3.431337, 3.754703, 3.652293, 3.85797, 
    4.084281, 3.821107, 4.116161, 3.854466, 3.920438, 3.579816, 3.757422, 
    6.07228, 3.640602, 4.422895, 3.821666, 4.082856, 3.770134, 3.966091, 
    21.26264,
  20.44768, 16.1873, 17.27027, 16.63962, 11.2657, 12.66232, 12.07111, 
    29.60023, 7.584904, 10.16815, 3.345697, 3.889911, 4.06545, 3.877009, 
    3.942673, 3.956659, 3.841271, 3.574344, 3.569604, 4.011981, 8.896669, 
    11.01674, 9.713631, 3.923651, 3.897095, 3.772776, 3.698681, 3.816121, 
    10.06392,
  5.819567, 3.979094, 5.33284, 21.90224, 1.618454, 11.986, 23.98764, 
    12.49476, 10.50791, 22.82114, 10.11723, 3.519705, 3.924908, 4.110197, 
    3.959261, 3.766245, 3.703685, 3.580501, 3.486065, 9.28066, 14.60048, 
    13.40509, 15.42212, 4.686903, 3.460612, 3.456538, 3.643784, 3.638644, 
    4.951267,
  4.46006, 17.64599, 19.80454, 26.09016, 25.67087, 25.65604, 10.51527, 
    26.13885, 11.2677, 6.029901, 9.281079, 16.93486, 3.377563, 3.14502, 
    3.498232, 3.350618, 3.421001, 3.566548, 3.787931, 21.26295, 18.95897, 
    22.50855, 17.02384, 20.5606, 9.398446, 3.213188, 3.221211, 3.395527, 
    3.674494,
  3.28493, 10.60896, 9.686433, 14.26786, 14.9195, 15.4171, 16.67404, 
    15.87479, 12.78058, 12.86592, 11.89554, 21.28938, 21.58181, 17.3119, 
    2.331954, 18.95504, 18.73707, 9.409877, 20.89851, 13.72099, 15.0461, 
    21.41998, 25.83009, 21.14217, 2.510523, 5.807779, 3.01138, 2.862548, 
    3.149322,
  0.2170782, 0.1998534, 1.60941, 0.2023845, 1.487759, 2.803855, 2.333739, 
    2.340957, 2.339506, 2.266188, 1.499686, 1.328582, 2.350045, 2.866114, 
    2.902692, 3.075826, 2.677449, 2.986262, 3.037555, 3.148364, 2.59273, 
    2.839533, 2.731728, 2.686438, 2.830736, 2.432736, 2.509262, 2.706268, 
    0.2339574,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  76.45917, 76.45917, 76.45917, 76.45917, 76.45917, 76.45917, 76.45917, 
    76.43328, 76.43328, 76.43328, 76.43328, 76.43328, 76.43328, 76.43328, 
    76.42191, 76.42191, 76.42191, 76.42191, 76.42191, 76.42191, 76.42191, 
    76.449, 76.449, 76.449, 76.449, 76.449, 76.449, 76.449, 76.45917,
  73.2886, 73.07695, 72.97181, 73.06145, 72.80318, 72.95871, 72.936, 
    72.87094, 72.98722, 73.16007, 72.89707, 73.16093, 73.2952, 73.66615, 
    73.70831, 72.95576, 73.75297, 73.02355, 73.13512, 73.86424, 74.08417, 
    74.02661, 73.99445, 73.5184, 74.90501, 73.0404, 74.13445, 73.61415, 
    73.41138,
  36.23158, 39.08492, 8.197051, 48.59606, 55.79223, 56.33447, 39.68078, 
    56.16028, 56.34244, 56.38931, 55.90307, 55.63747, 55.06417, 16.26642, 
    5.666276, 5.549684, 5.491557, 5.207502, 5.106162, 14.33389, 29.07833, 
    19.24171, 47.23975, 48.43013, 48.76183, 48.46383, 5.348134, 5.34516, 
    6.573974,
  4.405357, 4.704306, 4.566124, 4.492412, 4.321194, 4.636532, 4.404022, 
    4.263696, 4.073736, 4.115807, 4.098264, 4.086076, 4.105236, 4.314836, 
    4.372684, 4.356957, 4.550645, 4.292406, 4.530819, 4.595967, 4.777292, 
    4.868098, 4.973146, 4.670944, 4.466017, 4.309252, 4.309019, 4.496097, 
    4.204756,
  4.001403, 3.928081, 3.917543, 4.029042, 4.120102, 4.01884, 3.994899, 
    4.115098, 4.074612, 3.99983, 3.974346, 3.879889, 3.930383, 4.001359, 
    4.134026, 3.923068, 3.900476, 3.863004, 3.922684, 3.988853, 4.351483, 
    4.204781, 4.320621, 7.920043, 4.544635, 4.473603, 4.080145, 4.088374, 
    3.853456,
  3.944897, 3.861458, 4.030285, 3.937043, 3.976325, 3.873581, 3.963225, 
    3.957992, 3.817767, 3.795911, 3.726904, 3.865148, 4.098183, 4.076849, 
    9.451921, 3.811332, 3.668489, 3.811529, 3.618815, 3.782974, 3.872181, 
    3.915739, 4.050651, 9.510299, 4.46232, 3.959151, 3.881984, 3.932582, 
    3.851061,
  3.823867, 4.146844, 11.96496, 3.923861, 3.728617, 3.674473, 3.986218, 
    3.81689, 3.74832, 3.770288, 9.842348, 14.72773, 10.38958, 3.534102, 
    3.725843, 3.862411, 3.589865, 3.462924, 3.432689, 3.666065, 3.890041, 
    3.911281, 3.660732, 4.250847, 9.446749, 3.442542, 3.697413, 3.786202, 
    4.06009,
  3.462525, 9.714795, 12.34819, 3.437921, 3.407514, 3.463205, 3.749433, 
    3.433265, 3.819202, 3.377622, 12.11267, 11.52564, 3.518436, 3.70469, 
    3.669248, 3.676431, 3.308367, 3.495304, 3.334153, 3.693307, 3.763031, 
    3.741152, 3.47233, 3.162376, 8.896646, 9.289168, 4.127048, 3.718527, 
    3.967968,
  3.346734, 6.424582, 8.489165, 9.166639, 3.28045, 3.079649, 3.461074, 
    3.192868, 3.213534, 3.162419, 4.417192, 3.154662, 4.306151, 3.262828, 
    3.279814, 3.694389, 3.416149, 3.48554, 3.515137, 3.789929, 3.515477, 
    3.861778, 3.368286, 8.297206, 8.478291, 8.931256, 3.536549, 3.607129, 
    3.852432,
  3.190302, 8.748127, 8.598197, 9.784511, 3.306857, 3.426537, 3.280895, 
    3.2013, 8.491368, 8.233953, 3.303932, 3.289718, 3.312943, 3.309985, 
    3.40817, 3.631974, 3.579544, 3.657517, 3.539551, 3.718251, 3.643723, 
    3.485451, 3.403467, 8.430391, 8.407042, 3.246675, 3.387213, 3.413406, 
    3.102407,
  9.941072, 10.2034, 10.86059, 9.36496, 14.30751, 3.48508, 5.273398, 
    3.528155, 3.788224, 3.514122, 4.04993, 3.52584, 3.169337, 3.315392, 
    3.511275, 3.349547, 3.500227, 3.6294, 3.573085, 3.361885, 3.452937, 
    3.358069, 8.5172, 7.574263, 3.241806, 3.379826, 3.134778, 3.254349, 
    8.933478,
  17.04294, 19.18196, 20.89131, 3.811861, 21.14993, 3.781086, 10.54798, 
    4.116045, 9.222888, 3.502119, 3.480253, 3.639374, 3.788913, 3.684109, 
    3.66345, 3.887252, 3.751604, 3.659064, 3.91035, 3.453437, 4.024704, 
    6.2445, 3.715603, 4.350075, 3.829098, 3.926389, 3.599743, 3.695969, 
    21.5905,
  21.32687, 16.65648, 17.88854, 17.25213, 11.97403, 13.42809, 12.27196, 
    31.26753, 8.968997, 10.21701, 3.341084, 3.769291, 3.767126, 3.83973, 
    3.807955, 3.703246, 3.812414, 3.533507, 3.706733, 3.775363, 11.82451, 
    12.28015, 12.38632, 3.730866, 3.825301, 4.021869, 3.917362, 4.121207, 
    10.28849,
  6.420385, 4.216809, 6.005682, 14.42303, 1.753146, 13.27746, 27.98412, 
    13.09059, 11.34089, 21.25572, 8.939497, 3.627133, 3.531458, 3.678192, 
    3.864844, 3.744547, 3.218771, 3.511888, 3.667216, 11.27147, 20.65945, 
    16.26377, 14.17427, 4.469598, 3.405205, 3.5141, 3.479134, 3.645145, 
    4.798005,
  5.402888, 13.71243, 13.26558, 26.55079, 27.90294, 30.1681, 14.07335, 
    30.90282, 13.37775, 6.54888, 10.78616, 20.05787, 29.08957, 3.154229, 
    2.917741, 3.388083, 3.979062, 4.46939, 4.227643, 26.96186, 21.7495, 
    27.55103, 23.09704, 26.45032, 14.76512, 3.288174, 3.83193, 3.910752, 
    4.175916,
  4.258328, 14.99212, 17.48242, 20.09841, 21.55565, 22.24979, 23.88414, 
    23.3321, 19.42969, 19.09633, 17.72355, 29.15338, 29.5917, 24.76481, 
    3.189342, 33.67865, 26.04653, 13.68272, 29.26419, 20.08663, 21.70513, 
    29.47783, 35.08366, 29.12443, 2.59019, 8.414856, 4.320223, 3.93939, 
    4.319108,
  3.338975, 3.286114, 14.50453, 2.192807, 13.89081, 25.48105, 22.1773, 
    22.16393, 21.83546, 21.57184, 14.41854, 13.2157, 21.75819, 26.14826, 
    25.86154, 26.59015, 23.55722, 23.89894, 25.68204, 25.74167, 22.05218, 
    24.55587, 22.93271, 22.54877, 26.45882, 22.19027, 22.35586, 24.0005, 
    3.11839,
  2.36072, 2.232137, 2.486619, 2.568626, 2.344075, 2.295451, 2.471391, 
    2.382453, 2.390175, 2.345577, 2.262931, 2.175778, 2.368063, 2.521156, 
    2.585221, 2.532338, 2.521052, 2.771684, 2.892035, 2.651999, 2.768883, 
    2.525065, 2.293117, 2.531285, 2.242146, 2.339462, 2.09494, 2.267562, 
    2.641243,
  47.00509, 47.00509, 47.00509, 47.00509, 47.00509, 47.00509, 47.00509, 
    47.207, 47.207, 47.207, 47.207, 47.207, 47.207, 47.207, 47.35126, 
    47.35126, 47.35126, 47.35126, 47.35126, 47.35126, 47.35126, 47.26274, 
    47.26274, 47.26274, 47.26274, 47.26274, 47.26274, 47.26274, 47.00509,
  43.41802, 43.26198, 43.2297, 43.19894, 43.23173, 43.14181, 43.07385, 
    43.03705, 43.1942, 43.04394, 42.98541, 43.05552, 43.08139, 43.53246, 
    43.88158, 44.17169, 44.44234, 44.21972, 43.94145, 43.71065, 43.79564, 
    43.60255, 43.82034, 44.40745, 44.26767, 43.91338, 44.39358, 44.09753, 
    43.48222,
  34.31173, 17.62353, 7.772996, 35.78193, 41.48267, 41.49949, 42.89697, 
    41.43308, 41.38667, 41.66811, 41.67223, 41.46978, 41.72201, 7.964752, 
    4.785087, 4.777347, 4.552975, 4.312444, 4.382721, 6.166889, 12.59647, 
    14.4838, 44.47932, 40.36126, 42.29098, 39.57077, 4.762288, 3.9568, 
    24.16419,
  4.361288, 4.714728, 4.749916, 4.233894, 4.309018, 4.02312, 4.09586, 
    3.883536, 3.912441, 4.183074, 4.328512, 3.839681, 3.602955, 3.818161, 
    4.102726, 3.988666, 3.897598, 3.820446, 3.667719, 3.885858, 4.180392, 
    4.192776, 4.03876, 4.069193, 3.785183, 3.566906, 3.667979, 3.71048, 
    3.932217,
  3.591743, 3.731552, 3.659863, 3.834902, 3.847799, 3.910193, 3.903333, 
    3.874974, 3.960241, 3.846503, 3.732418, 3.839593, 3.784921, 3.652741, 
    4.020271, 3.605739, 3.727224, 3.545761, 3.606998, 3.794217, 3.81216, 
    4.024345, 3.820562, 7.248759, 4.330713, 4.037424, 3.706614, 3.601245, 
    3.536268,
  3.639362, 3.803677, 3.914585, 3.861439, 3.869304, 3.916616, 3.687128, 
    3.565039, 3.67272, 3.792469, 3.768072, 3.846053, 3.903736, 3.613356, 
    8.859904, 4.030863, 3.835163, 3.889855, 3.804514, 3.853976, 3.759839, 
    3.739673, 3.972824, 8.710025, 4.268406, 3.850047, 3.756501, 3.628733, 
    3.558794,
  3.671089, 4.012972, 11.63802, 3.773257, 3.66773, 3.494874, 3.502003, 
    3.623757, 3.70066, 3.757786, 9.382825, 14.00719, 9.895658, 3.623048, 
    3.670224, 3.940018, 3.559848, 3.396999, 3.415107, 3.631811, 3.625233, 
    3.726732, 3.706743, 4.309098, 8.966111, 3.797353, 3.649904, 3.680139, 
    3.799315,
  3.484785, 9.653737, 11.94688, 3.771977, 3.40637, 3.596052, 3.641788, 
    3.526633, 3.31628, 3.608676, 11.89484, 11.30811, 3.70166, 3.353507, 
    3.29592, 3.457842, 3.42501, 3.39677, 3.492682, 3.594455, 3.692969, 
    3.865273, 3.556261, 3.358956, 8.859101, 8.761039, 3.442259, 3.51239, 
    3.854824,
  3.298866, 6.160888, 8.434052, 8.926915, 3.27112, 3.409948, 3.379484, 
    3.249834, 3.138885, 3.299453, 4.56195, 3.130016, 4.316838, 3.343702, 
    3.536328, 3.426655, 3.295448, 3.444016, 3.354187, 3.55823, 3.596699, 
    3.687744, 3.449866, 8.325864, 8.281964, 8.604132, 3.512689, 3.510839, 
    3.646696,
  3.041514, 8.630935, 8.342789, 9.841524, 3.398857, 3.319081, 3.286037, 
    3.170005, 8.462026, 8.283673, 3.244136, 3.273758, 3.358891, 3.287982, 
    3.314742, 3.372326, 3.291441, 3.562221, 3.535237, 3.580569, 3.530737, 
    3.466143, 3.255036, 8.444114, 8.315844, 3.217355, 3.250921, 3.270492, 
    3.03652,
  10.03063, 10.37877, 10.55742, 9.63239, 14.9585, 3.395489, 5.15769, 
    3.258547, 3.664075, 3.342825, 4.16545, 3.409747, 3.364542, 3.420861, 
    3.397936, 3.285661, 3.449412, 3.496249, 3.350706, 3.437526, 3.366874, 
    3.430092, 8.831871, 7.36871, 3.390548, 3.266041, 3.21741, 3.21391, 
    9.033566,
  17.56821, 20.05806, 22.14445, 3.643493, 22.08451, 3.716119, 10.64469, 
    3.769943, 9.720462, 3.316581, 3.599488, 3.589075, 3.719428, 3.795307, 
    3.76674, 3.797487, 3.586294, 3.786657, 3.49191, 3.408953, 3.687326, 
    6.352117, 3.698886, 4.371268, 3.616202, 3.664411, 3.426768, 3.497861, 
    22.93208,
  22.77159, 18.51805, 19.69564, 18.36106, 12.26649, 13.97128, 12.31452, 
    30.01598, 9.159367, 10.28255, 3.414062, 3.532921, 3.539192, 3.488049, 
    3.601582, 3.506472, 3.601328, 3.524866, 3.597698, 3.849004, 12.64213, 
    11.30001, 9.084694, 3.547216, 3.576727, 3.602456, 3.416848, 3.681121, 
    10.99291,
  6.813754, 4.253103, 6.093978, 22.01879, 1.90161, 13.6763, 28.4531, 14.2811, 
    12.27043, 9.726168, 9.243841, 3.892117, 3.821793, 3.839948, 3.890555, 
    3.786743, 3.799345, 3.617912, 3.607546, 11.48324, 15.19301, 14.65386, 
    15.59088, 4.54654, 3.631999, 3.49895, 3.591216, 3.650815, 5.432932,
  5.655741, 14.3637, 15.24894, 14.63072, 21.88419, 33.955, 11.03448, 
    35.26326, 14.22122, 7.266745, 8.172451, 21.13739, 32.81843, 4.078194, 
    4.171196, 4.087504, 4.093245, 4.03052, 4.12637, 30.34744, 16.54679, 
    25.63973, 25.9432, 30.71552, 24.08567, 3.74632, 3.562862, 3.843323, 
    3.79351,
  4.211899, 16.28345, 20.03632, 26.58307, 28.04645, 26.72468, 29.96821, 
    29.91189, 25.72614, 26.39638, 24.8932, 37.90231, 38.57235, 35.27555, 
    4.175857, 41.35753, 32.13757, 15.87314, 35.62113, 25.71491, 27.53022, 
    36.97559, 45.36838, 38.39294, 4.107834, 10.68332, 4.57786, 4.02182, 
    4.280853,
  5.264061, 5.385809, 24.98239, 4.260882, 18.22739, 43.88689, 37.78481, 
    37.64494, 37.39049, 37.235, 25.55986, 22.91653, 37.35707, 43.94092, 
    43.67566, 44.6829, 39.97056, 40.23317, 43.28332, 43.10358, 37.31806, 
    41.18439, 38.52766, 37.98093, 44.75806, 37.98307, 37.85838, 41.38931, 
    4.842242,
  39.6379, 41.04997, 39.32433, 41.67879, 40.5295, 40.30993, 41.70043, 
    41.47575, 41.73232, 41.78044, 41.9758, 42.13523, 41.9308, 42.06394, 
    41.90507, 41.68589, 41.68418, 41.75086, 41.79604, 41.73426, 41.88638, 
    39.60005, 36.63077, 37.39766, 35.53342, 35.36537, 35.391, 35.95628, 
    41.8296,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  10.06781, 10.30963, 10.37245, 9.950179, 10.25171, 10.25342, 10.24704, 
    10.36679, 10.20778, 10.22712, 10.71072, 10.31766, 10.17462, 10.49983, 
    10.49558, 10.56847, 10.45121, 10.47752, 10.00297, 9.959476, 10.07948, 
    10.20749, 9.874797, 10.10994, 10.1636, 10.55846, 10.46031, 10.51081, 
    10.29923,
  21.33254, 17.54087, 10.77614, 17.36137, 27.60639, 27.63409, 30.17433, 
    27.7312, 27.79449, 27.92349, 27.54135, 27.32893, 27.61736, 5.812678, 
    2.980455, 3.123223, 3.283215, 3.197704, 3.123408, 4.887712, 21.70844, 
    19.20755, 28.5282, 28.42415, 29.72311, 29.8378, 15.6193, 2.993301, 
    28.01747,
  3.641266, 3.660086, 4.231604, 3.748159, 3.982475, 3.942498, 3.904545, 
    3.650586, 3.659087, 3.567922, 3.489419, 3.332066, 3.084815, 3.300662, 
    3.863025, 3.763938, 3.443957, 3.271327, 3.489348, 3.602946, 3.511353, 
    3.289782, 3.402983, 3.482747, 3.512392, 3.270386, 3.345474, 3.699584, 
    3.685734,
  3.414323, 3.789241, 3.498008, 3.779015, 3.852454, 3.527755, 3.680082, 
    3.633424, 3.874781, 3.672975, 3.660796, 3.548215, 3.57187, 3.762647, 
    3.784957, 3.68486, 3.601735, 3.918074, 3.714533, 3.698895, 3.513701, 
    3.451171, 3.670374, 6.92707, 3.754934, 4.027737, 3.826754, 3.673887, 
    3.555152,
  3.565046, 3.531621, 3.743589, 3.867813, 3.589109, 3.739125, 3.834466, 
    3.66626, 3.622496, 3.725603, 3.525759, 3.608027, 4.20938, 3.976595, 
    8.065894, 3.769532, 3.731821, 3.600407, 3.662379, 3.649263, 3.448509, 
    3.606586, 3.73553, 7.889583, 4.075655, 3.880592, 3.767508, 3.720715, 
    3.498325,
  3.942025, 3.940371, 11.27313, 3.897967, 3.934367, 3.784591, 3.664937, 
    3.882538, 3.613128, 3.929311, 8.859979, 13.3902, 9.462267, 3.876194, 
    3.70536, 3.72437, 3.829572, 3.669921, 3.562486, 3.562336, 3.64634, 
    3.962029, 3.886373, 4.348446, 8.274636, 3.671387, 3.53213, 3.842062, 
    3.678894,
  3.693393, 9.387356, 9.670104, 3.750037, 3.587999, 3.429611, 3.32776, 
    3.684697, 3.371006, 3.822074, 12.07596, 11.46374, 3.697133, 3.59508, 
    3.410365, 3.505252, 3.620275, 3.433203, 3.666055, 3.725376, 3.881763, 
    3.748379, 3.494147, 3.374702, 8.638007, 8.758164, 3.595792, 3.752937, 
    3.657124,
  3.353219, 6.389432, 8.540174, 8.494987, 3.364108, 3.341235, 3.255082, 
    3.505634, 3.236038, 3.404618, 4.607475, 3.655158, 4.107643, 3.289246, 
    3.474776, 3.263751, 3.336441, 3.444605, 3.403574, 3.617547, 3.713014, 
    3.385672, 3.178258, 8.663651, 8.093015, 8.734487, 3.635257, 3.36479, 
    3.465219,
  3.12014, 8.402856, 8.242336, 9.637259, 3.506828, 3.62834, 3.504736, 
    3.445772, 8.520418, 8.135445, 3.247473, 3.315686, 3.129511, 3.36816, 
    3.403229, 3.513544, 3.504243, 3.511133, 3.476398, 3.413405, 3.421702, 
    3.355357, 3.273948, 8.353836, 8.361552, 3.337653, 3.262424, 3.257322, 
    3.107685,
  10.15848, 10.56538, 10.53348, 9.797899, 15.11613, 3.248322, 5.283098, 
    3.363175, 3.692744, 3.385587, 4.554461, 3.357669, 3.368163, 3.259391, 
    3.218551, 3.42132, 3.288456, 3.36222, 3.324572, 3.319499, 3.151019, 
    3.361838, 8.883085, 7.65364, 3.545639, 3.225646, 3.059128, 3.208666, 
    8.863873,
  18.23812, 20.89123, 22.94378, 3.607815, 22.84093, 3.542257, 10.90097, 
    3.453624, 9.826267, 3.242689, 3.646268, 3.549084, 3.779115, 3.858719, 
    3.773204, 3.890577, 3.659426, 3.857513, 3.383864, 3.567827, 3.538277, 
    6.523942, 3.681404, 4.361062, 3.798398, 3.501698, 3.627276, 3.366014, 
    23.72788,
  24.09764, 20.42845, 21.06888, 19.59613, 12.79473, 14.39093, 12.6885, 
    17.96437, 8.374874, 10.22642, 3.469686, 3.516647, 3.461391, 3.530388, 
    3.681937, 3.618462, 3.571718, 3.774199, 3.471538, 3.973617, 10.57937, 
    11.82847, 9.29106, 3.527991, 3.699153, 3.516746, 3.775223, 3.621475, 
    11.43572,
  7.806798, 4.138757, 6.134325, 11.18061, 2.103832, 15.56828, 21.28419, 
    15.4277, 13.39498, 10.93934, 8.032671, 3.659639, 3.675356, 3.774322, 
    3.720161, 3.748963, 3.735933, 3.785663, 3.5605, 12.19872, 11.80634, 
    14.23763, 13.47598, 4.703897, 3.744191, 3.719102, 3.796106, 3.800264, 
    5.374824,
  6.207018, 12.36987, 15.22383, 16.20746, 13.67617, 22.61468, 9.644892, 
    39.04796, 13.20683, 8.620715, 8.044651, 13.64735, 18.47056, 4.116431, 
    4.043595, 3.977867, 4.166586, 4.090584, 4.302946, 30.34043, 11.90335, 
    12.09083, 19.66936, 29.90433, 10.53675, 3.717414, 4.029939, 4.296762, 
    4.278459,
  4.612814, 11.9985, 17.44275, 10.38926, 21.56886, 21.25337, 35.71466, 
    34.74107, 27.32059, 30.07104, 28.91668, 45.57052, 46.49475, 41.9038, 
    19.20038, 43.91259, 32.34013, 18.39344, 41.07797, 13.65606, 17.55307, 
    44.17083, 53.99283, 46.28572, 4.945357, 11.60767, 5.371981, 4.919231, 
    4.811394,
  5.49254, 5.651546, 29.62201, 5.200398, 35.4924, 51.78225, 50.90521, 
    52.06754, 51.98355, 51.26308, 37.30087, 33.33862, 51.85875, 61.14124, 
    60.68857, 61.44812, 54.18727, 52.66937, 57.91113, 57.32364, 51.71809, 
    57.29054, 53.37889, 52.64061, 62.23112, 52.61938, 52.39771, 58.84809, 
    5.826498,
  79.2588, 76.23703, 77.19462, 79.83168, 76.67937, 76.62772, 79.38733, 
    80.95038, 81.46128, 82.16718, 82.25, 82.31062, 82.07681, 81.92217, 
    82.06875, 82.25754, 82.22446, 81.97395, 81.88003, 81.93622, 81.79897, 
    77.49718, 72.02083, 72.92411, 69.42635, 68.81229, 69.17027, 70.47285, 
    81.91506,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  8.207256, 10.0288, 7.99017, 7.568598, 9.309444, 9.259027, 10.40392, 
    9.342898, 9.505941, 9.632073, 9.441983, 9.373121, 9.316809, 6.802946, 
    3.190262, 4.785258, 1.131119, 1.165537, 1.001179, 2.732987, 7.420048, 
    7.318288, 8.691492, 9.070669, 10.82669, 11.03732, 10.68446, 10.56755, 
    10.96981,
  3.717459, 3.347145, 3.275454, 3.400887, 2.97375, 3.337593, 2.966784, 
    3.605263, 3.407352, 3.071518, 3.067331, 3.049931, 2.621258, 3.064583, 
    3.151114, 2.893444, 3.225947, 3.399968, 3.467685, 3.846123, 3.377921, 
    3.474773, 3.029948, 2.744399, 2.55506, 9.647677, 14.49294, 3.034203, 
    3.278522,
  3.243275, 2.990554, 3.29349, 3.122252, 3.543504, 3.099396, 3.45611, 
    3.509915, 3.574297, 3.912737, 3.821485, 3.610381, 3.598147, 3.496101, 
    3.789952, 3.860787, 3.692404, 3.8653, 4.151141, 3.753389, 3.740206, 
    3.766736, 3.466482, 6.217369, 3.644935, 3.253769, 3.006925, 3.263073, 
    3.162447,
  3.294076, 3.908727, 3.877239, 3.661117, 3.495336, 3.692113, 3.312955, 
    3.659133, 3.960662, 3.892213, 3.935293, 3.885657, 3.879363, 3.935404, 
    7.388865, 3.905109, 3.862436, 3.91192, 3.662843, 3.428011, 3.511194, 
    3.95246, 3.866337, 7.34412, 4.3292, 3.906341, 3.964477, 3.749019, 3.459183,
  3.966131, 4.18679, 11.25269, 4.039012, 3.980976, 4.046475, 3.892925, 
    4.042104, 3.702626, 3.846639, 9.042244, 13.08361, 9.393846, 4.037091, 
    3.781149, 3.815426, 3.881052, 3.6226, 3.411772, 3.723072, 3.881524, 
    3.776348, 3.887493, 4.158095, 8.241242, 3.91399, 3.836318, 3.97145, 3.8913,
  3.695997, 9.334023, 10.83084, 3.79668, 3.562694, 3.791313, 3.7272, 
    3.896931, 3.479294, 3.912553, 11.44284, 11.59082, 3.943803, 3.718443, 
    3.665551, 3.734051, 3.747056, 3.543619, 3.864798, 3.711821, 4.086782, 
    3.868855, 3.615122, 3.844854, 8.744532, 8.938788, 3.775171, 4.073379, 
    3.592957,
  3.353571, 6.21144, 9.013899, 8.800789, 3.267844, 3.300543, 3.283633, 
    3.509015, 3.24568, 3.36619, 4.581576, 3.699583, 4.118513, 3.309355, 
    3.536814, 3.366899, 3.751721, 3.686109, 3.801296, 3.719811, 4.03373, 
    3.71311, 3.238358, 8.548631, 8.535704, 8.673987, 3.806253, 3.82039, 
    3.407928,
  3.23827, 8.319117, 8.121634, 9.993693, 3.593557, 3.657191, 3.549173, 
    3.49974, 8.608858, 8.139314, 3.48091, 3.473274, 3.65677, 3.638784, 
    3.585654, 3.650481, 3.63186, 3.75653, 3.693013, 3.738704, 3.640287, 
    3.546712, 3.20966, 8.164235, 8.375542, 3.356811, 3.437966, 3.327031, 
    3.302691,
  9.87033, 10.23562, 10.52158, 9.748078, 15.32731, 3.319685, 5.093399, 
    3.291493, 3.753616, 3.357207, 4.783806, 3.440593, 3.376664, 3.261026, 
    3.262197, 3.278097, 3.24708, 3.555046, 3.294425, 3.45071, 3.289405, 
    3.507437, 8.981514, 7.470119, 3.592278, 3.388705, 3.505288, 3.131666, 
    8.912589,
  18.79504, 21.36793, 23.58884, 3.440795, 23.77795, 3.549949, 11.25973, 
    3.290038, 9.47822, 3.360876, 3.717684, 3.497666, 3.593436, 3.710073, 
    3.77193, 3.818357, 3.758261, 3.898856, 3.528942, 3.522373, 3.912834, 
    6.803573, 3.762353, 4.310958, 3.572999, 3.760216, 3.928047, 3.601358, 
    24.5563,
  25.31771, 21.3885, 22.21191, 20.39403, 13.34363, 15.15663, 13.10202, 
    17.61603, 9.189785, 10.87638, 3.625542, 3.606702, 3.564163, 3.570833, 
    3.789462, 3.681687, 3.791456, 3.743671, 3.563538, 3.909212, 11.38967, 
    12.38427, 9.789193, 3.761185, 3.692599, 3.718527, 3.749333, 3.762103, 
    11.79674,
  8.395414, 4.137861, 6.379588, 11.0263, 2.249986, 15.83882, 10.55409, 
    16.61084, 14.29836, 11.68246, 8.145136, 3.989533, 3.869372, 3.776348, 
    3.731889, 3.765002, 3.79399, 3.689878, 3.856785, 13.09292, 11.89373, 
    14.74358, 13.71684, 4.750682, 3.831369, 4.006458, 3.858976, 4.172945, 
    5.34117,
  6.618307, 13.6469, 15.298, 16.0422, 14.82098, 12.84583, 9.074828, 23.78996, 
    9.981394, 8.268737, 8.157477, 8.203937, 4.175727, 4.217169, 4.290664, 
    4.207808, 4.081609, 4.184828, 4.259978, 11.78154, 11.36257, 10.98482, 
    7.924463, 10.06155, 5.862984, 4.153483, 4.353708, 4.25402, 4.35544,
  5.038737, 8.420995, 12.56352, 8.368599, 9.674547, 9.149107, 26.46828, 
    23.99571, 12.07325, 11.58191, 10.39726, 47.60344, 47.86214, 31.78186, 
    6.602672, 5.467993, 16.17012, 20.565, 32.74376, 8.537551, 8.350493, 
    33.77294, 49.47227, 42.1545, 5.20697, 10.30813, 4.573065, 4.914161, 
    4.858248,
  6.278323, 6.889002, 14.91238, 7.125478, 14.7873, 73.14732, 65.23597, 
    62.69674, 62.84936, 63.01077, 33.66816, 31.13625, 61.83462, 75.13591, 
    76.08392, 65.74132, 55.36371, 46.48162, 55.69169, 57.07106, 54.54035, 
    64.8662, 58.62131, 64.39354, 72.3419, 69.97951, 70.52843, 62.20162, 
    6.135671,
  68.74249, 70.39649, 75.34229, 80.95261, 79.26311, 81.17737, 82.98769, 
    81.48383, 82.01278, 81.73141, 81.46447, 80.54872, 79.22939, 75.26381, 
    74.80094, 75.28767, 73.63874, 72.42231, 73.32722, 73.13818, 72.79537, 
    70.16503, 72.04516, 75.82249, 74.40457, 76.41811, 76.54639, 71.75094, 
    71.32865,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  8.954749, 2.07305, 2.57466, 2.709603, 2.25497, 2.503206, 2.100795, 
    2.303388, 2.948401, 2.345654, 2.591513, 2.577687, 2.131613, 2.044556, 
    2.193775, 2.352979, 2.253003, 2.483256, 2.954404, 2.648228, 2.513153, 
    2.662241, 2.693469, 2.845018, 2.29283, 15.43419, 22.69668, 16.43883, 
    12.5816,
  3.079673, 3.361527, 3.359768, 3.404166, 3.244427, 3.157948, 3.038833, 
    3.419692, 3.582919, 3.376288, 3.432326, 3.431846, 3.496667, 3.330546, 
    3.482798, 3.06778, 3.099757, 3.299412, 3.305459, 3.093499, 3.250289, 
    3.301196, 3.558179, 8.886765, 4.224158, 3.722461, 3.196048, 3.518064, 
    3.30756,
  3.882203, 4.076994, 3.74076, 3.990009, 3.633744, 3.9717, 4.084915, 
    3.571853, 3.756551, 4.277793, 3.965776, 3.807415, 4.537826, 4.26976, 
    10.45502, 3.999001, 3.702674, 3.794469, 3.941078, 3.56096, 3.323897, 
    3.486602, 3.933547, 10.39358, 4.385761, 3.999719, 3.758258, 3.755826, 
    3.680813,
  3.744319, 4.401262, 11.56482, 4.356335, 4.011292, 3.855125, 4.20785, 
    4.086404, 4.314359, 4.332314, 8.354263, 12.18284, 9.457981, 4.193636, 
    3.961678, 3.844724, 3.933783, 4.058936, 3.694156, 3.619084, 3.639742, 
    4.042634, 3.882012, 4.261868, 8.222835, 3.621228, 3.884647, 4.144731, 
    4.22526,
  3.547275, 9.402644, 9.585195, 4.032499, 4.017748, 4.217079, 3.842115, 
    3.846157, 3.813982, 4.065452, 11.29434, 11.80803, 3.879341, 4.147933, 
    3.833889, 3.463091, 3.775755, 3.772486, 3.833218, 3.803063, 4.106861, 
    3.651666, 3.830302, 3.92455, 8.312923, 9.005594, 3.984306, 3.817648, 
    3.718852,
  3.660246, 6.51464, 9.22526, 9.151155, 3.741404, 3.59514, 3.511004, 
    3.617532, 3.311936, 3.736107, 4.685037, 3.703716, 4.351312, 3.430171, 
    3.335571, 3.262824, 3.440468, 3.609358, 4.084257, 3.872289, 3.969399, 
    3.619003, 3.332101, 8.578269, 8.904963, 9.090558, 3.82754, 4.023759, 
    3.482542,
  3.190102, 8.803493, 8.454676, 10.14264, 3.568033, 3.286018, 3.244746, 
    3.360569, 8.710108, 8.577391, 3.605627, 3.390007, 3.44909, 3.526023, 
    3.50042, 3.581457, 3.568253, 3.779721, 3.69309, 3.801732, 3.607781, 
    3.6493, 3.289777, 8.287563, 8.483267, 3.524786, 3.593329, 3.493928, 
    3.328434,
  9.750155, 10.29642, 10.58801, 9.934576, 15.17355, 3.271857, 5.029364, 
    3.089355, 3.693623, 3.264678, 4.441254, 3.43826, 3.301121, 3.378752, 
    3.448126, 3.422355, 3.275042, 3.771736, 3.405323, 3.494181, 3.470312, 
    3.321353, 8.997711, 7.659001, 3.381881, 3.219955, 3.325037, 3.114908, 
    8.919165,
  19.407, 21.77885, 23.57712, 3.539638, 24.29902, 3.128384, 11.07612, 
    3.215742, 9.131583, 3.406367, 3.534051, 3.467889, 3.896413, 3.677752, 
    3.627238, 3.961713, 3.777437, 3.813097, 3.570667, 3.777452, 3.695249, 
    6.705717, 3.444611, 4.096391, 3.835057, 3.633659, 3.627367, 3.510611, 
    24.5748,
  25.87362, 21.814, 22.70634, 20.94533, 13.99932, 15.94217, 12.93494, 
    10.85073, 8.750209, 10.93548, 3.631428, 3.680255, 3.706163, 3.68196, 
    3.718477, 3.877793, 4.149929, 3.93915, 3.810457, 3.814798, 11.61929, 
    12.28819, 9.97984, 3.742051, 3.709793, 4.079958, 3.920766, 3.987986, 
    11.98357,
  8.185322, 4.128829, 6.707524, 11.12386, 2.358731, 16.73757, 9.708811, 
    17.3283, 14.9468, 11.57462, 8.247165, 4.068477, 3.862055, 3.866282, 
    3.854724, 3.735801, 3.820976, 3.88736, 3.793909, 13.65651, 12.8303, 
    14.50419, 14.03579, 4.917433, 3.89262, 4.02083, 4.019463, 3.903403, 
    5.382471,
  6.96819, 14.3268, 15.28006, 16.59464, 15.24851, 13.51344, 9.621478, 
    12.9506, 9.158701, 8.159802, 7.894991, 7.495394, 4.22742, 4.204645, 
    4.10243, 4.22623, 4.139567, 4.328401, 4.404181, 10.35142, 11.51499, 
    11.27352, 7.94805, 7.698545, 6.001417, 4.575519, 4.492835, 4.491659, 
    4.623472,
  5.475673, 9.148862, 10.9201, 8.950768, 9.372644, 9.240079, 9.450485, 
    9.431724, 10.15784, 9.454295, 9.050331, 17.81958, 25.38977, 8.602552, 
    5.569464, 6.06113, 12.32584, 17.50919, 14.00767, 9.32409, 8.44162, 
    21.82711, 43.75837, 23.45077, 5.666492, 10.19251, 5.075019, 5.292585, 
    5.283402,
  6.190205, 7.239244, 11.84624, 7.086466, 7.145331, 59.70623, 43.59563, 
    47.21478, 36.46804, 35.86074, 17.23511, 14.78791, 29.94696, 59.01356, 
    58.16896, 59.48733, 34.62516, 34.18643, 51.18197, 55.30213, 29.55235, 
    49.74183, 36.45308, 56.67838, 46.5327, 68.29192, 74.0123, 37.76799, 
    6.518102,
  60.01873, 59.80387, 58.95005, 60.63799, 54.0267, 60.93587, 60.41843, 
    58.46654, 60.23501, 60.5098, 60.65059, 60.57858, 60.45856, 60.40287, 
    60.37328, 60.3328, 60.37081, 60.52739, 60.47021, 60.34467, 60.41519, 
    56.46355, 57.99541, 64.69775, 66.92129, 68.21605, 68.97215, 64.18209, 
    60.21944,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  3.937644, 4.059346, 4.093653, 3.796766, 3.408573, 3.431779, 3.745096, 
    3.323938, 3.482696, 3.529356, 3.343939, 3.22032, 3.372946, 4.092729, 
    4.173648, 4.276246, 4.449315, 3.769369, 0.3353124, 3.722301, 4.254342, 
    4.175943, 4.183346, 3.78994, 4.455185, 4.557441, 4.301361, 4.293293, 
    4.222141,
  25.89766, 23.12887, 2.648357, 3.164365, 3.235786, 3.135711, 21.7079, 
    2.690239, 3.192972, 3.539798, 3.313538, 2.835512, 3.029584, 3.054555, 
    3.138111, 2.945148, 2.734381, 2.543055, 2.768495, 3.018845, 2.851647, 
    2.793343, 2.922034, 2.529798, 13.36954, 25.29247, 26.029, 26.40083, 
    25.52853,
  3.15876, 3.00861, 2.887995, 2.946648, 2.993936, 3.507545, 3.587666, 
    3.802114, 3.483894, 3.443065, 3.277625, 3.606665, 3.454617, 3.658597, 
    3.492354, 3.706738, 3.854908, 3.460141, 3.492182, 3.65197, 3.708552, 
    3.727093, 4.002427, 9.955, 3.830147, 3.593657, 3.16708, 3.462798, 3.28865,
  3.65443, 3.930085, 4.056864, 3.860172, 3.80522, 3.76532, 3.971638, 
    3.877305, 3.936738, 4.021633, 4.177948, 4.015319, 4.357781, 4.259067, 
    11.62798, 4.358775, 4.07409, 4.066918, 3.753227, 3.586463, 3.500771, 
    3.598279, 3.826535, 9.860829, 4.266181, 3.698683, 3.786429, 3.631292, 
    3.894991,
  3.911689, 4.142035, 11.37072, 4.305263, 3.928467, 4.005132, 3.874589, 
    3.864589, 4.06596, 4.341518, 8.686159, 12.72344, 10.431, 4.309492, 
    3.980946, 4.115707, 3.868435, 3.943758, 3.836653, 3.942298, 4.007658, 
    4.246287, 3.744435, 4.392256, 8.550149, 3.736569, 3.88273, 4.209903, 
    4.024292,
  3.402113, 9.381686, 9.622629, 3.773943, 4.024459, 4.038765, 3.706077, 
    3.762275, 3.574021, 4.252287, 11.54507, 11.72849, 3.894633, 3.712766, 
    3.622651, 3.698479, 3.810027, 3.780233, 4.007181, 3.749032, 3.900777, 
    3.464803, 3.309209, 3.768842, 8.726899, 8.866632, 3.850883, 3.724762, 
    3.550537,
  3.29321, 6.262545, 9.219871, 9.050168, 3.692295, 3.643603, 3.381145, 
    3.379659, 3.386404, 3.803535, 4.740543, 3.725296, 4.203604, 3.217853, 
    3.281401, 3.401196, 3.830401, 3.748721, 4.050678, 3.797657, 3.915555, 
    3.521008, 3.328845, 8.864221, 8.896483, 9.14404, 3.775931, 4.041829, 
    3.546451,
  3.221054, 8.578339, 8.420505, 10.19775, 3.63319, 3.225121, 3.231062, 
    3.227568, 8.632911, 8.235376, 3.348819, 3.410092, 3.605053, 3.505699, 
    3.398328, 3.474182, 3.658822, 3.840991, 3.609741, 3.622594, 3.597298, 
    3.474097, 3.282867, 8.377344, 8.593021, 3.617082, 3.521437, 3.492408, 
    3.373537,
  9.675445, 10.16744, 9.974483, 9.479559, 15.07264, 3.281913, 5.027051, 
    3.022149, 3.593815, 3.242311, 4.267965, 3.304044, 3.346693, 3.42616, 
    3.356114, 3.498481, 3.470304, 3.663248, 3.376044, 3.397816, 3.237648, 
    3.229314, 9.03769, 7.589344, 3.297546, 3.136917, 3.216679, 3.162153, 
    8.596167,
  19.16027, 21.58859, 23.44779, 3.35374, 23.87273, 3.113803, 10.50242, 
    3.205509, 8.997926, 3.346938, 3.385014, 3.346428, 3.443252, 3.536772, 
    3.556845, 3.876737, 3.836796, 3.913261, 3.528102, 3.400731, 3.243321, 
    6.733939, 3.432934, 4.082909, 3.444126, 3.398406, 3.410426, 3.21179, 
    24.62262,
  25.34484, 21.59144, 22.66638, 20.60284, 13.61575, 15.89596, 12.50964, 
    9.89185, 7.236308, 10.65654, 3.56615, 3.852645, 3.601771, 3.737119, 
    4.204741, 4.069931, 4.09715, 3.856576, 3.671053, 3.925372, 11.78776, 
    12.04897, 9.525427, 3.621367, 3.661266, 4.088455, 4.040409, 3.703887, 
    11.63838,
  8.341124, 4.198357, 6.75784, 11.13409, 2.289093, 16.83676, 9.425503, 
    16.84243, 14.40416, 11.69723, 7.825489, 3.87232, 3.712683, 3.745603, 
    3.681738, 3.637065, 3.761827, 3.837428, 3.974648, 13.38368, 12.563, 
    14.66421, 13.65813, 4.614745, 3.80795, 3.940376, 4.048466, 4.039404, 
    5.641547,
  6.713972, 13.44479, 14.9993, 16.00343, 15.02882, 13.40419, 9.130196, 
    12.04097, 8.361918, 7.734684, 7.693208, 7.339312, 4.144758, 4.219711, 
    4.00974, 4.073275, 4.012276, 4.066431, 4.13551, 10.27823, 11.60113, 
    10.75518, 7.794538, 7.430983, 5.723678, 4.241274, 4.278132, 4.214406, 
    4.528553,
  5.093886, 8.450298, 9.947189, 8.526764, 8.947346, 8.818552, 8.846985, 
    8.863581, 9.113718, 8.989362, 8.581644, 13.18615, 13.15917, 8.073422, 
    5.060508, 4.959878, 11.50827, 15.9406, 12.70121, 8.767578, 7.884612, 
    13.77875, 5.230107, 13.23477, 5.336149, 10.24907, 5.058186, 4.879091, 
    4.818976,
  6.028561, 6.916415, 11.59007, 6.824832, 7.048464, 48.80408, 19.39706, 
    17.4463, 18.92422, 17.98593, 13.50359, 12.76028, 18.76376, 49.28145, 
    53.83068, 14.55631, 27.46205, 19.48911, 12.47585, 39.18582, 28.18076, 
    45.0043, 34.30557, 42.08452, 12.0874, 65.95777, 71.16652, 13.39094, 
    6.345264,
  60.06652, 49.63877, 48.94567, 50.07318, 29.84829, 52.32514, 59.37254, 
    14.16331, 59.7022, 60.14271, 60.23723, 60.15394, 60.13311, 60.14705, 
    60.15989, 60.18831, 60.2118, 60.33089, 60.37086, 60.35817, 60.46848, 
    51.4199, 52.35069, 61.93383, 71.22865, 66.34698, 72.34645, 60.49735, 
    60.1994,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  2.493829, 2.492429, 2.471442, 2.121521, 2.404775, 2.31636, 2.303638, 
    2.319246, 2.247494, 2.294985, 2.479152, 2.232728, 2.386821, 2.503096, 
    2.581967, 2.679867, 2.772909, 2.766962, 2.653347, 2.494684, 2.640127, 
    2.681441, 2.541608, 2.425219, 2.361829, 2.705937, 2.799138, 2.628233, 
    2.432264,
  25.31001, 25.43644, 26.39618, 24.62702, 22.29401, 22.23883, 24.42179, 
    22.20764, 22.19766, 22.25149, 22.28055, 22.30941, 22.43784, 26.35361, 
    26.54538, 26.4811, 26.41731, 26.36156, 9.725116, 25.16517, 25.21126, 
    25.51568, 26.25275, 24.506, 26.58585, 26.79025, 26.59775, 26.60295, 
    26.43914,
  32.34137, 33.31211, 3.197665, 3.655804, 3.828381, 4.19121, 33.64717, 
    4.166249, 3.350198, 4.188274, 3.91094, 3.851656, 3.005204, 3.385782, 
    3.43325, 3.552738, 3.108695, 3.343101, 3.670105, 4.002286, 4.255373, 
    4.054714, 4.087315, 4.173829, 29.23114, 31.94189, 32.45732, 32.66183, 
    33.08733,
  3.972982, 3.879125, 3.686785, 3.780803, 3.503103, 3.540745, 3.794511, 
    3.837054, 4.069533, 4.060327, 3.89285, 3.670757, 3.721102, 3.735834, 
    3.643999, 3.712911, 3.678112, 3.746373, 4.068103, 4.305541, 4.169703, 
    4.0704, 3.960535, 10.78808, 4.477331, 3.897174, 3.986733, 3.407463, 
    3.467773,
  3.635273, 3.850078, 3.921905, 3.625703, 3.574487, 3.567466, 3.656923, 
    3.769175, 3.735707, 4.154986, 3.943169, 3.984022, 4.273484, 4.032111, 
    12.51924, 4.06794, 4.148509, 3.938031, 4.049659, 3.834908, 3.88029, 
    3.774955, 3.665455, 10.77459, 4.234612, 3.734466, 3.693546, 3.748677, 
    3.532352,
  3.774355, 3.875211, 12.22545, 3.944428, 3.857469, 3.927598, 3.850542, 
    3.801685, 3.757984, 4.244765, 8.968526, 13.49369, 10.10252, 4.185449, 
    4.126674, 3.799822, 3.792712, 3.356117, 3.640818, 3.796725, 3.796721, 
    3.713194, 3.889997, 4.703434, 8.413291, 3.605881, 3.478864, 3.780583, 
    3.691799,
  3.259914, 9.512133, 9.80442, 3.826005, 3.690653, 3.767147, 3.874214, 
    3.903077, 3.538962, 4.269962, 11.55302, 11.26896, 3.833797, 3.699279, 
    3.445367, 3.5409, 3.636744, 3.492462, 4.131402, 3.676936, 3.810775, 
    3.44773, 3.15491, 3.734714, 9.104248, 8.98305, 3.628086, 4.015934, 
    3.405522,
  3.068291, 6.040157, 9.495571, 8.970817, 3.606194, 3.771368, 3.258763, 
    3.421397, 3.492193, 3.52643, 4.730158, 3.65137, 4.164867, 3.357155, 
    3.694999, 3.513344, 3.804169, 3.913147, 3.810285, 3.681695, 3.794073, 
    3.244341, 3.327145, 9.039392, 8.589607, 9.016556, 3.893803, 3.62863, 
    3.399747,
  3.133631, 8.421246, 8.424748, 10.00065, 3.496727, 3.108543, 3.075403, 
    3.148755, 8.493208, 8.136639, 3.073031, 3.174907, 3.185341, 3.442653, 
    3.487926, 3.564032, 3.563344, 3.700133, 3.576129, 3.600212, 3.546476, 
    3.284683, 3.23553, 8.562027, 8.713123, 3.42483, 3.482408, 3.337482, 
    3.200824,
  9.69042, 9.952655, 9.704674, 9.53069, 14.92811, 3.094155, 5.041256, 
    2.987249, 3.310392, 3.252799, 4.282717, 3.144106, 3.439252, 3.350933, 
    3.194822, 3.328511, 3.333667, 3.304145, 3.258198, 3.214577, 3.165806, 
    3.241184, 8.82091, 7.341235, 3.405256, 3.157803, 3.004761, 3.135985, 
    8.459505,
  18.1372, 20.99388, 23.23062, 3.178717, 23.26535, 3.07498, 10.15158, 
    3.117439, 9.028521, 3.142299, 3.301565, 3.27986, 3.154203, 3.267301, 
    3.325469, 3.518512, 3.55398, 3.896832, 3.298203, 3.419491, 3.378799, 
    6.165493, 3.369141, 4.135873, 3.316592, 3.278853, 3.315455, 3.061148, 
    23.88241,
  24.49442, 20.6781, 21.26427, 20.00345, 13.08182, 15.09585, 12.1964, 
    9.561179, 6.85343, 10.61206, 3.504281, 3.498742, 3.533332, 3.615898, 
    3.530036, 3.882113, 3.755616, 3.949048, 3.618906, 3.841248, 12.34305, 
    11.81472, 9.073066, 3.323836, 3.505931, 3.518508, 3.96582, 3.613935, 
    11.14605,
  6.676662, 4.276265, 6.411341, 10.60175, 2.14837, 15.69227, 8.990959, 
    15.75063, 13.56788, 11.15378, 7.464084, 3.885058, 3.847086, 3.529095, 
    3.847732, 3.638807, 3.699895, 3.956119, 3.8552, 12.6887, 11.4706, 
    13.9879, 13.00508, 4.479545, 3.729004, 3.838614, 3.854257, 3.887195, 
    5.360427,
  6.30231, 12.36273, 13.63856, 14.47003, 13.88133, 12.69853, 8.451757, 
    11.12163, 7.62409, 7.057515, 7.068615, 6.774438, 4.16987, 3.743387, 
    3.733598, 3.683196, 3.996392, 4.091352, 4.002153, 9.526365, 11.02099, 
    10.10777, 7.188038, 6.955253, 5.413029, 3.98207, 3.995911, 4.022892, 
    4.333362,
  4.845712, 7.441669, 8.747224, 7.343784, 7.995854, 7.623162, 7.717582, 
    7.876446, 7.809305, 7.765766, 7.634646, 11.30926, 11.84769, 7.139699, 
    4.927088, 4.813725, 9.829248, 15.09042, 10.97423, 7.910495, 6.977406, 
    11.6187, 4.819983, 11.53851, 4.174925, 8.772791, 4.158764, 4.347393, 
    4.486021,
  5.054276, 5.909121, 9.01218, 5.66084, 5.075035, 6.080107, 14.70819, 13.042, 
    13.9666, 14.06842, 10.19355, 10.01803, 13.9156, 10.07534, 19.13399, 
    5.147627, 10.4062, 10.85617, 6.88878, 8.737472, 21.56528, 19.82151, 
    19.29653, 29.13211, 5.396719, 52.01799, 56.30433, 9.183852, 4.950733,
  55.37937, 13.07278, 34.20408, 20.19646, 23.62682, 24.82287, 39.24474, 
    23.30175, 35.10054, 61.29577, 61.15277, 60.70659, 60.4595, 60.30219, 
    60.51845, 60.81598, 60.67836, 60.70415, 60.62838, 60.35335, 60.20845, 
    51.36092, 50.71568, 58.62269, 70.28262, 70.31542, 73.93369, 61.35513, 
    58.23784,
  20.90129, 20.90129, 20.90129, 20.90129, 20.90129, 20.90129, 20.90129, 
    21.08593, 21.08593, 21.08593, 21.08593, 21.08593, 21.08593, 21.08593, 
    20.77342, 20.77342, 20.77342, 20.77342, 20.77342, 20.77342, 20.77342, 
    20.7932, 20.7932, 20.7932, 20.7932, 20.7932, 20.7932, 20.7932, 20.90129,
  33.09964, 33.03193, 33.05904, 32.93226, 32.84799, 32.79695, 32.80107, 
    32.89754, 32.89782, 33.04958, 33.13911, 33.24326, 33.28473, 33.36491, 
    33.41805, 33.71605, 33.48211, 33.41721, 33.14462, 33.18063, 33.25198, 
    33.28024, 33.2229, 33.60783, 33.7056, 33.58025, 33.61534, 33.41937, 
    33.22408,
  41.64544, 41.62994, 43.15599, 40.20401, 36.5337, 36.49542, 39.96232, 
    36.56533, 36.61996, 36.71468, 36.6777, 36.64285, 36.93496, 43.02042, 
    43.30708, 43.14603, 43.2559, 43.13552, 42.07249, 41.60227, 40.69778, 
    39.49614, 39.07571, 37.90266, 43.09324, 43.27242, 43.38786, 43.44473, 
    43.34778,
  43.61283, 43.69456, 10.47307, 4.342847, 10.80238, 8.302503, 43.03923, 
    8.575305, 4.038308, 4.611137, 4.539783, 4.301235, 4.039899, 4.061869, 
    4.272611, 4.156531, 4.086718, 3.795734, 4.347197, 4.559931, 4.26293, 
    4.321833, 3.893597, 3.806245, 25.0619, 35.62947, 39.21054, 41.44508, 
    42.93018,
  3.819046, 3.990843, 3.950485, 3.927265, 3.922746, 3.823899, 3.808903, 
    3.990541, 3.949894, 4.112357, 4.022285, 3.938796, 3.986913, 3.780794, 
    3.891655, 4.026657, 4.015522, 3.985815, 4.05906, 3.926541, 3.846284, 
    3.986323, 3.798586, 8.057822, 4.339913, 3.651972, 3.641747, 3.445499, 
    3.746606,
  3.634842, 3.590599, 3.800956, 3.55193, 3.603643, 3.747187, 3.716654, 
    3.936337, 3.755795, 4.078915, 3.788451, 3.967173, 4.091709, 3.903577, 
    14.10535, 3.805816, 3.985785, 3.835906, 3.831385, 3.942745, 3.866541, 
    3.829321, 3.81178, 10.41127, 4.247932, 3.91557, 3.638119, 3.804725, 
    3.521243,
  3.66761, 3.773006, 12.72602, 3.51951, 3.618291, 3.681312, 3.821372, 
    3.810139, 3.63007, 4.061839, 9.488686, 14.00419, 11.35221, 3.881066, 
    3.720571, 3.558155, 3.768447, 3.699751, 3.373923, 3.377056, 3.74298, 
    3.585012, 3.554054, 4.445781, 8.791452, 3.524465, 3.547789, 3.457552, 
    3.586616,
  3.343278, 9.731485, 10.03323, 3.67545, 3.716024, 3.69691, 3.56251, 
    3.675848, 3.740429, 3.879701, 11.85861, 11.55573, 3.708889, 3.691036, 
    3.52657, 3.39075, 3.533785, 3.653764, 3.745188, 3.830686, 3.52587, 
    3.226712, 3.32978, 3.519117, 8.846123, 8.886536, 3.755616, 3.699037, 
    3.471109,
  3.156687, 6.091648, 9.017807, 9.150652, 3.64933, 3.597702, 3.276331, 
    3.300356, 3.423741, 3.52881, 4.858662, 3.561613, 4.307991, 3.159681, 
    3.187902, 3.32108, 3.600032, 3.837202, 3.655761, 3.798999, 3.580768, 
    3.284446, 3.332468, 8.609146, 8.507972, 11.83937, 3.657068, 3.419112, 
    3.247874,
  3.200632, 8.148125, 8.265129, 9.984423, 3.482576, 3.279022, 3.117794, 
    3.052537, 8.552002, 8.376835, 3.271375, 3.317401, 3.267097, 3.52293, 
    3.527341, 3.512039, 3.582831, 3.770384, 3.52225, 3.551509, 3.444216, 
    3.124511, 3.198072, 8.496183, 8.645205, 3.421478, 3.390983, 3.279215, 
    3.074495,
  9.597832, 9.847884, 9.772965, 9.33949, 14.61635, 3.309196, 4.931525, 
    3.12315, 3.182261, 3.150332, 4.039608, 3.104932, 3.263811, 3.247242, 
    3.189955, 3.250154, 3.337803, 3.479751, 3.506384, 3.214975, 3.148636, 
    3.141697, 8.59942, 7.369661, 3.454435, 3.151597, 3.033123, 3.131675, 
    8.5839,
  17.8673, 20.1948, 21.89411, 3.388096, 22.4759, 3.165919, 10.22369, 
    3.098615, 8.640246, 3.430589, 3.335502, 3.312146, 3.379266, 3.546149, 
    3.552728, 3.714237, 3.551233, 3.64214, 3.542567, 3.461562, 3.236046, 
    6.153461, 3.47058, 4.055276, 3.473653, 3.297194, 3.138513, 3.142396, 
    22.93318,
  22.98341, 19.29955, 20.09616, 18.87107, 12.64375, 14.52524, 11.8901, 
    9.986154, 6.819643, 9.802758, 3.427716, 3.539247, 3.617964, 3.554542, 
    3.789113, 3.683209, 3.635061, 3.753249, 3.525754, 3.828461, 11.96891, 
    11.93237, 8.691796, 3.597506, 3.628956, 3.487498, 3.694915, 3.721178, 
    10.42413,
  6.148839, 3.829409, 6.213335, 9.976778, 1.973944, 14.68624, 8.810743, 
    14.63238, 12.63992, 10.8413, 7.370614, 3.915973, 3.705724, 3.553941, 
    3.517221, 3.532708, 3.780565, 3.781206, 3.473422, 11.83168, 10.69566, 
    12.98729, 11.99576, 4.362588, 3.722741, 3.546784, 3.611377, 3.733143, 
    5.086323,
  6.035104, 11.11728, 12.05241, 12.57505, 12.09941, 11.27836, 7.590394, 
    11.66655, 8.83661, 6.760227, 6.597154, 6.16346, 3.749785, 3.661078, 
    3.835633, 3.737723, 3.720893, 4.057947, 4.131913, 8.549609, 10.07228, 
    9.330645, 6.442953, 6.153228, 4.989635, 3.597884, 3.649528, 4.078277, 
    4.161442,
  4.404262, 6.420896, 7.479022, 6.164582, 7.190842, 7.067245, 6.900622, 
    6.762216, 6.809305, 7.543815, 6.6517, 9.787057, 10.15287, 6.116961, 
    4.690738, 4.283021, 9.176804, 12.57676, 10.28384, 6.696338, 5.98974, 
    9.823442, 3.654905, 9.477062, 3.675352, 7.277973, 3.922466, 3.822765, 
    4.277844,
  4.151853, 4.754367, 6.999215, 4.42656, 4.226396, 5.125216, 11.63136, 
    12.11879, 13.63518, 12.04701, 9.019892, 7.894616, 10.85963, 5.226415, 
    21.77841, 4.664384, 9.99306, 15.29733, 9.544284, 6.84532, 17.29002, 
    10.80522, 14.04925, 24.11082, 4.988439, 41.65937, 43.01688, 8.080441, 
    4.215809,
  34.67865, 5.680239, 11.9314, 12.14448, 13.29152, 31.5202, 35.37904, 
    24.23923, 23.01473, 43.87937, 43.72669, 44.54483, 44.83745, 45.45209, 
    46.72717, 46.71783, 45.58794, 44.40288, 44.72347, 45.48284, 46.47599, 
    39.96976, 38.73441, 42.19539, 44.7522, 46.87964, 47.54099, 42.12761, 
    47.01162,
  76.34792, 76.34792, 76.34792, 76.34792, 76.34792, 76.34792, 76.34792, 
    76.29549, 76.29549, 76.29549, 76.29549, 76.29549, 76.29549, 76.29549, 
    76.1909, 76.1909, 76.1909, 76.1909, 76.1909, 76.1909, 76.1909, 76.33128, 
    76.33128, 76.33128, 76.33128, 76.33128, 76.33128, 76.33128, 76.34792,
  64.8836, 64.57207, 64.61784, 64.99524, 64.85411, 64.8848, 64.90484, 
    64.77013, 64.92882, 64.95878, 64.54097, 64.85989, 65.05613, 65.30067, 
    65.30379, 65.6069, 65.23344, 65.11444, 65.28864, 64.99837, 65.05997, 
    65.05544, 65.40359, 66.3326, 66.14386, 65.5992, 65.92085, 65.29882, 
    64.74574,
  57.14773, 57.26236, 59.44061, 55.34437, 50.38761, 50.4798, 55.41345, 
    50.51204, 50.3896, 50.49445, 50.36927, 50.42175, 50.73204, 59.16826, 
    59.40387, 58.27535, 56.2235, 57.23722, 57.98363, 58.07389, 55.20712, 
    52.11857, 47.70717, 46.60032, 51.54345, 50.50215, 50.72697, 51.77903, 
    57.41452,
  44.55904, 46.66686, 46.02581, 29.89131, 14.10824, 8.540816, 42.24285, 
    7.765872, 6.95402, 4.949214, 5.059228, 5.015715, 4.771024, 4.619771, 
    4.847534, 4.668594, 4.519419, 4.349875, 4.633832, 4.714952, 4.880421, 
    4.894166, 5.010652, 4.886749, 4.654101, 34.69159, 40.63885, 43.41626, 
    43.72532,
  3.912254, 3.81077, 3.826308, 3.876171, 4.05301, 4.030724, 4.068542, 
    4.131194, 4.184787, 4.044355, 4.1343, 4.02833, 4.169549, 4.13928, 
    4.163964, 4.023401, 3.833576, 3.980007, 3.923183, 4.028841, 4.17316, 
    4.217296, 4.13338, 7.934977, 4.46298, 3.929939, 3.825797, 4.07001, 
    3.987366,
  3.739376, 3.747684, 3.847212, 3.928405, 3.801199, 3.812694, 3.775181, 
    3.599036, 3.73538, 3.641643, 3.942143, 4.063015, 4.208814, 3.796031, 
    13.25613, 3.675733, 3.486383, 3.587488, 3.555808, 3.928852, 3.811433, 
    3.945117, 3.932839, 11.28014, 4.396631, 3.885188, 3.8827, 3.896135, 
    3.901909,
  3.497689, 3.947155, 12.41915, 3.681758, 3.658295, 3.540581, 3.787115, 
    3.54672, 3.858988, 3.929231, 9.924705, 14.97167, 10.68633, 3.855695, 
    3.587164, 3.757258, 3.607274, 3.796764, 3.380582, 3.691831, 3.659206, 
    3.79844, 3.803213, 4.51616, 9.221085, 3.569818, 3.602677, 3.489871, 
    3.613921,
  3.405143, 10.03319, 10.16408, 3.901414, 3.772617, 3.736023, 3.909662, 
    3.552707, 3.488516, 3.632147, 12.0702, 11.71833, 3.883914, 3.71501, 
    3.674783, 3.684717, 3.415746, 3.502274, 3.416227, 3.786545, 3.713336, 
    3.55746, 3.2184, 3.660077, 9.149323, 9.088811, 3.468332, 3.535538, 
    3.594057,
  3.175615, 6.05899, 8.6868, 9.368321, 3.46104, 3.353476, 3.569134, 3.335799, 
    3.40973, 3.437185, 4.80606, 3.265042, 4.524522, 3.414325, 3.145693, 
    3.518253, 3.342131, 3.615821, 3.607019, 3.807158, 3.577451, 3.650971, 
    3.200962, 8.334311, 8.813974, 11.90786, 3.629891, 3.41652, 3.388379,
  3.203526, 8.103395, 8.181146, 9.992857, 3.424624, 3.330621, 3.539443, 
    3.32143, 8.484052, 8.398689, 3.254187, 3.213645, 3.36041, 3.316066, 
    3.511811, 3.612092, 3.567742, 3.780416, 3.650619, 3.799321, 3.47945, 
    3.101351, 3.161267, 8.393649, 8.416717, 3.460916, 3.536686, 3.429475, 
    3.22228,
  9.387739, 10.04605, 10.31025, 9.081907, 14.59109, 3.570883, 4.964396, 
    3.321207, 3.327412, 3.262878, 3.98669, 3.199351, 3.022435, 3.176023, 
    3.247084, 3.109719, 3.168733, 3.436097, 3.313961, 3.432999, 3.421421, 
    3.034396, 8.324662, 7.39824, 3.147766, 3.204967, 3.049687, 2.966695, 
    8.693636,
  16.94649, 19.31001, 21.29592, 3.406748, 21.59598, 3.702733, 10.28362, 
    3.227338, 8.988012, 3.468667, 3.36557, 3.403026, 3.3912, 3.415849, 
    3.611377, 3.469244, 3.641126, 3.514956, 3.644757, 3.449636, 3.590362, 
    5.920456, 3.478851, 4.263922, 3.420608, 3.516079, 3.322428, 3.01893, 
    22.00011,
  21.53307, 17.99945, 18.7297, 17.61891, 12.02859, 13.8206, 11.59929, 
    9.998443, 10.53391, 10.06409, 3.516202, 3.722348, 3.533786, 3.668326, 
    3.634752, 3.59421, 3.866001, 3.78192, 3.702254, 4.032545, 11.49634, 
    11.06455, 8.72344, 3.734478, 3.417181, 3.836426, 3.508264, 3.834441, 
    9.774302,
  7.137391, 4.058389, 5.84375, 9.604799, 1.79822, 13.48337, 8.110905, 
    13.52328, 11.62199, 10.90083, 6.762012, 3.706711, 3.544802, 3.265991, 
    3.464738, 3.470135, 3.578688, 3.261449, 3.61293, 11.14855, 10.60005, 
    12.02816, 11.3733, 4.536029, 3.725235, 3.733176, 3.525459, 3.646761, 
    5.029325,
  5.018207, 9.678378, 10.76765, 11.32695, 10.60937, 10.06497, 6.717124, 
    12.75431, 7.388952, 6.719137, 6.618441, 8.19346, 3.541176, 3.852667, 
    3.715433, 3.745627, 3.799627, 3.660011, 3.536257, 7.801223, 8.857583, 
    8.204177, 7.376137, 6.533716, 4.5667, 3.441887, 3.443881, 3.356353, 
    3.532964,
  3.936877, 6.25112, 6.206897, 6.23612, 6.619791, 6.381757, 5.951904, 
    7.001349, 7.607394, 8.205813, 7.324815, 11.29995, 12.85331, 8.582529, 
    3.140881, 3.866322, 8.522807, 10.2372, 10.28791, 5.882853, 5.672953, 
    9.001056, 3.800046, 9.95096, 3.129219, 6.250645, 3.9175, 4.045475, 
    3.576432,
  3.800441, 4.152675, 8.62969, 3.496174, 3.225417, 3.850052, 11.68571, 
    12.72334, 17.63758, 25.05117, 12.94881, 8.190425, 10.7292, 27.8801, 
    31.26576, 3.522625, 20.67226, 19.57228, 15.23322, 5.985175, 17.96907, 
    23.36051, 21.68699, 22.38698, 3.157455, 28.7073, 28.50282, 16.20536, 
    3.273015,
  9.795769, 2.462685, 10.16049, 8.996198, 6.017338, 12.58445, 13.51844, 
    12.94057, 13.48582, 13.39214, 13.26702, 13.09277, 13.34129, 13.27341, 
    12.97331, 12.40372, 12.14484, 12.0119, 12.0934, 12.17131, 12.1664, 
    11.22708, 10.98061, 11.7254, 10.99343, 11.10572, 10.99553, 10.86483, 
    13.04578,
  76.27164, 76.27164, 76.27164, 76.27164, 76.27164, 76.27164, 76.27164, 
    76.27699, 76.27699, 76.27699, 76.27699, 76.27699, 76.27699, 76.27699, 
    76.2793, 76.2793, 76.2793, 76.2793, 76.2793, 76.2793, 76.2793, 76.31124, 
    76.31124, 76.31124, 76.31124, 76.31124, 76.31124, 76.31124, 76.27164,
  76.35242, 76.16932, 76.06711, 76.03042, 75.99735, 76.02655, 76.01499, 
    75.98363, 76.01456, 76.02307, 76.05218, 76.11053, 76.20306, 76.42274, 
    76.41149, 77.03011, 76.9541, 76.78632, 76.60933, 76.52366, 76.69807, 
    76.74238, 77.14258, 75.53281, 74.85128, 74.69977, 73.85787, 75.63739, 
    76.43199,
  67.68288, 65.99952, 74.47392, 69.74519, 68.26066, 68.23944, 60.80435, 
    67.74997, 67.47323, 67.71695, 67.68707, 67.65934, 68.14977, 78.42096, 
    77.30242, 73.7411, 70.80177, 71.81897, 71.12572, 69.0464, 66.53552, 
    44.25152, 59.31339, 59.27809, 62.20302, 64.34548, 63.27911, 63.52958, 
    66.61816,
  40.56993, 47.84757, 30.83875, 9.138043, 5.62297, 5.03018, 4.946997, 
    5.095215, 5.055817, 5.035543, 5.24988, 5.1634, 5.243423, 5.115674, 
    5.23986, 5.13573, 5.108906, 5.092359, 5.274127, 5.068138, 5.106168, 
    4.969546, 5.019871, 4.96153, 4.831969, 13.58893, 45.70667, 42.14108, 
    42.8769,
  4.083227, 4.417402, 4.463652, 4.524312, 4.498238, 4.409156, 4.377548, 
    4.492009, 4.556731, 4.497719, 4.402445, 4.330289, 4.42919, 4.088641, 
    4.258945, 4.582152, 4.517012, 4.354661, 4.35632, 4.23593, 4.199351, 
    4.297112, 4.266934, 8.726915, 4.702657, 4.366656, 4.206131, 4.122038, 
    4.276138,
  3.943547, 3.977809, 4.227108, 3.947287, 4.013211, 3.993726, 3.951106, 
    3.889347, 3.860957, 3.941604, 3.845921, 4.102917, 4.113184, 4.031137, 
    10.05186, 3.806201, 3.871399, 3.954737, 4.305062, 3.954795, 3.91937, 
    3.977437, 3.929244, 9.817687, 4.305885, 4.179577, 3.989821, 4.004017, 
    3.964952,
  3.944763, 4.045322, 12.92369, 3.782904, 3.846295, 3.797265, 3.913525, 
    3.829944, 3.748573, 4.062509, 10.21581, 15.83448, 11.017, 3.856991, 
    3.778453, 3.974533, 3.895796, 3.726755, 3.625791, 3.629362, 3.729891, 
    3.915893, 3.745347, 4.758852, 9.743622, 3.833191, 3.806345, 3.864904, 
    3.916213,
  3.29473, 10.51694, 10.50228, 3.592834, 3.644662, 3.739664, 3.782785, 
    3.772313, 3.861423, 3.736635, 12.45665, 12.18998, 3.69278, 3.734503, 
    3.717327, 3.831799, 3.63728, 3.572261, 3.509674, 3.988579, 3.921243, 
    3.75021, 3.374351, 3.566026, 9.410976, 9.390082, 3.805716, 3.588044, 
    3.689655,
  3.277909, 6.359814, 8.822883, 9.175161, 3.589143, 3.391065, 3.408422, 
    3.321093, 3.44991, 3.434615, 5.142993, 3.362371, 4.674433, 3.496783, 
    3.303743, 3.667776, 3.525543, 3.826428, 3.647396, 4.014215, 3.643505, 
    3.428507, 3.281067, 8.797507, 8.60709, 8.958352, 3.686894, 3.478005, 
    3.553292,
  3.154965, 8.509486, 8.271131, 9.676908, 3.477555, 3.498202, 3.53428, 
    3.381862, 8.411865, 8.215635, 3.279273, 3.451229, 3.304678, 3.451146, 
    3.468148, 3.582786, 3.620945, 3.789312, 3.589975, 3.797521, 3.453091, 
    3.219645, 3.423378, 8.40978, 8.392945, 3.432708, 3.495219, 3.497262, 
    3.33511,
  9.86727, 10.19926, 9.994411, 9.463506, 14.30549, 3.44985, 5.135857, 
    3.582154, 3.439611, 3.235509, 4.081657, 3.483027, 3.203094, 3.236126, 
    3.41261, 3.298735, 3.539014, 3.299747, 3.503453, 3.147183, 3.222244, 
    3.292617, 8.565457, 7.450588, 3.589347, 3.587792, 3.17352, 3.611574, 
    8.882711,
  16.58678, 18.71688, 20.60765, 3.752549, 20.75314, 3.94874, 10.49597, 
    3.935206, 8.776859, 3.483607, 3.205182, 3.365786, 3.660974, 3.860899, 
    4.040407, 3.826321, 4.010668, 3.714398, 3.599426, 3.643984, 4.013387, 
    5.806623, 3.458697, 4.303502, 3.688161, 3.675039, 3.563061, 3.623378, 
    21.21563,
  20.57167, 17.22454, 17.77888, 16.51601, 11.56951, 12.80246, 11.02453, 
    18.51127, 7.841946, 9.601162, 3.674597, 3.73408, 3.902867, 3.814044, 
    3.66318, 3.828666, 3.648663, 3.929135, 3.537109, 4.15015, 9.199241, 
    10.70751, 8.263031, 3.735389, 3.739969, 3.63305, 3.932399, 3.908388, 
    9.593773,
  6.029313, 4.386253, 5.540312, 9.291282, 1.637772, 12.1817, 11.68852, 
    12.2715, 10.93843, 10.46407, 7.057492, 3.493027, 4.097932, 3.882261, 
    3.832399, 3.992466, 3.376299, 3.293329, 3.661782, 9.736567, 9.545227, 
    11.32651, 10.12375, 4.234021, 3.470152, 3.560719, 3.55562, 3.904268, 
    4.902585,
  5.200981, 8.798709, 9.658195, 10.12296, 8.997507, 8.898866, 6.614154, 
    23.58991, 8.429526, 6.652975, 5.989398, 13.83663, 3.307596, 3.582465, 
    3.770773, 3.370727, 3.248988, 3.253174, 3.037222, 7.247458, 8.999235, 
    10.64048, 11.31876, 16.03565, 4.708081, 3.563449, 3.441991, 3.342852, 
    3.744542,
  3.634066, 10.39025, 6.751377, 8.584142, 7.016211, 9.086443, 6.584736, 
    10.30195, 10.16471, 10.49056, 7.651548, 20.9822, 23.64075, 11.34961, 
    2.242072, 3.039124, 11.63584, 10.00803, 19.44252, 7.331436, 9.957579, 
    22.2292, 3.192827, 22.19687, 3.056976, 4.88958, 3.144429, 3.223058, 
    3.081795,
  1.0364, 0.8928514, 3.837065, 0.8798878, 0.863392, 1.933193, 7.958504, 
    7.991439, 7.816866, 7.933673, 4.620799, 3.07819, 7.239893, 9.514277, 
    9.287303, 3.032434, 8.151765, 8.155948, 8.676926, 7.803829, 7.231671, 
    8.468578, 7.660348, 7.915191, 0.7866554, 7.945049, 7.969198, 7.98115, 
    0.9593921,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  76.13555, 76.13555, 76.13555, 76.13555, 76.13555, 76.13555, 76.13555, 
    76.16167, 76.16167, 76.16167, 76.16167, 76.16167, 76.16167, 76.16167, 
    76.20033, 76.20033, 76.20033, 76.20033, 76.20033, 76.20033, 76.20033, 
    76.18402, 76.18402, 76.18402, 76.18402, 76.18402, 76.18402, 76.18402, 
    76.13555,
  76.35452, 76.19527, 76.0992, 76.00932, 75.96207, 75.90783, 75.88535, 
    75.89178, 75.93999, 76.01354, 76.11885, 76.12794, 76.3341, 69.87098, 
    68.34055, 67.0013, 66.90444, 67.60623, 69.87836, 74.96468, 76.21087, 
    76.4316, 75.95966, 64.94259, 65.62067, 64.78209, 64.64643, 67.53224, 
    76.27279,
  46.66751, 40.14297, 63.61326, 65.48601, 76.34853, 76.73755, 56.03942, 
    75.99763, 75.86828, 75.86781, 75.9255, 75.9981, 72.26419, 71.03369, 
    51.40993, 28.35418, 25.06566, 60.26761, 52.76725, 60.77001, 47.95707, 
    37.22901, 61.19368, 63.48392, 64.68018, 60.53158, 44.86546, 38.2002, 
    46.03336,
  4.92067, 44.76322, 4.830221, 4.803882, 4.75036, 4.702308, 4.854949, 
    5.105814, 5.218238, 5.410077, 5.430798, 5.228028, 4.969777, 5.191349, 
    5.395777, 5.129903, 5.267948, 5.10267, 5.129266, 5.154373, 5.361742, 
    5.294181, 5.217529, 5.124929, 5.044704, 8.795198, 33.29396, 12.49164, 
    10.40916,
  4.316248, 4.409105, 4.280708, 4.398264, 4.432966, 4.347757, 4.465708, 
    4.394874, 4.337368, 4.42209, 4.593459, 4.458628, 4.462576, 4.33088, 
    4.499528, 4.551941, 4.309874, 4.502297, 4.363528, 4.701666, 4.5089, 
    4.519996, 4.449102, 8.88013, 5.197481, 4.755109, 4.497812, 4.227966, 
    4.365754,
  4.192708, 4.173234, 4.503735, 4.074657, 4.217872, 4.19254, 3.833158, 
    4.100229, 4.024463, 4.10667, 3.972231, 4.331143, 4.203409, 4.178179, 
    10.35894, 3.896481, 4.004969, 4.153093, 3.930152, 3.917884, 4.087285, 
    3.934559, 4.113989, 10.30507, 4.273955, 4.244535, 4.139349, 4.066302, 
    4.126666,
  3.805301, 4.152401, 13.13804, 3.649227, 3.917532, 4.115233, 3.750492, 
    4.096236, 3.812405, 4.210562, 10.47775, 16.23137, 10.94638, 4.168949, 
    3.957705, 3.850651, 4.137971, 3.820354, 3.509146, 3.662467, 4.060136, 
    3.95551, 3.973168, 4.900866, 9.677895, 3.851726, 3.792713, 3.929389, 
    3.947605,
  3.540888, 10.28622, 10.42877, 3.838864, 3.705942, 3.703078, 3.964645, 
    3.84033, 3.641634, 4.051556, 12.27944, 11.73181, 3.959391, 3.745161, 
    3.586811, 3.627119, 3.483611, 3.526035, 3.855895, 4.105494, 3.873019, 
    4.04405, 3.386294, 3.408751, 9.753648, 9.456862, 3.980017, 4.006966, 
    3.757917,
  3.233804, 6.676659, 9.000182, 9.283442, 3.459512, 3.506742, 3.303633, 
    3.408353, 3.597164, 3.304155, 4.888968, 3.512861, 4.531201, 3.331307, 
    3.319286, 3.587328, 3.507357, 3.842682, 3.574599, 4.000473, 3.68909, 
    3.660137, 3.353565, 8.928036, 8.574518, 8.910154, 3.800139, 3.577587, 
    3.737529,
  3.168326, 8.868134, 8.469222, 9.715761, 3.596029, 3.593704, 3.465655, 
    3.421366, 8.628778, 8.186518, 3.478569, 3.448586, 3.178027, 3.434965, 
    3.519555, 3.697637, 3.733233, 3.892927, 3.774205, 3.876055, 3.762301, 
    3.235647, 3.305473, 8.464889, 8.551067, 3.44493, 3.337162, 3.518698, 
    3.323592,
  10.06523, 10.38361, 10.35662, 9.324317, 13.99603, 3.472922, 5.653937, 
    3.951053, 3.390982, 3.592128, 4.250901, 3.447018, 3.466069, 3.5316, 
    3.428101, 3.534483, 3.735986, 3.267154, 3.712708, 3.392942, 3.431848, 
    3.649763, 8.481645, 7.159072, 3.453278, 3.61817, 3.151664, 3.467304, 
    8.997998,
  15.67493, 18.40475, 20.68396, 3.844038, 20.35705, 3.920913, 10.40217, 
    4.194667, 9.088999, 3.358753, 3.548091, 3.811486, 3.870946, 4.006296, 
    4.275704, 3.997265, 3.997861, 3.639422, 3.506804, 3.394515, 4.059182, 
    5.838926, 4.04731, 4.908596, 3.784641, 3.99811, 3.893771, 3.873172, 
    20.84708,
  20.04106, 16.56619, 17.03666, 16.0916, 10.75092, 12.03941, 10.94081, 
    20.17916, 10.68482, 9.593909, 3.514697, 3.754733, 4.100675, 3.971699, 
    3.918983, 3.783, 3.585099, 3.811981, 3.419732, 3.851769, 8.454815, 
    10.17857, 8.004357, 3.634355, 3.82267, 3.570081, 4.003907, 4.082883, 
    9.614446,
  5.246389, 4.197029, 4.96362, 11.39095, 1.5245, 11.27416, 16.30254, 
    12.56195, 10.251, 19.89279, 9.924774, 3.462151, 4.310572, 4.071455, 
    3.715486, 3.569047, 3.11763, 3.153113, 3.887731, 11.62304, 17.25614, 
    12.05905, 10.44522, 3.765343, 3.406249, 3.392457, 3.32948, 3.807827, 
    4.268058,
  4.22495, 7.949425, 10.9591, 15.06866, 15.35563, 17.33369, 9.934199, 
    22.58436, 10.27222, 5.911169, 5.263299, 15.50613, 3.446767, 4.018446, 
    3.574628, 3.218309, 3.363861, 3.65958, 4.054349, 11.57522, 12.45622, 
    19.55111, 14.85919, 19.90637, 5.09614, 3.338633, 3.385429, 3.608537, 
    3.49331,
  2.404103, 11.39395, 5.953698, 9.697238, 7.977333, 9.724386, 7.787672, 
    11.28488, 10.12462, 10.63467, 8.23129, 17.28834, 18.56227, 12.86236, 
    2.095158, 2.625715, 13.73327, 8.215582, 18.17134, 8.274078, 11.55905, 
    18.75428, 22.08476, 18.44226, 2.258399, 5.454312, 2.836203, 2.752644, 
    2.789562,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0 ;

 lat = -89.5, -79.5, -69.5, -59.5, -49.5, -39.5, -29.5, -19.5, -9.5, 0.5, 
    10.5, 20.5, 30.5, 40.5, 50.5, 60.5, 70.5, 80.5 ;

 lat_bnds =
  -90, -89,
  -80, -79,
  -70, -69,
  -60, -59,
  -50, -49,
  -40, -39,
  -30, -29,
  -20, -19,
  -10, -9,
  0, 1,
  10, 11,
  20, 21,
  30, 31,
  40, 41,
  50, 51,
  60, 61,
  70, 71,
  80, 81 ;

 lon = 0.625, 13.125, 25.625, 38.125, 50.625, 63.125, 75.625, 88.125, 
    100.625, 113.125, 125.625, 138.125, 150.625, 163.125, 175.625, 188.125, 
    200.625, 213.125, 225.625, 238.125, 250.625, 263.125, 275.625, 288.125, 
    300.625, 313.125, 325.625, 338.125, 350.625 ;

 lon_bnds =
  0, 1.25,
  12.5, 13.75,
  25, 26.25,
  37.5, 38.75,
  50, 51.25,
  62.5, 63.75,
  75, 76.25,
  87.5, 88.75,
  100, 101.25,
  112.5, 113.75,
  125, 126.25,
  137.5, 138.75,
  150, 151.25,
  162.5, 163.75,
  175, 176.25,
  187.5, 188.75,
  200, 201.25,
  212.5, 213.75,
  225, 226.25,
  237.5, 238.75,
  250, 251.25,
  262.5, 263.75,
  275, 276.25,
  287.5, 288.75,
  300, 301.25,
  312.5, 313.75,
  325, 326.25,
  337.5, 338.75,
  350, 351.25 ;

 time = 380.5, 410.5, 440.5, 471, 501.5, 532, 562.5, 593.5, 624, 654.5, 685, 
    715.5 ;

 time_bnds =
  365, 396,
  396, 425,
  425, 456,
  456, 486,
  486, 517,
  517, 547,
  547, 578,
  578, 609,
  609, 639,
  639, 670,
  670, 700,
  700, 731 ;
}
