netcdf LUmip_refined.185001-185412.gppLut {
dimensions:
	time = UNLIMITED ; // (60 currently)
	bnds = 2 ;
	landuse = 4 ;
	lat = 2 ;
	lon = 2 ;
variables:
	double average_DT(time) ;
		average_DT:long_name = "Length of average period" ;
		average_DT:units = "days" ;
		average_DT:missing_value = 1.e+20 ;
		average_DT:_FillValue = 1.e+20 ;
	double average_T1(time) ;
		average_T1:long_name = "Start time for average period" ;
		average_T1:units = "days since 1850-01-01 00:00:00" ;
		average_T1:missing_value = 1.e+20 ;
		average_T1:_FillValue = 1.e+20 ;
	double average_T2(time) ;
		average_T2:long_name = "End time for average period" ;
		average_T2:units = "days since 1850-01-01 00:00:00" ;
		average_T2:missing_value = 1.e+20 ;
		average_T2:_FillValue = 1.e+20 ;
	double bnds(bnds) ;
		bnds:long_name = "vertex number" ;
	float gppLut(time, landuse, lat, lon) ;
		gppLut:_FillValue = -1.f ;
		gppLut:long_name = "Gross Primary Productivity on Land Use Tile" ;
		gppLut:units = "kg m-2 s-1" ;
		gppLut:missing_value = -1.f ;
		gppLut:cell_methods = "area: mean time: mean" ;
		gppLut:cell_measures = "area: area" ;
		gppLut:time_avg_info = "average_T1,average_T2,average_DT" ;
		gppLut:standard_name = "gross_primary_productivity_of_biomass_expressed_as_carbon" ;
		gppLut:interp_method = "conserve_order1" ;
	int landuse(landuse) ;
		landuse:long_name = "Land use type" ;
		landuse:standard_name = "area_type" ;
		landuse:flag_values = 0, 1, 2, 3 ;
		landuse:flag_meanings = "psl pst crp urb" ;
	double lat(lat) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_N" ;
		lat:axis = "Y" ;
		lat:bounds = "lat_bnds" ;
	double lat_bnds(lat, bnds) ;
		lat_bnds:long_name = "latitude bounds" ;
		lat_bnds:units = "degrees_N" ;
		lat_bnds:axis = "Y" ;
	double lon(lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_E" ;
		lon:axis = "X" ;
		lon:bounds = "lon_bnds" ;
	double lon_bnds(lon, bnds) ;
		lon_bnds:long_name = "longitude bounds" ;
		lon_bnds:units = "degrees_E" ;
		lon_bnds:axis = "X" ;
	double time(time) ;
		time:long_name = "time" ;
		time:units = "days since 1850-01-01 00:00:00" ;
		time:axis = "T" ;
		time:calendar_type = "NOLEAP" ;
		time:calendar = "noleap" ;
		time:bounds = "time_bnds" ;
	double time_bnds(time, bnds) ;
		time_bnds:long_name = "time axis boundaries" ;
		time_bnds:units = "days since 1850-01-01 00:00:00" ;
		time_bnds:missing_value = 1.e+20 ;
		time_bnds:_FillValue = 1.e+20 ;

// global attributes:
		:filename = "LUmip_refined.185001-185412.gppLut.nc" ;
		:NumFilesInSet = 40 ;
		:title = "ESM4_historical_D1" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
		:history = "fregrid --standard_dimension --input_mosaic C96_mosaic.nc --input_file 18540101.lumip_refined --interp_method conserve_order1 --remap_file .fregrid_remap_file_288_by_180.nc --nlon 288 --nlat 180 --scalar_field time_bnds,geolat_t,geolon_t,area,gppLut,raLut,nppLut,rhLut,tasLut,tslsiLut,hussLut,hflsLut,hfssLut,rsusLut,rlusLut,laiLut,mrsosLut,mrroLut,mrsoLut,mrs1mLut,fracLut,cell_area --output_file out.nc" ;
		:code_version = "$Name: bronx-10_performance_z1l $" ;
		:external_variables = "area" ;
data:

 average_DT = 31, 28, 31, 30, 31, 30, 31, 31, 30, 31, 30, 31, 31, 28, 31, 30, 
    31, 30, 31, 31, 30, 31, 30, 31, 31, 28, 31, 30, 31, 30, 31, 31, 30, 31, 
    30, 31, 31, 28, 31, 30, 31, 30, 31, 31, 30, 31, 30, 31, 31, 28, 31, 30, 
    31, 30, 31, 31, 30, 31, 30, 31 ;

 average_T1 = 0, 31, 59, 90, 120, 151, 181, 212, 243, 273, 304, 334, 365, 
    396, 424, 455, 485, 516, 546, 577, 608, 638, 669, 699, 730, 761, 789, 
    820, 850, 881, 911, 942, 973, 1003, 1034, 1064, 1095, 1126, 1154, 1185, 
    1215, 1246, 1276, 1307, 1338, 1368, 1399, 1429, 1460, 1491, 1519, 1550, 
    1580, 1611, 1641, 1672, 1703, 1733, 1764, 1794 ;

 average_T2 = 31, 59, 90, 120, 151, 181, 212, 243, 273, 304, 334, 365, 396, 
    424, 455, 485, 516, 546, 577, 608, 638, 669, 699, 730, 761, 789, 820, 
    850, 881, 911, 942, 973, 1003, 1034, 1064, 1095, 1126, 1154, 1185, 1215, 
    1246, 1276, 1307, 1338, 1368, 1399, 1429, 1460, 1491, 1519, 1550, 1580, 
    1611, 1641, 1672, 1703, 1733, 1764, 1794, 1825 ;

 bnds = 1, 2 ;

 gppLut =
    2.47952e-08, 3.095144e-08, 3.532048e-08, 2.326242e-08, 3.522679e-08, 0, 
    3.018852e-09, 2.775054e-08, 1.807339e-08, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 0, 0, 1.179804e-10, 
    2.677578e-10, 0, 0, _, _, _, _, _, _, _, _, _, _, _, 0, 0, 0, 0, _, 0, 0, 
    0, 0, 0, 0, _, _, _, _, _, 5.878042e-08, 2.102753e-09, 0, 0, 0, 
    4.119591e-08, 2.277574e-08, 4.580447e-08, 3.790088e-08, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
    2.47952e-08, 3.095144e-08, 3.532048e-08, 2.326242e-08, 3.522679e-08, 0, 
    3.018852e-09, 2.775054e-08, 1.807339e-08, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 0, 0, 1.179804e-10, 
    2.677578e-10, 0, 0, _, _, _, _, _, _, _, _, _, _, _, 0, 0, 0, 0, _, 0, 0, 
    0, 0, 0, 0, _, _, _, _, _, 5.878042e-08, 2.102753e-09, 0, 0, 0, 
    4.119591e-08, 2.277574e-08, 4.580447e-08, 3.790088e-08, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
    2.47952e-08, 3.095144e-08, 3.532048e-08, 2.326242e-08, 3.522679e-08, 0, 
    3.018852e-09, 2.775054e-08, 1.807339e-08, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 0, 0, 1.179804e-10, 
    2.677578e-10, 0, 0, _, _, _, _, _, _, _, _, _, _, _, 0, 0, 0, 0, _, 0, 0, 
    0, 0, 0, 0, _, _, _, _, _, 5.878042e-08, 2.102753e-09, 0, 0, 0, 
    4.119591e-08, 2.277574e-08, 4.580447e-08, 3.790088e-08, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
    2.47952e-08, 3.095144e-08, 3.532048e-08, 2.326242e-08, 3.522679e-08, 0, 
    3.018852e-09, 2.775054e-08, 1.807339e-08, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 0, 0, 1.179804e-10, 
    2.677578e-10, 0, 0, _, _, _, _, _, _, _, _, _, _, _, 0, 0, 0, 0, _, 0, 0, 
    0, 0, 0, 0, _, _, _, _, _, 5.878042e-08, 2.102753e-09, 0, 0, 0, 
    4.119591e-08, 2.277574e-08, 4.580447e-08, 3.790088e-08, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
    2.47952e-08, 3.095144e-08, 3.532048e-08, 2.326242e-08, 3.522679e-08, 0, 
    3.018852e-09, 2.775054e-08, 1.807339e-08, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 0, 0, 1.179804e-10, 
    2.677578e-10, 0, 0, _, _, _, _, _, _, _, _, _, _, _, 0, 0, 0, 0, _, 0, 0, 
    0, 0, 0, 0, _, _, _, _, _, 5.878042e-08, 2.102753e-09, 0, 0, 0, 
    4.119591e-08, 2.277574e-08, 4.580447e-08, 3.790088e-08, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
    2.47952e-08, 3.095144e-08, 3.532048e-08, 2.326242e-08, 3.522679e-08, 0, 
    3.018852e-09, 2.775054e-08, 1.807339e-08, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 0, 0, 1.179804e-10, 
    2.677578e-10, 0, 0, _, _, _, _, _, _, _, _, _, _, _, 0, 0, 0, 0, _, 0, 0, 
    0, 0, 0, 0, _, _, _, _, _, 5.878042e-08, 2.102753e-09, 0, 0, 0, 
    4.119591e-08, 2.277574e-08, 4.580447e-08, 3.790088e-08, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
    2.47952e-08, 3.095144e-08, 3.532048e-08, 2.326242e-08, 3.522679e-08, 0, 
    3.018852e-09, 2.775054e-08, 1.807339e-08, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 0, 0, 1.179804e-10, 
    2.677578e-10, 0, 0, _, _, _, _, _, _, _, _, _, _, _, 0, 0, 0, 0, _, 0, 0, 
    0, 0, 0, 0, _, _, _, _, _, 5.878042e-08, 2.102753e-09, 0, 0, 0, 
    4.119591e-08, 2.277574e-08, 4.580447e-08, 3.790088e-08, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
    2.47952e-08, 3.095144e-08, 3.532048e-08, 2.326242e-08, 3.522679e-08, 0, 
    3.018852e-09, 2.775054e-08, 1.807339e-08, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 0, 0, 1.179804e-10, 
    2.677578e-10, 0, 0, _, _, _, _, _, _, _, _, _, _, _, 0, 0, 0, 0, _, 0, 0, 
    0, 0, 0, 0, _, _, _, _, _, 5.878042e-08, 2.102753e-09, 0, 0, 0, 
    4.119591e-08, 2.277574e-08, 4.580447e-08, 3.790088e-08, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _;


 landuse = 0, 1, 2, 3 ;

 lat = -89.5, -88.5;

 lat_bnds =
  -90, -89,
  -89, -88;

 lon = 0.625, 1.875;

 lon_bnds =
  0, 1.25,
  1.25, 2.5;

 time = 15.5, 45, 74.5, 105, 135.5, 166, 196.5, 227.5, 258, 288.5, 319, 
    349.5, 380.5, 410, 439.5, 470, 500.5, 531, 561.5, 592.5, 623, 653.5, 684, 
    714.5, 745.5, 775, 804.5, 835, 865.5, 896, 926.5, 957.5, 988, 1018.5, 
    1049, 1079.5, 1110.5, 1140, 1169.5, 1200, 1230.5, 1261, 1291.5, 1322.5, 
    1353, 1383.5, 1414, 1444.5, 1475.5, 1505, 1534.5, 1565, 1595.5, 1626, 
    1656.5, 1687.5, 1718, 1748.5, 1779, 1809.5 ;

 time_bnds =
  0, 31,
  31, 59,
  59, 90,
  90, 120,
  120, 151,
  151, 181,
  181, 212,
  212, 243,
  243, 273,
  273, 304,
  304, 334,
  334, 365,
  365, 396,
  396, 424,
  424, 455,
  455, 485,
  485, 516,
  516, 546,
  546, 577,
  577, 608,
  608, 638,
  638, 669,
  669, 699,
  699, 730,
  730, 761,
  761, 789,
  789, 820,
  820, 850,
  850, 881,
  881, 911,
  911, 942,
  942, 973,
  973, 1003,
  1003, 1034,
  1034, 1064,
  1064, 1095,
  1095, 1126,
  1126, 1154,
  1154, 1185,
  1185, 1215,
  1215, 1246,
  1246, 1276,
  1276, 1307,
  1307, 1338,
  1338, 1368,
  1368, 1399,
  1399, 1429,
  1429, 1460,
  1460, 1491,
  1491, 1519,
  1519, 1550,
  1550, 1580,
  1580, 1611,
  1611, 1641,
  1641, 1672,
  1672, 1703,
  1703, 1733,
  1733, 1764,
  1764, 1794,
  1794, 1825 ;
}


















