netcdf atmos_plev39_cmip.185001-185412.ta {
dimensions:
	time = UNLIMITED ; // (60 currently)
	bnds = 2 ;
	lat = 2 ;
	plev39 = 39 ;
variables:
	double average_DT(time) ;
		average_DT:long_name = "Length of average period" ;
		average_DT:units = "days" ;
		average_DT:missing_value = 1.e+20 ;
		average_DT:_FillValue = 1.e+20 ;
	double average_T1(time) ;
		average_T1:long_name = "Start time for average period" ;
		average_T1:units = "days since 1850-01-01 00:00:00" ;
		average_T1:missing_value = 1.e+20 ;
		average_T1:_FillValue = 1.e+20 ;
	double average_T2(time) ;
		average_T2:long_name = "End time for average period" ;
		average_T2:units = "days since 1850-01-01 00:00:00" ;
		average_T2:missing_value = 1.e+20 ;
		average_T2:_FillValue = 1.e+20 ;
	double bnds(bnds) ;
		bnds:long_name = "vertex number" ;
	double lat(lat) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_N" ;
		lat:axis = "Y" ;
		lat:bounds = "lat_bnds" ;
	double lat_bnds(lat, bnds) ;
		lat_bnds:long_name = "latitude bounds" ;
		lat_bnds:units = "degrees_N" ;
		lat_bnds:axis = "Y" ;
	double plev39(plev39) ;
		plev39:long_name = "pressure" ;
		plev39:units = "Pa" ;
		plev39:axis = "Z" ;
		plev39:positive = "down" ;
	float ta(time, plev39, lat) ;
		ta:long_name = "Air Temperature" ;
		ta:units = "K" ;
		ta:missing_value = 1.e+20f ;
		ta:cell_methods = "time: mean" ;
		ta:cell_measures = "area: area" ;
		ta:time_avg_info = "average_T1,average_T2,average_DT" ;
		ta:standard_name = "air_temperature" ;
		ta:interp_method = "conserve_order2" ;
		ta:_FillValue = 1.e+20f ;
	double time(time) ;
		time:long_name = "time" ;
		time:units = "days since 1850-01-01 00:00:00" ;
		time:axis = "T" ;
		time:calendar_type = "NOLEAP" ;
		time:calendar = "noleap" ;
		time:bounds = "time_bnds" ;
	double time_bnds(time, bnds) ;
		time_bnds:long_name = "time axis boundaries" ;
		time_bnds:units = "days since 1850-01-01 00:00:00" ;
		time_bnds:missing_value = 1.e+20 ;
		time_bnds:_FillValue = 1.e+20 ;

// global attributes:
		:filename = "atmos_plev39_cmip.185001-185412.ta.nc" ;
		:title = "ESM4_historical_D1" ;
		:associated_files = "area: 18540101.grid_spec.nc" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
		:history = "fregrid --standard_dimension --input_mosaic C96_mosaic.nc --input_file 18540101.atmos_month_plev39_refined --interp_method conserve_order2 --remap_file .fregrid_remap_file_288_by_180.nc --nlon 288 --nlat 180 --scalar_field time_bnds,bry,ch4,cly,hcl,hno3,ho2,meanage,n2o,noy,o3,oh,ta,ua,va,zg,tntmp,tntrl,tntrs,tntrlcs,tntrscs,tntc,tntscp,tntogw,tntnogw,utendogw,utendnogw --output_file out.nc" ;
		:code_version = "$Name: bronx-10_performance_z1l $" ;
		:external_variables = "area" ;
data:

 average_DT = 31, 28, 31, 30, 31, 30, 31, 31, 30, 31, 30, 31, 31, 28, 31, 30, 
    31, 30, 31, 31, 30, 31, 30, 31, 31, 28, 31, 30, 31, 30, 31, 31, 30, 31, 
    30, 31, 31, 28, 31, 30, 31, 30, 31, 31, 30, 31, 30, 31, 31, 28, 31, 30, 
    31, 30, 31, 31, 30, 31, 30, 31 ;

 average_T1 = 0, 31, 59, 90, 120, 151, 181, 212, 243, 273, 304, 334, 365, 
    396, 424, 455, 485, 516, 546, 577, 608, 638, 669, 699, 730, 761, 789, 
    820, 850, 881, 911, 942, 973, 1003, 1034, 1064, 1095, 1126, 1154, 1185, 
    1215, 1246, 1276, 1307, 1338, 1368, 1399, 1429, 1460, 1491, 1519, 1550, 
    1580, 1611, 1641, 1672, 1703, 1733, 1764, 1794 ;

 average_T2 = 31, 59, 90, 120, 151, 181, 212, 243, 273, 304, 334, 365, 396, 
    424, 455, 485, 516, 546, 577, 608, 638, 669, 699, 730, 761, 789, 820, 
    850, 881, 911, 942, 973, 1003, 1034, 1064, 1095, 1126, 1154, 1185, 1215, 
    1246, 1276, 1307, 1338, 1368, 1399, 1429, 1460, 1491, 1519, 1550, 1580, 
    1611, 1641, 1672, 1703, 1733, 1764, 1794, 1825 ;

 bnds = 1, 2 ;

 lat = -89.5, -88.5;

 lat_bnds =
  -90, -89,
  -89, -88;

 plev39 = 100000, 92500, 85000, 70000, 60000, 50000, 40000, 30000, 25000, 
    20000, 17000, 15000, 13000, 11500, 10000, 9000, 8000, 7000, 5000, 3000, 
    2000, 1500, 1000, 700, 500, 300, 200, 150, 100, 70, 50, 40, 30, 20, 15, 
    10, 7, 5, 3 ;

 ta =
    283.519, 284.2079, 284.8589, 285.5298, 286.2316, 286.9749, 287.7004, 
    288.4397, 288.9764, 289.7086, 290.403, 291.0512, 291.598, 292.0377, 
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793, 
    295.5613, 295.9263, 296.2113, 296.4967, 296.8282, 297.1194, 297.4232, 
    297.662, 297.9678, 298.1667, 298.4066, 298.5545, 298.7012, 298.8887,
	298.9477, 298.9558, 298.9343, 298.8975, 283.519, 284.2079, 284.8589,
	285.5298, 286.2316, 286.9749, 287.7004, 288.4397, 288.9764, 289.7086,
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793,
	290.403, 291.0512, 291.598, 292.0377, 
    283.519, 284.2079, 284.8589, 285.5298, 286.2316, 286.9749, 287.7004, 
    288.4397, 288.9764, 289.7086, 290.403, 291.0512, 291.598, 292.0377, 
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793, 
    295.5613, 295.9263, 296.2113, 296.4967, 296.8282, 297.1194, 297.4232, 
    297.662, 297.9678, 298.1667, 298.4066, 298.5545, 298.7012, 298.8887,
	298.9477, 298.9558, 298.9343, 298.8975, 283.519, 284.2079, 284.8589,
	285.5298, 286.2316, 286.9749, 287.7004, 288.4397, 288.9764, 289.7086,
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793,
	290.403, 291.0512, 291.598, 292.0377,

    283.519, 284.2079, 284.8589, 285.5298, 286.2316, 286.9749, 287.7004, 
    288.4397, 288.9764, 289.7086, 290.403, 291.0512, 291.598, 292.0377, 
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793, 
    295.5613, 295.9263, 296.2113, 296.4967, 296.8282, 297.1194, 297.4232, 
    297.662, 297.9678, 298.1667, 298.4066, 298.5545, 298.7012, 298.8887,
	298.9477, 298.9558, 298.9343, 298.8975, 283.519, 284.2079, 284.8589,
	285.5298, 286.2316, 286.9749, 287.7004, 288.4397, 288.9764, 289.7086,
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793,
	290.403, 291.0512, 291.598, 292.0377, 
    283.519, 284.2079, 284.8589, 285.5298, 286.2316, 286.9749, 287.7004, 
    288.4397, 288.9764, 289.7086, 290.403, 291.0512, 291.598, 292.0377, 
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793, 
    295.5613, 295.9263, 296.2113, 296.4967, 296.8282, 297.1194, 297.4232, 
    297.662, 297.9678, 298.1667, 298.4066, 298.5545, 298.7012, 298.8887,
	298.9477, 298.9558, 298.9343, 298.8975, 283.519, 284.2079, 284.8589,
	285.5298, 286.2316, 286.9749, 287.7004, 288.4397, 288.9764, 289.7086,
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793,
	290.403, 291.0512, 291.598, 292.0377,

    283.519, 284.2079, 284.8589, 285.5298, 286.2316, 286.9749, 287.7004, 
    288.4397, 288.9764, 289.7086, 290.403, 291.0512, 291.598, 292.0377, 
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793, 
    295.5613, 295.9263, 296.2113, 296.4967, 296.8282, 297.1194, 297.4232, 
    297.662, 297.9678, 298.1667, 298.4066, 298.5545, 298.7012, 298.8887,
	298.9477, 298.9558, 298.9343, 298.8975, 283.519, 284.2079, 284.8589,
	285.5298, 286.2316, 286.9749, 287.7004, 288.4397, 288.9764, 289.7086,
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793,
	290.403, 291.0512, 291.598, 292.0377, 
    283.519, 284.2079, 284.8589, 285.5298, 286.2316, 286.9749, 287.7004, 
    288.4397, 288.9764, 289.7086, 290.403, 291.0512, 291.598, 292.0377, 
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793, 
    295.5613, 295.9263, 296.2113, 296.4967, 296.8282, 297.1194, 297.4232, 
    297.662, 297.9678, 298.1667, 298.4066, 298.5545, 298.7012, 298.8887,
	298.9477, 298.9558, 298.9343, 298.8975, 283.519, 284.2079, 284.8589,
	285.5298, 286.2316, 286.9749, 287.7004, 288.4397, 288.9764, 289.7086,
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793,
	290.403, 291.0512, 291.598, 292.0377,

    283.519, 284.2079, 284.8589, 285.5298, 286.2316, 286.9749, 287.7004, 
    288.4397, 288.9764, 289.7086, 290.403, 291.0512, 291.598, 292.0377, 
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793, 
    295.5613, 295.9263, 296.2113, 296.4967, 296.8282, 297.1194, 297.4232, 
    297.662, 297.9678, 298.1667, 298.4066, 298.5545, 298.7012, 298.8887,
	298.9477, 298.9558, 298.9343, 298.8975, 283.519, 284.2079, 284.8589,
	285.5298, 286.2316, 286.9749, 287.7004, 288.4397, 288.9764, 289.7086,
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793,
	290.403, 291.0512, 291.598, 292.0377, 
    283.519, 284.2079, 284.8589, 285.5298, 286.2316, 286.9749, 287.7004, 
    288.4397, 288.9764, 289.7086, 290.403, 291.0512, 291.598, 292.0377, 
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793, 
    295.5613, 295.9263, 296.2113, 296.4967, 296.8282, 297.1194, 297.4232, 
    297.662, 297.9678, 298.1667, 298.4066, 298.5545, 298.7012, 298.8887,
	298.9477, 298.9558, 298.9343, 298.8975, 283.519, 284.2079, 284.8589,
	285.5298, 286.2316, 286.9749, 287.7004, 288.4397, 288.9764, 289.7086,
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793,
	290.403, 291.0512, 291.598, 292.0377,

    283.519, 284.2079, 284.8589, 285.5298, 286.2316, 286.9749, 287.7004, 
    288.4397, 288.9764, 289.7086, 290.403, 291.0512, 291.598, 292.0377, 
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793, 
    295.5613, 295.9263, 296.2113, 296.4967, 296.8282, 297.1194, 297.4232, 
    297.662, 297.9678, 298.1667, 298.4066, 298.5545, 298.7012, 298.8887,
	298.9477, 298.9558, 298.9343, 298.8975, 283.519, 284.2079, 284.8589,
	285.5298, 286.2316, 286.9749, 287.7004, 288.4397, 288.9764, 289.7086,
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793,
	290.403, 291.0512, 291.598, 292.0377, 
    283.519, 284.2079, 284.8589, 285.5298, 286.2316, 286.9749, 287.7004, 
    288.4397, 288.9764, 289.7086, 290.403, 291.0512, 291.598, 292.0377, 
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793, 
    295.5613, 295.9263, 296.2113, 296.4967, 296.8282, 297.1194, 297.4232, 
    297.662, 297.9678, 298.1667, 298.4066, 298.5545, 298.7012, 298.8887,
	298.9477, 298.9558, 298.9343, 298.8975, 283.519, 284.2079, 284.8589,
	285.5298, 286.2316, 286.9749, 287.7004, 288.4397, 288.9764, 289.7086,
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793,
	290.403, 291.0512, 291.598, 292.0377,

    283.519, 284.2079, 284.8589, 285.5298, 286.2316, 286.9749, 287.7004, 
    288.4397, 288.9764, 289.7086, 290.403, 291.0512, 291.598, 292.0377, 
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793, 
    295.5613, 295.9263, 296.2113, 296.4967, 296.8282, 297.1194, 297.4232, 
    297.662, 297.9678, 298.1667, 298.4066, 298.5545, 298.7012, 298.8887,
	298.9477, 298.9558, 298.9343, 298.8975, 283.519, 284.2079, 284.8589,
	285.5298, 286.2316, 286.9749, 287.7004, 288.4397, 288.9764, 289.7086,
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793,
	290.403, 291.0512, 291.598, 292.0377, 
    283.519, 284.2079, 284.8589, 285.5298, 286.2316, 286.9749, 287.7004, 
    288.4397, 288.9764, 289.7086, 290.403, 291.0512, 291.598, 292.0377, 
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793, 
    295.5613, 295.9263, 296.2113, 296.4967, 296.8282, 297.1194, 297.4232, 
    297.662, 297.9678, 298.1667, 298.4066, 298.5545, 298.7012, 298.8887,
	298.9477, 298.9558, 298.9343, 298.8975, 283.519, 284.2079, 284.8589,
	285.5298, 286.2316, 286.9749, 287.7004, 288.4397, 288.9764, 289.7086,
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793,
	290.403, 291.0512, 291.598, 292.0377,

    283.519, 284.2079, 284.8589, 285.5298, 286.2316, 286.9749, 287.7004, 
    288.4397, 288.9764, 289.7086, 290.403, 291.0512, 291.598, 292.0377, 
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793, 
    295.5613, 295.9263, 296.2113, 296.4967, 296.8282, 297.1194, 297.4232, 
    297.662, 297.9678, 298.1667, 298.4066, 298.5545, 298.7012, 298.8887,
	298.9477, 298.9558, 298.9343, 298.8975, 283.519, 284.2079, 284.8589,
	285.5298, 286.2316, 286.9749, 287.7004, 288.4397, 288.9764, 289.7086,
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793,
	290.403, 291.0512, 291.598, 292.0377, 
    283.519, 284.2079, 284.8589, 285.5298, 286.2316, 286.9749, 287.7004, 
    288.4397, 288.9764, 289.7086, 290.403, 291.0512, 291.598, 292.0377, 
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793, 
    295.5613, 295.9263, 296.2113, 296.4967, 296.8282, 297.1194, 297.4232, 
    297.662, 297.9678, 298.1667, 298.4066, 298.5545, 298.7012, 298.8887,
	298.9477, 298.9558, 298.9343, 298.8975, 283.519, 284.2079, 284.8589,
	285.5298, 286.2316, 286.9749, 287.7004, 288.4397, 288.9764, 289.7086,
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793,
	290.403, 291.0512, 291.598, 292.0377,

    283.519, 284.2079, 284.8589, 285.5298, 286.2316, 286.9749, 287.7004, 
    288.4397, 288.9764, 289.7086, 290.403, 291.0512, 291.598, 292.0377, 
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793, 
    295.5613, 295.9263, 296.2113, 296.4967, 296.8282, 297.1194, 297.4232, 
    297.662, 297.9678, 298.1667, 298.4066, 298.5545, 298.7012, 298.8887,
	298.9477, 298.9558, 298.9343, 298.8975, 283.519, 284.2079, 284.8589,
	285.5298, 286.2316, 286.9749, 287.7004, 288.4397, 288.9764, 289.7086,
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793,
	290.403, 291.0512, 291.598, 292.0377, 
    283.519, 284.2079, 284.8589, 285.5298, 286.2316, 286.9749, 287.7004, 
    288.4397, 288.9764, 289.7086, 290.403, 291.0512, 291.598, 292.0377, 
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793, 
    295.5613, 295.9263, 296.2113, 296.4967, 296.8282, 297.1194, 297.4232, 
    297.662, 297.9678, 298.1667, 298.4066, 298.5545, 298.7012, 298.8887,
	298.9477, 298.9558, 298.9343, 298.8975, 283.519, 284.2079, 284.8589,
	285.5298, 286.2316, 286.9749, 287.7004, 288.4397, 288.9764, 289.7086,
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793,
	290.403, 291.0512, 291.598, 292.0377,

    283.519, 284.2079, 284.8589, 285.5298, 286.2316, 286.9749, 287.7004, 
    288.4397, 288.9764, 289.7086, 290.403, 291.0512, 291.598, 292.0377, 
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793, 
    295.5613, 295.9263, 296.2113, 296.4967, 296.8282, 297.1194, 297.4232, 
    297.662, 297.9678, 298.1667, 298.4066, 298.5545, 298.7012, 298.8887,
	298.9477, 298.9558, 298.9343, 298.8975, 283.519, 284.2079, 284.8589,
	285.5298, 286.2316, 286.9749, 287.7004, 288.4397, 288.9764, 289.7086,
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793,
	290.403, 291.0512, 291.598, 292.0377, 
    283.519, 284.2079, 284.8589, 285.5298, 286.2316, 286.9749, 287.7004, 
    288.4397, 288.9764, 289.7086, 290.403, 291.0512, 291.598, 292.0377, 
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793, 
    295.5613, 295.9263, 296.2113, 296.4967, 296.8282, 297.1194, 297.4232, 
    297.662, 297.9678, 298.1667, 298.4066, 298.5545, 298.7012, 298.8887,
	298.9477, 298.9558, 298.9343, 298.8975, 283.519, 284.2079, 284.8589,
	285.5298, 286.2316, 286.9749, 287.7004, 288.4397, 288.9764, 289.7086,
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793,
	290.403, 291.0512, 291.598, 292.0377,

    283.519, 284.2079, 284.8589, 285.5298, 286.2316, 286.9749, 287.7004, 
    288.4397, 288.9764, 289.7086, 290.403, 291.0512, 291.598, 292.0377, 
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793, 
    295.5613, 295.9263, 296.2113, 296.4967, 296.8282, 297.1194, 297.4232, 
    297.662, 297.9678, 298.1667, 298.4066, 298.5545, 298.7012, 298.8887,
	298.9477, 298.9558, 298.9343, 298.8975, 283.519, 284.2079, 284.8589,
	285.5298, 286.2316, 286.9749, 287.7004, 288.4397, 288.9764, 289.7086,
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793,
	290.403, 291.0512, 291.598, 292.0377, 
    283.519, 284.2079, 284.8589, 285.5298, 286.2316, 286.9749, 287.7004, 
    288.4397, 288.9764, 289.7086, 290.403, 291.0512, 291.598, 292.0377, 
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793, 
    295.5613, 295.9263, 296.2113, 296.4967, 296.8282, 297.1194, 297.4232, 
    297.662, 297.9678, 298.1667, 298.4066, 298.5545, 298.7012, 298.8887,
	298.9477, 298.9558, 298.9343, 298.8975, 283.519, 284.2079, 284.8589,
	285.5298, 286.2316, 286.9749, 287.7004, 288.4397, 288.9764, 289.7086,
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793,
	290.403, 291.0512, 291.598, 292.0377,

    283.519, 284.2079, 284.8589, 285.5298, 286.2316, 286.9749, 287.7004, 
    288.4397, 288.9764, 289.7086, 290.403, 291.0512, 291.598, 292.0377, 
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793, 
    295.5613, 295.9263, 296.2113, 296.4967, 296.8282, 297.1194, 297.4232, 
    297.662, 297.9678, 298.1667, 298.4066, 298.5545, 298.7012, 298.8887,
	298.9477, 298.9558, 298.9343, 298.8975, 283.519, 284.2079, 284.8589,
	285.5298, 286.2316, 286.9749, 287.7004, 288.4397, 288.9764, 289.7086,
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793,
	290.403, 291.0512, 291.598, 292.0377, 
    283.519, 284.2079, 284.8589, 285.5298, 286.2316, 286.9749, 287.7004, 
    288.4397, 288.9764, 289.7086, 290.403, 291.0512, 291.598, 292.0377, 
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793, 
    295.5613, 295.9263, 296.2113, 296.4967, 296.8282, 297.1194, 297.4232, 
    297.662, 297.9678, 298.1667, 298.4066, 298.5545, 298.7012, 298.8887,
	298.9477, 298.9558, 298.9343, 298.8975, 283.519, 284.2079, 284.8589,
	285.5298, 286.2316, 286.9749, 287.7004, 288.4397, 288.9764, 289.7086,
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793,
	290.403, 291.0512, 291.598, 292.0377,

    283.519, 284.2079, 284.8589, 285.5298, 286.2316, 286.9749, 287.7004, 
    288.4397, 288.9764, 289.7086, 290.403, 291.0512, 291.598, 292.0377, 
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793, 
    295.5613, 295.9263, 296.2113, 296.4967, 296.8282, 297.1194, 297.4232, 
    297.662, 297.9678, 298.1667, 298.4066, 298.5545, 298.7012, 298.8887,
	298.9477, 298.9558, 298.9343, 298.8975, 283.519, 284.2079, 284.8589,
	285.5298, 286.2316, 286.9749, 287.7004, 288.4397, 288.9764, 289.7086,
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793,
	290.403, 291.0512, 291.598, 292.0377, 
    283.519, 284.2079, 284.8589, 285.5298, 286.2316, 286.9749, 287.7004, 
    288.4397, 288.9764, 289.7086, 290.403, 291.0512, 291.598, 292.0377, 
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793, 
    295.5613, 295.9263, 296.2113, 296.4967, 296.8282, 297.1194, 297.4232, 
    297.662, 297.9678, 298.1667, 298.4066, 298.5545, 298.7012, 298.8887,
	298.9477, 298.9558, 298.9343, 298.8975, 283.519, 284.2079, 284.8589,
	285.5298, 286.2316, 286.9749, 287.7004, 288.4397, 288.9764, 289.7086,
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793,
	290.403, 291.0512, 291.598, 292.0377,

    283.519, 284.2079, 284.8589, 285.5298, 286.2316, 286.9749, 287.7004, 
    288.4397, 288.9764, 289.7086, 290.403, 291.0512, 291.598, 292.0377, 
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793, 
    295.5613, 295.9263, 296.2113, 296.4967, 296.8282, 297.1194, 297.4232, 
    297.662, 297.9678, 298.1667, 298.4066, 298.5545, 298.7012, 298.8887,
	298.9477, 298.9558, 298.9343, 298.8975, 283.519, 284.2079, 284.8589,
	285.5298, 286.2316, 286.9749, 287.7004, 288.4397, 288.9764, 289.7086,
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793,
	290.403, 291.0512, 291.598, 292.0377, 
    283.519, 284.2079, 284.8589, 285.5298, 286.2316, 286.9749, 287.7004, 
    288.4397, 288.9764, 289.7086, 290.403, 291.0512, 291.598, 292.0377, 
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793, 
    295.5613, 295.9263, 296.2113, 296.4967, 296.8282, 297.1194, 297.4232, 
    297.662, 297.9678, 298.1667, 298.4066, 298.5545, 298.7012, 298.8887,
	298.9477, 298.9558, 298.9343, 298.8975, 283.519, 284.2079, 284.8589,
	285.5298, 286.2316, 286.9749, 287.7004, 288.4397, 288.9764, 289.7086,
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793,
	290.403, 291.0512, 291.598, 292.0377,

    283.519, 284.2079, 284.8589, 285.5298, 286.2316, 286.9749, 287.7004, 
    288.4397, 288.9764, 289.7086, 290.403, 291.0512, 291.598, 292.0377, 
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793, 
    295.5613, 295.9263, 296.2113, 296.4967, 296.8282, 297.1194, 297.4232, 
    297.662, 297.9678, 298.1667, 298.4066, 298.5545, 298.7012, 298.8887,
	298.9477, 298.9558, 298.9343, 298.8975, 283.519, 284.2079, 284.8589,
	285.5298, 286.2316, 286.9749, 287.7004, 288.4397, 288.9764, 289.7086,
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793,
	290.403, 291.0512, 291.598, 292.0377, 
    283.519, 284.2079, 284.8589, 285.5298, 286.2316, 286.9749, 287.7004, 
    288.4397, 288.9764, 289.7086, 290.403, 291.0512, 291.598, 292.0377, 
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793, 
    295.5613, 295.9263, 296.2113, 296.4967, 296.8282, 297.1194, 297.4232, 
    297.662, 297.9678, 298.1667, 298.4066, 298.5545, 298.7012, 298.8887,
	298.9477, 298.9558, 298.9343, 298.8975, 283.519, 284.2079, 284.8589,
	285.5298, 286.2316, 286.9749, 287.7004, 288.4397, 288.9764, 289.7086,
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793,
	290.403, 291.0512, 291.598, 292.0377,

    283.519, 284.2079, 284.8589, 285.5298, 286.2316, 286.9749, 287.7004, 
    288.4397, 288.9764, 289.7086, 290.403, 291.0512, 291.598, 292.0377, 
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793, 
    295.5613, 295.9263, 296.2113, 296.4967, 296.8282, 297.1194, 297.4232, 
    297.662, 297.9678, 298.1667, 298.4066, 298.5545, 298.7012, 298.8887,
	298.9477, 298.9558, 298.9343, 298.8975, 283.519, 284.2079, 284.8589,
	285.5298, 286.2316, 286.9749, 287.7004, 288.4397, 288.9764, 289.7086,
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793,
	290.403, 291.0512, 291.598, 292.0377, 
    283.519, 284.2079, 284.8589, 285.5298, 286.2316, 286.9749, 287.7004, 
    288.4397, 288.9764, 289.7086, 290.403, 291.0512, 291.598, 292.0377, 
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793, 
    295.5613, 295.9263, 296.2113, 296.4967, 296.8282, 297.1194, 297.4232, 
    297.662, 297.9678, 298.1667, 298.4066, 298.5545, 298.7012, 298.8887,
	298.9477, 298.9558, 298.9343, 298.8975, 283.519, 284.2079, 284.8589,
	285.5298, 286.2316, 286.9749, 287.7004, 288.4397, 288.9764, 289.7086,
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793,
	290.403, 291.0512, 291.598, 292.0377,

    283.519, 284.2079, 284.8589, 285.5298, 286.2316, 286.9749, 287.7004, 
    288.4397, 288.9764, 289.7086, 290.403, 291.0512, 291.598, 292.0377, 
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793, 
    295.5613, 295.9263, 296.2113, 296.4967, 296.8282, 297.1194, 297.4232, 
    297.662, 297.9678, 298.1667, 298.4066, 298.5545, 298.7012, 298.8887,
	298.9477, 298.9558, 298.9343, 298.8975, 283.519, 284.2079, 284.8589,
	285.5298, 286.2316, 286.9749, 287.7004, 288.4397, 288.9764, 289.7086,
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793,
	290.403, 291.0512, 291.598, 292.0377, 
    283.519, 284.2079, 284.8589, 285.5298, 286.2316, 286.9749, 287.7004, 
    288.4397, 288.9764, 289.7086, 290.403, 291.0512, 291.598, 292.0377, 
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793, 
    295.5613, 295.9263, 296.2113, 296.4967, 296.8282, 297.1194, 297.4232, 
    297.662, 297.9678, 298.1667, 298.4066, 298.5545, 298.7012, 298.8887,
	298.9477, 298.9558, 298.9343, 298.8975, 283.519, 284.2079, 284.8589,
	285.5298, 286.2316, 286.9749, 287.7004, 288.4397, 288.9764, 289.7086,
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793,
	290.403, 291.0512, 291.598, 292.0377,

    283.519, 284.2079, 284.8589, 285.5298, 286.2316, 286.9749, 287.7004, 
    288.4397, 288.9764, 289.7086, 290.403, 291.0512, 291.598, 292.0377, 
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793, 
    295.5613, 295.9263, 296.2113, 296.4967, 296.8282, 297.1194, 297.4232, 
    297.662, 297.9678, 298.1667, 298.4066, 298.5545, 298.7012, 298.8887,
	298.9477, 298.9558, 298.9343, 298.8975, 283.519, 284.2079, 284.8589,
	285.5298, 286.2316, 286.9749, 287.7004, 288.4397, 288.9764, 289.7086,
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793,
	290.403, 291.0512, 291.598, 292.0377, 
    283.519, 284.2079, 284.8589, 285.5298, 286.2316, 286.9749, 287.7004, 
    288.4397, 288.9764, 289.7086, 290.403, 291.0512, 291.598, 292.0377, 
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793, 
    295.5613, 295.9263, 296.2113, 296.4967, 296.8282, 297.1194, 297.4232, 
    297.662, 297.9678, 298.1667, 298.4066, 298.5545, 298.7012, 298.8887,
	298.9477, 298.9558, 298.9343, 298.8975, 283.519, 284.2079, 284.8589,
	285.5298, 286.2316, 286.9749, 287.7004, 288.4397, 288.9764, 289.7086,
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793,
	290.403, 291.0512, 291.598, 292.0377,

    283.519, 284.2079, 284.8589, 285.5298, 286.2316, 286.9749, 287.7004, 
    288.4397, 288.9764, 289.7086, 290.403, 291.0512, 291.598, 292.0377, 
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793, 
    295.5613, 295.9263, 296.2113, 296.4967, 296.8282, 297.1194, 297.4232, 
    297.662, 297.9678, 298.1667, 298.4066, 298.5545, 298.7012, 298.8887,
	298.9477, 298.9558, 298.9343, 298.8975, 283.519, 284.2079, 284.8589,
	285.5298, 286.2316, 286.9749, 287.7004, 288.4397, 288.9764, 289.7086,
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793,
	290.403, 291.0512, 291.598, 292.0377, 
    283.519, 284.2079, 284.8589, 285.5298, 286.2316, 286.9749, 287.7004, 
    288.4397, 288.9764, 289.7086, 290.403, 291.0512, 291.598, 292.0377, 
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793, 
    295.5613, 295.9263, 296.2113, 296.4967, 296.8282, 297.1194, 297.4232, 
    297.662, 297.9678, 298.1667, 298.4066, 298.5545, 298.7012, 298.8887,
	298.9477, 298.9558, 298.9343, 298.8975, 283.519, 284.2079, 284.8589,
	285.5298, 286.2316, 286.9749, 287.7004, 288.4397, 288.9764, 289.7086,
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793,
	290.403, 291.0512, 291.598, 292.0377,

    283.519, 284.2079, 284.8589, 285.5298, 286.2316, 286.9749, 287.7004, 
    288.4397, 288.9764, 289.7086, 290.403, 291.0512, 291.598, 292.0377, 
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793, 
    295.5613, 295.9263, 296.2113, 296.4967, 296.8282, 297.1194, 297.4232, 
    297.662, 297.9678, 298.1667, 298.4066, 298.5545, 298.7012, 298.8887,
	298.9477, 298.9558, 298.9343, 298.8975, 283.519, 284.2079, 284.8589,
	285.5298, 286.2316, 286.9749, 287.7004, 288.4397, 288.9764, 289.7086,
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793,
	290.403, 291.0512, 291.598, 292.0377, 
    283.519, 284.2079, 284.8589, 285.5298, 286.2316, 286.9749, 287.7004, 
    288.4397, 288.9764, 289.7086, 290.403, 291.0512, 291.598, 292.0377, 
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793, 
    295.5613, 295.9263, 296.2113, 296.4967, 296.8282, 297.1194, 297.4232, 
    297.662, 297.9678, 298.1667, 298.4066, 298.5545, 298.7012, 298.8887,
	298.9477, 298.9558, 298.9343, 298.8975, 283.519, 284.2079, 284.8589,
	285.5298, 286.2316, 286.9749, 287.7004, 288.4397, 288.9764, 289.7086,
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793,
	290.403, 291.0512, 291.598, 292.0377,

    283.519, 284.2079, 284.8589, 285.5298, 286.2316, 286.9749, 287.7004, 
    288.4397, 288.9764, 289.7086, 290.403, 291.0512, 291.598, 292.0377, 
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793, 
    295.5613, 295.9263, 296.2113, 296.4967, 296.8282, 297.1194, 297.4232, 
    297.662, 297.9678, 298.1667, 298.4066, 298.5545, 298.7012, 298.8887,
	298.9477, 298.9558, 298.9343, 298.8975, 283.519, 284.2079, 284.8589,
	285.5298, 286.2316, 286.9749, 287.7004, 288.4397, 288.9764, 289.7086,
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793,
	290.403, 291.0512, 291.598, 292.0377, 
    283.519, 284.2079, 284.8589, 285.5298, 286.2316, 286.9749, 287.7004, 
    288.4397, 288.9764, 289.7086, 290.403, 291.0512, 291.598, 292.0377, 
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793, 
    295.5613, 295.9263, 296.2113, 296.4967, 296.8282, 297.1194, 297.4232, 
    297.662, 297.9678, 298.1667, 298.4066, 298.5545, 298.7012, 298.8887,
	298.9477, 298.9558, 298.9343, 298.8975, 283.519, 284.2079, 284.8589,
	285.5298, 286.2316, 286.9749, 287.7004, 288.4397, 288.9764, 289.7086,
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793,
	290.403, 291.0512, 291.598, 292.0377,

    283.519, 284.2079, 284.8589, 285.5298, 286.2316, 286.9749, 287.7004, 
    288.4397, 288.9764, 289.7086, 290.403, 291.0512, 291.598, 292.0377, 
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793, 
    295.5613, 295.9263, 296.2113, 296.4967, 296.8282, 297.1194, 297.4232, 
    297.662, 297.9678, 298.1667, 298.4066, 298.5545, 298.7012, 298.8887,
	298.9477, 298.9558, 298.9343, 298.8975, 283.519, 284.2079, 284.8589,
	285.5298, 286.2316, 286.9749, 287.7004, 288.4397, 288.9764, 289.7086,
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793,
	290.403, 291.0512, 291.598, 292.0377, 
    283.519, 284.2079, 284.8589, 285.5298, 286.2316, 286.9749, 287.7004, 
    288.4397, 288.9764, 289.7086, 290.403, 291.0512, 291.598, 292.0377, 
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793, 
    295.5613, 295.9263, 296.2113, 296.4967, 296.8282, 297.1194, 297.4232, 
    297.662, 297.9678, 298.1667, 298.4066, 298.5545, 298.7012, 298.8887,
	298.9477, 298.9558, 298.9343, 298.8975, 283.519, 284.2079, 284.8589,
	285.5298, 286.2316, 286.9749, 287.7004, 288.4397, 288.9764, 289.7086,
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793,
	290.403, 291.0512, 291.598, 292.0377,

    283.519, 284.2079, 284.8589, 285.5298, 286.2316, 286.9749, 287.7004, 
    288.4397, 288.9764, 289.7086, 290.403, 291.0512, 291.598, 292.0377, 
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793, 
    295.5613, 295.9263, 296.2113, 296.4967, 296.8282, 297.1194, 297.4232, 
    297.662, 297.9678, 298.1667, 298.4066, 298.5545, 298.7012, 298.8887,
	298.9477, 298.9558, 298.9343, 298.8975, 283.519, 284.2079, 284.8589,
	285.5298, 286.2316, 286.9749, 287.7004, 288.4397, 288.9764, 289.7086,
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793,
	290.403, 291.0512, 291.598, 292.0377, 
    283.519, 284.2079, 284.8589, 285.5298, 286.2316, 286.9749, 287.7004, 
    288.4397, 288.9764, 289.7086, 290.403, 291.0512, 291.598, 292.0377, 
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793, 
    295.5613, 295.9263, 296.2113, 296.4967, 296.8282, 297.1194, 297.4232, 
    297.662, 297.9678, 298.1667, 298.4066, 298.5545, 298.7012, 298.8887,
	298.9477, 298.9558, 298.9343, 298.8975, 283.519, 284.2079, 284.8589,
	285.5298, 286.2316, 286.9749, 287.7004, 288.4397, 288.9764, 289.7086,
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793,
	290.403, 291.0512, 291.598, 292.0377,

    283.519, 284.2079, 284.8589, 285.5298, 286.2316, 286.9749, 287.7004, 
    288.4397, 288.9764, 289.7086, 290.403, 291.0512, 291.598, 292.0377, 
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793, 
    295.5613, 295.9263, 296.2113, 296.4967, 296.8282, 297.1194, 297.4232, 
    297.662, 297.9678, 298.1667, 298.4066, 298.5545, 298.7012, 298.8887,
	298.9477, 298.9558, 298.9343, 298.8975, 283.519, 284.2079, 284.8589,
	285.5298, 286.2316, 286.9749, 287.7004, 288.4397, 288.9764, 289.7086,
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793,
	290.403, 291.0512, 291.598, 292.0377, 
    283.519, 284.2079, 284.8589, 285.5298, 286.2316, 286.9749, 287.7004, 
    288.4397, 288.9764, 289.7086, 290.403, 291.0512, 291.598, 292.0377, 
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793, 
    295.5613, 295.9263, 296.2113, 296.4967, 296.8282, 297.1194, 297.4232, 
    297.662, 297.9678, 298.1667, 298.4066, 298.5545, 298.7012, 298.8887,
	298.9477, 298.9558, 298.9343, 298.8975, 283.519, 284.2079, 284.8589,
	285.5298, 286.2316, 286.9749, 287.7004, 288.4397, 288.9764, 289.7086,
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793,
	290.403, 291.0512, 291.598, 292.0377,

    283.519, 284.2079, 284.8589, 285.5298, 286.2316, 286.9749, 287.7004, 
    288.4397, 288.9764, 289.7086, 290.403, 291.0512, 291.598, 292.0377, 
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793, 
    295.5613, 295.9263, 296.2113, 296.4967, 296.8282, 297.1194, 297.4232, 
    297.662, 297.9678, 298.1667, 298.4066, 298.5545, 298.7012, 298.8887,
	298.9477, 298.9558, 298.9343, 298.8975, 283.519, 284.2079, 284.8589,
	285.5298, 286.2316, 286.9749, 287.7004, 288.4397, 288.9764, 289.7086,
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793,
	290.403, 291.0512, 291.598, 292.0377, 
    283.519, 284.2079, 284.8589, 285.5298, 286.2316, 286.9749, 287.7004, 
    288.4397, 288.9764, 289.7086, 290.403, 291.0512, 291.598, 292.0377, 
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793, 
    295.5613, 295.9263, 296.2113, 296.4967, 296.8282, 297.1194, 297.4232, 
    297.662, 297.9678, 298.1667, 298.4066, 298.5545, 298.7012, 298.8887,
	298.9477, 298.9558, 298.9343, 298.8975, 283.519, 284.2079, 284.8589,
	285.5298, 286.2316, 286.9749, 287.7004, 288.4397, 288.9764, 289.7086,
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793,
	290.403, 291.0512, 291.598, 292.0377,

    283.519, 284.2079, 284.8589, 285.5298, 286.2316, 286.9749, 287.7004, 
    288.4397, 288.9764, 289.7086, 290.403, 291.0512, 291.598, 292.0377, 
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793, 
    295.5613, 295.9263, 296.2113, 296.4967, 296.8282, 297.1194, 297.4232, 
    297.662, 297.9678, 298.1667, 298.4066, 298.5545, 298.7012, 298.8887,
	298.9477, 298.9558, 298.9343, 298.8975, 283.519, 284.2079, 284.8589,
	285.5298, 286.2316, 286.9749, 287.7004, 288.4397, 288.9764, 289.7086,
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793,
	290.403, 291.0512, 291.598, 292.0377, 
    283.519, 284.2079, 284.8589, 285.5298, 286.2316, 286.9749, 287.7004, 
    288.4397, 288.9764, 289.7086, 290.403, 291.0512, 291.598, 292.0377, 
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793, 
    295.5613, 295.9263, 296.2113, 296.4967, 296.8282, 297.1194, 297.4232, 
    297.662, 297.9678, 298.1667, 298.4066, 298.5545, 298.7012, 298.8887,
	298.9477, 298.9558, 298.9343, 298.8975, 283.519, 284.2079, 284.8589,
	285.5298, 286.2316, 286.9749, 287.7004, 288.4397, 288.9764, 289.7086,
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793,
	290.403, 291.0512, 291.598, 292.0377,

    283.519, 284.2079, 284.8589, 285.5298, 286.2316, 286.9749, 287.7004, 
    288.4397, 288.9764, 289.7086, 290.403, 291.0512, 291.598, 292.0377, 
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793, 
    295.5613, 295.9263, 296.2113, 296.4967, 296.8282, 297.1194, 297.4232, 
    297.662, 297.9678, 298.1667, 298.4066, 298.5545, 298.7012, 298.8887,
	298.9477, 298.9558, 298.9343, 298.8975, 283.519, 284.2079, 284.8589,
	285.5298, 286.2316, 286.9749, 287.7004, 288.4397, 288.9764, 289.7086,
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793,
	290.403, 291.0512, 291.598, 292.0377, 
    283.519, 284.2079, 284.8589, 285.5298, 286.2316, 286.9749, 287.7004, 
    288.4397, 288.9764, 289.7086, 290.403, 291.0512, 291.598, 292.0377, 
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793, 
    295.5613, 295.9263, 296.2113, 296.4967, 296.8282, 297.1194, 297.4232, 
    297.662, 297.9678, 298.1667, 298.4066, 298.5545, 298.7012, 298.8887,
	298.9477, 298.9558, 298.9343, 298.8975, 283.519, 284.2079, 284.8589,
	285.5298, 286.2316, 286.9749, 287.7004, 288.4397, 288.9764, 289.7086,
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793,
	290.403, 291.0512, 291.598, 292.0377,

    283.519, 284.2079, 284.8589, 285.5298, 286.2316, 286.9749, 287.7004, 
    288.4397, 288.9764, 289.7086, 290.403, 291.0512, 291.598, 292.0377, 
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793, 
    295.5613, 295.9263, 296.2113, 296.4967, 296.8282, 297.1194, 297.4232, 
    297.662, 297.9678, 298.1667, 298.4066, 298.5545, 298.7012, 298.8887,
	298.9477, 298.9558, 298.9343, 298.8975, 283.519, 284.2079, 284.8589,
	285.5298, 286.2316, 286.9749, 287.7004, 288.4397, 288.9764, 289.7086,
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793,
	290.403, 291.0512, 291.598, 292.0377, 
    283.519, 284.2079, 284.8589, 285.5298, 286.2316, 286.9749, 287.7004, 
    288.4397, 288.9764, 289.7086, 290.403, 291.0512, 291.598, 292.0377, 
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793, 
    295.5613, 295.9263, 296.2113, 296.4967, 296.8282, 297.1194, 297.4232, 
    297.662, 297.9678, 298.1667, 298.4066, 298.5545, 298.7012, 298.8887,
	298.9477, 298.9558, 298.9343, 298.8975, 283.519, 284.2079, 284.8589,
	285.5298, 286.2316, 286.9749, 287.7004, 288.4397, 288.9764, 289.7086,
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793,
	290.403, 291.0512, 291.598, 292.0377,

    283.519, 284.2079, 284.8589, 285.5298, 286.2316, 286.9749, 287.7004, 
    288.4397, 288.9764, 289.7086, 290.403, 291.0512, 291.598, 292.0377, 
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793, 
    295.5613, 295.9263, 296.2113, 296.4967, 296.8282, 297.1194, 297.4232, 
    297.662, 297.9678, 298.1667, 298.4066, 298.5545, 298.7012, 298.8887,
	298.9477, 298.9558, 298.9343, 298.8975, 283.519, 284.2079, 284.8589,
	285.5298, 286.2316, 286.9749, 287.7004, 288.4397, 288.9764, 289.7086,
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793,
	290.403, 291.0512, 291.598, 292.0377, 
    283.519, 284.2079, 284.8589, 285.5298, 286.2316, 286.9749, 287.7004, 
    288.4397, 288.9764, 289.7086, 290.403, 291.0512, 291.598, 292.0377, 
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793, 
    295.5613, 295.9263, 296.2113, 296.4967, 296.8282, 297.1194, 297.4232, 
    297.662, 297.9678, 298.1667, 298.4066, 298.5545, 298.7012, 298.8887,
	298.9477, 298.9558, 298.9343, 298.8975, 283.519, 284.2079, 284.8589,
	285.5298, 286.2316, 286.9749, 287.7004, 288.4397, 288.9764, 289.7086,
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793,
	290.403, 291.0512, 291.598, 292.0377,

    283.519, 284.2079, 284.8589, 285.5298, 286.2316, 286.9749, 287.7004, 
    288.4397, 288.9764, 289.7086, 290.403, 291.0512, 291.598, 292.0377, 
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793, 
    295.5613, 295.9263, 296.2113, 296.4967, 296.8282, 297.1194, 297.4232, 
    297.662, 297.9678, 298.1667, 298.4066, 298.5545, 298.7012, 298.8887,
	298.9477, 298.9558, 298.9343, 298.8975, 283.519, 284.2079, 284.8589,
	285.5298, 286.2316, 286.9749, 287.7004, 288.4397, 288.9764, 289.7086,
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793,
	290.403, 291.0512, 291.598, 292.0377, 
    283.519, 284.2079, 284.8589, 285.5298, 286.2316, 286.9749, 287.7004, 
    288.4397, 288.9764, 289.7086, 290.403, 291.0512, 291.598, 292.0377, 
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793, 
    295.5613, 295.9263, 296.2113, 296.4967, 296.8282, 297.1194, 297.4232, 
    297.662, 297.9678, 298.1667, 298.4066, 298.5545, 298.7012, 298.8887,
	298.9477, 298.9558, 298.9343, 298.8975, 283.519, 284.2079, 284.8589,
	285.5298, 286.2316, 286.9749, 287.7004, 288.4397, 288.9764, 289.7086,
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793,
	290.403, 291.0512, 291.598, 292.0377,

    283.519, 284.2079, 284.8589, 285.5298, 286.2316, 286.9749, 287.7004, 
    288.4397, 288.9764, 289.7086, 290.403, 291.0512, 291.598, 292.0377, 
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793, 
    295.5613, 295.9263, 296.2113, 296.4967, 296.8282, 297.1194, 297.4232, 
    297.662, 297.9678, 298.1667, 298.4066, 298.5545, 298.7012, 298.8887,
	298.9477, 298.9558, 298.9343, 298.8975, 283.519, 284.2079, 284.8589,
	285.5298, 286.2316, 286.9749, 287.7004, 288.4397, 288.9764, 289.7086,
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793,
	290.403, 291.0512, 291.598, 292.0377, 
    283.519, 284.2079, 284.8589, 285.5298, 286.2316, 286.9749, 287.7004, 
    288.4397, 288.9764, 289.7086, 290.403, 291.0512, 291.598, 292.0377, 
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793, 
    295.5613, 295.9263, 296.2113, 296.4967, 296.8282, 297.1194, 297.4232, 
    297.662, 297.9678, 298.1667, 298.4066, 298.5545, 298.7012, 298.8887,
	298.9477, 298.9558, 298.9343, 298.8975, 283.519, 284.2079, 284.8589,
	285.5298, 286.2316, 286.9749, 287.7004, 288.4397, 288.9764, 289.7086,
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793,
	290.403, 291.0512, 291.598, 292.0377,

    283.519, 284.2079, 284.8589, 285.5298, 286.2316, 286.9749, 287.7004, 
    288.4397, 288.9764, 289.7086, 290.403, 291.0512, 291.598, 292.0377, 
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793, 
    295.5613, 295.9263, 296.2113, 296.4967, 296.8282, 297.1194, 297.4232, 
    297.662, 297.9678, 298.1667, 298.4066, 298.5545, 298.7012, 298.8887,
	298.9477, 298.9558, 298.9343, 298.8975, 283.519, 284.2079, 284.8589,
	285.5298, 286.2316, 286.9749, 287.7004, 288.4397, 288.9764, 289.7086,
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793,
	290.403, 291.0512, 291.598, 292.0377, 
    283.519, 284.2079, 284.8589, 285.5298, 286.2316, 286.9749, 287.7004, 
    288.4397, 288.9764, 289.7086, 290.403, 291.0512, 291.598, 292.0377, 
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793, 
    295.5613, 295.9263, 296.2113, 296.4967, 296.8282, 297.1194, 297.4232, 
    297.662, 297.9678, 298.1667, 298.4066, 298.5545, 298.7012, 298.8887,
	298.9477, 298.9558, 298.9343, 298.8975, 283.519, 284.2079, 284.8589,
	285.5298, 286.2316, 286.9749, 287.7004, 288.4397, 288.9764, 289.7086,
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793,
	290.403, 291.0512, 291.598, 292.0377,

    283.519, 284.2079, 284.8589, 285.5298, 286.2316, 286.9749, 287.7004, 
    288.4397, 288.9764, 289.7086, 290.403, 291.0512, 291.598, 292.0377, 
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793, 
    295.5613, 295.9263, 296.2113, 296.4967, 296.8282, 297.1194, 297.4232, 
    297.662, 297.9678, 298.1667, 298.4066, 298.5545, 298.7012, 298.8887,
	298.9477, 298.9558, 298.9343, 298.8975, 283.519, 284.2079, 284.8589,
	285.5298, 286.2316, 286.9749, 287.7004, 288.4397, 288.9764, 289.7086,
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793,
	290.403, 291.0512, 291.598, 292.0377, 
    283.519, 284.2079, 284.8589, 285.5298, 286.2316, 286.9749, 287.7004, 
    288.4397, 288.9764, 289.7086, 290.403, 291.0512, 291.598, 292.0377, 
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793, 
    295.5613, 295.9263, 296.2113, 296.4967, 296.8282, 297.1194, 297.4232, 
    297.662, 297.9678, 298.1667, 298.4066, 298.5545, 298.7012, 298.8887,
	298.9477, 298.9558, 298.9343, 298.8975, 283.519, 284.2079, 284.8589,
	285.5298, 286.2316, 286.9749, 287.7004, 288.4397, 288.9764, 289.7086,
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793,
	290.403, 291.0512, 291.598, 292.0377,

    283.519, 284.2079, 284.8589, 285.5298, 286.2316, 286.9749, 287.7004, 
    288.4397, 288.9764, 289.7086, 290.403, 291.0512, 291.598, 292.0377, 
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793, 
    295.5613, 295.9263, 296.2113, 296.4967, 296.8282, 297.1194, 297.4232, 
    297.662, 297.9678, 298.1667, 298.4066, 298.5545, 298.7012, 298.8887,
	298.9477, 298.9558, 298.9343, 298.8975, 283.519, 284.2079, 284.8589,
	285.5298, 286.2316, 286.9749, 287.7004, 288.4397, 288.9764, 289.7086,
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793,
	290.403, 291.0512, 291.598, 292.0377, 
    283.519, 284.2079, 284.8589, 285.5298, 286.2316, 286.9749, 287.7004, 
    288.4397, 288.9764, 289.7086, 290.403, 291.0512, 291.598, 292.0377, 
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793, 
    295.5613, 295.9263, 296.2113, 296.4967, 296.8282, 297.1194, 297.4232, 
    297.662, 297.9678, 298.1667, 298.4066, 298.5545, 298.7012, 298.8887,
	298.9477, 298.9558, 298.9343, 298.8975, 283.519, 284.2079, 284.8589,
	285.5298, 286.2316, 286.9749, 287.7004, 288.4397, 288.9764, 289.7086,
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793,
	290.403, 291.0512, 291.598, 292.0377,

    283.519, 284.2079, 284.8589, 285.5298, 286.2316, 286.9749, 287.7004, 
    288.4397, 288.9764, 289.7086, 290.403, 291.0512, 291.598, 292.0377, 
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793, 
    295.5613, 295.9263, 296.2113, 296.4967, 296.8282, 297.1194, 297.4232, 
    297.662, 297.9678, 298.1667, 298.4066, 298.5545, 298.7012, 298.8887,
	298.9477, 298.9558, 298.9343, 298.8975, 283.519, 284.2079, 284.8589,
	285.5298, 286.2316, 286.9749, 287.7004, 288.4397, 288.9764, 289.7086,
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793,
	290.403, 291.0512, 291.598, 292.0377, 
    283.519, 284.2079, 284.8589, 285.5298, 286.2316, 286.9749, 287.7004, 
    288.4397, 288.9764, 289.7086, 290.403, 291.0512, 291.598, 292.0377, 
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793, 
    295.5613, 295.9263, 296.2113, 296.4967, 296.8282, 297.1194, 297.4232, 
    297.662, 297.9678, 298.1667, 298.4066, 298.5545, 298.7012, 298.8887,
	298.9477, 298.9558, 298.9343, 298.8975, 283.519, 284.2079, 284.8589,
	285.5298, 286.2316, 286.9749, 287.7004, 288.4397, 288.9764, 289.7086,
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793,
	290.403, 291.0512, 291.598, 292.0377,

    283.519, 284.2079, 284.8589, 285.5298, 286.2316, 286.9749, 287.7004, 
    288.4397, 288.9764, 289.7086, 290.403, 291.0512, 291.598, 292.0377, 
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793, 
    295.5613, 295.9263, 296.2113, 296.4967, 296.8282, 297.1194, 297.4232, 
    297.662, 297.9678, 298.1667, 298.4066, 298.5545, 298.7012, 298.8887,
	298.9477, 298.9558, 298.9343, 298.8975, 283.519, 284.2079, 284.8589,
	285.5298, 286.2316, 286.9749, 287.7004, 288.4397, 288.9764, 289.7086,
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793,
	290.403, 291.0512, 291.598, 292.0377, 
    283.519, 284.2079, 284.8589, 285.5298, 286.2316, 286.9749, 287.7004, 
    288.4397, 288.9764, 289.7086, 290.403, 291.0512, 291.598, 292.0377, 
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793, 
    295.5613, 295.9263, 296.2113, 296.4967, 296.8282, 297.1194, 297.4232, 
    297.662, 297.9678, 298.1667, 298.4066, 298.5545, 298.7012, 298.8887,
	298.9477, 298.9558, 298.9343, 298.8975, 283.519, 284.2079, 284.8589,
	285.5298, 286.2316, 286.9749, 287.7004, 288.4397, 288.9764, 289.7086,
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793,
	290.403, 291.0512, 291.598, 292.0377,

    283.519, 284.2079, 284.8589, 285.5298, 286.2316, 286.9749, 287.7004, 
    288.4397, 288.9764, 289.7086, 290.403, 291.0512, 291.598, 292.0377, 
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793, 
    295.5613, 295.9263, 296.2113, 296.4967, 296.8282, 297.1194, 297.4232, 
    297.662, 297.9678, 298.1667, 298.4066, 298.5545, 298.7012, 298.8887,
	298.9477, 298.9558, 298.9343, 298.8975, 283.519, 284.2079, 284.8589,
	285.5298, 286.2316, 286.9749, 287.7004, 288.4397, 288.9764, 289.7086,
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793,
	290.403, 291.0512, 291.598, 292.0377, 
    283.519, 284.2079, 284.8589, 285.5298, 286.2316, 286.9749, 287.7004, 
    288.4397, 288.9764, 289.7086, 290.403, 291.0512, 291.598, 292.0377, 
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793, 
    295.5613, 295.9263, 296.2113, 296.4967, 296.8282, 297.1194, 297.4232, 
    297.662, 297.9678, 298.1667, 298.4066, 298.5545, 298.7012, 298.8887,
	298.9477, 298.9558, 298.9343, 298.8975, 283.519, 284.2079, 284.8589,
	285.5298, 286.2316, 286.9749, 287.7004, 288.4397, 288.9764, 289.7086,
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793,
	290.403, 291.0512, 291.598, 292.0377,

    283.519, 284.2079, 284.8589, 285.5298, 286.2316, 286.9749, 287.7004, 
    288.4397, 288.9764, 289.7086, 290.403, 291.0512, 291.598, 292.0377, 
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793, 
    295.5613, 295.9263, 296.2113, 296.4967, 296.8282, 297.1194, 297.4232, 
    297.662, 297.9678, 298.1667, 298.4066, 298.5545, 298.7012, 298.8887,
	298.9477, 298.9558, 298.9343, 298.8975, 283.519, 284.2079, 284.8589,
	285.5298, 286.2316, 286.9749, 287.7004, 288.4397, 288.9764, 289.7086,
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793,
	290.403, 291.0512, 291.598, 292.0377, 
    283.519, 284.2079, 284.8589, 285.5298, 286.2316, 286.9749, 287.7004, 
    288.4397, 288.9764, 289.7086, 290.403, 291.0512, 291.598, 292.0377, 
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793, 
    295.5613, 295.9263, 296.2113, 296.4967, 296.8282, 297.1194, 297.4232, 
    297.662, 297.9678, 298.1667, 298.4066, 298.5545, 298.7012, 298.8887,
	298.9477, 298.9558, 298.9343, 298.8975, 283.519, 284.2079, 284.8589,
	285.5298, 286.2316, 286.9749, 287.7004, 288.4397, 288.9764, 289.7086,
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793,
	290.403, 291.0512, 291.598, 292.0377,

    283.519, 284.2079, 284.8589, 285.5298, 286.2316, 286.9749, 287.7004, 
    288.4397, 288.9764, 289.7086, 290.403, 291.0512, 291.598, 292.0377, 
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793, 
    295.5613, 295.9263, 296.2113, 296.4967, 296.8282, 297.1194, 297.4232, 
    297.662, 297.9678, 298.1667, 298.4066, 298.5545, 298.7012, 298.8887,
	298.9477, 298.9558, 298.9343, 298.8975, 283.519, 284.2079, 284.8589,
	285.5298, 286.2316, 286.9749, 287.7004, 288.4397, 288.9764, 289.7086,
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793,
	290.403, 291.0512, 291.598, 292.0377, 
    283.519, 284.2079, 284.8589, 285.5298, 286.2316, 286.9749, 287.7004, 
    288.4397, 288.9764, 289.7086, 290.403, 291.0512, 291.598, 292.0377, 
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793, 
    295.5613, 295.9263, 296.2113, 296.4967, 296.8282, 297.1194, 297.4232, 
    297.662, 297.9678, 298.1667, 298.4066, 298.5545, 298.7012, 298.8887,
	298.9477, 298.9558, 298.9343, 298.8975, 283.519, 284.2079, 284.8589,
	285.5298, 286.2316, 286.9749, 287.7004, 288.4397, 288.9764, 289.7086,
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793,
	290.403, 291.0512, 291.598, 292.0377,

    283.519, 284.2079, 284.8589, 285.5298, 286.2316, 286.9749, 287.7004, 
    288.4397, 288.9764, 289.7086, 290.403, 291.0512, 291.598, 292.0377, 
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793, 
    295.5613, 295.9263, 296.2113, 296.4967, 296.8282, 297.1194, 297.4232, 
    297.662, 297.9678, 298.1667, 298.4066, 298.5545, 298.7012, 298.8887,
	298.9477, 298.9558, 298.9343, 298.8975, 283.519, 284.2079, 284.8589,
	285.5298, 286.2316, 286.9749, 287.7004, 288.4397, 288.9764, 289.7086,
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793,
	290.403, 291.0512, 291.598, 292.0377, 
    283.519, 284.2079, 284.8589, 285.5298, 286.2316, 286.9749, 287.7004, 
    288.4397, 288.9764, 289.7086, 290.403, 291.0512, 291.598, 292.0377, 
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793, 
    295.5613, 295.9263, 296.2113, 296.4967, 296.8282, 297.1194, 297.4232, 
    297.662, 297.9678, 298.1667, 298.4066, 298.5545, 298.7012, 298.8887,
	298.9477, 298.9558, 298.9343, 298.8975, 283.519, 284.2079, 284.8589,
	285.5298, 286.2316, 286.9749, 287.7004, 288.4397, 288.9764, 289.7086,
    292.5377, 293.0864, 293.6501, 294.1322, 294.6041, 295.0236, 295.2793,
	290.403, 291.0512, 291.598, 292.0377 ;

 time = 15.5, 45, 74.5, 105, 135.5, 166, 196.5, 227.5, 258, 288.5, 319, 
    349.5, 380.5, 410, 439.5, 470, 500.5, 531, 561.5, 592.5, 623, 653.5, 684, 
    714.5, 745.5, 775, 804.5, 835, 865.5, 896, 926.5, 957.5, 988, 1018.5, 
    1049, 1079.5, 1110.5, 1140, 1169.5, 1200, 1230.5, 1261, 1291.5, 1322.5, 
    1353, 1383.5, 1414, 1444.5, 1475.5, 1505, 1534.5, 1565, 1595.5, 1626, 
    1656.5, 1687.5, 1718, 1748.5, 1779, 1809.5 ;

 time_bnds =
  0, 31,
  31, 59,
  59, 90,
  90, 120,
  120, 151,
  151, 181,
  181, 212,
  212, 243,
  243, 273,
  273, 304,
  304, 334,
  334, 365,
  365, 396,
  396, 424,
  424, 455,
  455, 485,
  485, 516,
  516, 546,
  546, 577,
  577, 608,
  608, 638,
  638, 669,
  669, 699,
  699, 730,
  730, 761,
  761, 789,
  789, 820,
  820, 850,
  850, 881,
  881, 911,
  911, 942,
  942, 973,
  973, 1003,
  1003, 1034,
  1034, 1064,
  1064, 1095,
  1095, 1126,
  1126, 1154,
  1154, 1185,
  1185, 1215,
  1215, 1246,
  1246, 1276,
  1276, 1307,
  1307, 1338,
  1338, 1368,
  1368, 1399,
  1399, 1429,
  1429, 1460,
  1460, 1491,
  1491, 1519,
  1519, 1550,
  1550, 1580,
  1580, 1611,
  1611, 1641,
  1641, 1672,
  1672, 1703,
  1703, 1733,
  1733, 1764,
  1764, 1794,
  1794, 1825 ;
}
