netcdf atmos.1980-1981.alb_sfc.11 {
dimensions:
	time = UNLIMITED ; // (1 currently)
	lat = 18 ;
	lon = 29 ;
	bnds = 2 ;
variables:
	float alb_sfc(time, lat, lon) ;
		alb_sfc:long_name = "Surface Albedo for  Flux" ;
		alb_sfc:units = "percent" ;
		alb_sfc:_FillValue = 1.e+20f ;
		alb_sfc:missing_value = 1.e+20f ;
		alb_sfc:cell_measures = "area: area" ;
		alb_sfc:interp_method = "conserve_order1" ;
		alb_sfc:cell_methods = "time: mean within months time: mean over years" ;
		alb_sfc:time_avg_info = "average_T1,average_T2,average_DT" ;
	double average_DT(time) ;
		average_DT:long_name = "Length of average period" ;
		average_DT:units = "days" ;
	double average_T1(time) ;
		average_T1:long_name = "Start time for average period" ;
		average_T1:units = "days since 1979-01-01 00:00:00" ;
	double average_T2(time) ;
		average_T2:long_name = "End time for average period" ;
		average_T2:units = "days since 1979-01-01 00:00:00" ;
	double climatology_bounds(time, bnds) ;
	double lat(lat) ;
		lat:standard_name = "latitude" ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_N" ;
		lat:axis = "Y" ;
		lat:bounds = "lat_bnds" ;
	double lat_bnds(lat, bnds) ;
	double lon(lon) ;
		lon:standard_name = "longitude" ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_E" ;
		lon:axis = "X" ;
		lon:bounds = "lon_bnds" ;
	double lon_bnds(lon, bnds) ;
	double time(time) ;
		time:standard_name = "time" ;
		time:long_name = "time" ;
		time:climatology = "climatology_bounds" ;
		time:units = "days since 1979-01-01 00:00:00" ;
		time:calendar = "standard" ;
		time:axis = "T" ;

// global attributes:
		:CDI = "Climate Data Interface version 2.4.4 (https://mpimet.mpg.de/cdi)" ;
		:Conventions = "CF-1.6" ;
		:title = "c96L65_am5f9d8r0_amip" ;
		:associated_files = "area: 19800101.grid_spec.nc" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
		:code_release_version = "2024.05" ;
		:git_hash = "5d306c05d9fe755cab04eedc8fd3de0d3c8355a0" ;
		:creationtime = "Mon Aug 25 14:09:46 2025" ;
		:hostname = "pp050" ;
		:history = "Mon Aug 25 13:32:22 2025: ncks -d lat,,,10 -d lon,,,10 atmos.1980-1981.alb_sfc.11.nc reduced/atmos.1980-1981.alb_sfc.11.nc\n",
			"Mon Aug 25 14:40:09 2025: cdo -O -s -select,month=11 merged_output.nc monthly_nc_files/all_years.11.nc\n",
			"Mon Aug 25 14:40:01 2025: cdo -O -s -mergetime /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/shards/ts/regrid-xy/180_288.conserve_order2/atmos_month/P1M/P1Y/atmos_month.198001-198012.alb_sfc.nc /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/shards/ts/regrid-xy/180_288.conserve_order2/atmos_month/P1M/P1Y/atmos_month.198101-198112.alb_sfc.nc merged_output.nc\n",
			"Mon Aug 25 14:12:17 2025: cdo --history splitname 19800101.atmos_month.nc /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/cycle/19800101T0000Z/split/regrid-xy/180_288.conserve_order2/19800101.atmos_month.\n",
			"fregrid --debug --standard_dimension --input_mosaic C96_mosaic.nc --input_dir /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/cycle/19800101T0000Z/history/native --input_file 19800101.atmos_month --associated_file_dir /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/cycle/19800101T0000Z/history/native --interp_method conserve_order2 --remap_file fregrid_remap_file_288_by_180.nc --nlon 288 --nlat 180 --scalar_field (**please see the field list in this file**) --output_file 19800101.atmos_month.nc" ;
		:CDO = "Climate Data Operators version 2.4.4 (https://mpimet.mpg.de/cdo)" ;
		:comment = "FMS time averaging, version 3.0, precision=double" ;
		:NCO = "netCDF Operators version 5.2.4 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco, Citation = 10.1016/j.envsoft.2008.03.004)" ;
data:

 alb_sfc =
  76.28321, 76.28321, 76.28321, 76.28321, 76.28321, 76.28321, 76.28321, 
    76.27275, 76.27275, 76.27275, 76.27275, 76.27275, 76.27275, 76.27275, 
    76.26085, 76.26085, 76.26085, 76.26085, 76.26085, 76.26085, 76.26085, 
    76.30629, 76.30629, 76.30629, 76.30629, 76.30629, 76.30629, 76.30629, 
    76.28321,
  76.33073, 76.21892, 76.12687, 76.08855, 76.0436, 76.05582, 76.04623, 
    76.00616, 76.01494, 76.03448, 76.06387, 76.13065, 76.21382, 76.52481, 
    76.5704, 76.69276, 76.4317, 76.48534, 76.5417, 76.5211, 76.61867, 
    76.60396, 77.12971, 75.07339, 74.12468, 74.492, 74.04332, 76.05251, 
    76.3915,
  65.19052, 51.79762, 69.10509, 68.80449, 68.13489, 68.14877, 64.6349, 
    67.73249, 67.44228, 67.58685, 67.63368, 67.57153, 67.7093, 76.76891, 
    75.76566, 73.66827, 71.37943, 71.98882, 71.36288, 70.99538, 69.53935, 
    57.35296, 61.86291, 60.45116, 63.49646, 63.12741, 61.11821, 61.73548, 
    63.4162,
  42.9173, 47.09008, 35.32267, 7.009246, 5.145768, 4.890486, 8.231593, 
    4.96782, 6.935204, 4.979663, 4.980195, 4.938543, 4.937977, 4.935597, 
    5.093824, 4.91185, 4.805215, 4.791977, 5.047561, 5.044189, 5.106452, 
    5.064185, 5.088437, 5.006056, 4.825216, 10.43241, 33.53594, 35.90094, 
    42.75307,
  4.142395, 4.284228, 4.388851, 4.418045, 4.41597, 4.352337, 4.3191, 
    4.385942, 4.38787, 4.384038, 4.387404, 4.398344, 4.452306, 4.244187, 
    4.362875, 4.377433, 4.355393, 4.258412, 4.183645, 4.264458, 4.205622, 
    4.293778, 4.155342, 8.690409, 4.799713, 4.417268, 4.224765, 4.218978, 
    4.271422,
  3.942469, 3.994837, 4.299252, 4.020767, 4.044106, 4.026037, 3.96878, 
    3.98288, 3.820512, 4.000469, 3.85624, 4.096023, 4.218265, 4.108027, 
    10.00251, 3.879276, 3.920696, 3.862439, 4.058027, 3.911481, 3.845759, 
    3.894607, 3.955948, 9.882301, 4.324738, 4.091618, 3.814946, 3.950861, 
    3.852124,
  3.910253, 4.05676, 12.90845, 3.751325, 3.793828, 3.773717, 3.840524, 
    3.817252, 3.720776, 4.158886, 10.24454, 15.8526, 11.1237, 3.818633, 
    3.804595, 3.922285, 3.853743, 3.787419, 3.786406, 3.652873, 3.747263, 
    3.93185, 3.758221, 4.774544, 9.745634, 3.838506, 3.769886, 3.83898, 
    3.86746,
  3.313769, 10.43597, 10.55423, 3.704276, 3.688191, 3.779661, 3.866831, 
    3.73739, 3.812957, 3.727036, 12.59037, 12.19861, 3.672113, 3.64335, 
    3.687149, 3.805719, 3.58829, 3.630629, 3.475151, 4.024055, 3.850879, 
    3.676029, 3.354238, 3.594729, 9.375131, 9.329957, 3.783937, 3.561587, 
    3.613341,
  3.22937, 6.190372, 8.831119, 9.187737, 3.53105, 3.358895, 3.503801, 
    3.393708, 3.46354, 3.401496, 4.983201, 3.355683, 4.565188, 3.443879, 
    3.352483, 3.577514, 3.47636, 3.784834, 3.640507, 3.975571, 3.605827, 
    3.469147, 3.287411, 8.771511, 8.680509, 8.993187, 3.689122, 3.495514, 
    3.623564,
  3.195363, 8.314839, 8.219286, 9.613474, 3.472168, 3.458517, 3.526326, 
    3.367467, 8.435708, 8.32423, 3.233224, 3.370108, 3.245116, 3.468582, 
    3.543793, 3.635197, 3.688558, 3.798904, 3.632118, 3.802565, 3.462997, 
    3.214236, 3.408481, 8.417072, 8.406038, 3.460675, 3.386421, 3.467225, 
    3.381497,
  9.831889, 10.11974, 9.913081, 9.345377, 14.2288, 3.451887, 5.17906, 
    3.491068, 3.45395, 3.293067, 4.043437, 3.441373, 3.152276, 3.172021, 
    3.364024, 3.316625, 3.527467, 3.269423, 3.536421, 3.218539, 3.403562, 
    3.322315, 8.567595, 7.361147, 3.513149, 3.584383, 3.169573, 3.445986, 
    8.827256,
  16.55211, 18.70415, 20.50001, 3.764664, 20.67388, 3.813122, 10.5044, 
    3.824242, 8.743545, 3.578709, 3.311585, 3.555695, 3.697256, 3.796683, 
    3.92872, 3.759367, 3.854741, 3.656994, 3.620532, 3.514278, 3.920097, 
    5.975677, 3.667953, 4.297356, 3.657661, 3.731857, 3.466843, 3.644318, 
    21.14793,
  20.52013, 17.15657, 17.68227, 16.45034, 11.23848, 12.84089, 10.99735, 
    17.9341, 8.815908, 9.652834, 3.578817, 3.746892, 3.88652, 3.828691, 
    3.63179, 3.770017, 3.752579, 3.869717, 3.622046, 4.21103, 9.149229, 
    10.67795, 8.240385, 3.779605, 3.75184, 3.595713, 3.904256, 3.978267, 
    9.623957,
  5.888193, 4.19626, 5.521075, 8.964939, 1.644011, 12.25978, 10.1837, 
    12.29495, 10.94318, 10.41779, 7.062436, 3.535761, 3.707375, 3.558279, 
    3.695022, 3.791929, 3.392071, 3.368127, 3.575197, 9.972665, 9.898775, 
    11.45455, 10.2675, 4.281878, 3.603737, 3.543788, 3.63715, 3.723872, 
    4.781573,
  4.903425, 8.637146, 9.367579, 9.796785, 8.968102, 8.808298, 6.473489, 
    25.63412, 11.47304, 6.612338, 8.035072, 11.02518, 3.474778, 3.56885, 
    3.866337, 3.735358, 3.565325, 3.412671, 3.26757, 8.31568, 9.047657, 
    9.819481, 9.363935, 16.09324, 4.478539, 3.521692, 3.533371, 3.62005, 
    3.928103,
  3.6887, 9.049425, 6.119119, 8.472935, 7.086675, 8.556673, 9.324328, 
    12.48832, 11.6236, 10.23409, 7.944249, 22.04226, 23.37843, 11.00023, 
    2.64938, 3.474224, 14.27784, 10.0872, 20.85916, 7.595808, 9.395947, 
    21.70179, 2.834043, 21.90183, 2.860404, 5.128787, 3.225574, 3.265324, 
    3.422497,
  1.163998, 0.9130338, 3.19914, 0.838528, 0.8111365, 1.519564, 8.09005, 
    8.069554, 7.69157, 7.666807, 4.734021, 3.102786, 7.372371, 9.536769, 
    9.320639, 4.321461, 8.188543, 8.316654, 8.225592, 7.114708, 7.544911, 
    8.623745, 7.853431, 7.846618, 1.144613, 7.947784, 8.019742, 8.051539, 
    1.044186,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0 ;

 average_DT = 730 ;

 average_T1 = 320 ;

 average_T2 = 1050 ;

 climatology_bounds =
  320, 1050 ;

 lat = -89.5, -79.5, -69.5, -59.5, -49.5, -39.5, -29.5, -19.5, -9.5, 0.5, 
    10.5, 20.5, 30.5, 40.5, 50.5, 60.5, 70.5, 80.5 ;

 lat_bnds =
  -90, -89,
  -80, -79,
  -70, -69,
  -60, -59,
  -50, -49,
  -40, -39,
  -30, -29,
  -20, -19,
  -10, -9,
  0, 1,
  10, 11,
  20, 21,
  30, 31,
  40, 41,
  50, 51,
  60, 61,
  70, 71,
  80, 81 ;

 lon = 0.625, 13.125, 25.625, 38.125, 50.625, 63.125, 75.625, 88.125, 
    100.625, 113.125, 125.625, 138.125, 150.625, 163.125, 175.625, 188.125, 
    200.625, 213.125, 225.625, 238.125, 250.625, 263.125, 275.625, 288.125, 
    300.625, 313.125, 325.625, 338.125, 350.625 ;

 lon_bnds =
  0, 1.25,
  12.5, 13.75,
  25, 26.25,
  37.5, 38.75,
  50, 51.25,
  62.5, 63.75,
  75, 76.25,
  87.5, 88.75,
  100, 101.25,
  112.5, 113.75,
  125, 126.25,
  137.5, 138.75,
  150, 151.25,
  162.5, 163.75,
  175, 176.25,
  187.5, 188.75,
  200, 201.25,
  212.5, 213.75,
  225, 226.25,
  237.5, 238.75,
  250, 251.25,
  262.5, 263.75,
  275, 276.25,
  287.5, 288.75,
  300, 301.25,
  312.5, 313.75,
  325, 326.25,
  337.5, 338.75,
  350, 351.25 ;

 time = 0 ;
}
