netcdf \00010101.ocean_static {
dimensions:
	yq = 15 ;
	xq = 15 ;
	yh = 10 ;
	xh = 15 ;
	time = UNLIMITED ; // (1 currently)
variables:
	float Coriolis(yq, xq) ;
		Coriolis:_FillValue = 1.e+20f ;
		Coriolis:missing_value = 1.e+20f ;
		Coriolis:units = "s-1" ;
		Coriolis:long_name = "Coriolis parameter at corner (Bu) points" ;
		Coriolis:cell_methods = "time: point" ;
		Coriolis:interp_method = "none" ;
	float areacello(yh, xh) ;
		areacello:_FillValue = 1.e+20f ;
		areacello:missing_value = 1.e+20f ;
		areacello:units = "m2" ;
		areacello:long_name = "Ocean Grid-Cell Area" ;
		areacello:cell_methods = "area:sum yh:sum xh:sum time: point" ;
		areacello:standard_name = "cell_area" ;
	float areacello_bu(yq, xq) ;
		areacello_bu:_FillValue = 1.e+20f ;
		areacello_bu:missing_value = 1.e+20f ;
		areacello_bu:units = "m2" ;
		areacello_bu:long_name = "Ocean Grid-Cell Area" ;
		areacello_bu:cell_methods = "area:sum yq:sum xq:sum time: point" ;
		areacello_bu:standard_name = "cell_area" ;
	float areacello_cu(yh, xq) ;
		areacello_cu:_FillValue = 1.e+20f ;
		areacello_cu:missing_value = 1.e+20f ;
		areacello_cu:units = "m2" ;
		areacello_cu:long_name = "Ocean Grid-Cell Area" ;
		areacello_cu:cell_methods = "area:sum yh:sum xq:sum time: point" ;
		areacello_cu:standard_name = "cell_area" ;
	float areacello_cv(yq, xh) ;
		areacello_cv:_FillValue = 1.e+20f ;
		areacello_cv:missing_value = 1.e+20f ;
		areacello_cv:units = "m2" ;
		areacello_cv:long_name = "Ocean Grid-Cell Area" ;
		areacello_cv:cell_methods = "area:sum yq:sum xh:sum time: point" ;
		areacello_cv:standard_name = "cell_area" ;
	float deptho(yh, xh) ;
		deptho:_FillValue = 1.e+20f ;
		deptho:missing_value = 1.e+20f ;
		deptho:units = "m" ;
		deptho:long_name = "Sea Floor Depth" ;
		deptho:cell_methods = "area:mean yh:mean xh:mean time: point" ;
		deptho:cell_measures = "area: areacello" ;
		deptho:standard_name = "sea_floor_depth_below_geoid" ;
	float dxCu(yh, xq) ;
		dxCu:_FillValue = 1.e+20f ;
		dxCu:missing_value = 1.e+20f ;
		dxCu:units = "m" ;
		dxCu:long_name = "Delta(x) at u points (meter)" ;
		dxCu:cell_methods = "time: point" ;
		dxCu:interp_method = "none" ;
	float dxCv(yq, xh) ;
		dxCv:_FillValue = 1.e+20f ;
		dxCv:missing_value = 1.e+20f ;
		dxCv:units = "m" ;
		dxCv:long_name = "Delta(x) at v points (meter)" ;
		dxCv:cell_methods = "time: point" ;
		dxCv:interp_method = "none" ;
	float dxt(yh, xh) ;
		dxt:_FillValue = 1.e+20f ;
		dxt:missing_value = 1.e+20f ;
		dxt:units = "m" ;
		dxt:long_name = "Delta(x) at thickness/tracer points (meter)" ;
		dxt:cell_methods = "time: point" ;
		dxt:interp_method = "none" ;
	float dyCu(yh, xq) ;
		dyCu:_FillValue = 1.e+20f ;
		dyCu:missing_value = 1.e+20f ;
		dyCu:units = "m" ;
		dyCu:long_name = "Delta(y) at u points (meter)" ;
		dyCu:cell_methods = "time: point" ;
		dyCu:interp_method = "none" ;
	float dyCv(yq, xh) ;
		dyCv:_FillValue = 1.e+20f ;
		dyCv:missing_value = 1.e+20f ;
		dyCv:units = "m" ;
		dyCv:long_name = "Delta(y) at v points (meter)" ;
		dyCv:cell_methods = "time: point" ;
		dyCv:interp_method = "none" ;
	float dyt(yh, xh) ;
		dyt:_FillValue = 1.e+20f ;
		dyt:missing_value = 1.e+20f ;
		dyt:units = "m" ;
		dyt:long_name = "Delta(y) at thickness/tracer points (meter)" ;
		dyt:cell_methods = "time: point" ;
		dyt:interp_method = "none" ;
	float geolat(yh, xh) ;
		geolat:_FillValue = 1.e+20f ;
		geolat:missing_value = 1.e+20f ;
		geolat:units = "degrees_north" ;
		geolat:long_name = "Latitude of tracer (T) points" ;
		geolat:cell_methods = "time: point" ;
	float geolat_c(yq, xq) ;
		geolat_c:_FillValue = 1.e+20f ;
		geolat_c:missing_value = 1.e+20f ;
		geolat_c:units = "degrees_north" ;
		geolat_c:long_name = "Latitude of corner (Bu) points" ;
		geolat_c:cell_methods = "time: point" ;
		geolat_c:interp_method = "none" ;
	float geolat_u(yh, xq) ;
		geolat_u:_FillValue = 1.e+20f ;
		geolat_u:missing_value = 1.e+20f ;
		geolat_u:units = "degrees_north" ;
		geolat_u:long_name = "Latitude of zonal velocity (Cu) points" ;
		geolat_u:cell_methods = "time: point" ;
		geolat_u:interp_method = "none" ;
	float geolat_v(yq, xh) ;
		geolat_v:_FillValue = 1.e+20f ;
		geolat_v:missing_value = 1.e+20f ;
		geolat_v:units = "degrees_north" ;
		geolat_v:long_name = "Latitude of meridional velocity (Cv) points" ;
		geolat_v:cell_methods = "time: point" ;
		geolat_v:interp_method = "none" ;
	float geolon(yh, xh) ;
		geolon:_FillValue = 1.e+20f ;
		geolon:missing_value = 1.e+20f ;
		geolon:units = "degrees_east" ;
		geolon:long_name = "Longitude of tracer (T) points" ;
		geolon:cell_methods = "time: point" ;
	float geolon_c(yq, xq) ;
		geolon_c:_FillValue = 1.e+20f ;
		geolon_c:missing_value = 1.e+20f ;
		geolon_c:units = "degrees_east" ;
		geolon_c:long_name = "Longitude of corner (Bu) points" ;
		geolon_c:cell_methods = "time: point" ;
		geolon_c:interp_method = "none" ;
	float geolon_u(yh, xq) ;
		geolon_u:_FillValue = 1.e+20f ;
		geolon_u:missing_value = 1.e+20f ;
		geolon_u:units = "degrees_east" ;
		geolon_u:long_name = "Longitude of zonal velocity (Cu) points" ;
		geolon_u:cell_methods = "time: point" ;
		geolon_u:interp_method = "none" ;
	float geolon_v(yq, xh) ;
		geolon_v:_FillValue = 1.e+20f ;
		geolon_v:missing_value = 1.e+20f ;
		geolon_v:units = "degrees_east" ;
		geolon_v:long_name = "Longitude of meridional velocity (Cv) points" ;
		geolon_v:cell_methods = "time: point" ;
		geolon_v:interp_method = "none" ;
	float hfgeou(yh, xh) ;
		hfgeou:_FillValue = 1.e+20f ;
		hfgeou:missing_value = 1.e+20f ;
		hfgeou:units = "W m-2" ;
		hfgeou:long_name = "Upward geothermal heat flux at sea floor" ;
		hfgeou:cell_methods = "area:mean yh:mean xh:mean time: point" ;
		hfgeou:standard_name = "upward_geothermal_heat_flux_at_sea_floor" ;
	float sftof(yh, xh) ;
		sftof:_FillValue = 1.e+20f ;
		sftof:missing_value = 1.e+20f ;
		sftof:units = "%" ;
		sftof:long_name = "Sea Area Fraction" ;
		sftof:cell_methods = "area:mean yh:mean xh:mean time: point" ;
		sftof:standard_name = "SeaAreaFraction" ;
	double time(time) ;
		time:units = "days since 0001-01-01 00:00:00" ;
		time:long_name = "time" ;
		time:axis = "T" ;
		time:calendar_type = "NOLEAP" ;
		time:calendar = "noleap" ;
	float wet(yh, xh) ;
		wet:_FillValue = 1.e+20f ;
		wet:missing_value = 1.e+20f ;
		wet:long_name = "0 if land, 1 if ocean at tracer points" ;
		wet:cell_methods = "time: point" ;
		wet:cell_measures = "area: areacello" ;
	float wet_c(yq, xq) ;
		wet_c:_FillValue = 1.e+20f ;
		wet_c:missing_value = 1.e+20f ;
		wet_c:long_name = "0 if land, 1 if ocean at corner (Bu) points" ;
		wet_c:cell_methods = "time: point" ;
		wet_c:interp_method = "none" ;
	float wet_u(yh, xq) ;
		wet_u:_FillValue = 1.e+20f ;
		wet_u:missing_value = 1.e+20f ;
		wet_u:long_name = "0 if land, 1 if ocean at zonal velocity (Cu) points" ;
		wet_u:cell_methods = "time: point" ;
		wet_u:interp_method = "none" ;
	float wet_v(yq, xh) ;
		wet_v:_FillValue = 1.e+20f ;
		wet_v:missing_value = 1.e+20f ;
		wet_v:long_name = "0 if land, 1 if ocean at meridional velocity (Cv) points" ;
		wet_v:cell_methods = "time: point" ;
		wet_v:interp_method = "none" ;
	double xh(xh) ;
		xh:units = "degrees_east" ;
		xh:long_name = "h point nominal longitude" ;
		xh:axis = "X" ;
	double xq(xq) ;
		xq:units = "degrees_east" ;
		xq:long_name = "q point nominal longitude" ;
		xq:axis = "X" ;
	double yh(yh) ;
		yh:units = "degrees_north" ;
		yh:long_name = "h point nominal latitude" ;
		yh:axis = "Y" ;
	double yq(yq) ;
		yq:units = "degrees_north" ;
		yq:long_name = "q point nominal latitude" ;
		yq:axis = "Y" ;

// global attributes:
		:title = "cm5_c96_am5f7c1r0_b06_piC_galb_noiceinit_alb" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
		:history = "Tue May 27 16:22:52 2025: ncks -d xh,0,14 -d yh,0,9 -d xq,0,14 -d yq,0,14 /home/cew/Code/cmip7-sprint/testfiles/input/00010101.ocean_static.nc -O /home/cew/Code/cmip7-sprint/testfiles/00010101.ocean_static.nc" ;
		:NCO = "netCDF Operators version 5.1.9 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco, Citation = 10.1016/j.envsoft.2008.03.004)" ;
data:

 Coriolis =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 areacello =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 areacello_bu =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 areacello_cu =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 areacello_cv =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 deptho =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 dxCu =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 dxCv =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 dxt =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 dyCu =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 dyCv =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 dyt =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 geolat =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 geolat_c =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 geolat_u =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 geolat_v =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 geolon =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 geolon_c =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 geolon_u =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 geolon_v =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 hfgeou =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 sftof =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 time = 0 ;

 wet =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 wet_c =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 wet_u =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 wet_v =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 xh = -299.875, -299.625, -299.375, -299.125, -298.875, -298.625, -298.375, 
    -298.125, -297.875, -297.625, -297.375, -297.125, -296.875, -296.625, 
    -296.375 ;

 xq = -300, -299.75, -299.5, -299.25, -299, -298.75, -298.5, -298.25, -298, 
    -297.75, -297.5, -297.25, -297, -296.75, -296.5 ;

 yh = -88.5208813286133, -88.4226439858398, -88.3244066430664, 
    -88.2261693002929, -88.1279319575195, -88.029694614746, 
    -87.9314572719726, -87.8332199291991, -87.7349825864257, -87.6367452436523 ;

 yq = -88.57, -88.4717626572265, -88.3735253144531, -88.2752879716797, 
    -88.1770506289062, -88.0788132861328, -87.9805759433593, 
    -87.8823386005859, -87.7841012578124, -87.685863915039, 
    -87.5876265722655, -87.4893892294921, -87.3911518867186, 
    -87.2929145439452, -87.1946772011717 ;
}
