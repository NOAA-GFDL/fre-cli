netcdf atmos_month.198101-198112.alb_sfc {
dimensions:
	time = UNLIMITED ; // (12 currently)
	lat = 18 ;
	lon = 29 ;
	bnds = 2 ;
variables:
	float alb_sfc(time, lat, lon) ;
		alb_sfc:long_name = "Surface Albedo for  Flux" ;
		alb_sfc:units = "percent" ;
		alb_sfc:_FillValue = 1.e+20f ;
		alb_sfc:missing_value = 1.e+20f ;
		alb_sfc:cell_methods = "time: mean" ;
		alb_sfc:cell_measures = "area: area" ;
		alb_sfc:interp_method = "conserve_order1" ;
	double lat(lat) ;
		lat:standard_name = "latitude" ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_N" ;
		lat:axis = "Y" ;
		lat:bounds = "lat_bnds" ;
	double lat_bnds(lat, bnds) ;
	double lon(lon) ;
		lon:standard_name = "longitude" ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_E" ;
		lon:axis = "X" ;
		lon:bounds = "lon_bnds" ;
	double lon_bnds(lon, bnds) ;
	double time(time) ;
		time:standard_name = "time" ;
		time:long_name = "time" ;
		time:bounds = "time_bnds" ;
		time:units = "days since 1979-01-01 00:00:00" ;
		time:calendar = "standard" ;
		time:axis = "T" ;
	double time_bnds(time, bnds) ;

// global attributes:
		:CDI = "Climate Data Interface version 2.4.4 (https://mpimet.mpg.de/cdi)" ;
		:Conventions = "CF-1.6" ;
		:title = "c96L65_am5f9d8r0_amip" ;
		:associated_files = "area: 19810101.grid_spec.nc" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
		:code_release_version = "2024.05" ;
		:git_hash = "5d306c05d9fe755cab04eedc8fd3de0d3c8355a0" ;
		:creationtime = "Mon Aug 11 19:59:00 2025" ;
		:hostname = "pp030" ;
		:history = "Mon Aug 11 16:16:23 2025: ncks -d lat,,,10 -d lon,,,10 atmos_month.198101-198112.alb_sfc.nc reduced/atmos_month.198101-198112.alb_sfc.nc\n",
			"Mon Aug 11 20:01:59 2025: cdo --history splitname 19810101.atmos_month.nc /home/Chris.Blanton/cylc-run/c96L65_am5f9d8r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run1/share/cycle/19810101T0000Z/split/regrid-xy/180_288.conserve_order2/19810101.atmos_month.\n",
			"fregrid --debug --standard_dimension --input_mosaic C96_mosaic.nc --input_dir /home/Chris.Blanton/cylc-run/c96L65_am5f9d8r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run1/share/cycle/19810101T0000Z/history/native --input_file 19810101.atmos_month --associated_file_dir /home/Chris.Blanton/cylc-run/c96L65_am5f9d8r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run1/share/cycle/19810101T0000Z/history/native --interp_method conserve_order2 --remap_file fregrid_remap_file_288_by_180.nc --nlon 288 --nlat 180 --scalar_field (**please see the field list in this file**) --output_file 19810101.atmos_month.nc" ;
		:CDO = "Climate Data Operators version 2.4.4 (https://mpimet.mpg.de/cdo)" ;
		:NCO = "netCDF Operators version 5.2.4 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco, Citation = 10.1016/j.envsoft.2008.03.004)" ;
data:

 alb_sfc =
  76.25285, 76.25285, 76.25285, 76.25285, 76.25285, 76.25285, 76.25285, 
    76.25897, 76.25897, 76.25897, 76.25897, 76.25897, 76.25897, 76.25897, 
    76.24693, 76.24693, 76.24693, 76.24693, 76.24693, 76.24693, 76.24693, 
    76.27441, 76.27441, 76.27441, 76.27441, 76.27441, 76.27441, 76.27441, 
    76.25285,
  76.44437, 76.19061, 76.10728, 76.03162, 76.02551, 76.04452, 76.02316, 
    76.02529, 76.07803, 76.17192, 76.2251, 76.33382, 76.38404, 76.72162, 
    77.61076, 74.43082, 76.99693, 72.19584, 67.54581, 73.11387, 75.10155, 
    76.1926, 74.58293, 68.24023, 75.52526, 66.1054, 74.86777, 69.23141, 
    76.51962,
  28.50309, 24.33908, 50.42044, 64.34027, 72.01418, 72.00896, 47.81725, 
    72.62207, 72.56776, 71.69529, 72.38673, 72.76912, 67.12334, 60.87822, 
    6.322688, 5.9809, 6.582986, 6.815576, 6.37846, 21.82946, 9.001003, 
    18.95372, 56.81915, 60.97662, 61.21234, 13.32665, 6.244976, 6.660918, 
    7.287549,
  4.62552, 4.729858, 4.944829, 4.697002, 4.679885, 4.614884, 4.769694, 
    4.555934, 4.72069, 4.641797, 4.762366, 4.648767, 4.550398, 4.819422, 
    4.937311, 4.889597, 4.622276, 4.741107, 4.810156, 5.127718, 5.094404, 
    5.162316, 5.103305, 5.040258, 4.68521, 4.503845, 4.626632, 4.79687, 
    4.605134,
  4.186664, 4.317166, 4.253982, 4.457397, 4.329167, 4.314857, 4.309872, 
    4.192106, 4.188114, 4.281168, 4.51259, 4.353054, 4.375732, 4.524392, 
    4.42281, 4.22637, 4.194461, 4.34935, 4.364345, 4.467135, 4.447765, 
    4.480952, 4.397642, 8.589765, 4.88754, 4.370362, 4.252131, 4.175511, 
    4.238363,
  4.030228, 4.017932, 4.396855, 4.220715, 4.090051, 4.037546, 4.015064, 
    3.891837, 3.850593, 4.004006, 3.979544, 4.26432, 4.157741, 3.916245, 
    10.10682, 3.979578, 4.139743, 4.018028, 3.941245, 3.824202, 3.923378, 
    4.00177, 4.018346, 10.01776, 4.546876, 4.170698, 3.920205, 3.899943, 
    3.910404,
  3.973957, 3.976381, 12.54141, 3.895043, 4.089889, 3.898044, 3.797119, 
    3.967796, 3.762332, 4.120789, 10.42475, 16.04226, 10.42725, 3.939613, 
    4.165726, 3.877569, 3.917168, 3.781408, 3.631483, 3.949666, 4.072561, 
    4.175301, 3.837363, 4.599521, 9.660911, 3.805533, 3.69835, 3.956614, 
    3.988466,
  3.638758, 10.09365, 12.24548, 3.55879, 3.49978, 3.341087, 3.606533, 
    3.587746, 3.66411, 3.468076, 12.20152, 11.09819, 3.551778, 3.6474, 
    3.614573, 3.596542, 3.366595, 3.623096, 3.68731, 4.076787, 3.956673, 
    3.828458, 3.366333, 3.301217, 9.224553, 9.545017, 3.955695, 3.992986, 
    4.019764,
  3.448313, 6.498559, 8.795625, 9.331126, 3.299385, 3.375395, 3.537181, 
    3.47185, 3.588164, 3.24944, 4.617576, 3.271331, 4.36395, 3.393754, 
    3.40133, 3.621265, 3.463986, 3.7496, 3.578741, 3.973477, 3.621236, 
    3.674351, 3.449006, 8.752406, 8.622976, 8.862894, 3.84174, 3.603243, 
    3.67109,
  3.212863, 8.847048, 8.667336, 9.959523, 3.4798, 3.344474, 3.176226, 
    3.269013, 8.738402, 8.242429, 3.20764, 3.217577, 3.184929, 3.335654, 
    3.49186, 3.725949, 3.737191, 3.901747, 3.829139, 3.990755, 3.646087, 
    3.363367, 3.362743, 8.482767, 8.490137, 3.138422, 3.359119, 3.466349, 
    3.170737,
  10.1605, 10.20571, 10.58627, 9.518259, 14.22514, 3.411071, 5.477973, 
    3.591974, 3.489619, 3.599905, 4.178845, 3.321407, 3.33167, 3.600458, 
    3.636446, 3.574635, 3.823971, 3.534467, 3.801881, 3.497605, 3.551521, 
    3.620317, 8.583489, 7.248289, 3.535151, 3.625779, 3.302197, 3.64899, 
    9.00752,
  16.19405, 18.68271, 20.70156, 3.654742, 20.67924, 4.112761, 10.10409, 
    4.042687, 9.035423, 3.249509, 3.692606, 3.787453, 3.69267, 4.116786, 
    4.045927, 3.724722, 3.861744, 3.821295, 3.776413, 3.398991, 3.935206, 
    6.209273, 3.900632, 4.669007, 3.829282, 4.02164, 3.573931, 3.562109, 
    21.1219,
  20.53044, 16.34159, 17.11703, 16.58839, 11.25486, 12.74166, 12.41082, 
    21.42238, 11.88453, 10.45427, 3.453351, 3.576255, 3.993596, 3.838589, 
    3.789434, 3.847592, 3.853415, 3.629769, 3.937521, 4.005362, 9.518476, 
    11.08754, 9.671306, 3.517058, 4.017105, 3.898309, 3.800087, 4.08324, 
    9.876928,
  5.734525, 4.369344, 5.639949, 21.29601, 1.619299, 12.19106, 20.12887, 
    15.48073, 10.39243, 24.40797, 12.21084, 3.67704, 4.066605, 4.122468, 
    3.867066, 3.775214, 3.357579, 3.497929, 3.588675, 13.28588, 28.14277, 
    23.84485, 16.60576, 4.959707, 3.574054, 3.478571, 3.573528, 3.429143, 
    4.788535,
  4.305625, 13.1902, 16.90124, 21.3148, 25.39365, 26.22113, 14.24677, 
    25.07507, 12.0619, 6.294494, 5.517313, 19.02976, 3.690831, 4.284812, 
    3.494217, 3.357742, 3.040316, 3.186808, 3.57993, 15.95235, 15.42676, 
    22.88089, 18.80218, 22.60502, 6.709063, 3.649329, 4.217072, 3.713891, 
    3.390046,
  3.079972, 15.78787, 10.24107, 14.76607, 13.05266, 14.36469, 13.92672, 
    15.51315, 13.11488, 13.60625, 10.80467, 20.16291, 21.60268, 17.35262, 
    2.253484, 20.5484, 17.69775, 9.012324, 20.81408, 12.31257, 14.79779, 
    21.6341, 26.01353, 22.05828, 2.126907, 5.843377, 3.076459, 3.15899, 
    3.165395,
  0.2413161, 0.2188116, 1.978713, 0.2684774, 0.9168655, 3.137789, 2.81116, 
    2.770568, 2.58713, 2.514809, 1.782062, 1.440114, 2.58055, 3.285434, 
    3.192125, 3.514523, 2.955585, 3.285028, 3.393564, 3.490463, 2.886969, 
    3.258077, 3.040147, 3.001601, 3.180703, 2.797944, 2.839205, 3.350022, 
    0.2942657,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  76.47349, 76.47349, 76.47349, 76.47349, 76.47349, 76.47349, 76.47349, 
    76.46885, 76.46885, 76.46885, 76.46885, 76.46885, 76.46885, 76.46885, 
    76.46272, 76.46272, 76.46272, 76.46272, 76.46272, 76.46272, 76.46272, 
    76.51137, 76.51137, 76.51137, 76.51137, 76.51137, 76.51137, 76.51137, 
    76.47349,
  73.38937, 73.0288, 72.95197, 73.06375, 72.88479, 72.92987, 72.85201, 
    72.84698, 73.00648, 72.99537, 72.78703, 73.31318, 73.35129, 73.63771, 
    74.05005, 73.25165, 74.23699, 72.93342, 73.60738, 73.87808, 74.08434, 
    74.27706, 74.08244, 73.94949, 74.34531, 71.2145, 73.02779, 73.33174, 
    73.55668,
  23.68905, 19.22613, 7.555005, 45.89272, 55.90423, 55.29077, 46.16449, 
    55.35531, 55.35733, 55.78025, 55.45878, 55.49192, 55.65055, 30.94169, 
    5.616188, 5.393435, 5.653991, 5.101903, 5.123664, 5.076049, 5.43658, 
    11.23932, 43.55555, 47.11147, 46.63531, 5.308214, 5.236366, 5.124593, 
    5.305081,
  4.542045, 4.202247, 4.455595, 4.116914, 4.055612, 4.002218, 4.12833, 
    4.592474, 4.614058, 4.669598, 4.800887, 4.390934, 4.320484, 4.384887, 
    4.566933, 4.485081, 4.287245, 4.233551, 4.612134, 4.628309, 4.59808, 
    4.808796, 4.484952, 4.345573, 4.137033, 4.078397, 4.145028, 4.41147, 
    4.253036,
  4.045811, 3.981613, 4.024312, 4.009115, 4.011377, 4.066682, 3.895648, 
    4.082625, 4.103643, 4.164188, 4.197336, 4.229297, 4.166733, 4.168899, 
    4.027658, 3.926782, 4.091369, 3.929942, 4.227895, 4.137807, 4.257522, 
    4.004555, 4.095086, 7.86202, 4.548726, 4.069358, 3.997149, 4.021692, 
    3.785915,
  3.824169, 3.946234, 4.002593, 3.928079, 3.735591, 3.73566, 3.712724, 
    3.502936, 3.595342, 3.816068, 3.997175, 4.019819, 4.038631, 3.992, 
    9.304639, 3.574995, 3.901952, 3.701087, 3.848388, 3.885811, 3.810099, 
    3.891664, 3.72386, 9.538174, 4.321431, 3.845592, 3.672635, 3.87425, 
    3.849491,
  3.933947, 4.205045, 11.94157, 3.856716, 3.725211, 3.463316, 3.893256, 
    3.725722, 3.905588, 4.059326, 9.689536, 14.59482, 10.31497, 3.897257, 
    3.577773, 3.635252, 3.524714, 3.62618, 3.585831, 3.8431, 3.7784, 4.01124, 
    3.769807, 4.16202, 9.40954, 3.434255, 3.887748, 3.788271, 4.119768,
  3.42633, 9.744349, 12.25169, 3.670028, 3.270532, 3.634238, 3.811703, 
    3.593475, 3.703417, 3.275148, 11.84588, 11.33382, 3.803502, 3.558307, 
    3.331904, 3.486379, 3.371178, 3.683268, 3.462898, 3.813497, 3.804553, 
    3.708179, 3.438823, 3.534403, 8.973072, 8.768469, 3.763811, 3.569672, 
    3.914507,
  3.296974, 6.313697, 8.427731, 9.145274, 3.414996, 3.396683, 3.677496, 
    3.552946, 3.39261, 3.304254, 4.592828, 3.127028, 4.335747, 3.13157, 
    3.031756, 3.449894, 3.431673, 3.556704, 3.547427, 3.836514, 3.562861, 
    3.809493, 3.479173, 8.358654, 8.393641, 8.737321, 3.504572, 3.469503, 
    3.659154,
  3.092581, 8.687326, 8.511052, 9.861168, 3.285424, 3.127158, 3.247306, 
    3.229949, 8.669594, 8.481945, 3.200342, 3.282953, 3.236895, 3.137813, 
    3.266041, 3.530599, 3.602223, 3.779, 3.65051, 3.740967, 3.578296, 
    3.396876, 3.357579, 8.693338, 8.441473, 3.134681, 3.160415, 3.264361, 
    3.057022,
  9.951073, 10.1648, 10.8296, 9.336568, 14.27404, 3.517084, 5.359812, 
    3.615214, 3.757757, 3.378586, 3.911884, 3.403492, 3.241949, 3.403089, 
    3.607373, 3.423151, 3.610794, 3.44924, 3.330248, 3.212582, 3.408447, 
    3.431586, 8.548915, 7.690048, 3.409532, 3.553764, 3.212499, 3.31555, 
    9.025295,
  17.17299, 19.24684, 20.98844, 3.770304, 21.16425, 3.788384, 10.67969, 
    4.14293, 9.152899, 3.380504, 3.226138, 3.577653, 3.761951, 3.754867, 
    3.67754, 3.792931, 3.961147, 3.502704, 3.679859, 3.298177, 3.745206, 
    6.274539, 3.788821, 4.496214, 3.924277, 4.031633, 3.573115, 3.894007, 
    21.86384,
  21.32451, 16.6807, 17.80998, 17.25264, 11.82918, 13.47122, 12.33112, 
    19.7534, 10.94252, 11.02758, 3.219759, 3.544452, 3.796863, 3.76445, 
    3.716333, 3.322585, 3.721414, 3.350798, 3.643692, 4.139328, 11.99729, 
    12.45723, 12.11444, 3.391979, 3.586865, 3.630364, 3.606144, 3.466739, 
    10.11079,
  5.441322, 4.263473, 6.195023, 16.24177, 1.745014, 12.59807, 25.24848, 
    13.49161, 11.4486, 23.89228, 10.09495, 3.706543, 3.658422, 4.004444, 
    3.904898, 3.7628, 3.393523, 3.429749, 3.868484, 11.55112, 31.38688, 
    20.96553, 24.33289, 4.92922, 3.399285, 3.390161, 3.588398, 3.799552, 
    4.801128,
  4.930236, 13.34633, 13.83937, 27.03154, 29.84692, 31.23927, 17.26562, 
    29.58057, 14.12615, 6.566063, 6.105516, 22.29372, 3.91268, 4.037742, 
    4.179052, 4.434782, 3.702923, 3.429086, 3.570111, 21.59432, 18.39, 
    27.40141, 23.28908, 27.86168, 10.42874, 3.681109, 3.85862, 3.831404, 
    3.484537,
  3.447603, 21.83692, 16.81063, 21.95956, 20.8015, 20.77264, 21.03954, 
    22.70031, 19.15129, 19.67199, 16.16232, 27.71015, 29.27386, 25.9633, 
    3.293368, 32.77077, 25.36459, 12.48012, 28.4809, 18.40113, 20.78348, 
    29.33702, 35.18491, 29.62201, 3.013771, 8.086734, 3.999071, 3.640182, 
    3.499787,
  2.77061, 2.599666, 15.2395, 2.776066, 12.51746, 26.23814, 22.15353, 
    22.19633, 21.89847, 21.8501, 15.19132, 12.38034, 21.76487, 26.25883, 
    26.07509, 26.7859, 23.93197, 23.9042, 25.85169, 26.03227, 21.99245, 
    24.62457, 22.72041, 22.6867, 26.74351, 22.75857, 22.73637, 25.10599, 
    2.971133,
  2.347429, 2.28148, 2.50774, 2.489999, 2.331524, 2.116885, 2.359385, 
    2.386973, 2.347938, 2.132972, 2.142857, 2.117281, 2.199756, 2.476933, 
    2.378642, 2.319304, 2.491861, 2.707309, 2.880671, 2.679748, 2.725112, 
    2.544869, 2.257616, 2.48093, 2.15655, 2.199329, 2.057053, 2.09281, 
    2.556672,
  47.86325, 47.86325, 47.86325, 47.86325, 47.86325, 47.86325, 47.86325, 
    47.9864, 47.9864, 47.9864, 47.9864, 47.9864, 47.9864, 47.9864, 47.88717, 
    47.88717, 47.88717, 47.88717, 47.88717, 47.88717, 47.88717, 47.66661, 
    47.66661, 47.66661, 47.66661, 47.66661, 47.66661, 47.66661, 47.86325,
  43.60559, 43.56427, 43.51102, 43.64766, 43.46303, 43.40103, 43.36587, 
    43.29021, 43.13161, 43.11645, 43.22464, 43.29139, 43.46806, 43.94561, 
    44.1, 44.53913, 44.12061, 44.00351, 43.80995, 44.3302, 44.47427, 
    44.31205, 44.0598, 44.22716, 44.25876, 44.0233, 43.8876, 43.85018, 
    43.58686,
  19.13547, 15.21168, 8.159559, 35.79597, 42.11032, 42.00614, 44.69871, 
    41.86934, 41.54436, 41.61552, 41.60257, 41.78421, 42.02669, 13.27865, 
    4.428499, 4.379848, 4.495051, 4.303891, 4.467598, 4.404344, 3.975779, 
    8.574464, 22.07154, 38.01693, 44.161, 4.688285, 4.321562, 4.572248, 
    4.775513,
  4.458996, 4.321667, 4.589545, 4.165012, 4.007765, 4.052714, 3.882623, 
    3.753137, 3.896985, 4.261047, 4.618036, 4.308486, 3.777787, 4.034236, 
    4.213739, 4.08694, 3.948004, 3.784545, 4.03844, 4.325053, 4.250377, 
    4.359186, 4.082337, 4.054464, 3.762205, 3.791435, 3.861564, 4.001741, 
    4.528336,
  3.688109, 3.927964, 4.009128, 3.949556, 3.680764, 3.805731, 3.73416, 
    3.78597, 3.841884, 3.908787, 3.856374, 3.935338, 3.766527, 3.774638, 
    3.849305, 3.836555, 3.811591, 3.983771, 4.133485, 4.059247, 4.066262, 
    4.001992, 3.943551, 7.216831, 4.377115, 3.927748, 3.634935, 3.420948, 
    3.663777,
  3.643287, 3.774722, 4.038914, 3.767598, 3.714923, 3.848742, 3.743246, 
    3.550682, 3.674261, 3.747315, 3.797193, 3.859452, 4.05143, 3.555408, 
    8.700632, 3.691863, 3.78288, 3.677866, 3.631777, 3.680036, 3.593408, 
    3.421868, 3.837591, 8.896569, 4.387879, 3.70465, 3.648818, 3.581098, 
    3.746436,
  3.819831, 3.954465, 11.39918, 3.641202, 3.754565, 3.560645, 3.543408, 
    3.637597, 3.584126, 3.886977, 9.559267, 14.14689, 9.789516, 3.876059, 
    3.733354, 3.623034, 3.601084, 3.597252, 3.520065, 3.859849, 3.788543, 
    4.046131, 3.763992, 4.329397, 8.939814, 3.666645, 3.500868, 3.777254, 
    3.999557,
  3.530055, 9.687468, 11.4823, 3.446306, 3.32619, 3.270144, 3.607909, 
    3.478441, 3.648197, 3.657271, 12.18188, 11.2819, 3.561635, 3.522341, 
    3.318063, 3.436456, 3.423648, 3.503818, 3.552208, 3.821551, 3.541161, 
    3.769471, 3.37883, 3.28507, 8.907555, 8.722985, 3.549581, 3.632228, 
    3.882436,
  3.343881, 6.243426, 8.473501, 9.03372, 3.347484, 3.47118, 3.402011, 
    3.261284, 3.32978, 3.26004, 4.741865, 3.386581, 4.161629, 3.175197, 
    3.118029, 3.425899, 3.192819, 3.389931, 3.393841, 3.516606, 3.517272, 
    3.700892, 3.447294, 8.406621, 8.305228, 8.582374, 3.422557, 3.569338, 
    3.580556,
  3.032411, 8.583547, 8.253314, 9.844931, 3.237589, 3.260622, 3.178483, 
    3.311226, 8.484381, 8.004576, 3.33273, 3.186717, 3.201923, 3.209167, 
    3.167309, 3.281495, 3.465244, 3.721592, 3.5209, 3.561671, 3.399062, 
    3.461138, 3.221265, 8.4309, 8.444202, 3.079857, 3.183247, 3.237569, 
    3.055395,
  9.936267, 10.3758, 10.4497, 9.511047, 14.96278, 3.321997, 5.296031, 
    3.519904, 3.699653, 3.437191, 4.403192, 3.434813, 3.307281, 3.445473, 
    3.42362, 3.443806, 3.477342, 3.375141, 3.37443, 3.409642, 3.183667, 
    3.38012, 8.705035, 7.393296, 3.377709, 3.270824, 3.140347, 3.138105, 
    8.938948,
  17.54675, 19.97657, 22.06772, 3.355389, 22.15116, 3.694685, 10.62347, 
    3.727415, 9.631269, 3.247338, 3.469681, 3.588007, 3.587141, 3.71011, 
    3.72732, 3.638066, 3.626317, 3.710674, 3.31276, 3.551157, 3.702705, 
    6.095897, 3.713453, 4.495441, 3.764348, 3.594611, 3.358636, 3.193894, 
    22.81223,
  22.69071, 18.48763, 19.76144, 18.43981, 12.31849, 13.98708, 12.12571, 
    20.77826, 9.783124, 10.23105, 3.43657, 3.526586, 3.561235, 3.492108, 
    3.433186, 3.521192, 3.575243, 3.578695, 3.522346, 3.933529, 12.53056, 
    11.27386, 8.969935, 3.560365, 3.473804, 3.595534, 3.49794, 3.488692, 
    11.10925,
  6.911561, 4.239717, 6.104644, 21.97217, 1.914341, 13.87077, 26.11742, 
    14.23802, 12.24114, 9.978435, 10.09568, 3.71858, 3.702274, 3.762507, 
    3.722198, 3.640781, 3.57287, 3.414088, 3.522391, 12.08503, 28.11846, 
    15.39535, 15.52871, 4.664992, 3.563662, 3.589667, 3.672574, 3.712969, 
    5.711269,
  5.764884, 14.28816, 15.10825, 15.08293, 18.25835, 31.7608, 12.38274, 
    33.24897, 14.07794, 8.719583, 7.598753, 26.03641, 4.230794, 3.920293, 
    3.835678, 3.967264, 3.468098, 3.418922, 3.628094, 21.76154, 15.44891, 
    30.85045, 28.21659, 33.07829, 12.505, 3.736768, 3.75719, 3.866677, 
    3.871763,
  4.258918, 24.43213, 19.03308, 28.24267, 26.65698, 25.58398, 25.1888, 
    27.88618, 24.23011, 25.07871, 21.42915, 36.19353, 37.99911, 34.10403, 
    5.123603, 39.10859, 33.15577, 15.88712, 36.0847, 25.83543, 26.8081, 
    37.6773, 45.43743, 38.32676, 3.606916, 15.28094, 4.68666, 4.615879, 
    4.42591,
  4.64036, 4.496507, 26.49236, 3.753574, 40.07278, 41.52692, 36.99358, 
    37.25118, 37.39013, 37.20338, 26.67743, 21.91695, 36.85708, 43.78579, 
    43.5141, 44.55828, 39.65234, 39.41783, 43.1633, 43.03728, 36.64069, 
    40.92839, 37.88924, 37.70203, 44.70045, 37.8121, 37.62402, 42.34515, 
    4.654528,
  40.45809, 41.46996, 39.06857, 41.36221, 40.28374, 39.8233, 41.39633, 
    41.09312, 41.31589, 41.54827, 41.6129, 41.53643, 41.66534, 41.64058, 
    41.63769, 41.49719, 41.45634, 41.44926, 41.48461, 41.55274, 41.46035, 
    39.10433, 36.1328, 36.97921, 35.14833, 34.9593, 34.98283, 35.66399, 
    41.59682,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  10.2823, 10.3841, 10.42082, 10.13789, 10.49899, 10.3605, 10.49905, 
    10.62477, 10.44701, 10.40105, 10.84681, 10.39646, 10.54596, 10.63387, 
    10.65538, 10.67723, 10.66201, 10.5154, 10.21663, 10.19349, 10.11368, 
    10.2536, 10.01198, 10.12654, 10.01575, 10.64864, 10.71651, 10.67458, 
    10.36253,
  16.68602, 26.36262, 23.26848, 29.56888, 27.71469, 27.61427, 30.32085, 
    27.81997, 27.69191, 27.78355, 27.4902, 27.40155, 27.72713, 27.49432, 
    13.36353, 9.111379, 9.316815, 3.530072, 3.093677, 2.7488, 6.863021, 
    7.774731, 22.34785, 28.59387, 32.22757, 25.79162, 15.73503, 8.648671, 
    10.06623,
  3.657752, 3.762981, 4.065264, 3.864401, 3.860222, 3.563244, 3.574946, 
    3.983171, 3.657056, 3.804006, 4.339695, 3.510604, 3.287935, 3.804054, 
    3.977929, 3.822574, 3.598054, 3.482534, 3.562351, 3.632492, 3.721176, 
    3.586183, 3.285668, 3.858269, 3.046769, 3.513323, 3.148836, 3.524644, 
    3.711871,
  3.435922, 3.297428, 3.481202, 3.655682, 3.570048, 3.480334, 3.770097, 
    3.85387, 3.733075, 3.675462, 3.511822, 3.741722, 3.711176, 3.708241, 
    3.785329, 3.880292, 3.944672, 3.538287, 3.478637, 3.571687, 3.332803, 
    3.471545, 3.701307, 6.419241, 4.149329, 3.649121, 3.777497, 3.710568, 
    3.537232,
  3.769923, 3.652518, 3.892305, 3.680295, 3.69354, 3.748533, 3.699768, 
    3.702356, 3.652145, 3.667692, 3.737045, 3.820895, 4.154766, 4.068425, 
    8.116899, 3.795965, 3.8204, 3.489031, 3.866335, 3.635876, 3.893694, 
    3.865578, 3.786244, 8.09507, 4.115847, 3.898019, 3.892253, 3.956658, 
    3.589979,
  3.903672, 3.811388, 11.33152, 3.631394, 3.722037, 3.840865, 3.592829, 
    3.843861, 3.465478, 4.119938, 9.109232, 13.55053, 9.611348, 4.071254, 
    3.985947, 3.607096, 3.634933, 3.470713, 3.803634, 3.562391, 3.494386, 
    3.842924, 3.840994, 4.245013, 8.624439, 3.975048, 3.561342, 3.840764, 
    3.745887,
  3.515443, 9.56234, 9.826855, 3.550074, 3.469092, 3.639843, 3.545595, 
    3.712024, 3.523921, 3.867049, 12.10823, 11.40595, 3.646642, 3.705272, 
    3.532951, 3.389792, 3.481561, 3.496129, 3.814245, 3.726813, 3.870294, 
    3.713054, 3.421106, 3.506603, 8.734684, 8.953725, 3.737519, 3.958822, 
    3.696936,
  3.271075, 6.538677, 8.858203, 8.635196, 3.456529, 3.339016, 3.17222, 
    3.360709, 3.26179, 3.263445, 4.434933, 3.225948, 4.091791, 3.346676, 
    3.384546, 3.137582, 3.473373, 3.781934, 3.616079, 3.6603, 3.676176, 
    3.520726, 3.280417, 8.591984, 8.225548, 8.841343, 3.842262, 3.523408, 
    3.517268,
  3.050037, 8.405201, 8.133167, 9.779788, 3.46048, 3.43335, 3.511436, 
    3.320469, 8.701575, 8.214864, 3.316143, 3.294436, 3.186212, 3.476882, 
    3.324012, 3.409436, 3.412533, 3.544314, 3.470723, 3.489922, 3.494511, 
    3.487345, 3.249383, 8.048944, 8.290181, 3.309446, 3.136048, 3.23063, 
    3.072796,
  10.09554, 10.34316, 10.413, 9.911973, 14.89494, 3.252333, 5.350966, 
    3.359843, 3.525831, 3.389397, 4.420576, 3.230442, 3.46165, 3.293792, 
    3.222665, 3.297614, 3.253946, 3.260309, 3.341802, 3.434858, 3.294699, 
    3.508016, 8.875221, 7.450827, 3.505873, 3.336764, 3.199981, 3.216482, 
    8.831358,
  18.11437, 20.77784, 22.80289, 3.525267, 22.71027, 3.508467, 10.97071, 
    3.476373, 10.01117, 3.305715, 3.564311, 3.669705, 3.74422, 3.744949, 
    3.735702, 3.865381, 3.531675, 3.745332, 3.327504, 3.541386, 3.728203, 
    6.566255, 3.776703, 4.381808, 3.927527, 3.500829, 3.560474, 3.518139, 
    23.6546,
  24.04209, 20.23202, 20.96905, 19.43071, 12.52403, 14.31042, 12.53258, 
    19.1592, 9.196596, 10.10672, 3.464012, 3.425197, 3.362109, 3.459697, 
    3.582243, 3.509008, 3.480688, 3.856695, 3.510452, 3.883758, 10.43557, 
    11.87629, 9.447504, 3.635334, 3.908524, 3.675807, 3.767608, 3.688599, 
    11.39904,
  7.723964, 4.034106, 5.892714, 10.63053, 2.083908, 15.33471, 14.35986, 
    15.45729, 13.49847, 11.05388, 8.272856, 3.963526, 3.825073, 3.805083, 
    3.705377, 3.618259, 3.650476, 3.825672, 3.694233, 12.2094, 11.59688, 
    14.60992, 13.69412, 4.398408, 3.817233, 3.863486, 3.760123, 3.745281, 
    5.22649,
  5.927563, 12.75562, 15.07015, 16.07172, 13.4171, 13.44447, 8.557118, 
    35.95807, 9.348412, 8.132102, 8.362915, 24.70223, 3.890318, 4.08754, 
    4.177126, 4.466231, 4.019747, 3.973223, 4.11716, 12.20696, 11.56637, 
    18.62702, 22.45228, 34.49789, 9.831541, 3.888309, 3.998572, 4.421502, 
    4.211093,
  4.860225, 15.57729, 15.5633, 26.31043, 21.73938, 16.39543, 19.12786, 
    33.81788, 30.27572, 30.3998, 23.83459, 44.69674, 45.89076, 38.74989, 
    4.384302, 17.46636, 39.101, 18.39072, 41.11026, 15.33483, 19.51368, 
    44.22225, 52.94443, 46.3211, 4.140852, 11.75031, 5.009665, 4.852435, 
    4.723929,
  4.9528, 6.093573, 34.59067, 6.246111, 56.09219, 60.14931, 51.99076, 
    52.06572, 52.17702, 51.59848, 37.50103, 31.75468, 51.68705, 60.98213, 
    60.55804, 62.0252, 55.71251, 55.42488, 60.22522, 59.84231, 51.22786, 
    56.88989, 52.98647, 52.69043, 59.16868, 52.55598, 52.44607, 55.47049, 
    5.370459,
  74.78991, 70.48125, 70.88749, 74.39713, 75.89007, 77.97993, 81.33638, 
    81.22336, 81.46358, 82.073, 82, 81.99393, 81.88242, 81.67651, 81.80884, 
    81.94019, 81.92454, 81.66813, 81.50029, 81.6239, 81.65494, 76.94597, 
    71.53992, 72.72562, 69.36823, 69.05082, 69.29929, 70.80599, 80.0174,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  10.4232, 10.66378, 11.0925, 10.3434, 9.441807, 9.431978, 10.42794, 
    9.478423, 9.675533, 9.697056, 9.604809, 9.410529, 9.430476, 11.1859, 
    10.19321, 7.149058, 10.37973, 8.566884, 5.287404, 9.082601, 9.36251, 
    7.434439, 9.500381, 9.185423, 11.0356, 11.20379, 10.05745, 10.77281, 
    11.00603,
  2.737919, 3.406557, 3.750786, 3.589836, 3.198654, 3.00509, 2.878663, 
    2.963968, 2.976619, 3.261252, 3.099189, 2.901306, 2.918248, 2.6566, 
    2.997812, 2.909362, 2.958345, 3.145292, 3.11168, 3.201442, 3.281427, 
    3.187022, 3.288355, 2.825517, 2.67851, 2.812316, 2.798754, 2.649971, 
    2.722737,
  3.692113, 3.535609, 3.796281, 3.590552, 3.310591, 3.616301, 3.22162, 
    3.454179, 3.501966, 3.501212, 3.509827, 3.224519, 3.397851, 3.305832, 
    3.131092, 3.386782, 3.656504, 3.597195, 3.835471, 3.809779, 3.894062, 
    3.946064, 3.158932, 6.158599, 3.999078, 3.337545, 3.364511, 3.579407, 
    3.570997,
  3.504381, 3.896251, 3.966372, 3.729223, 3.911295, 3.910284, 3.965196, 
    3.76421, 3.665496, 3.900346, 4.115698, 4.09838, 4.184096, 3.799531, 
    7.389039, 3.856648, 3.528082, 3.606489, 3.587971, 3.787832, 3.547339, 
    3.427481, 3.609859, 7.738131, 3.875213, 3.735732, 4.104619, 3.767625, 
    3.744976,
  3.678461, 4.104763, 11.1795, 3.978556, 3.982644, 3.942193, 4.052356, 
    4.005466, 4.006149, 4.267581, 9.154458, 13.212, 9.520465, 4.130663, 
    4.001759, 3.507063, 3.607414, 3.798941, 3.501741, 3.514313, 3.588105, 
    3.872707, 3.854005, 4.320979, 8.395721, 3.947547, 3.997191, 3.942077, 
    3.844327,
  3.761771, 9.390458, 10.87209, 4.004695, 3.874057, 3.763717, 3.767859, 
    4.003623, 3.646869, 4.224083, 11.32798, 11.69181, 3.979162, 3.592889, 
    3.750282, 3.631039, 3.836272, 3.585665, 3.888454, 3.783914, 3.957422, 
    3.922023, 3.531223, 3.849338, 8.656506, 8.6977, 3.545544, 4.203999, 
    3.579089,
  3.534266, 6.343275, 9.039492, 8.915622, 3.498135, 3.445469, 3.448263, 
    3.442595, 3.321507, 3.470936, 4.296668, 3.383607, 4.271377, 3.242501, 
    3.618202, 3.665243, 3.839926, 3.825007, 4.004071, 3.786164, 3.829327, 
    3.516105, 3.20495, 8.656515, 8.555301, 8.757083, 3.849654, 3.797588, 
    3.469767,
  3.24389, 8.3931, 8.137314, 9.757134, 3.441632, 3.209482, 3.287992, 
    3.250447, 8.601323, 8.400973, 3.31124, 3.396881, 3.599487, 3.518656, 
    3.379457, 3.481494, 3.538258, 3.635646, 3.598418, 3.780856, 3.671923, 
    3.768071, 3.148979, 8.283686, 8.49495, 3.41376, 3.491836, 3.417027, 
    3.284626,
  9.912714, 10.46082, 10.72436, 9.949521, 15.34627, 3.313577, 5.155846, 
    3.17882, 3.488288, 3.18223, 4.220709, 3.188723, 3.340144, 3.31947, 
    3.374011, 3.378586, 3.314257, 3.571228, 3.398951, 3.578348, 3.333654, 
    3.232614, 9.011678, 7.399442, 3.553965, 3.302969, 3.290559, 3.15291, 
    9.018363,
  18.82865, 21.61217, 23.64423, 3.49488, 23.96092, 3.624819, 11.23171, 
    3.327998, 9.419011, 3.372988, 3.72691, 3.702123, 3.575365, 3.650487, 
    3.726664, 3.757225, 3.605601, 3.786683, 3.386598, 3.842465, 3.97668, 
    6.749997, 3.604721, 4.039994, 3.563851, 3.482942, 3.77642, 3.647016, 
    24.58926,
  25.31614, 21.34241, 22.21624, 20.46692, 13.40833, 15.26431, 13.26155, 
    17.68552, 9.975374, 10.76912, 3.659368, 3.55358, 3.543811, 3.74603, 
    3.778268, 3.653555, 3.807941, 3.772186, 3.774717, 3.978642, 11.24806, 
    12.2783, 9.959605, 3.77776, 3.715867, 3.742874, 3.716936, 3.735712, 
    11.79764,
  8.313829, 3.980488, 6.46824, 10.84984, 2.252835, 15.93054, 10.24387, 
    16.6604, 14.39943, 11.69016, 8.180788, 4.111171, 3.959324, 3.811295, 
    3.740052, 3.775197, 3.866387, 3.785929, 3.736854, 13.03179, 12.09779, 
    14.78621, 13.92286, 4.844381, 3.908955, 3.903589, 4.013534, 4.317868, 
    5.245015,
  6.443024, 13.54856, 15.23941, 15.88912, 14.73211, 13.06655, 9.178881, 
    23.77223, 9.979302, 8.4163, 8.148265, 9.034524, 4.282784, 4.389501, 
    4.101119, 4.113883, 4.158012, 4.367456, 4.35952, 10.24662, 11.74794, 
    10.97176, 7.646235, 14.66767, 5.57172, 3.979575, 4.288142, 4.396487, 
    4.41933,
  5.443273, 9.223376, 10.98321, 8.944587, 10.14637, 10.25516, 9.081723, 
    17.20312, 12.542, 12.19896, 9.38532, 39.78866, 48.25568, 31.72913, 
    4.913126, 5.612537, 23.25904, 20.9513, 36.81985, 8.656455, 8.792933, 
    37.55586, 47.29005, 38.68701, 4.713165, 10.18047, 4.514663, 4.644034, 
    5.17561,
  6.397051, 7.638515, 41.04818, 6.892959, 66.37019, 72.70956, 65.02373, 
    65.62538, 65.86261, 65.21964, 42.63134, 32.73222, 64.29359, 68.53593, 
    66.77146, 67.87492, 64.37669, 59.94524, 66.35417, 63.89745, 65.30217, 
    65.12147, 57.81121, 63.64092, 55.16029, 68.9875, 70.49863, 63.15816, 
    6.344803,
  80.03839, 78.25382, 79.95118, 86.21111, 77.07464, 84.75726, 86.04649, 
    82.08135, 80.90128, 80.72463, 81.73735, 81.41127, 81.22662, 81.55504, 
    81.31358, 80.26396, 78.57015, 77.81126, 77.90018, 78.43227, 78.14822, 
    74.34625, 71.93066, 74.74102, 73.22122, 76.18527, 76.41434, 73.42256, 
    81.2297,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  3.263511, 2.871547, 3.068769, 2.57056, 2.73269, 2.376283, 2.028909, 
    2.238716, 2.151823, 1.968595, 2.13811, 2.184833, 2.147407, 2.162898, 
    2.439598, 2.308298, 2.099518, 2.77752, 2.550699, 2.676296, 2.88038, 
    2.923593, 3.093461, 2.655603, 2.539268, 9.024633, 8.603427, 4.242791, 
    15.3846,
  3.375126, 3.772299, 3.64349, 3.941743, 3.843183, 3.999619, 3.692043, 
    3.643797, 3.662182, 3.596931, 3.540162, 3.801683, 3.699805, 3.486027, 
    2.940073, 3.325436, 3.17168, 2.744081, 2.982688, 3.262203, 3.56422, 
    3.715354, 3.690225, 6.682123, 4.032764, 3.484746, 2.775695, 3.072027, 
    3.40358,
  3.883566, 3.920665, 3.831119, 3.926497, 3.514178, 3.667463, 3.94953, 
    3.605897, 3.500216, 3.82802, 3.960593, 3.706436, 4.232745, 3.892069, 
    10.36085, 4.281847, 3.928047, 3.493215, 3.569869, 3.726625, 3.703248, 
    3.901162, 3.766456, 8.395045, 4.101943, 3.719264, 3.482977, 3.642318, 
    4.006248,
  4.129162, 4.320088, 11.34565, 4.142805, 3.900762, 3.880364, 4.197795, 
    3.868919, 4.210166, 4.443914, 8.608879, 12.47732, 9.711339, 4.192898, 
    3.963542, 4.107327, 3.931527, 3.792522, 3.575509, 3.537056, 3.892575, 
    4.120211, 3.829014, 4.029256, 8.445096, 3.916228, 4.207069, 4.225374, 
    3.970522,
  3.552503, 9.473972, 9.532101, 3.773272, 4.145745, 4.266947, 3.91959, 
    4.109857, 3.873394, 4.291677, 11.63893, 12.03733, 3.940695, 3.62879, 
    3.701909, 3.802103, 3.8874, 3.651448, 3.852399, 3.939101, 4.134181, 
    3.839121, 3.541822, 3.880651, 8.468306, 8.875341, 3.846882, 3.784984, 
    3.663264,
  3.323679, 6.460494, 9.233714, 8.970462, 3.527218, 3.666316, 3.680627, 
    3.539894, 3.297183, 3.765352, 4.592725, 3.651731, 4.18259, 3.514647, 
    3.518247, 3.718238, 4.063127, 3.81191, 4.145193, 3.886687, 3.896607, 
    3.51206, 3.337671, 8.589912, 8.833002, 9.04817, 3.731555, 4.02777, 
    3.428335,
  3.245783, 8.69947, 8.486801, 10.10091, 3.579259, 3.562538, 3.203916, 
    3.210117, 8.613183, 8.617889, 3.338706, 3.352777, 3.256126, 3.44677, 
    3.397043, 3.525545, 3.622299, 3.722323, 3.667889, 3.790951, 3.685432, 
    3.616921, 3.299768, 8.274657, 8.532505, 3.574447, 3.512349, 3.448248, 
    3.288983,
  9.862949, 10.28637, 10.50127, 10.0743, 15.23599, 3.430345, 5.092399, 
    3.020758, 3.4208, 3.148396, 4.116941, 3.221134, 3.203755, 3.378935, 
    3.572417, 3.462322, 3.30362, 3.580242, 3.335833, 3.555261, 3.529677, 
    3.367766, 8.992569, 7.84314, 3.400465, 3.267994, 3.478723, 3.111313, 
    8.896255,
  19.47336, 21.78134, 23.60131, 3.576867, 24.277, 3.240448, 11.2632, 
    3.198735, 9.330683, 3.383981, 3.421008, 3.469214, 3.83172, 3.865665, 
    3.745772, 3.937711, 3.855377, 3.93339, 3.770758, 3.713422, 3.745214, 
    7.157488, 3.509474, 4.016141, 3.766808, 3.704838, 3.67332, 3.428144, 
    24.68721,
  25.8821, 21.88877, 22.79087, 20.88961, 13.85859, 15.88787, 13.38695, 
    10.82006, 8.169576, 11.14356, 3.618793, 3.607252, 3.563813, 3.813328, 
    3.656165, 3.647125, 3.882546, 3.976109, 3.88458, 3.862215, 11.65398, 
    12.56013, 9.834899, 3.742311, 3.581003, 4.125137, 3.922454, 3.935769, 
    11.98001,
  8.343321, 4.29432, 6.857409, 10.98879, 2.347787, 16.7195, 9.930901, 
    17.28986, 15.04951, 11.77565, 8.13041, 3.911289, 3.697823, 3.816411, 
    3.975359, 3.779339, 3.926732, 3.838076, 3.904479, 13.62941, 12.78611, 
    14.90687, 14.1657, 4.955834, 3.872963, 4.010866, 4.114388, 4.080603, 
    5.490836,
  6.799867, 13.89786, 15.28787, 16.58183, 15.54438, 13.44357, 9.464064, 
    12.82403, 8.609111, 8.172264, 7.971641, 7.7271, 4.301348, 4.365732, 
    4.146388, 4.234674, 4.222887, 4.20106, 4.465114, 10.24579, 11.7159, 
    11.38736, 8.089664, 7.590556, 6.079084, 4.430407, 4.373153, 4.321528, 
    4.748059,
  5.374411, 9.165045, 10.84608, 8.912563, 9.355453, 9.229032, 9.299223, 
    9.38324, 9.460958, 9.583862, 9.271997, 16.27015, 24.94757, 8.859853, 
    5.409078, 5.912062, 12.0257, 16.97542, 14.03381, 9.393799, 8.414137, 
    21.41707, 46.6626, 23.0479, 5.575336, 9.896134, 5.164502, 5.051294, 
    5.227304,
  6.43579, 6.835717, 12.51027, 7.02615, 14.3982, 59.88136, 43.08378, 
    41.04231, 34.49965, 33.69981, 17.20938, 15.30407, 33.17641, 58.88225, 
    58.30133, 54.94777, 37.31762, 35.04766, 52.86144, 18.66801, 35.24426, 
    48.52745, 35.72696, 50.14744, 27.48733, 69.51991, 74.656, 41.79357, 
    6.996423,
  60.89682, 57.11327, 56.84207, 60.40711, 43.83316, 58.52504, 60.40191, 
    59.89787, 60.01779, 60.29117, 60.42509, 60.63473, 60.65119, 60.79604, 
    60.66422, 60.52024, 60.41507, 60.523, 60.91508, 60.52288, 60.63238, 
    56.62858, 58.12341, 64.67667, 65.4202, 69.8543, 69.8737, 64.36972, 
    61.53412,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  3.849893, 3.856283, 3.876297, 3.722874, 3.312477, 3.303909, 3.728273, 
    3.271839, 3.404781, 3.456355, 3.315954, 3.216712, 3.217213, 3.979126, 
    4.067082, 4.12159, 4.292443, 4.25784, 4.043362, 4.088735, 4.206679, 
    4.139745, 3.941573, 3.650811, 4.270883, 4.339611, 4.129677, 4.173456, 
    4.11991,
  23.3913, 21.10123, 2.384663, 2.738321, 2.825331, 2.662113, 19.72605, 
    7.915842, 3.079172, 2.974945, 2.963715, 2.85387, 2.528532, 2.573021, 
    2.486332, 2.571714, 2.502167, 2.793546, 3.164559, 3.342665, 3.497552, 
    3.41118, 3.365852, 3.163154, 3.130959, 11.98952, 23.35816, 22.89286, 
    24.6501,
  3.378531, 2.953474, 3.242178, 3.110556, 3.257246, 3.378793, 3.477828, 
    4.037461, 3.990792, 3.864687, 4.04198, 3.742432, 3.57092, 3.773334, 
    3.453762, 3.615848, 3.763057, 3.640034, 3.907608, 3.400746, 3.747702, 
    3.555107, 3.321162, 6.382054, 3.734557, 3.742974, 3.305307, 3.465575, 
    3.282292,
  3.450989, 3.847913, 3.911248, 4.018094, 3.833026, 3.907627, 4.074425, 
    3.796141, 4.055058, 3.81418, 4.105705, 4.078651, 4.345757, 3.985118, 
    11.32582, 3.831229, 3.755456, 3.785145, 3.721199, 3.812036, 3.615114, 
    3.415135, 3.426016, 8.919117, 4.264057, 3.88468, 4.136335, 3.552783, 
    3.626698,
  4.0069, 4.28548, 11.58804, 4.11476, 4.076484, 3.958518, 4.007677, 3.613632, 
    3.982361, 4.3216, 8.783336, 12.74564, 10.93033, 4.248031, 3.976979, 
    3.862868, 3.842033, 3.751975, 3.70548, 3.541082, 3.761027, 4.017263, 
    3.579243, 4.299872, 8.528915, 4.067359, 4.048556, 3.931433, 3.905582,
  3.375264, 9.45883, 9.837132, 3.880792, 4.143943, 4.162468, 3.734957, 
    4.075751, 3.534219, 4.211858, 11.50331, 11.81786, 3.991126, 3.747541, 
    3.708467, 3.523463, 4.031811, 3.700854, 4.061032, 3.885763, 3.945246, 
    3.34333, 3.168113, 3.929471, 8.861012, 8.835147, 3.808527, 3.614073, 
    3.302133,
  3.318061, 6.23445, 9.393153, 9.185542, 3.713145, 3.694351, 3.499408, 
    3.543348, 3.500188, 3.765476, 4.678342, 3.610532, 4.049887, 3.383706, 
    3.619837, 3.695357, 4.014354, 3.784348, 4.012377, 3.752182, 3.752322, 
    3.40899, 3.431316, 8.917912, 8.802418, 9.150582, 3.86287, 4.01437, 
    3.529638,
  3.161242, 8.697525, 8.604968, 10.14865, 3.414701, 3.277946, 3.106585, 
    3.155272, 8.759369, 8.663495, 3.288543, 3.19271, 3.466063, 3.339281, 
    3.467445, 3.685304, 3.692217, 3.771382, 3.686859, 3.817103, 3.710386, 
    3.556711, 3.535718, 8.557709, 8.691965, 3.514397, 3.585006, 3.415441, 
    3.44202,
  9.784891, 10.24779, 9.976641, 9.295855, 14.96083, 3.111283, 5.009281, 
    3.02579, 3.463272, 3.099203, 4.215755, 3.193274, 3.242134, 3.30835, 
    3.361334, 3.386925, 3.369128, 3.485404, 3.240921, 3.412645, 3.253392, 
    3.228375, 8.81122, 7.650157, 3.368878, 3.217982, 3.178265, 3.101236, 
    8.80668,
  19.22267, 21.60826, 23.52611, 3.338216, 23.94795, 3.072971, 9.989408, 
    3.321576, 8.694997, 3.321878, 3.448324, 3.337141, 3.498293, 3.541253, 
    3.543709, 3.75351, 3.680443, 3.725989, 3.478187, 3.473844, 3.462271, 
    6.661892, 3.427514, 4.061265, 3.537899, 3.410243, 3.425969, 3.196785, 
    24.72017,
  25.36008, 21.49814, 22.59903, 20.63654, 13.53841, 15.82099, 12.61559, 
    10.37165, 7.683127, 10.83131, 3.689949, 3.787359, 3.420891, 3.647969, 
    3.902458, 3.636904, 3.915183, 3.865264, 3.799143, 3.928563, 11.88778, 
    12.17339, 9.500583, 3.66592, 3.675743, 3.925926, 3.92686, 3.699883, 
    11.71703,
  8.169175, 4.076253, 6.748446, 11.17791, 2.289379, 16.78876, 9.549583, 
    16.95436, 14.5035, 11.31938, 7.862218, 3.964858, 3.729162, 3.711964, 
    3.65044, 3.675449, 3.825419, 3.835011, 3.962104, 13.52691, 12.50951, 
    14.72277, 13.83352, 4.728748, 3.912308, 3.935472, 3.871082, 3.948413, 
    5.441088,
  6.575819, 13.68782, 15.24972, 15.68476, 14.95733, 13.67452, 9.135143, 
    11.64115, 8.331523, 8.041239, 7.795383, 7.292559, 4.094804, 4.116693, 
    4.004654, 3.996922, 3.990916, 4.04765, 4.190957, 10.43866, 11.87364, 
    11.01475, 7.708714, 7.455135, 5.668116, 4.197755, 4.393662, 4.134894, 
    4.560749,
  5.169791, 8.841509, 10.22076, 8.399336, 8.952921, 8.826251, 8.781018, 
    8.72908, 8.911089, 8.906417, 8.898951, 13.24638, 13.35855, 8.029644, 
    4.979704, 5.01109, 11.43125, 17.001, 12.86888, 8.891726, 8.065603, 
    13.92177, 6.374236, 13.20597, 5.60521, 10.18694, 4.989675, 5.126527, 
    4.832425,
  6.24145, 6.204876, 11.30593, 7.485038, 6.726289, 48.20478, 19.89283, 
    18.10007, 18.50454, 18.63955, 13.58515, 12.43399, 17.80441, 20.52042, 
    54.84818, 15.30902, 26.05787, 29.62769, 27.20374, 11.69455, 28.39441, 
    45.23884, 33.15934, 41.78193, 7.385835, 67.25801, 71.84697, 18.19055, 
    6.546476,
  60.07401, 43.80394, 48.32499, 55.75319, 35.60721, 52.76728, 59.96224, 
    58.50709, 59.74198, 60.18441, 60.20528, 60.21327, 60.2471, 60.25859, 
    60.2449, 60.25675, 60.31661, 60.29691, 60.48621, 60.64716, 60.14647, 
    51.25051, 52.23624, 58.10523, 69.70419, 65.57051, 73.06789, 60.31311, 
    44.12394,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  2.23983, 2.443991, 2.369467, 2.061352, 2.231854, 2.199944, 2.20608, 
    2.189638, 2.097535, 2.098871, 2.3531, 2.086133, 2.039821, 2.318063, 
    2.385066, 2.538923, 2.478305, 2.616679, 2.471617, 2.344972, 2.532229, 
    2.439283, 2.412121, 2.334194, 2.196361, 2.605808, 2.638407, 2.487885, 
    2.414575,
  25.21568, 25.38106, 26.26929, 24.3962, 22.1197, 22.12864, 24.32268, 
    22.13681, 22.21647, 22.34777, 22.2838, 22.31196, 22.61312, 26.23935, 
    26.30697, 26.22862, 26.19667, 26.23034, 26.08508, 26.00303, 26.31087, 
    25.8761, 25.92479, 24.37402, 26.44881, 26.64913, 26.54453, 26.41795, 
    26.32568,
  33.94374, 34.05513, 3.567151, 3.743794, 3.680321, 3.648973, 33.28426, 
    28.60334, 5.229125, 3.768654, 3.433515, 3.495399, 3.140697, 2.972671, 
    2.992865, 2.988852, 2.847082, 2.904128, 3.202813, 3.47594, 4.258402, 
    4.429258, 3.89246, 4.226138, 3.50216, 22.47453, 32.12323, 33.56538, 
    33.98292,
  3.986871, 4.270828, 3.962986, 3.7876, 3.54119, 3.481346, 3.856209, 
    3.818406, 3.958141, 4.172368, 3.84959, 3.958691, 3.805797, 3.899226, 
    3.477826, 3.817496, 3.699108, 3.566858, 3.574215, 3.658361, 3.555261, 
    3.915254, 3.910434, 8.117191, 4.188196, 3.827264, 3.5369, 3.87921, 3.96026,
  3.655027, 3.768519, 4.046415, 3.772287, 3.887514, 3.878178, 4.028559, 
    4.077557, 3.800567, 4.011391, 3.911467, 4.058834, 4.275026, 4.039367, 
    12.62784, 3.699128, 3.761713, 3.644035, 3.783242, 3.78049, 3.648092, 
    3.601111, 3.749682, 10.48611, 4.500976, 3.967303, 3.685591, 3.588793, 
    3.576775,
  3.77985, 3.6988, 12.45261, 3.985422, 3.892268, 4.03973, 3.855812, 4.0346, 
    3.863726, 4.212935, 9.077677, 13.52706, 10.32984, 3.924035, 4.089614, 
    3.863557, 3.777445, 3.623222, 3.756045, 3.646693, 3.929814, 3.795756, 
    3.943604, 4.593791, 8.499731, 3.741817, 3.628763, 3.739041, 3.68416,
  3.360407, 9.540145, 9.860668, 3.907832, 3.822461, 3.82277, 3.782165, 
    3.693602, 3.45107, 4.394618, 11.54702, 11.45898, 3.88114, 3.536068, 
    3.706231, 3.769371, 3.788575, 3.639736, 4.028832, 3.701462, 3.775473, 
    3.465806, 3.339548, 3.6957, 9.15306, 9.169831, 3.747611, 4.005865, 
    3.326907,
  3.248349, 6.060346, 9.453049, 9.052529, 3.520314, 3.568033, 3.233526, 
    3.374818, 3.485114, 3.496161, 4.733906, 3.557626, 4.044427, 3.411057, 
    3.604439, 3.422251, 3.69981, 3.961051, 3.835346, 3.729769, 3.813331, 
    3.287973, 3.302269, 9.054506, 8.70335, 9.105979, 3.919947, 3.747223, 
    3.354568,
  3.122762, 8.55567, 8.355515, 9.973453, 3.378729, 3.236324, 3.238411, 
    3.178522, 8.565884, 8.219251, 3.215302, 3.225085, 3.285427, 3.378826, 
    3.478092, 3.561123, 3.581481, 3.747563, 3.647296, 3.632422, 3.46284, 
    3.275675, 3.268298, 8.629727, 8.742919, 3.475494, 3.512121, 3.327066, 
    3.217284,
  9.555881, 9.858054, 9.483795, 9.106402, 14.87067, 3.284304, 5.066569, 
    3.062972, 3.314403, 3.186854, 4.178864, 3.126484, 3.259096, 3.403163, 
    3.180083, 3.408219, 3.235415, 3.221657, 3.240705, 3.321643, 3.138992, 
    3.251199, 8.816936, 7.305283, 3.255131, 3.083033, 2.956294, 3.112124, 
    8.507084,
  18.10869, 20.90464, 23.11588, 3.030486, 22.99694, 3.1357, 9.917166, 
    3.151852, 8.793662, 3.187633, 3.317825, 3.312697, 3.218035, 3.342903, 
    3.425536, 3.631901, 3.579019, 3.875694, 3.294317, 3.436236, 3.231664, 
    6.221606, 3.387435, 4.132294, 3.278371, 3.287123, 3.341487, 3.047742, 
    23.92474,
  24.53785, 20.70071, 21.31325, 19.87343, 12.95154, 15.00467, 12.09935, 
    9.990979, 7.163763, 10.37748, 3.631232, 3.547702, 3.702656, 3.639263, 
    3.541899, 3.930404, 3.852043, 4.097413, 3.71733, 3.946666, 12.31873, 
    12.02222, 9.268805, 3.40761, 3.711939, 3.769091, 4.069635, 3.596241, 
    11.26148,
  6.698274, 4.234491, 6.355492, 10.6562, 2.140969, 15.76149, 9.034671, 
    15.93241, 13.6342, 11.29838, 7.360078, 3.746908, 3.539001, 3.698002, 
    3.57632, 3.610885, 3.555323, 3.754485, 3.753139, 12.69716, 11.70098, 
    13.82215, 12.97426, 4.381145, 3.687301, 3.702881, 3.898651, 4.023606, 
    5.257266,
  6.113511, 12.57968, 14.0047, 14.60622, 13.79177, 12.70931, 8.372281, 
    11.4504, 7.765956, 7.147082, 7.110018, 6.958457, 3.905505, 3.824898, 
    3.736065, 3.666218, 3.805678, 3.806703, 4.222828, 9.444231, 10.93531, 
    9.989761, 7.042933, 6.854623, 5.361516, 4.172703, 4.123868, 4.255902, 
    3.898669,
  4.403711, 7.684649, 8.728783, 7.2373, 7.716644, 7.61562, 7.614408, 
    7.691447, 7.842656, 7.800129, 7.696713, 11.7016, 11.85282, 6.789203, 
    4.290509, 4.501255, 9.926376, 15.47871, 11.3439, 7.688498, 7.074048, 
    11.8417, 4.843839, 11.54759, 4.421161, 8.920911, 4.256143, 4.254754, 
    4.204268,
  4.902468, 5.356794, 8.584962, 5.182193, 4.990663, 5.959644, 13.45371, 
    13.23414, 13.93448, 13.77028, 10.48293, 10.05518, 13.44768, 5.727123, 
    22.71744, 5.045751, 10.6288, 10.26272, 6.977019, 8.426332, 25.44161, 
    20.3479, 18.82711, 29.10439, 5.707048, 52.92152, 56.82689, 8.719672, 
    4.964287,
  46.44859, 8.624842, 33.5353, 38.29524, 29.6681, 25.47851, 60.32549, 
    58.76976, 60.0569, 60.48402, 60.96387, 60.74286, 61.35557, 61.58157, 
    62.03634, 62.57771, 62.88708, 63.0727, 62.76698, 61.4595, 61.33596, 
    52.38147, 52.7865, 59.35516, 71.28531, 71.3038, 75.68409, 59.36493, 
    27.36596,
  20.42517, 20.42517, 20.42517, 20.42517, 20.42517, 20.42517, 20.42517, 
    20.09119, 20.09119, 20.09119, 20.09119, 20.09119, 20.09119, 20.09119, 
    20.08523, 20.08523, 20.08523, 20.08523, 20.08523, 20.08523, 20.08523, 
    20.22404, 20.22404, 20.22404, 20.22404, 20.22404, 20.22404, 20.22404, 
    20.42517,
  32.94125, 32.81193, 32.7462, 32.62016, 32.60735, 32.53995, 32.55154, 
    32.60879, 32.63617, 32.75629, 32.89869, 32.8534, 32.93066, 32.98158, 
    32.9904, 33.3036, 33.1595, 33.18209, 33.08523, 33.03173, 32.95968, 
    33.09716, 33.1664, 33.41994, 33.28544, 33.45037, 33.7359, 33.31431, 
    33.07684,
  41.40041, 41.49811, 43.02742, 40.09346, 36.54895, 36.48399, 39.82904, 
    36.51166, 36.56657, 36.69514, 36.67208, 36.65713, 37.04079, 42.89258, 
    43.07217, 41.98176, 41.53115, 42.28184, 42.39245, 42.49495, 42.80083, 
    42.0033, 42.42709, 39.5406, 42.0658, 43.13004, 43.20388, 43.27909, 
    43.22318,
  43.34626, 43.84412, 7.245405, 4.107951, 5.041785, 24.19967, 42.5238, 
    42.84676, 37.33493, 4.475881, 4.353141, 4.424299, 4.003063, 4.149846, 
    4.319924, 3.876502, 3.632577, 3.517452, 3.694416, 3.972339, 4.125613, 
    4.139646, 4.374284, 4.262466, 4.13805, 24.07879, 38.38928, 40.54487, 
    42.65262,
  3.824639, 3.737813, 3.852404, 3.687712, 3.893946, 3.991609, 3.946618, 
    4.100024, 4.196376, 4.026991, 4.008016, 4.01666, 3.919827, 4.156059, 
    3.909164, 3.821612, 3.651886, 3.473112, 3.713415, 3.675363, 3.917446, 
    3.937159, 3.801884, 8.744837, 4.108849, 3.953249, 3.754754, 3.710914, 
    3.700302,
  3.769916, 3.899818, 3.759683, 3.636419, 3.621782, 3.674057, 3.755948, 
    3.830639, 3.749517, 3.832144, 3.816481, 3.986923, 4.03429, 3.712, 
    13.58318, 3.648126, 3.924413, 3.673778, 3.428505, 3.615889, 3.824427, 
    3.960303, 3.854511, 11.54646, 4.417253, 3.875874, 3.655298, 3.665133, 
    3.660108,
  3.663294, 3.698711, 12.74467, 3.706316, 3.848587, 3.626447, 3.727762, 
    3.860199, 3.864508, 4.164116, 9.472161, 14.21188, 11.51188, 3.699133, 
    3.666499, 3.685274, 3.679271, 3.496044, 3.312791, 3.567279, 3.765356, 
    3.728959, 3.57938, 4.610554, 8.89137, 3.513083, 3.588584, 3.606128, 
    3.629589,
  3.211739, 9.627126, 10.16239, 3.791265, 3.777721, 3.815249, 3.685612, 
    3.596207, 3.57436, 3.77978, 11.98766, 11.84783, 3.708216, 3.492156, 
    3.585597, 3.522187, 3.631813, 3.723169, 3.767975, 3.830483, 3.604028, 
    3.308804, 3.222849, 3.668372, 8.989523, 9.204117, 3.843618, 3.676141, 
    3.516706,
  3.005261, 6.073549, 9.06297, 9.060443, 3.60012, 3.586196, 3.269781, 
    3.298595, 3.451119, 3.487191, 4.628163, 3.334808, 4.110469, 3.330947, 
    3.391282, 3.363851, 3.527205, 3.710023, 3.617498, 3.665666, 3.555247, 
    3.252955, 3.31916, 8.872885, 8.67463, 12.1769, 3.786543, 3.414071, 
    3.232029,
  3.21147, 8.193237, 8.145697, 9.871732, 3.427397, 3.198226, 3.101713, 
    3.100278, 8.561978, 8.101552, 3.349819, 3.430828, 3.445236, 3.422158, 
    3.483327, 3.570497, 3.549356, 3.713785, 3.49914, 3.528497, 3.328302, 
    3.229834, 3.147955, 8.456, 8.51399, 3.425318, 3.451754, 3.316885, 3.232519,
  9.472232, 9.751119, 9.683608, 9.38919, 14.58545, 3.225212, 4.99315, 
    3.033324, 3.197616, 3.115312, 3.961886, 3.144968, 3.267263, 3.157135, 
    3.186447, 3.270558, 3.253317, 3.394457, 3.269204, 3.237173, 3.154395, 
    3.133573, 8.584388, 7.294443, 3.427665, 3.222716, 3.159964, 3.094719, 
    8.360596,
  17.80005, 20.15772, 21.78689, 3.383359, 22.42377, 3.095594, 10.15558, 
    3.088015, 8.617355, 3.283748, 3.306589, 3.253113, 3.39214, 3.426768, 
    3.37475, 3.652326, 3.697832, 3.806445, 3.424033, 3.433588, 3.145402, 
    5.981155, 3.356054, 3.957218, 3.358468, 3.240247, 3.164384, 3.163117, 
    22.89814,
  23.05764, 19.41514, 20.09536, 18.86579, 12.588, 14.48705, 11.82205, 
    9.881642, 7.513378, 10.07812, 3.55706, 3.596499, 3.829221, 3.786097, 
    3.637519, 3.79669, 3.722465, 3.955158, 3.531701, 3.696517, 11.88948, 
    11.89851, 8.850475, 3.458386, 3.531002, 3.62397, 3.68233, 3.521421, 
    10.73441,
  6.227854, 3.89501, 6.177783, 9.957928, 1.979744, 14.75507, 8.627841, 
    14.61809, 12.65156, 10.96726, 7.199634, 3.675231, 3.522413, 3.572904, 
    3.695084, 3.467112, 3.391214, 3.470338, 3.703646, 11.74969, 10.68325, 
    12.73934, 12.2229, 4.338383, 3.777027, 3.840066, 3.873803, 3.780555, 
    5.245914,
  5.647316, 11.0129, 12.38766, 13.05047, 12.52302, 11.23402, 7.478331, 
    11.49345, 7.499798, 7.00538, 7.036828, 6.237599, 3.906703, 4.055851, 
    4.053195, 4.174885, 3.783634, 3.774828, 3.688944, 8.377676, 9.83066, 
    9.301428, 6.303364, 6.235791, 5.015049, 4.053378, 3.804047, 3.765507, 
    4.006456,
  4.391366, 6.472799, 7.523004, 6.216074, 6.466147, 6.503433, 6.538387, 
    6.722376, 6.729311, 7.07069, 6.813744, 11.89696, 10.96997, 6.351046, 
    3.964693, 4.27127, 8.861506, 12.84572, 9.849312, 7.302434, 6.03785, 
    11.35029, 3.91993, 10.46148, 4.040409, 7.975544, 4.582049, 4.642265, 
    4.44525,
  4.058449, 4.476113, 6.878038, 3.813162, 3.976066, 4.715731, 10.74337, 
    11.32191, 11.41297, 12.13756, 12.40652, 10.78269, 13.0156, 4.597189, 
    13.23346, 3.809593, 8.500738, 8.734775, 5.679147, 6.968148, 18.11316, 
    11.77869, 16.19608, 31.67456, 3.95826, 43.13771, 43.30083, 9.660636, 
    4.306415,
  13.56715, 5.160811, 10.48074, 11.97082, 16.8765, 21.0169, 43.48619, 
    43.55082, 44.19431, 44.87406, 44.93296, 46.32714, 46.88927, 46.42255, 
    46.39574, 46.27839, 45.83002, 45.13892, 44.89439, 45.91873, 47.12955, 
    46.08286, 41.01465, 46.908, 47.14761, 47.55635, 47.77073, 45.6171, 
    15.97072,
  76.32105, 76.32105, 76.32105, 76.32105, 76.32105, 76.32105, 76.32105, 
    76.26913, 76.26913, 76.26913, 76.26913, 76.26913, 76.26913, 76.26913, 
    76.28025, 76.28025, 76.28025, 76.28025, 76.28025, 76.28025, 76.28025, 
    76.33347, 76.33347, 76.33347, 76.33347, 76.33347, 76.33347, 76.33347, 
    76.32105,
  64.90369, 64.6298, 64.63443, 64.83301, 64.60438, 64.77776, 64.71052, 
    64.61693, 64.6462, 64.64974, 64.30616, 64.62667, 64.61202, 64.64821, 
    64.71255, 65.20638, 64.75205, 64.60986, 64.72108, 64.61427, 64.43154, 
    64.38303, 64.76843, 65.12057, 65.37663, 64.97582, 64.90881, 64.89304, 
    64.90021,
  55.46278, 56.32965, 59.34335, 55.24179, 50.3285, 50.47661, 55.33776, 
    50.47486, 50.2331, 50.42131, 50.47485, 50.2812, 50.76092, 59.0295, 
    59.42395, 58.79338, 58.38962, 58.24303, 58.40985, 58.65955, 58.74493, 
    59.22123, 58.74757, 53.72588, 57.0346, 55.81038, 53.18273, 53.08663, 
    55.35767,
  42.74674, 45.07474, 37.85433, 4.844555, 6.726536, 27.37482, 45.47479, 
    35.14567, 40.49166, 4.468805, 4.787293, 4.93224, 4.755197, 4.766776, 
    4.954597, 4.746784, 4.448916, 4.27868, 4.436535, 4.554966, 4.836428, 
    4.893676, 4.728329, 4.619895, 4.494048, 24.14004, 38.83576, 40.21775, 
    41.48883,
  3.759887, 4.124198, 4.102218, 4.042541, 4.047965, 4.171541, 4.080013, 
    4.047744, 3.918811, 3.918705, 3.975539, 4.040512, 4.217172, 4.272469, 
    4.353305, 4.128162, 3.913845, 3.942405, 3.881875, 3.990181, 4.057024, 
    4.104878, 4.093611, 9.022662, 4.761724, 4.04408, 3.751832, 3.964305, 
    3.711627,
  3.597251, 3.861883, 3.98396, 4.010903, 3.974269, 3.805978, 3.746219, 
    3.784802, 3.724791, 3.776561, 3.838946, 3.90498, 4.093378, 3.880047, 
    13.29206, 3.82261, 3.667262, 3.905445, 3.671196, 3.808156, 3.5578, 
    3.762915, 3.792232, 11.42567, 4.227711, 3.921521, 3.84165, 3.944218, 
    3.926139,
  3.453191, 3.769577, 12.44823, 3.635506, 3.718819, 3.570599, 3.806918, 
    3.610323, 3.568839, 3.998961, 9.999844, 14.93241, 10.75942, 3.847121, 
    3.793644, 3.727141, 3.608136, 3.802898, 3.535383, 3.788461, 3.57925, 
    3.650622, 3.505897, 4.613866, 9.256697, 3.443614, 3.705482, 3.734038, 
    3.691552,
  3.40959, 10.04336, 10.31814, 3.903711, 3.651334, 3.695894, 3.898786, 
    3.591596, 3.722478, 3.720148, 12.26171, 11.45577, 3.630054, 3.762288, 
    3.641325, 3.609985, 3.456588, 3.638541, 3.514789, 3.84078, 3.579578, 
    3.61583, 3.365269, 3.746, 9.247554, 9.009339, 3.547721, 3.459064, 3.583747,
  3.151502, 6.117112, 8.841331, 9.552134, 3.543856, 3.226698, 3.409431, 
    3.453269, 3.47725, 3.381563, 4.723243, 3.084631, 4.400764, 3.31239, 
    3.28071, 3.649858, 3.417897, 3.60295, 3.603931, 3.788716, 3.459665, 
    3.531705, 3.227995, 8.41416, 8.820116, 11.91147, 3.580215, 3.399566, 
    3.272576,
  3.355619, 8.005797, 8.086666, 9.973727, 3.474389, 3.536972, 3.432515, 
    3.287076, 8.420215, 8.444087, 3.187692, 3.197689, 3.268533, 3.390196, 
    3.464622, 3.689172, 3.631422, 3.715518, 3.619369, 3.739494, 3.475422, 
    3.136345, 3.283118, 8.476778, 8.514912, 3.50335, 3.596057, 3.421993, 
    3.47837,
  9.414896, 9.912844, 10.257, 9.036853, 14.64171, 3.569959, 4.932691, 
    3.468506, 3.447018, 3.144296, 3.931025, 3.139849, 3.041277, 3.16235, 
    3.174126, 2.994262, 3.295756, 3.197782, 3.23338, 3.291637, 3.22328, 
    3.085449, 8.601447, 7.418859, 3.267622, 3.246141, 3.098917, 3.064136, 
    8.668287,
  16.93372, 19.39404, 21.33942, 3.360438, 21.46722, 3.555222, 10.3599, 
    3.608676, 9.011078, 3.546573, 3.264677, 3.318602, 3.306113, 3.548603, 
    3.6917, 3.574667, 3.792122, 3.570747, 3.612278, 3.283613, 3.576888, 
    5.962729, 3.423355, 4.153275, 3.377117, 3.740672, 3.506525, 3.520546, 
    21.9014,
  21.70075, 18.03231, 18.83429, 17.46478, 11.81038, 13.65395, 11.62505, 
    9.458474, 8.352261, 10.01765, 3.379685, 3.303967, 3.538415, 3.69253, 
    3.648841, 3.480973, 3.782424, 3.608298, 3.725628, 3.446829, 11.12496, 
    11.01906, 8.683892, 3.572111, 3.381171, 3.911537, 3.899033, 4.180006, 
    9.879284,
  6.795138, 3.663016, 5.853401, 9.415535, 1.801388, 13.43976, 8.889196, 
    13.9995, 11.60817, 10.73502, 6.91687, 4.144278, 3.567039, 3.557197, 
    3.560689, 3.676418, 3.738649, 3.316923, 3.485469, 10.90593, 9.860681, 
    12.23584, 11.25569, 4.652129, 3.599483, 3.707473, 3.698868, 3.912867, 
    4.880559,
  5.383226, 9.84245, 10.9893, 11.40605, 10.66375, 9.853643, 7.602111, 
    15.64213, 9.81413, 6.983168, 9.442024, 7.068858, 3.863439, 3.933296, 
    4.053083, 3.638697, 3.593762, 3.209559, 3.585823, 7.802095, 8.617135, 
    8.31904, 6.973976, 8.467867, 4.685915, 3.45572, 3.53631, 4.001267, 
    4.131925,
  3.90865, 5.162776, 5.713617, 4.792522, 5.629866, 5.691249, 7.173501, 
    9.412261, 9.386623, 8.347288, 8.294571, 14.94284, 11.7121, 7.036501, 
    3.297727, 3.553821, 7.118531, 10.16525, 8.933929, 7.209597, 5.866919, 
    9.635096, 4.285679, 12.56851, 3.496054, 6.549919, 3.932243, 3.938029, 
    4.112247,
  2.853425, 3.414564, 5.4924, 3.225325, 3.134174, 4.178444, 11.87287, 
    12.38258, 17.76958, 23.88107, 15.04493, 7.321695, 8.730595, 24.01825, 
    29.05392, 3.113914, 19.46789, 15.97541, 4.35999, 5.696687, 24.51343, 
    22.21526, 23.66739, 25.38987, 3.455673, 28.37093, 28.48327, 19.81969, 
    2.5725,
  8.358735, 1.2442, 8.2303, 6.755699, 3.732956, 10.47798, 13.59545, 13.52574, 
    13.64481, 13.31298, 12.6013, 12.01397, 12.54815, 13.01806, 12.99609, 
    12.92617, 12.83615, 13.04976, 13.15103, 13.14319, 12.82171, 12.26593, 
    11.3403, 11.86761, 11.40641, 11.37071, 11.21965, 11.38273, 13.30919,
  76.29478, 76.29478, 76.29478, 76.29478, 76.29478, 76.29478, 76.29478, 
    76.26852, 76.26852, 76.26852, 76.26852, 76.26852, 76.26852, 76.26852, 
    76.24239, 76.24239, 76.24239, 76.24239, 76.24239, 76.24239, 76.24239, 
    76.30133, 76.30133, 76.30133, 76.30133, 76.30133, 76.30133, 76.30133, 
    76.29478,
  76.30904, 76.26852, 76.18663, 76.14668, 76.08985, 76.0851, 76.07748, 
    76.0287, 76.01533, 76.04591, 76.07558, 76.15076, 76.22458, 76.62688, 
    76.72932, 76.35542, 75.90929, 76.18436, 76.47408, 76.51854, 76.53927, 
    76.46555, 77.11685, 74.61399, 73.39807, 74.28423, 74.22876, 76.46761, 
    76.35101,
  62.69817, 37.59571, 63.73626, 67.86379, 68.00912, 68.05811, 68.46545, 
    67.71501, 67.41134, 67.45674, 67.58029, 67.48372, 67.26883, 75.11686, 
    74.22889, 73.59544, 71.9571, 72.15868, 71.60004, 72.94436, 72.54318, 
    70.4544, 64.41242, 61.62423, 64.78989, 61.90934, 58.9573, 59.94139, 
    60.21424,
  45.26468, 46.33259, 39.80659, 4.880448, 4.668566, 4.750793, 11.51619, 
    4.840425, 8.81459, 4.923784, 4.710509, 4.713686, 4.632531, 4.755519, 
    4.947788, 4.68797, 4.501524, 4.491595, 4.820996, 5.020241, 5.106737, 
    5.158825, 5.157003, 5.050581, 4.818464, 7.275883, 21.36522, 29.6608, 
    42.62926,
  4.201563, 4.151055, 4.31405, 4.311779, 4.333702, 4.295519, 4.260652, 
    4.279875, 4.219009, 4.270357, 4.372364, 4.466399, 4.475421, 4.399734, 
    4.466805, 4.172714, 4.193775, 4.162163, 4.010971, 4.292985, 4.211893, 
    4.290444, 4.04375, 8.653903, 4.896769, 4.467879, 4.243398, 4.315917, 
    4.266707,
  3.94139, 4.011866, 4.371395, 4.094247, 4.075, 4.058349, 3.986454, 4.076413, 
    3.780067, 4.059334, 3.86656, 4.089129, 4.323344, 4.184918, 9.953151, 
    3.952351, 3.969993, 3.770141, 3.810992, 3.868167, 3.772148, 3.811777, 
    3.982652, 9.946915, 4.343589, 4.003659, 3.64007, 3.897705, 3.739297,
  3.875742, 4.068198, 12.89322, 3.719746, 3.74136, 3.750169, 3.767522, 
    3.80456, 3.692979, 4.255264, 10.27328, 15.87072, 11.23041, 3.780274, 
    3.830738, 3.870037, 3.811691, 3.848084, 3.947021, 3.676383, 3.764634, 
    3.947807, 3.771096, 4.790236, 9.747645, 3.843821, 3.733427, 3.813056, 
    3.818707,
  3.332808, 10.355, 10.60618, 3.815717, 3.731721, 3.819657, 3.950878, 
    3.702467, 3.764491, 3.717438, 12.72409, 12.20723, 3.651446, 3.552197, 
    3.656971, 3.77964, 3.539301, 3.688996, 3.440627, 4.05953, 3.780515, 
    3.601847, 3.334125, 3.623432, 9.339285, 9.269832, 3.762157, 3.53513, 
    3.537027,
  3.180831, 6.020929, 8.839355, 9.200312, 3.472956, 3.326724, 3.599181, 
    3.466324, 3.477169, 3.368377, 4.823409, 3.348995, 4.455943, 3.390975, 
    3.401223, 3.487251, 3.427177, 3.743241, 3.633617, 3.936927, 3.568148, 
    3.509787, 3.293755, 8.745516, 8.753927, 9.028022, 3.69135, 3.513023, 
    3.693835,
  3.235761, 8.120193, 8.167442, 9.55004, 3.466782, 3.418832, 3.518373, 
    3.353072, 8.459551, 8.432825, 3.187175, 3.288986, 3.185555, 3.486019, 
    3.619438, 3.687609, 3.756171, 3.808496, 3.67426, 3.80761, 3.472903, 
    3.208827, 3.393583, 8.424366, 8.419132, 3.488642, 3.277623, 3.437188, 
    3.427883,
  9.796509, 10.04021, 9.831751, 9.227248, 14.15211, 3.453925, 5.222262, 
    3.399982, 3.46829, 3.350626, 4.005218, 3.39972, 3.101459, 3.107916, 
    3.315438, 3.334515, 3.515921, 3.239099, 3.569389, 3.289895, 3.584881, 
    3.352013, 8.569733, 7.271706, 3.43695, 3.580975, 3.165626, 3.280397, 
    8.771801,
  16.51744, 18.69143, 20.39238, 3.776779, 20.59461, 3.677503, 10.51283, 
    3.713278, 8.71023, 3.673811, 3.417988, 3.745603, 3.733539, 3.732467, 
    3.817034, 3.692412, 3.698813, 3.599589, 3.641639, 3.384573, 3.826808, 
    6.144732, 3.877209, 4.291211, 3.627161, 3.788675, 3.370625, 3.665258, 
    21.08022,
  20.46859, 17.0886, 17.58566, 16.38467, 10.90745, 12.87932, 10.97016, 
    17.35693, 9.789871, 9.704507, 3.483038, 3.759705, 3.870174, 3.843338, 
    3.6004, 3.711369, 3.856496, 3.810298, 3.706984, 4.271911, 9.099217, 
    10.64838, 8.217738, 3.82382, 3.763711, 3.558376, 3.876113, 4.048146, 
    9.65414,
  5.747074, 4.006268, 5.501839, 8.638597, 1.65025, 12.33786, 8.678884, 
    12.3184, 10.94792, 10.37151, 7.06738, 3.578495, 3.316818, 3.234298, 
    3.557645, 3.591391, 3.407844, 3.442925, 3.488613, 10.20876, 10.25232, 
    11.5826, 10.41125, 4.329733, 3.737321, 3.526857, 3.718681, 3.543477, 
    4.660561,
  4.605869, 8.475582, 9.076962, 9.47061, 8.938696, 8.717731, 6.332824, 
    27.67833, 14.51656, 6.571701, 10.08075, 8.213726, 3.64196, 3.555236, 
    3.961901, 4.099989, 3.881661, 3.572167, 3.497919, 9.383901, 9.09608, 
    8.998482, 7.409111, 16.15083, 4.248996, 3.479935, 3.624752, 3.897249, 
    4.111664,
  3.743334, 7.708599, 5.486861, 8.361729, 7.157138, 8.026904, 12.06392, 
    14.67469, 13.0825, 9.977619, 8.236951, 23.10231, 23.11611, 10.65085, 
    3.056688, 3.909323, 16.91984, 10.16638, 22.2758, 7.86018, 8.834314, 
    21.17439, 2.475259, 21.60678, 2.663831, 5.367994, 3.306719, 3.30759, 
    3.763198,
  1.291596, 0.9332163, 2.561215, 0.7971681, 0.7588809, 1.105934, 8.221596, 
    8.14767, 7.566274, 7.399941, 4.847243, 3.127383, 7.504849, 9.55926, 
    9.353975, 5.610487, 8.225322, 8.47736, 7.774258, 6.425588, 7.858152, 
    8.778911, 8.046515, 7.778044, 1.502571, 7.950519, 8.070286, 8.121929, 
    1.128979,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  76.07452, 76.07452, 76.07452, 76.07452, 76.07452, 76.07452, 76.07452, 
    76.00054, 76.00054, 76.00054, 76.00054, 76.00054, 76.00054, 76.00054, 
    75.99906, 75.99906, 75.99906, 75.99906, 75.99906, 75.99906, 75.99906, 
    76.03716, 76.03716, 76.03716, 76.03716, 76.03716, 76.03716, 76.03716, 
    76.07452,
  76.23776, 76.06744, 75.97851, 75.93897, 75.93933, 75.96429, 75.93755, 
    75.9159, 75.93393, 75.95274, 75.96122, 76.07576, 76.21194, 74.26964, 
    68.83714, 66.3562, 67.03481, 67.30183, 71.08145, 75.5315, 76.10185, 
    76.10247, 75.96873, 64.99692, 65.36275, 65.31129, 64.52369, 67.46635, 
    76.14603,
  47.08821, 39.78064, 65.17686, 67.06091, 75.39043, 75.62454, 54.02661, 
    76.28989, 75.92274, 75.67311, 75.77917, 75.83623, 72.31573, 70.41719, 
    67.30744, 63.81781, 60.51402, 62.70388, 62.79856, 63.08656, 64.12659, 
    56.74884, 63.06895, 63.94172, 62.46814, 62.30279, 46.9643, 62.07563, 
    65.29506,
  28.70593, 24.29932, 5.277404, 4.664639, 4.733109, 4.740892, 4.712512, 
    4.933883, 4.723403, 5.195364, 4.863607, 5.131938, 4.87483, 5.037911, 
    5.217434, 5.140977, 4.973939, 4.822694, 5.080806, 5.114286, 5.077697, 
    4.996029, 5.008913, 4.972516, 4.86502, 4.792601, 4.877259, 5.121644, 
    12.98983,
  4.242709, 4.477846, 4.294391, 4.488003, 4.357565, 4.338476, 4.446472, 
    4.390183, 4.360558, 4.408836, 4.546145, 4.411483, 4.437038, 4.52511, 
    4.588255, 4.485234, 4.425212, 4.546773, 4.422399, 4.574793, 4.428821, 
    4.426642, 4.49695, 8.935439, 5.102932, 4.47962, 4.352555, 4.394399, 
    4.31924,
  4.098804, 4.198433, 4.449523, 4.097005, 4.076146, 4.286565, 3.934423, 
    4.09562, 4.029839, 3.877523, 3.965692, 4.479001, 4.151289, 4.015486, 
    10.35105, 3.922551, 4.218702, 4.150631, 3.862169, 3.932716, 4.129335, 
    4.04199, 4.2734, 10.22346, 4.441556, 4.373238, 4.121648, 4.090972, 
    4.135964,
  3.799037, 4.181551, 13.122, 3.751425, 3.922001, 4.028002, 3.687085, 
    3.914338, 3.908565, 4.102907, 10.39286, 16.10341, 10.87443, 3.962623, 
    3.945045, 3.729527, 3.972012, 3.647161, 3.494816, 3.76027, 4.089788, 
    4.043815, 3.952126, 4.859788, 9.687916, 3.941732, 3.778603, 3.785552, 
    3.765045,
  3.622912, 10.14244, 10.3128, 3.867978, 3.530591, 3.436364, 3.921525, 
    3.841564, 3.823227, 4.102831, 12.51932, 11.68597, 3.862648, 3.637559, 
    3.448077, 3.686473, 3.61252, 3.639603, 3.882136, 4.104214, 3.957531, 
    3.893538, 3.315006, 3.330784, 9.600559, 9.133184, 3.779639, 3.998035, 
    3.798149,
  3.332698, 6.781849, 8.950177, 9.335812, 3.323235, 3.42967, 3.561319, 
    3.412487, 3.695856, 3.343009, 4.94712, 3.316008, 4.531771, 3.700585, 
    3.637039, 3.73866, 3.600437, 3.875443, 3.696248, 3.970558, 3.781482, 
    3.769193, 3.387362, 9.030635, 8.611618, 9.098142, 4.085333, 3.62775, 
    3.722712,
  3.226397, 8.863524, 8.44458, 9.837615, 3.393033, 3.319263, 3.32145, 
    3.244461, 8.550245, 8.21362, 3.318355, 3.421618, 3.307756, 3.593971, 
    3.586608, 3.706766, 3.862183, 3.992337, 3.819756, 3.93947, 3.708955, 
    3.313099, 3.509924, 8.525232, 8.511231, 3.397391, 3.302927, 3.442458, 
    3.324693,
  10.15579, 10.30067, 10.27834, 9.530962, 14.23251, 3.497124, 5.580375, 
    3.773961, 3.494882, 3.444101, 3.971205, 3.308688, 3.445687, 3.560337, 
    3.384125, 3.4559, 3.818717, 3.291538, 3.496067, 3.266223, 3.291957, 
    3.448824, 8.504575, 7.272306, 3.578774, 3.734716, 3.161728, 3.756382, 
    9.166369,
  15.87409, 18.47683, 20.7076, 3.649283, 20.40932, 3.998232, 10.29874, 
    3.877515, 9.137363, 3.268897, 3.27869, 3.878571, 3.864924, 4.041171, 
    4.186173, 3.669262, 3.985262, 3.824546, 3.569679, 3.433971, 3.961447, 
    6.000515, 3.868928, 4.85245, 3.943801, 4.243917, 3.738083, 3.567279, 
    21.03829,
  20.07133, 16.46431, 16.99092, 16.12315, 10.76974, 12.59963, 11.23757, 
    22.38011, 16.87654, 9.544673, 3.381925, 3.788702, 4.119921, 3.816537, 
    3.515094, 3.704862, 3.718484, 3.97688, 3.851808, 3.923357, 8.550056, 
    10.18563, 8.113522, 3.488494, 3.902388, 3.823717, 4.091905, 3.791627, 
    9.709495,
  5.574897, 4.423749, 5.452045, 11.50318, 1.533152, 10.90562, 16.86831, 
    12.27624, 10.12835, 12.47072, 7.53353, 3.573075, 3.743525, 3.755694, 
    3.727368, 3.76037, 3.161195, 3.272928, 3.577691, 10.42197, 15.32513, 
    11.7495, 10.20657, 4.132444, 3.66544, 3.518038, 3.891251, 3.97131, 
    4.699478,
  3.826842, 7.969535, 11.62514, 15.42164, 12.25134, 15.7647, 9.899959, 
    25.54912, 14.56804, 6.937693, 11.18779, 11.23886, 3.539949, 3.755506, 
    4.003037, 3.359331, 3.57896, 3.228468, 3.513859, 12.04069, 11.82376, 
    15.23148, 10.29594, 20.54312, 5.637074, 3.43277, 3.26886, 3.248068, 
    3.125845,
  2.491312, 12.81094, 7.388693, 12.31697, 8.81054, 9.459171, 12.4113, 
    13.81019, 12.87046, 10.82043, 8.736136, 18.45498, 18.26361, 12.66025, 
    2.359894, 4.170528, 16.18436, 7.71747, 17.95869, 9.912076, 11.25335, 
    18.51919, 19.1211, 18.4709, 2.127753, 5.513164, 2.406839, 2.451899, 
    2.142247,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0 ;

 lat = -89.5, -79.5, -69.5, -59.5, -49.5, -39.5, -29.5, -19.5, -9.5, 0.5, 
    10.5, 20.5, 30.5, 40.5, 50.5, 60.5, 70.5, 80.5 ;

 lat_bnds =
  -90, -89,
  -80, -79,
  -70, -69,
  -60, -59,
  -50, -49,
  -40, -39,
  -30, -29,
  -20, -19,
  -10, -9,
  0, 1,
  10, 11,
  20, 21,
  30, 31,
  40, 41,
  50, 51,
  60, 61,
  70, 71,
  80, 81 ;

 lon = 0.625, 13.125, 25.625, 38.125, 50.625, 63.125, 75.625, 88.125, 
    100.625, 113.125, 125.625, 138.125, 150.625, 163.125, 175.625, 188.125, 
    200.625, 213.125, 225.625, 238.125, 250.625, 263.125, 275.625, 288.125, 
    300.625, 313.125, 325.625, 338.125, 350.625 ;

 lon_bnds =
  0, 1.25,
  12.5, 13.75,
  25, 26.25,
  37.5, 38.75,
  50, 51.25,
  62.5, 63.75,
  75, 76.25,
  87.5, 88.75,
  100, 101.25,
  112.5, 113.75,
  125, 126.25,
  137.5, 138.75,
  150, 151.25,
  162.5, 163.75,
  175, 176.25,
  187.5, 188.75,
  200, 201.25,
  212.5, 213.75,
  225, 226.25,
  237.5, 238.75,
  250, 251.25,
  262.5, 263.75,
  275, 276.25,
  287.5, 288.75,
  300, 301.25,
  312.5, 313.75,
  325, 326.25,
  337.5, 338.75,
  350, 351.25 ;

 time = 746.5, 776, 805.5, 836, 866.5, 897, 927.5, 958.5, 989, 1019.5, 1050, 
    1080.5 ;

 time_bnds =
  731, 762,
  762, 790,
  790, 821,
  821, 851,
  851, 882,
  882, 912,
  912, 943,
  943, 974,
  974, 1004,
  1004, 1035,
  1035, 1065,
  1065, 1096 ;
}
