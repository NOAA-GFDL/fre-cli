netcdf \20030101.grid_spec.tile5 {
dimensions:
	grid_x = 97 ;
	grid_y = 97 ;
	time = UNLIMITED ; // (1 currently)
	grid_xt = 96 ;
	grid_yt = 96 ;
	phalf = 50 ;
variables:
	double grid_x(grid_x) ;
		grid_x:units = "degrees_E" ;
		grid_x:long_name = "cell corner longitude" ;
		grid_x:axis = "X" ;
	double grid_y(grid_y) ;
		grid_y:units = "degrees_N" ;
		grid_y:long_name = "cell corner latitude" ;
		grid_y:axis = "Y" ;
	double time(time) ;
		time:units = "days since 1870-01-01 00:00:00" ;
		time:long_name = "time" ;
		time:axis = "T" ;
		time:calendar_type = "JULIAN" ;
		time:calendar = "julian" ;
	double grid_xt(grid_xt) ;
		grid_xt:units = "degrees_E" ;
		grid_xt:long_name = "T-cell longitude" ;
		grid_xt:axis = "X" ;
	double grid_yt(grid_yt) ;
		grid_yt:units = "degrees_N" ;
		grid_yt:long_name = "T-cell latitude" ;
		grid_yt:axis = "Y" ;
	double phalf(phalf) ;
		phalf:units = "mb" ;
		phalf:long_name = "ref half pressure level" ;
		phalf:axis = "Z" ;
		phalf:positive = "down" ;
	float grid_lon(grid_y, grid_x) ;
		grid_lon:_FillValue = 1.e+20f ;
		grid_lon:missing_value = 1.e+20f ;
		grid_lon:units = "degrees_E" ;
		grid_lon:long_name = "longitude" ;
		grid_lon:cell_methods = "time: point" ;
	float grid_lat(grid_y, grid_x) ;
		grid_lat:_FillValue = 1.e+20f ;
		grid_lat:missing_value = 1.e+20f ;
		grid_lat:units = "degrees_N" ;
		grid_lat:long_name = "latitude" ;
		grid_lat:cell_methods = "time: point" ;
	float grid_lont(grid_yt, grid_xt) ;
		grid_lont:_FillValue = 1.e+20f ;
		grid_lont:missing_value = 1.e+20f ;
		grid_lont:units = "degrees_E" ;
		grid_lont:long_name = "longitude" ;
		grid_lont:cell_methods = "time: point" ;
	float grid_latt(grid_yt, grid_xt) ;
		grid_latt:_FillValue = 1.e+20f ;
		grid_latt:missing_value = 1.e+20f ;
		grid_latt:units = "degrees_N" ;
		grid_latt:long_name = "latitude" ;
		grid_latt:cell_methods = "time: point" ;
	float area(grid_yt, grid_xt) ;
		area:_FillValue = 1.e+20f ;
		area:missing_value = 1.e+20f ;
		area:units = "m**2" ;
		area:long_name = "cell area" ;
		area:cell_methods = "time: point" ;
	float bk(phalf) ;
		bk:_FillValue = 1.e+20f ;
		bk:missing_value = 1.e+20f ;
		bk:long_name = "vertical coordinate sigma value" ;
		bk:cell_methods = "time: point" ;
	float pk(phalf) ;
		pk:_FillValue = 1.e+20f ;
		pk:missing_value = 1.e+20f ;
		pk:units = "pascal" ;
		pk:long_name = "pressure part of the hybrid coordinate" ;
		pk:cell_methods = "time: point" ;
	float sftlf(grid_yt, grid_xt) ;
		sftlf:_FillValue = 1.e+20f ;
		sftlf:missing_value = 1.e+20f ;
		sftlf:units = "1.0" ;
		sftlf:long_name = "Fraction of the Grid Cell Occupied by Land" ;
		sftlf:cell_methods = "time: point" ;
		sftlf:cell_measures = "area: area" ;
		sftlf:standard_name = "land_area_fraction" ;
		sftlf:interp_method = "conserve_order1" ;
	float orog(grid_yt, grid_xt) ;
		orog:_FillValue = 1.e+20f ;
		orog:missing_value = 1.e+20f ;
		orog:units = "m" ;
		orog:long_name = "Surface Altitude" ;
		orog:cell_methods = "time: point" ;
		orog:cell_measures = "area: area" ;
		orog:standard_name = "surface_altitude" ;
		orog:interp_method = "conserve_order1" ;
	float land_mask(grid_yt, grid_xt) ;
		land_mask:_FillValue = 1.e+20f ;
		land_mask:missing_value = 1.e+20f ;
		land_mask:valid_range = -0.01f, 1.01f ;
		land_mask:long_name = "fractional amount of land" ;
		land_mask:cell_methods = "time: point" ;
		land_mask:interp_method = "conserve_order1" ;
	float zsurf(grid_yt, grid_xt) ;
		zsurf:_FillValue = 1.e+20f ;
		zsurf:missing_value = 1.e+20f ;
		zsurf:units = "m" ;
		zsurf:long_name = "surface height" ;
		zsurf:cell_methods = "time: point" ;

// global attributes:
		:title = "ESM4_longamip_D1_am4p2_proto7b_whiteCapsAlbedo_salt_SIS2" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
data:

 grid_x = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19, 
    20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 37, 
    38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 54, 55, 
    56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 72, 73, 
    74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 90, 91, 
    92, 93, 94, 95, 96, 97 ;

 grid_y = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19, 
    20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 37, 
    38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 54, 55, 
    56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 72, 73, 
    74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 90, 91, 
    92, 93, 94, 95, 96, 97 ;

 time = 0 ;

 grid_xt = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19, 
    20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 37, 
    38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 54, 55, 
    56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 72, 73, 
    74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 90, 91, 
    92, 93, 94, 95, 96 ;

 grid_yt = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19, 
    20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 37, 
    38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 54, 55, 
    56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 72, 73, 
    74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 90, 91, 
    92, 93, 94, 95, 96 ;

 phalf = 0.01, 0.0269722, 0.0517136, 0.0889455, 0.142479, 0.2207157, 
    0.3361283, 0.5048096, 0.7479993, 1.0940055, 1.580046, 2.2544108, 
    3.178956, 4.431935, 6.1111558, 8.3374392, 11.2583405, 15.0520759, 
    19.9315829, 26.1486254, 33.997842, 43.820624, 56.0087014, 71.0073115, 
    89.3178242, 111.4997021, 138.1716841, 170.012093, 207.7581856, 
    252.2033875, 304.1464563, 363.9522552, 430.6429622, 501.015122, 
    570.6113482, 635.806353, 694.8286462, 747.1992533, 793.0044191, 
    832.5750255, 866.4443202, 895.1917865, 919.4060705, 939.6860264, 
    956.4664631, 970.1833931, 981.1347983, 989.68, 995.9, 1000 ;

 grid_lon =
  215, 215, 215, 215, 215, 215, 215, 215, 215, 215, 215, 215, 215, 215, 215, 
    215, 215, 215, 215, 215, 215, 215, 215, 215, 215, 215, 215, 215, 215, 
    215, 215, 215, 215, 215, 215, 215, 215, 215, 215, 215, 215, 215, 215, 
    215, 215, 215, 215, 215, 215, 215, 215, 215, 215, 215, 215, 215, 215, 
    215, 215, 215, 215, 215, 215, 215, 215, 215, 215, 215, 215, 215, 215, 
    215, 215, 215, 215, 215, 215, 215, 215, 215, 215, 215, 215, 215, 215, 
    215, 215, 215, 215, 215, 215, 215, 215, 215, 215, 215, 215,
  215.7828, 215.7828, 215.7828, 215.7828, 215.7828, 215.7828, 215.7828, 
    215.7828, 215.7828, 215.7828, 215.7828, 215.7828, 215.7828, 215.7828, 
    215.7828, 215.7828, 215.7828, 215.7828, 215.7828, 215.7828, 215.7828, 
    215.7828, 215.7828, 215.7828, 215.7828, 215.7828, 215.7828, 215.7828, 
    215.7828, 215.7828, 215.7828, 215.7828, 215.7828, 215.7828, 215.7828, 
    215.7828, 215.7828, 215.7828, 215.7828, 215.7828, 215.7828, 215.7828, 
    215.7828, 215.7828, 215.7828, 215.7828, 215.7828, 215.7828, 215.7828, 
    215.7828, 215.7828, 215.7828, 215.7828, 215.7828, 215.7828, 215.7828, 
    215.7828, 215.7828, 215.7828, 215.7828, 215.7828, 215.7828, 215.7828, 
    215.7828, 215.7828, 215.7828, 215.7828, 215.7828, 215.7828, 215.7828, 
    215.7828, 215.7828, 215.7828, 215.7828, 215.7828, 215.7828, 215.7828, 
    215.7828, 215.7828, 215.7828, 215.7828, 215.7828, 215.7828, 215.7828, 
    215.7828, 215.7828, 215.7828, 215.7828, 215.7828, 215.7828, 215.7828, 
    215.7828, 215.7828, 215.7828, 215.7828, 215.7828, 215.7828,
  216.5727, 216.5727, 216.5727, 216.5727, 216.5727, 216.5727, 216.5727, 
    216.5727, 216.5727, 216.5727, 216.5727, 216.5727, 216.5727, 216.5727, 
    216.5727, 216.5727, 216.5727, 216.5727, 216.5727, 216.5727, 216.5727, 
    216.5727, 216.5727, 216.5727, 216.5727, 216.5727, 216.5727, 216.5727, 
    216.5727, 216.5727, 216.5727, 216.5727, 216.5727, 216.5727, 216.5727, 
    216.5727, 216.5727, 216.5727, 216.5727, 216.5727, 216.5727, 216.5727, 
    216.5727, 216.5727, 216.5727, 216.5727, 216.5727, 216.5727, 216.5727, 
    216.5727, 216.5727, 216.5727, 216.5727, 216.5727, 216.5727, 216.5727, 
    216.5727, 216.5727, 216.5727, 216.5727, 216.5727, 216.5727, 216.5727, 
    216.5727, 216.5727, 216.5727, 216.5727, 216.5727, 216.5727, 216.5727, 
    216.5727, 216.5727, 216.5727, 216.5727, 216.5727, 216.5727, 216.5727, 
    216.5727, 216.5727, 216.5727, 216.5727, 216.5727, 216.5727, 216.5727, 
    216.5727, 216.5727, 216.5727, 216.5727, 216.5727, 216.5727, 216.5727, 
    216.5727, 216.5727, 216.5727, 216.5727, 216.5727, 216.5727,
  217.3698, 217.3698, 217.3698, 217.3698, 217.3698, 217.3698, 217.3698, 
    217.3698, 217.3698, 217.3698, 217.3698, 217.3698, 217.3698, 217.3698, 
    217.3698, 217.3698, 217.3698, 217.3698, 217.3698, 217.3698, 217.3698, 
    217.3698, 217.3698, 217.3698, 217.3698, 217.3698, 217.3698, 217.3698, 
    217.3698, 217.3698, 217.3698, 217.3698, 217.3698, 217.3698, 217.3698, 
    217.3698, 217.3698, 217.3698, 217.3698, 217.3698, 217.3698, 217.3698, 
    217.3698, 217.3698, 217.3698, 217.3698, 217.3698, 217.3698, 217.3698, 
    217.3698, 217.3698, 217.3698, 217.3698, 217.3698, 217.3698, 217.3698, 
    217.3698, 217.3698, 217.3698, 217.3698, 217.3698, 217.3698, 217.3698, 
    217.3698, 217.3698, 217.3698, 217.3698, 217.3698, 217.3698, 217.3698, 
    217.3698, 217.3698, 217.3698, 217.3698, 217.3698, 217.3698, 217.3698, 
    217.3698, 217.3698, 217.3698, 217.3698, 217.3698, 217.3698, 217.3698, 
    217.3698, 217.3698, 217.3698, 217.3698, 217.3698, 217.3698, 217.3698, 
    217.3698, 217.3698, 217.3698, 217.3698, 217.3698, 217.3698,
  218.1741, 218.1741, 218.1741, 218.1741, 218.1741, 218.1741, 218.1741, 
    218.1741, 218.1741, 218.1741, 218.1741, 218.1741, 218.1741, 218.1741, 
    218.1741, 218.1741, 218.1741, 218.1741, 218.1741, 218.1741, 218.1741, 
    218.1741, 218.1741, 218.1741, 218.1741, 218.1741, 218.1741, 218.1741, 
    218.1741, 218.1741, 218.1741, 218.1741, 218.1741, 218.1741, 218.1741, 
    218.1741, 218.1741, 218.1741, 218.1741, 218.1741, 218.1741, 218.1741, 
    218.1741, 218.1741, 218.1741, 218.1741, 218.1741, 218.1741, 218.1741, 
    218.1741, 218.1741, 218.1741, 218.1741, 218.1741, 218.1741, 218.1741, 
    218.1741, 218.1741, 218.1741, 218.1741, 218.1741, 218.1741, 218.1741, 
    218.1741, 218.1741, 218.1741, 218.1741, 218.1741, 218.1741, 218.1741, 
    218.1741, 218.1741, 218.1741, 218.1741, 218.1741, 218.1741, 218.1741, 
    218.1741, 218.1741, 218.1741, 218.1741, 218.1741, 218.1741, 218.1741, 
    218.1741, 218.1741, 218.1741, 218.1741, 218.1741, 218.1741, 218.1741, 
    218.1741, 218.1741, 218.1741, 218.1741, 218.1741, 218.1741,
  218.9857, 218.9857, 218.9857, 218.9857, 218.9857, 218.9857, 218.9857, 
    218.9857, 218.9857, 218.9857, 218.9857, 218.9857, 218.9857, 218.9857, 
    218.9857, 218.9857, 218.9857, 218.9857, 218.9857, 218.9857, 218.9857, 
    218.9857, 218.9857, 218.9857, 218.9857, 218.9857, 218.9857, 218.9857, 
    218.9857, 218.9857, 218.9857, 218.9857, 218.9857, 218.9857, 218.9857, 
    218.9857, 218.9857, 218.9857, 218.9857, 218.9857, 218.9857, 218.9857, 
    218.9857, 218.9857, 218.9857, 218.9857, 218.9857, 218.9857, 218.9857, 
    218.9857, 218.9857, 218.9857, 218.9857, 218.9857, 218.9857, 218.9857, 
    218.9857, 218.9857, 218.9857, 218.9857, 218.9857, 218.9857, 218.9857, 
    218.9857, 218.9857, 218.9857, 218.9857, 218.9857, 218.9857, 218.9857, 
    218.9857, 218.9857, 218.9857, 218.9857, 218.9857, 218.9857, 218.9857, 
    218.9857, 218.9857, 218.9857, 218.9857, 218.9857, 218.9857, 218.9857, 
    218.9857, 218.9857, 218.9857, 218.9857, 218.9857, 218.9857, 218.9857, 
    218.9857, 218.9857, 218.9857, 218.9857, 218.9857, 218.9857,
  219.8047, 219.8047, 219.8047, 219.8047, 219.8047, 219.8047, 219.8047, 
    219.8047, 219.8047, 219.8047, 219.8047, 219.8047, 219.8047, 219.8047, 
    219.8047, 219.8047, 219.8047, 219.8047, 219.8047, 219.8047, 219.8047, 
    219.8047, 219.8047, 219.8047, 219.8047, 219.8047, 219.8047, 219.8047, 
    219.8047, 219.8047, 219.8047, 219.8047, 219.8047, 219.8047, 219.8047, 
    219.8047, 219.8047, 219.8047, 219.8047, 219.8047, 219.8047, 219.8047, 
    219.8047, 219.8047, 219.8047, 219.8047, 219.8047, 219.8047, 219.8047, 
    219.8047, 219.8047, 219.8047, 219.8047, 219.8047, 219.8047, 219.8047, 
    219.8047, 219.8047, 219.8047, 219.8047, 219.8047, 219.8047, 219.8047, 
    219.8047, 219.8047, 219.8047, 219.8047, 219.8047, 219.8047, 219.8047, 
    219.8047, 219.8047, 219.8047, 219.8047, 219.8047, 219.8047, 219.8047, 
    219.8047, 219.8047, 219.8047, 219.8047, 219.8047, 219.8047, 219.8047, 
    219.8047, 219.8047, 219.8047, 219.8047, 219.8047, 219.8047, 219.8047, 
    219.8047, 219.8047, 219.8047, 219.8047, 219.8047, 219.8047,
  220.6309, 220.6309, 220.6309, 220.6309, 220.6309, 220.6309, 220.6309, 
    220.6309, 220.6309, 220.6309, 220.6309, 220.6309, 220.6309, 220.6309, 
    220.6309, 220.6309, 220.6309, 220.6309, 220.6309, 220.6309, 220.6309, 
    220.6309, 220.6309, 220.6309, 220.6309, 220.6309, 220.6309, 220.6309, 
    220.6309, 220.6309, 220.6309, 220.6309, 220.6309, 220.6309, 220.6309, 
    220.6309, 220.6309, 220.6309, 220.6309, 220.6309, 220.6309, 220.6309, 
    220.6309, 220.6309, 220.6309, 220.6309, 220.6309, 220.6309, 220.6309, 
    220.6309, 220.6309, 220.6309, 220.6309, 220.6309, 220.6309, 220.6309, 
    220.6309, 220.6309, 220.6309, 220.6309, 220.6309, 220.6309, 220.6309, 
    220.6309, 220.6309, 220.6309, 220.6309, 220.6309, 220.6309, 220.6309, 
    220.6309, 220.6309, 220.6309, 220.6309, 220.6309, 220.6309, 220.6309, 
    220.6309, 220.6309, 220.6309, 220.6309, 220.6309, 220.6309, 220.6309, 
    220.6309, 220.6309, 220.6309, 220.6309, 220.6309, 220.6309, 220.6309, 
    220.6309, 220.6309, 220.6309, 220.6309, 220.6309, 220.6309,
  221.4646, 221.4646, 221.4646, 221.4646, 221.4646, 221.4646, 221.4646, 
    221.4646, 221.4646, 221.4646, 221.4646, 221.4646, 221.4646, 221.4646, 
    221.4646, 221.4646, 221.4646, 221.4646, 221.4646, 221.4646, 221.4646, 
    221.4646, 221.4646, 221.4646, 221.4646, 221.4646, 221.4646, 221.4646, 
    221.4646, 221.4646, 221.4646, 221.4646, 221.4646, 221.4646, 221.4646, 
    221.4646, 221.4646, 221.4646, 221.4646, 221.4646, 221.4646, 221.4646, 
    221.4646, 221.4646, 221.4646, 221.4646, 221.4646, 221.4646, 221.4646, 
    221.4646, 221.4646, 221.4646, 221.4646, 221.4646, 221.4646, 221.4646, 
    221.4646, 221.4646, 221.4646, 221.4646, 221.4646, 221.4646, 221.4646, 
    221.4646, 221.4646, 221.4646, 221.4646, 221.4646, 221.4646, 221.4646, 
    221.4646, 221.4646, 221.4646, 221.4646, 221.4646, 221.4646, 221.4646, 
    221.4646, 221.4646, 221.4646, 221.4646, 221.4646, 221.4646, 221.4646, 
    221.4646, 221.4646, 221.4646, 221.4646, 221.4646, 221.4646, 221.4646, 
    221.4646, 221.4646, 221.4646, 221.4646, 221.4646, 221.4646,
  222.3056, 222.3056, 222.3056, 222.3056, 222.3056, 222.3056, 222.3056, 
    222.3056, 222.3056, 222.3056, 222.3056, 222.3056, 222.3056, 222.3056, 
    222.3056, 222.3056, 222.3056, 222.3056, 222.3056, 222.3056, 222.3056, 
    222.3056, 222.3056, 222.3056, 222.3056, 222.3056, 222.3056, 222.3056, 
    222.3056, 222.3056, 222.3056, 222.3056, 222.3056, 222.3056, 222.3056, 
    222.3056, 222.3056, 222.3056, 222.3056, 222.3056, 222.3056, 222.3056, 
    222.3056, 222.3056, 222.3056, 222.3056, 222.3056, 222.3056, 222.3056, 
    222.3056, 222.3056, 222.3056, 222.3056, 222.3056, 222.3056, 222.3056, 
    222.3056, 222.3056, 222.3056, 222.3056, 222.3056, 222.3056, 222.3056, 
    222.3056, 222.3056, 222.3056, 222.3056, 222.3056, 222.3056, 222.3056, 
    222.3056, 222.3056, 222.3056, 222.3056, 222.3056, 222.3056, 222.3056, 
    222.3056, 222.3056, 222.3056, 222.3056, 222.3056, 222.3056, 222.3056, 
    222.3056, 222.3056, 222.3056, 222.3056, 222.3056, 222.3056, 222.3056, 
    222.3056, 222.3056, 222.3056, 222.3056, 222.3056, 222.3056,
  223.1541, 223.1541, 223.1541, 223.1541, 223.1541, 223.1541, 223.1541, 
    223.1541, 223.1541, 223.1541, 223.1541, 223.1541, 223.1541, 223.1541, 
    223.1541, 223.1541, 223.1541, 223.1541, 223.1541, 223.1541, 223.1541, 
    223.1541, 223.1541, 223.1541, 223.1541, 223.1541, 223.1541, 223.1541, 
    223.1541, 223.1541, 223.1541, 223.1541, 223.1541, 223.1541, 223.1541, 
    223.1541, 223.1541, 223.1541, 223.1541, 223.1541, 223.1541, 223.1541, 
    223.1541, 223.1541, 223.1541, 223.1541, 223.1541, 223.1541, 223.1541, 
    223.1541, 223.1541, 223.1541, 223.1541, 223.1541, 223.1541, 223.1541, 
    223.1541, 223.1541, 223.1541, 223.1541, 223.1541, 223.1541, 223.1541, 
    223.1541, 223.1541, 223.1541, 223.1541, 223.1541, 223.1541, 223.1541, 
    223.1541, 223.1541, 223.1541, 223.1541, 223.1541, 223.1541, 223.1541, 
    223.1541, 223.1541, 223.1541, 223.1541, 223.1541, 223.1541, 223.1541, 
    223.1541, 223.1541, 223.1541, 223.1541, 223.1541, 223.1541, 223.1541, 
    223.1541, 223.1541, 223.1541, 223.1541, 223.1541, 223.1541,
  224.01, 224.01, 224.01, 224.01, 224.01, 224.01, 224.01, 224.01, 224.01, 
    224.01, 224.01, 224.01, 224.01, 224.01, 224.01, 224.01, 224.01, 224.01, 
    224.01, 224.01, 224.01, 224.01, 224.01, 224.01, 224.01, 224.01, 224.01, 
    224.01, 224.01, 224.01, 224.01, 224.01, 224.01, 224.01, 224.01, 224.01, 
    224.01, 224.01, 224.01, 224.01, 224.01, 224.01, 224.01, 224.01, 224.01, 
    224.01, 224.01, 224.01, 224.01, 224.01, 224.01, 224.01, 224.01, 224.01, 
    224.01, 224.01, 224.01, 224.01, 224.01, 224.01, 224.01, 224.01, 224.01, 
    224.01, 224.01, 224.01, 224.01, 224.01, 224.01, 224.01, 224.01, 224.01, 
    224.01, 224.01, 224.01, 224.01, 224.01, 224.01, 224.01, 224.01, 224.01, 
    224.01, 224.01, 224.01, 224.01, 224.01, 224.01, 224.01, 224.01, 224.01, 
    224.01, 224.01, 224.01, 224.01, 224.01, 224.01, 224.01,
  224.8733, 224.8733, 224.8733, 224.8733, 224.8733, 224.8733, 224.8733, 
    224.8733, 224.8733, 224.8733, 224.8733, 224.8733, 224.8733, 224.8733, 
    224.8733, 224.8733, 224.8733, 224.8733, 224.8733, 224.8733, 224.8733, 
    224.8733, 224.8733, 224.8733, 224.8733, 224.8733, 224.8733, 224.8733, 
    224.8733, 224.8733, 224.8733, 224.8733, 224.8733, 224.8733, 224.8733, 
    224.8733, 224.8733, 224.8733, 224.8733, 224.8733, 224.8733, 224.8733, 
    224.8733, 224.8733, 224.8733, 224.8733, 224.8733, 224.8733, 224.8733, 
    224.8733, 224.8733, 224.8733, 224.8733, 224.8733, 224.8733, 224.8733, 
    224.8733, 224.8733, 224.8733, 224.8733, 224.8733, 224.8733, 224.8733, 
    224.8733, 224.8733, 224.8733, 224.8733, 224.8733, 224.8733, 224.8733, 
    224.8733, 224.8733, 224.8733, 224.8733, 224.8733, 224.8733, 224.8733, 
    224.8733, 224.8733, 224.8733, 224.8733, 224.8733, 224.8733, 224.8733, 
    224.8733, 224.8733, 224.8733, 224.8733, 224.8733, 224.8733, 224.8733, 
    224.8733, 224.8733, 224.8733, 224.8733, 224.8733, 224.8733,
  225.744, 225.744, 225.744, 225.744, 225.744, 225.744, 225.744, 225.744, 
    225.744, 225.744, 225.744, 225.744, 225.744, 225.744, 225.744, 225.744, 
    225.744, 225.744, 225.744, 225.744, 225.744, 225.744, 225.744, 225.744, 
    225.744, 225.744, 225.744, 225.744, 225.744, 225.744, 225.744, 225.744, 
    225.744, 225.744, 225.744, 225.744, 225.744, 225.744, 225.744, 225.744, 
    225.744, 225.744, 225.744, 225.744, 225.744, 225.744, 225.744, 225.744, 
    225.744, 225.744, 225.744, 225.744, 225.744, 225.744, 225.744, 225.744, 
    225.744, 225.744, 225.744, 225.744, 225.744, 225.744, 225.744, 225.744, 
    225.744, 225.744, 225.744, 225.744, 225.744, 225.744, 225.744, 225.744, 
    225.744, 225.744, 225.744, 225.744, 225.744, 225.744, 225.744, 225.744, 
    225.744, 225.744, 225.744, 225.744, 225.744, 225.744, 225.744, 225.744, 
    225.744, 225.744, 225.744, 225.744, 225.744, 225.744, 225.744, 225.744, 
    225.744,
  226.6221, 226.6221, 226.6221, 226.6221, 226.6221, 226.6221, 226.6221, 
    226.6221, 226.6221, 226.6221, 226.6221, 226.6221, 226.6221, 226.6221, 
    226.6221, 226.6221, 226.6221, 226.6221, 226.6221, 226.6221, 226.6221, 
    226.6221, 226.6221, 226.6221, 226.6221, 226.6221, 226.6221, 226.6221, 
    226.6221, 226.6221, 226.6221, 226.6221, 226.6221, 226.6221, 226.6221, 
    226.6221, 226.6221, 226.6221, 226.6221, 226.6221, 226.6221, 226.6221, 
    226.6221, 226.6221, 226.6221, 226.6221, 226.6221, 226.6221, 226.6221, 
    226.6221, 226.6221, 226.6221, 226.6221, 226.6221, 226.6221, 226.6221, 
    226.6221, 226.6221, 226.6221, 226.6221, 226.6221, 226.6221, 226.6221, 
    226.6221, 226.6221, 226.6221, 226.6221, 226.6221, 226.6221, 226.6221, 
    226.6221, 226.6221, 226.6221, 226.6221, 226.6221, 226.6221, 226.6221, 
    226.6221, 226.6221, 226.6221, 226.6221, 226.6221, 226.6221, 226.6221, 
    226.6221, 226.6221, 226.6221, 226.6221, 226.6221, 226.6221, 226.6221, 
    226.6221, 226.6221, 226.6221, 226.6221, 226.6221, 226.6221,
  227.5075, 227.5075, 227.5075, 227.5075, 227.5075, 227.5075, 227.5075, 
    227.5075, 227.5075, 227.5075, 227.5075, 227.5075, 227.5075, 227.5075, 
    227.5075, 227.5075, 227.5075, 227.5075, 227.5075, 227.5075, 227.5075, 
    227.5075, 227.5075, 227.5075, 227.5075, 227.5075, 227.5075, 227.5075, 
    227.5075, 227.5075, 227.5075, 227.5075, 227.5075, 227.5075, 227.5075, 
    227.5075, 227.5075, 227.5075, 227.5075, 227.5075, 227.5075, 227.5075, 
    227.5075, 227.5075, 227.5075, 227.5075, 227.5075, 227.5075, 227.5075, 
    227.5075, 227.5075, 227.5075, 227.5075, 227.5075, 227.5075, 227.5075, 
    227.5075, 227.5075, 227.5075, 227.5075, 227.5075, 227.5075, 227.5075, 
    227.5075, 227.5075, 227.5075, 227.5075, 227.5075, 227.5075, 227.5075, 
    227.5075, 227.5075, 227.5075, 227.5075, 227.5075, 227.5075, 227.5075, 
    227.5075, 227.5075, 227.5075, 227.5075, 227.5075, 227.5075, 227.5075, 
    227.5075, 227.5075, 227.5075, 227.5075, 227.5075, 227.5075, 227.5075, 
    227.5075, 227.5075, 227.5075, 227.5075, 227.5075, 227.5075,
  228.4002, 228.4002, 228.4002, 228.4002, 228.4002, 228.4002, 228.4002, 
    228.4002, 228.4002, 228.4002, 228.4002, 228.4002, 228.4002, 228.4002, 
    228.4002, 228.4002, 228.4002, 228.4002, 228.4002, 228.4002, 228.4002, 
    228.4002, 228.4002, 228.4002, 228.4002, 228.4002, 228.4002, 228.4002, 
    228.4002, 228.4002, 228.4002, 228.4002, 228.4002, 228.4002, 228.4002, 
    228.4002, 228.4002, 228.4002, 228.4002, 228.4002, 228.4002, 228.4002, 
    228.4002, 228.4002, 228.4002, 228.4002, 228.4002, 228.4002, 228.4002, 
    228.4002, 228.4002, 228.4002, 228.4002, 228.4002, 228.4002, 228.4002, 
    228.4002, 228.4002, 228.4002, 228.4002, 228.4002, 228.4002, 228.4002, 
    228.4002, 228.4002, 228.4002, 228.4002, 228.4002, 228.4002, 228.4002, 
    228.4002, 228.4002, 228.4002, 228.4002, 228.4002, 228.4002, 228.4002, 
    228.4002, 228.4002, 228.4002, 228.4002, 228.4002, 228.4002, 228.4002, 
    228.4002, 228.4002, 228.4002, 228.4002, 228.4002, 228.4002, 228.4002, 
    228.4002, 228.4002, 228.4002, 228.4002, 228.4002, 228.4002,
  229.3002, 229.3002, 229.3002, 229.3002, 229.3002, 229.3002, 229.3002, 
    229.3002, 229.3002, 229.3002, 229.3002, 229.3002, 229.3002, 229.3002, 
    229.3002, 229.3002, 229.3002, 229.3002, 229.3002, 229.3002, 229.3002, 
    229.3002, 229.3002, 229.3002, 229.3002, 229.3002, 229.3002, 229.3002, 
    229.3002, 229.3002, 229.3002, 229.3002, 229.3002, 229.3002, 229.3002, 
    229.3002, 229.3002, 229.3002, 229.3002, 229.3002, 229.3002, 229.3002, 
    229.3002, 229.3002, 229.3002, 229.3002, 229.3002, 229.3002, 229.3002, 
    229.3002, 229.3002, 229.3002, 229.3002, 229.3002, 229.3002, 229.3002, 
    229.3002, 229.3002, 229.3002, 229.3002, 229.3002, 229.3002, 229.3002, 
    229.3002, 229.3002, 229.3002, 229.3002, 229.3002, 229.3002, 229.3002, 
    229.3002, 229.3002, 229.3002, 229.3002, 229.3002, 229.3002, 229.3002, 
    229.3002, 229.3002, 229.3002, 229.3002, 229.3002, 229.3002, 229.3002, 
    229.3002, 229.3002, 229.3002, 229.3002, 229.3002, 229.3002, 229.3002, 
    229.3002, 229.3002, 229.3002, 229.3002, 229.3002, 229.3002,
  230.2074, 230.2074, 230.2074, 230.2074, 230.2074, 230.2074, 230.2074, 
    230.2074, 230.2074, 230.2074, 230.2074, 230.2074, 230.2074, 230.2074, 
    230.2074, 230.2074, 230.2074, 230.2074, 230.2074, 230.2074, 230.2074, 
    230.2074, 230.2074, 230.2074, 230.2074, 230.2074, 230.2074, 230.2074, 
    230.2074, 230.2074, 230.2074, 230.2074, 230.2074, 230.2074, 230.2074, 
    230.2074, 230.2074, 230.2074, 230.2074, 230.2074, 230.2074, 230.2074, 
    230.2074, 230.2074, 230.2074, 230.2074, 230.2074, 230.2074, 230.2074, 
    230.2074, 230.2074, 230.2074, 230.2074, 230.2074, 230.2074, 230.2074, 
    230.2074, 230.2074, 230.2074, 230.2074, 230.2074, 230.2074, 230.2074, 
    230.2074, 230.2074, 230.2074, 230.2074, 230.2074, 230.2074, 230.2074, 
    230.2074, 230.2074, 230.2074, 230.2074, 230.2074, 230.2074, 230.2074, 
    230.2074, 230.2074, 230.2074, 230.2074, 230.2074, 230.2074, 230.2074, 
    230.2074, 230.2074, 230.2074, 230.2074, 230.2074, 230.2074, 230.2074, 
    230.2074, 230.2074, 230.2074, 230.2074, 230.2074, 230.2074,
  231.1216, 231.1216, 231.1216, 231.1216, 231.1216, 231.1216, 231.1216, 
    231.1216, 231.1216, 231.1216, 231.1216, 231.1216, 231.1216, 231.1216, 
    231.1216, 231.1216, 231.1216, 231.1216, 231.1216, 231.1216, 231.1216, 
    231.1216, 231.1216, 231.1216, 231.1216, 231.1216, 231.1216, 231.1216, 
    231.1216, 231.1216, 231.1216, 231.1216, 231.1216, 231.1216, 231.1216, 
    231.1216, 231.1216, 231.1216, 231.1216, 231.1216, 231.1216, 231.1216, 
    231.1216, 231.1216, 231.1216, 231.1216, 231.1216, 231.1216, 231.1216, 
    231.1216, 231.1216, 231.1216, 231.1216, 231.1216, 231.1216, 231.1216, 
    231.1216, 231.1216, 231.1216, 231.1216, 231.1216, 231.1216, 231.1216, 
    231.1216, 231.1216, 231.1216, 231.1216, 231.1216, 231.1216, 231.1216, 
    231.1216, 231.1216, 231.1216, 231.1216, 231.1216, 231.1216, 231.1216, 
    231.1216, 231.1216, 231.1216, 231.1216, 231.1216, 231.1216, 231.1216, 
    231.1216, 231.1216, 231.1216, 231.1216, 231.1216, 231.1216, 231.1216, 
    231.1216, 231.1216, 231.1216, 231.1216, 231.1216, 231.1216,
  232.043, 232.043, 232.043, 232.043, 232.043, 232.043, 232.043, 232.043, 
    232.043, 232.043, 232.043, 232.043, 232.043, 232.043, 232.043, 232.043, 
    232.043, 232.043, 232.043, 232.043, 232.043, 232.043, 232.043, 232.043, 
    232.043, 232.043, 232.043, 232.043, 232.043, 232.043, 232.043, 232.043, 
    232.043, 232.043, 232.043, 232.043, 232.043, 232.043, 232.043, 232.043, 
    232.043, 232.043, 232.043, 232.043, 232.043, 232.043, 232.043, 232.043, 
    232.043, 232.043, 232.043, 232.043, 232.043, 232.043, 232.043, 232.043, 
    232.043, 232.043, 232.043, 232.043, 232.043, 232.043, 232.043, 232.043, 
    232.043, 232.043, 232.043, 232.043, 232.043, 232.043, 232.043, 232.043, 
    232.043, 232.043, 232.043, 232.043, 232.043, 232.043, 232.043, 232.043, 
    232.043, 232.043, 232.043, 232.043, 232.043, 232.043, 232.043, 232.043, 
    232.043, 232.043, 232.043, 232.043, 232.043, 232.043, 232.043, 232.043, 
    232.043,
  232.9712, 232.9712, 232.9712, 232.9712, 232.9712, 232.9712, 232.9712, 
    232.9712, 232.9712, 232.9712, 232.9712, 232.9712, 232.9712, 232.9712, 
    232.9712, 232.9712, 232.9712, 232.9712, 232.9712, 232.9712, 232.9712, 
    232.9712, 232.9712, 232.9712, 232.9712, 232.9712, 232.9712, 232.9712, 
    232.9712, 232.9712, 232.9712, 232.9712, 232.9712, 232.9712, 232.9712, 
    232.9712, 232.9712, 232.9712, 232.9712, 232.9712, 232.9712, 232.9712, 
    232.9712, 232.9712, 232.9712, 232.9712, 232.9712, 232.9712, 232.9712, 
    232.9712, 232.9712, 232.9712, 232.9712, 232.9712, 232.9712, 232.9712, 
    232.9712, 232.9712, 232.9712, 232.9712, 232.9712, 232.9712, 232.9712, 
    232.9712, 232.9712, 232.9712, 232.9712, 232.9712, 232.9712, 232.9712, 
    232.9712, 232.9712, 232.9712, 232.9712, 232.9712, 232.9712, 232.9712, 
    232.9712, 232.9712, 232.9712, 232.9712, 232.9712, 232.9712, 232.9712, 
    232.9712, 232.9712, 232.9712, 232.9712, 232.9712, 232.9712, 232.9712, 
    232.9712, 232.9712, 232.9712, 232.9712, 232.9712, 232.9712,
  233.9063, 233.9063, 233.9063, 233.9063, 233.9063, 233.9063, 233.9063, 
    233.9063, 233.9063, 233.9063, 233.9063, 233.9063, 233.9063, 233.9063, 
    233.9063, 233.9063, 233.9063, 233.9063, 233.9063, 233.9063, 233.9063, 
    233.9063, 233.9063, 233.9063, 233.9063, 233.9063, 233.9063, 233.9063, 
    233.9063, 233.9063, 233.9063, 233.9063, 233.9063, 233.9063, 233.9063, 
    233.9063, 233.9063, 233.9063, 233.9063, 233.9063, 233.9063, 233.9063, 
    233.9063, 233.9063, 233.9063, 233.9063, 233.9063, 233.9063, 233.9063, 
    233.9063, 233.9063, 233.9063, 233.9063, 233.9063, 233.9063, 233.9063, 
    233.9063, 233.9063, 233.9063, 233.9063, 233.9063, 233.9063, 233.9063, 
    233.9063, 233.9063, 233.9063, 233.9063, 233.9063, 233.9063, 233.9063, 
    233.9063, 233.9063, 233.9063, 233.9063, 233.9063, 233.9063, 233.9063, 
    233.9063, 233.9063, 233.9063, 233.9063, 233.9063, 233.9063, 233.9063, 
    233.9063, 233.9063, 233.9063, 233.9063, 233.9063, 233.9063, 233.9063, 
    233.9063, 233.9063, 233.9063, 233.9063, 233.9063, 233.9063,
  234.8482, 234.8482, 234.8482, 234.8482, 234.8482, 234.8482, 234.8482, 
    234.8482, 234.8482, 234.8482, 234.8482, 234.8482, 234.8482, 234.8482, 
    234.8482, 234.8482, 234.8482, 234.8482, 234.8482, 234.8482, 234.8482, 
    234.8482, 234.8482, 234.8482, 234.8482, 234.8482, 234.8482, 234.8482, 
    234.8482, 234.8482, 234.8482, 234.8482, 234.8482, 234.8482, 234.8482, 
    234.8482, 234.8482, 234.8482, 234.8482, 234.8482, 234.8482, 234.8482, 
    234.8482, 234.8482, 234.8482, 234.8482, 234.8482, 234.8482, 234.8482, 
    234.8482, 234.8482, 234.8482, 234.8482, 234.8482, 234.8482, 234.8482, 
    234.8482, 234.8482, 234.8482, 234.8482, 234.8482, 234.8482, 234.8482, 
    234.8482, 234.8482, 234.8482, 234.8482, 234.8482, 234.8482, 234.8482, 
    234.8482, 234.8482, 234.8482, 234.8482, 234.8482, 234.8482, 234.8482, 
    234.8482, 234.8482, 234.8482, 234.8482, 234.8482, 234.8482, 234.8482, 
    234.8482, 234.8482, 234.8482, 234.8482, 234.8482, 234.8482, 234.8482, 
    234.8482, 234.8482, 234.8482, 234.8482, 234.8482, 234.8482,
  235.7966, 235.7966, 235.7966, 235.7966, 235.7966, 235.7966, 235.7966, 
    235.7966, 235.7966, 235.7966, 235.7966, 235.7966, 235.7966, 235.7966, 
    235.7966, 235.7966, 235.7966, 235.7966, 235.7966, 235.7966, 235.7966, 
    235.7966, 235.7966, 235.7966, 235.7966, 235.7966, 235.7966, 235.7966, 
    235.7966, 235.7966, 235.7966, 235.7966, 235.7966, 235.7966, 235.7966, 
    235.7966, 235.7966, 235.7966, 235.7966, 235.7966, 235.7966, 235.7966, 
    235.7966, 235.7966, 235.7966, 235.7966, 235.7966, 235.7966, 235.7966, 
    235.7966, 235.7966, 235.7966, 235.7966, 235.7966, 235.7966, 235.7966, 
    235.7966, 235.7966, 235.7966, 235.7966, 235.7966, 235.7966, 235.7966, 
    235.7966, 235.7966, 235.7966, 235.7966, 235.7966, 235.7966, 235.7966, 
    235.7966, 235.7966, 235.7966, 235.7966, 235.7966, 235.7966, 235.7966, 
    235.7966, 235.7966, 235.7966, 235.7966, 235.7966, 235.7966, 235.7966, 
    235.7966, 235.7966, 235.7966, 235.7966, 235.7966, 235.7966, 235.7966, 
    235.7966, 235.7966, 235.7966, 235.7966, 235.7966, 235.7966,
  236.7514, 236.7514, 236.7514, 236.7514, 236.7514, 236.7514, 236.7514, 
    236.7514, 236.7514, 236.7514, 236.7514, 236.7514, 236.7514, 236.7514, 
    236.7514, 236.7514, 236.7514, 236.7514, 236.7514, 236.7514, 236.7514, 
    236.7514, 236.7514, 236.7514, 236.7514, 236.7514, 236.7514, 236.7514, 
    236.7514, 236.7514, 236.7514, 236.7514, 236.7514, 236.7514, 236.7514, 
    236.7514, 236.7514, 236.7514, 236.7514, 236.7514, 236.7514, 236.7514, 
    236.7514, 236.7514, 236.7514, 236.7514, 236.7514, 236.7514, 236.7514, 
    236.7514, 236.7514, 236.7514, 236.7514, 236.7514, 236.7514, 236.7514, 
    236.7514, 236.7514, 236.7514, 236.7514, 236.7514, 236.7514, 236.7514, 
    236.7514, 236.7514, 236.7514, 236.7514, 236.7514, 236.7514, 236.7514, 
    236.7514, 236.7514, 236.7514, 236.7514, 236.7514, 236.7514, 236.7514, 
    236.7514, 236.7514, 236.7514, 236.7514, 236.7514, 236.7514, 236.7514, 
    236.7514, 236.7514, 236.7514, 236.7514, 236.7514, 236.7514, 236.7514, 
    236.7514, 236.7514, 236.7514, 236.7514, 236.7514, 236.7514,
  237.7126, 237.7126, 237.7126, 237.7126, 237.7126, 237.7126, 237.7126, 
    237.7126, 237.7126, 237.7126, 237.7126, 237.7126, 237.7126, 237.7126, 
    237.7126, 237.7126, 237.7126, 237.7126, 237.7126, 237.7126, 237.7126, 
    237.7126, 237.7126, 237.7126, 237.7126, 237.7126, 237.7126, 237.7126, 
    237.7126, 237.7126, 237.7126, 237.7126, 237.7126, 237.7126, 237.7126, 
    237.7126, 237.7126, 237.7126, 237.7126, 237.7126, 237.7126, 237.7126, 
    237.7126, 237.7126, 237.7126, 237.7126, 237.7126, 237.7126, 237.7126, 
    237.7126, 237.7126, 237.7126, 237.7126, 237.7126, 237.7126, 237.7126, 
    237.7126, 237.7126, 237.7126, 237.7126, 237.7126, 237.7126, 237.7126, 
    237.7126, 237.7126, 237.7126, 237.7126, 237.7126, 237.7126, 237.7126, 
    237.7126, 237.7126, 237.7126, 237.7126, 237.7126, 237.7126, 237.7126, 
    237.7126, 237.7126, 237.7126, 237.7126, 237.7126, 237.7126, 237.7126, 
    237.7126, 237.7126, 237.7126, 237.7126, 237.7126, 237.7126, 237.7126, 
    237.7126, 237.7126, 237.7126, 237.7126, 237.7126, 237.7126,
  238.6799, 238.6799, 238.6799, 238.6799, 238.6799, 238.6799, 238.6799, 
    238.6799, 238.6799, 238.6799, 238.6799, 238.6799, 238.6799, 238.6799, 
    238.6799, 238.6799, 238.6799, 238.6799, 238.6799, 238.6799, 238.6799, 
    238.6799, 238.6799, 238.6799, 238.6799, 238.6799, 238.6799, 238.6799, 
    238.6799, 238.6799, 238.6799, 238.6799, 238.6799, 238.6799, 238.6799, 
    238.6799, 238.6799, 238.6799, 238.6799, 238.6799, 238.6799, 238.6799, 
    238.6799, 238.6799, 238.6799, 238.6799, 238.6799, 238.6799, 238.6799, 
    238.6799, 238.6799, 238.6799, 238.6799, 238.6799, 238.6799, 238.6799, 
    238.6799, 238.6799, 238.6799, 238.6799, 238.6799, 238.6799, 238.6799, 
    238.6799, 238.6799, 238.6799, 238.6799, 238.6799, 238.6799, 238.6799, 
    238.6799, 238.6799, 238.6799, 238.6799, 238.6799, 238.6799, 238.6799, 
    238.6799, 238.6799, 238.6799, 238.6799, 238.6799, 238.6799, 238.6799, 
    238.6799, 238.6799, 238.6799, 238.6799, 238.6799, 238.6799, 238.6799, 
    238.6799, 238.6799, 238.6799, 238.6799, 238.6799, 238.6799,
  239.6532, 239.6532, 239.6532, 239.6532, 239.6532, 239.6532, 239.6532, 
    239.6532, 239.6532, 239.6532, 239.6532, 239.6532, 239.6532, 239.6532, 
    239.6532, 239.6532, 239.6532, 239.6532, 239.6532, 239.6532, 239.6532, 
    239.6532, 239.6532, 239.6532, 239.6532, 239.6532, 239.6532, 239.6532, 
    239.6532, 239.6532, 239.6532, 239.6532, 239.6532, 239.6532, 239.6532, 
    239.6532, 239.6532, 239.6532, 239.6532, 239.6532, 239.6532, 239.6532, 
    239.6532, 239.6532, 239.6532, 239.6532, 239.6532, 239.6532, 239.6532, 
    239.6532, 239.6532, 239.6532, 239.6532, 239.6532, 239.6532, 239.6532, 
    239.6532, 239.6532, 239.6532, 239.6532, 239.6532, 239.6532, 239.6532, 
    239.6532, 239.6532, 239.6532, 239.6532, 239.6532, 239.6532, 239.6532, 
    239.6532, 239.6532, 239.6532, 239.6532, 239.6532, 239.6532, 239.6532, 
    239.6532, 239.6532, 239.6532, 239.6532, 239.6532, 239.6532, 239.6532, 
    239.6532, 239.6532, 239.6532, 239.6532, 239.6532, 239.6532, 239.6532, 
    239.6532, 239.6532, 239.6532, 239.6532, 239.6532, 239.6532,
  240.6322, 240.6322, 240.6322, 240.6322, 240.6322, 240.6322, 240.6322, 
    240.6322, 240.6322, 240.6322, 240.6322, 240.6322, 240.6322, 240.6322, 
    240.6322, 240.6322, 240.6322, 240.6322, 240.6322, 240.6322, 240.6322, 
    240.6322, 240.6322, 240.6322, 240.6322, 240.6322, 240.6322, 240.6322, 
    240.6322, 240.6322, 240.6322, 240.6322, 240.6322, 240.6322, 240.6322, 
    240.6322, 240.6322, 240.6322, 240.6322, 240.6322, 240.6322, 240.6322, 
    240.6322, 240.6322, 240.6322, 240.6322, 240.6322, 240.6322, 240.6322, 
    240.6322, 240.6322, 240.6322, 240.6322, 240.6322, 240.6322, 240.6322, 
    240.6322, 240.6322, 240.6322, 240.6322, 240.6322, 240.6322, 240.6322, 
    240.6322, 240.6322, 240.6322, 240.6322, 240.6322, 240.6322, 240.6322, 
    240.6322, 240.6322, 240.6322, 240.6322, 240.6322, 240.6322, 240.6322, 
    240.6322, 240.6322, 240.6322, 240.6322, 240.6322, 240.6322, 240.6322, 
    240.6322, 240.6322, 240.6322, 240.6322, 240.6322, 240.6322, 240.6322, 
    240.6322, 240.6322, 240.6322, 240.6322, 240.6322, 240.6322,
  241.6168, 241.6168, 241.6168, 241.6168, 241.6168, 241.6168, 241.6168, 
    241.6168, 241.6168, 241.6168, 241.6168, 241.6168, 241.6168, 241.6168, 
    241.6168, 241.6168, 241.6168, 241.6168, 241.6168, 241.6168, 241.6168, 
    241.6168, 241.6168, 241.6168, 241.6168, 241.6168, 241.6168, 241.6168, 
    241.6168, 241.6168, 241.6168, 241.6168, 241.6168, 241.6168, 241.6168, 
    241.6168, 241.6168, 241.6168, 241.6168, 241.6168, 241.6168, 241.6168, 
    241.6168, 241.6168, 241.6168, 241.6168, 241.6168, 241.6168, 241.6168, 
    241.6168, 241.6168, 241.6168, 241.6168, 241.6168, 241.6168, 241.6168, 
    241.6168, 241.6168, 241.6168, 241.6168, 241.6168, 241.6168, 241.6168, 
    241.6168, 241.6168, 241.6168, 241.6168, 241.6168, 241.6168, 241.6168, 
    241.6168, 241.6168, 241.6168, 241.6168, 241.6168, 241.6168, 241.6168, 
    241.6168, 241.6168, 241.6168, 241.6168, 241.6168, 241.6168, 241.6168, 
    241.6168, 241.6168, 241.6168, 241.6168, 241.6168, 241.6168, 241.6168, 
    241.6168, 241.6168, 241.6168, 241.6168, 241.6168, 241.6168,
  242.6068, 242.6068, 242.6068, 242.6068, 242.6068, 242.6068, 242.6068, 
    242.6068, 242.6068, 242.6068, 242.6068, 242.6068, 242.6068, 242.6068, 
    242.6068, 242.6068, 242.6068, 242.6068, 242.6068, 242.6068, 242.6068, 
    242.6068, 242.6068, 242.6068, 242.6068, 242.6068, 242.6068, 242.6068, 
    242.6068, 242.6068, 242.6068, 242.6068, 242.6068, 242.6068, 242.6068, 
    242.6068, 242.6068, 242.6068, 242.6068, 242.6068, 242.6068, 242.6068, 
    242.6068, 242.6068, 242.6068, 242.6068, 242.6068, 242.6068, 242.6068, 
    242.6068, 242.6068, 242.6068, 242.6068, 242.6068, 242.6068, 242.6068, 
    242.6068, 242.6068, 242.6068, 242.6068, 242.6068, 242.6068, 242.6068, 
    242.6068, 242.6068, 242.6068, 242.6068, 242.6068, 242.6068, 242.6068, 
    242.6068, 242.6068, 242.6068, 242.6068, 242.6068, 242.6068, 242.6068, 
    242.6068, 242.6068, 242.6068, 242.6068, 242.6068, 242.6068, 242.6068, 
    242.6068, 242.6068, 242.6068, 242.6068, 242.6068, 242.6068, 242.6068, 
    242.6068, 242.6068, 242.6068, 242.6068, 242.6068, 242.6068,
  243.6019, 243.6019, 243.6019, 243.6019, 243.6019, 243.6019, 243.6019, 
    243.6019, 243.6019, 243.6019, 243.6019, 243.6019, 243.6019, 243.6019, 
    243.6019, 243.6019, 243.6019, 243.6019, 243.6019, 243.6019, 243.6019, 
    243.6019, 243.6019, 243.6019, 243.6019, 243.6019, 243.6019, 243.6019, 
    243.6019, 243.6019, 243.6019, 243.6019, 243.6019, 243.6019, 243.6019, 
    243.6019, 243.6019, 243.6019, 243.6019, 243.6019, 243.6019, 243.6019, 
    243.6019, 243.6019, 243.6019, 243.6019, 243.6019, 243.6019, 243.6019, 
    243.6019, 243.6019, 243.6019, 243.6019, 243.6019, 243.6019, 243.6019, 
    243.6019, 243.6019, 243.6019, 243.6019, 243.6019, 243.6019, 243.6019, 
    243.6019, 243.6019, 243.6019, 243.6019, 243.6019, 243.6019, 243.6019, 
    243.6019, 243.6019, 243.6019, 243.6019, 243.6019, 243.6019, 243.6019, 
    243.6019, 243.6019, 243.6019, 243.6019, 243.6019, 243.6019, 243.6019, 
    243.6019, 243.6019, 243.6019, 243.6019, 243.6019, 243.6019, 243.6019, 
    243.6019, 243.6019, 243.6019, 243.6019, 243.6019, 243.6019,
  244.6019, 244.6019, 244.6019, 244.6019, 244.6019, 244.6019, 244.6019, 
    244.6019, 244.6019, 244.6019, 244.6019, 244.6019, 244.6019, 244.6019, 
    244.6019, 244.6019, 244.6019, 244.6019, 244.6019, 244.6019, 244.6019, 
    244.6019, 244.6019, 244.6019, 244.6019, 244.6019, 244.6019, 244.6019, 
    244.6019, 244.6019, 244.6019, 244.6019, 244.6019, 244.6019, 244.6019, 
    244.6019, 244.6019, 244.6019, 244.6019, 244.6019, 244.6019, 244.6019, 
    244.6019, 244.6019, 244.6019, 244.6019, 244.6019, 244.6019, 244.6019, 
    244.6019, 244.6019, 244.6019, 244.6019, 244.6019, 244.6019, 244.6019, 
    244.6019, 244.6019, 244.6019, 244.6019, 244.6019, 244.6019, 244.6019, 
    244.6019, 244.6019, 244.6019, 244.6019, 244.6019, 244.6019, 244.6019, 
    244.6019, 244.6019, 244.6019, 244.6019, 244.6019, 244.6019, 244.6019, 
    244.6019, 244.6019, 244.6019, 244.6019, 244.6019, 244.6019, 244.6019, 
    244.6019, 244.6019, 244.6019, 244.6019, 244.6019, 244.6019, 244.6019, 
    244.6019, 244.6019, 244.6019, 244.6019, 244.6019, 244.6019,
  245.6065, 245.6065, 245.6065, 245.6065, 245.6065, 245.6065, 245.6065, 
    245.6065, 245.6065, 245.6065, 245.6065, 245.6065, 245.6065, 245.6065, 
    245.6065, 245.6065, 245.6065, 245.6065, 245.6065, 245.6065, 245.6065, 
    245.6065, 245.6065, 245.6065, 245.6065, 245.6065, 245.6065, 245.6065, 
    245.6065, 245.6065, 245.6065, 245.6065, 245.6065, 245.6065, 245.6065, 
    245.6065, 245.6065, 245.6065, 245.6065, 245.6065, 245.6065, 245.6065, 
    245.6065, 245.6065, 245.6065, 245.6065, 245.6065, 245.6065, 245.6065, 
    245.6065, 245.6065, 245.6065, 245.6065, 245.6065, 245.6065, 245.6065, 
    245.6065, 245.6065, 245.6065, 245.6065, 245.6065, 245.6065, 245.6065, 
    245.6065, 245.6065, 245.6065, 245.6065, 245.6065, 245.6065, 245.6065, 
    245.6065, 245.6065, 245.6065, 245.6065, 245.6065, 245.6065, 245.6065, 
    245.6065, 245.6065, 245.6065, 245.6065, 245.6065, 245.6065, 245.6065, 
    245.6065, 245.6065, 245.6065, 245.6065, 245.6065, 245.6065, 245.6065, 
    245.6065, 245.6065, 245.6065, 245.6065, 245.6065, 245.6065,
  246.6156, 246.6156, 246.6156, 246.6156, 246.6156, 246.6156, 246.6156, 
    246.6156, 246.6156, 246.6156, 246.6156, 246.6156, 246.6156, 246.6156, 
    246.6156, 246.6156, 246.6156, 246.6156, 246.6156, 246.6156, 246.6156, 
    246.6156, 246.6156, 246.6156, 246.6156, 246.6156, 246.6156, 246.6156, 
    246.6156, 246.6156, 246.6156, 246.6156, 246.6156, 246.6156, 246.6156, 
    246.6156, 246.6156, 246.6156, 246.6156, 246.6156, 246.6156, 246.6156, 
    246.6156, 246.6156, 246.6156, 246.6156, 246.6156, 246.6156, 246.6156, 
    246.6156, 246.6156, 246.6156, 246.6156, 246.6156, 246.6156, 246.6156, 
    246.6156, 246.6156, 246.6156, 246.6156, 246.6156, 246.6156, 246.6156, 
    246.6156, 246.6156, 246.6156, 246.6156, 246.6156, 246.6156, 246.6156, 
    246.6156, 246.6156, 246.6156, 246.6156, 246.6156, 246.6156, 246.6156, 
    246.6156, 246.6156, 246.6156, 246.6156, 246.6156, 246.6156, 246.6156, 
    246.6156, 246.6156, 246.6156, 246.6156, 246.6156, 246.6156, 246.6156, 
    246.6156, 246.6156, 246.6156, 246.6156, 246.6156, 246.6156,
  247.6287, 247.6287, 247.6287, 247.6287, 247.6287, 247.6287, 247.6287, 
    247.6287, 247.6287, 247.6287, 247.6287, 247.6287, 247.6287, 247.6287, 
    247.6287, 247.6287, 247.6287, 247.6287, 247.6287, 247.6287, 247.6287, 
    247.6287, 247.6287, 247.6287, 247.6287, 247.6287, 247.6287, 247.6287, 
    247.6287, 247.6287, 247.6287, 247.6287, 247.6287, 247.6287, 247.6287, 
    247.6287, 247.6287, 247.6287, 247.6287, 247.6287, 247.6287, 247.6287, 
    247.6287, 247.6287, 247.6287, 247.6287, 247.6287, 247.6287, 247.6287, 
    247.6287, 247.6287, 247.6287, 247.6287, 247.6287, 247.6287, 247.6287, 
    247.6287, 247.6287, 247.6287, 247.6287, 247.6287, 247.6287, 247.6287, 
    247.6287, 247.6287, 247.6287, 247.6287, 247.6287, 247.6287, 247.6287, 
    247.6287, 247.6287, 247.6287, 247.6287, 247.6287, 247.6287, 247.6287, 
    247.6287, 247.6287, 247.6287, 247.6287, 247.6287, 247.6287, 247.6287, 
    247.6287, 247.6287, 247.6287, 247.6287, 247.6287, 247.6287, 247.6287, 
    247.6287, 247.6287, 247.6287, 247.6287, 247.6287, 247.6287,
  248.6458, 248.6458, 248.6458, 248.6458, 248.6458, 248.6458, 248.6458, 
    248.6458, 248.6458, 248.6458, 248.6458, 248.6458, 248.6458, 248.6458, 
    248.6458, 248.6458, 248.6458, 248.6458, 248.6458, 248.6458, 248.6458, 
    248.6458, 248.6458, 248.6458, 248.6458, 248.6458, 248.6458, 248.6458, 
    248.6458, 248.6458, 248.6458, 248.6458, 248.6458, 248.6458, 248.6458, 
    248.6458, 248.6458, 248.6458, 248.6458, 248.6458, 248.6458, 248.6458, 
    248.6458, 248.6458, 248.6458, 248.6458, 248.6458, 248.6458, 248.6458, 
    248.6458, 248.6458, 248.6458, 248.6458, 248.6458, 248.6458, 248.6458, 
    248.6458, 248.6458, 248.6458, 248.6458, 248.6458, 248.6458, 248.6458, 
    248.6458, 248.6458, 248.6458, 248.6458, 248.6458, 248.6458, 248.6458, 
    248.6458, 248.6458, 248.6458, 248.6458, 248.6458, 248.6458, 248.6458, 
    248.6458, 248.6458, 248.6458, 248.6458, 248.6458, 248.6458, 248.6458, 
    248.6458, 248.6458, 248.6458, 248.6458, 248.6458, 248.6458, 248.6458, 
    248.6458, 248.6458, 248.6458, 248.6458, 248.6458, 248.6458,
  249.6663, 249.6663, 249.6663, 249.6663, 249.6663, 249.6663, 249.6663, 
    249.6663, 249.6663, 249.6663, 249.6663, 249.6663, 249.6663, 249.6663, 
    249.6663, 249.6663, 249.6663, 249.6663, 249.6663, 249.6663, 249.6663, 
    249.6663, 249.6663, 249.6663, 249.6663, 249.6663, 249.6663, 249.6663, 
    249.6663, 249.6663, 249.6663, 249.6663, 249.6663, 249.6663, 249.6663, 
    249.6663, 249.6663, 249.6663, 249.6663, 249.6663, 249.6663, 249.6663, 
    249.6663, 249.6663, 249.6663, 249.6663, 249.6663, 249.6663, 249.6663, 
    249.6663, 249.6663, 249.6663, 249.6663, 249.6663, 249.6663, 249.6663, 
    249.6663, 249.6663, 249.6663, 249.6663, 249.6663, 249.6663, 249.6663, 
    249.6663, 249.6663, 249.6663, 249.6663, 249.6663, 249.6663, 249.6663, 
    249.6663, 249.6663, 249.6663, 249.6663, 249.6663, 249.6663, 249.6663, 
    249.6663, 249.6663, 249.6663, 249.6663, 249.6663, 249.6663, 249.6663, 
    249.6663, 249.6663, 249.6663, 249.6663, 249.6663, 249.6663, 249.6663, 
    249.6663, 249.6663, 249.6663, 249.6663, 249.6663, 249.6663,
  250.6902, 250.6902, 250.6902, 250.6902, 250.6902, 250.6902, 250.6902, 
    250.6902, 250.6902, 250.6902, 250.6902, 250.6902, 250.6902, 250.6902, 
    250.6902, 250.6902, 250.6902, 250.6902, 250.6902, 250.6902, 250.6902, 
    250.6902, 250.6902, 250.6902, 250.6902, 250.6902, 250.6902, 250.6902, 
    250.6902, 250.6902, 250.6902, 250.6902, 250.6902, 250.6902, 250.6902, 
    250.6902, 250.6902, 250.6902, 250.6902, 250.6902, 250.6902, 250.6902, 
    250.6902, 250.6902, 250.6902, 250.6902, 250.6902, 250.6902, 250.6902, 
    250.6902, 250.6902, 250.6902, 250.6902, 250.6902, 250.6902, 250.6902, 
    250.6902, 250.6902, 250.6902, 250.6902, 250.6902, 250.6902, 250.6902, 
    250.6902, 250.6902, 250.6902, 250.6902, 250.6902, 250.6902, 250.6902, 
    250.6902, 250.6902, 250.6902, 250.6902, 250.6902, 250.6902, 250.6902, 
    250.6902, 250.6902, 250.6902, 250.6902, 250.6902, 250.6902, 250.6902, 
    250.6902, 250.6902, 250.6902, 250.6902, 250.6902, 250.6902, 250.6902, 
    250.6902, 250.6902, 250.6902, 250.6902, 250.6902, 250.6902,
  251.717, 251.717, 251.717, 251.717, 251.717, 251.717, 251.717, 251.717, 
    251.717, 251.717, 251.717, 251.717, 251.717, 251.717, 251.717, 251.717, 
    251.717, 251.717, 251.717, 251.717, 251.717, 251.717, 251.717, 251.717, 
    251.717, 251.717, 251.717, 251.717, 251.717, 251.717, 251.717, 251.717, 
    251.717, 251.717, 251.717, 251.717, 251.717, 251.717, 251.717, 251.717, 
    251.717, 251.717, 251.717, 251.717, 251.717, 251.717, 251.717, 251.717, 
    251.717, 251.717, 251.717, 251.717, 251.717, 251.717, 251.717, 251.717, 
    251.717, 251.717, 251.717, 251.717, 251.717, 251.717, 251.717, 251.717, 
    251.717, 251.717, 251.717, 251.717, 251.717, 251.717, 251.717, 251.717, 
    251.717, 251.717, 251.717, 251.717, 251.717, 251.717, 251.717, 251.717, 
    251.717, 251.717, 251.717, 251.717, 251.717, 251.717, 251.717, 251.717, 
    251.717, 251.717, 251.717, 251.717, 251.717, 251.717, 251.717, 251.717, 
    251.717,
  252.7465, 252.7465, 252.7465, 252.7465, 252.7465, 252.7465, 252.7465, 
    252.7465, 252.7465, 252.7465, 252.7465, 252.7465, 252.7465, 252.7465, 
    252.7465, 252.7465, 252.7465, 252.7465, 252.7465, 252.7465, 252.7465, 
    252.7465, 252.7465, 252.7465, 252.7465, 252.7465, 252.7465, 252.7465, 
    252.7465, 252.7465, 252.7465, 252.7465, 252.7465, 252.7465, 252.7465, 
    252.7465, 252.7465, 252.7465, 252.7465, 252.7465, 252.7465, 252.7465, 
    252.7465, 252.7465, 252.7465, 252.7465, 252.7465, 252.7465, 252.7465, 
    252.7465, 252.7465, 252.7465, 252.7465, 252.7465, 252.7465, 252.7465, 
    252.7465, 252.7465, 252.7465, 252.7465, 252.7465, 252.7465, 252.7465, 
    252.7465, 252.7465, 252.7465, 252.7465, 252.7465, 252.7465, 252.7465, 
    252.7465, 252.7465, 252.7465, 252.7465, 252.7465, 252.7465, 252.7465, 
    252.7465, 252.7465, 252.7465, 252.7465, 252.7465, 252.7465, 252.7465, 
    252.7465, 252.7465, 252.7465, 252.7465, 252.7465, 252.7465, 252.7465, 
    252.7465, 252.7465, 252.7465, 252.7465, 252.7465, 252.7465,
  253.7783, 253.7783, 253.7783, 253.7783, 253.7783, 253.7783, 253.7783, 
    253.7783, 253.7783, 253.7783, 253.7783, 253.7783, 253.7783, 253.7783, 
    253.7783, 253.7783, 253.7783, 253.7783, 253.7783, 253.7783, 253.7783, 
    253.7783, 253.7783, 253.7783, 253.7783, 253.7783, 253.7783, 253.7783, 
    253.7783, 253.7783, 253.7783, 253.7783, 253.7783, 253.7783, 253.7783, 
    253.7783, 253.7783, 253.7783, 253.7783, 253.7783, 253.7783, 253.7783, 
    253.7783, 253.7783, 253.7783, 253.7783, 253.7783, 253.7783, 253.7783, 
    253.7783, 253.7783, 253.7783, 253.7783, 253.7783, 253.7783, 253.7783, 
    253.7783, 253.7783, 253.7783, 253.7783, 253.7783, 253.7783, 253.7783, 
    253.7783, 253.7783, 253.7783, 253.7783, 253.7783, 253.7783, 253.7783, 
    253.7783, 253.7783, 253.7783, 253.7783, 253.7783, 253.7783, 253.7783, 
    253.7783, 253.7783, 253.7783, 253.7783, 253.7783, 253.7783, 253.7783, 
    253.7783, 253.7783, 253.7783, 253.7783, 253.7783, 253.7783, 253.7783, 
    253.7783, 253.7783, 253.7783, 253.7783, 253.7783, 253.7783,
  254.8122, 254.8122, 254.8122, 254.8122, 254.8122, 254.8122, 254.8122, 
    254.8122, 254.8122, 254.8122, 254.8122, 254.8122, 254.8122, 254.8122, 
    254.8122, 254.8122, 254.8122, 254.8122, 254.8122, 254.8122, 254.8122, 
    254.8122, 254.8122, 254.8122, 254.8122, 254.8122, 254.8122, 254.8122, 
    254.8122, 254.8122, 254.8122, 254.8122, 254.8122, 254.8122, 254.8122, 
    254.8122, 254.8122, 254.8122, 254.8122, 254.8122, 254.8122, 254.8122, 
    254.8122, 254.8122, 254.8122, 254.8122, 254.8122, 254.8122, 254.8122, 
    254.8122, 254.8122, 254.8122, 254.8122, 254.8122, 254.8122, 254.8122, 
    254.8122, 254.8122, 254.8122, 254.8122, 254.8122, 254.8122, 254.8122, 
    254.8122, 254.8122, 254.8122, 254.8122, 254.8122, 254.8122, 254.8122, 
    254.8122, 254.8122, 254.8122, 254.8122, 254.8122, 254.8122, 254.8122, 
    254.8122, 254.8122, 254.8122, 254.8122, 254.8122, 254.8122, 254.8122, 
    254.8122, 254.8122, 254.8122, 254.8122, 254.8122, 254.8122, 254.8122, 
    254.8122, 254.8122, 254.8122, 254.8122, 254.8122, 254.8122,
  255.8477, 255.8477, 255.8477, 255.8477, 255.8477, 255.8477, 255.8477, 
    255.8477, 255.8477, 255.8477, 255.8477, 255.8477, 255.8477, 255.8477, 
    255.8477, 255.8477, 255.8477, 255.8477, 255.8477, 255.8477, 255.8477, 
    255.8477, 255.8477, 255.8477, 255.8477, 255.8477, 255.8477, 255.8477, 
    255.8477, 255.8477, 255.8477, 255.8477, 255.8477, 255.8477, 255.8477, 
    255.8477, 255.8477, 255.8477, 255.8477, 255.8477, 255.8477, 255.8477, 
    255.8477, 255.8477, 255.8477, 255.8477, 255.8477, 255.8477, 255.8477, 
    255.8477, 255.8477, 255.8477, 255.8477, 255.8477, 255.8477, 255.8477, 
    255.8477, 255.8477, 255.8477, 255.8477, 255.8477, 255.8477, 255.8477, 
    255.8477, 255.8477, 255.8477, 255.8477, 255.8477, 255.8477, 255.8477, 
    255.8477, 255.8477, 255.8477, 255.8477, 255.8477, 255.8477, 255.8477, 
    255.8477, 255.8477, 255.8477, 255.8477, 255.8477, 255.8477, 255.8477, 
    255.8477, 255.8477, 255.8477, 255.8477, 255.8477, 255.8477, 255.8477, 
    255.8477, 255.8477, 255.8477, 255.8477, 255.8477, 255.8477,
  256.8846, 256.8846, 256.8846, 256.8846, 256.8846, 256.8846, 256.8846, 
    256.8846, 256.8846, 256.8846, 256.8846, 256.8846, 256.8846, 256.8846, 
    256.8846, 256.8846, 256.8846, 256.8846, 256.8846, 256.8846, 256.8846, 
    256.8846, 256.8846, 256.8846, 256.8846, 256.8846, 256.8846, 256.8846, 
    256.8846, 256.8846, 256.8846, 256.8846, 256.8846, 256.8846, 256.8846, 
    256.8846, 256.8846, 256.8846, 256.8846, 256.8846, 256.8846, 256.8846, 
    256.8846, 256.8846, 256.8846, 256.8846, 256.8846, 256.8846, 256.8846, 
    256.8846, 256.8846, 256.8846, 256.8846, 256.8846, 256.8846, 256.8846, 
    256.8846, 256.8846, 256.8846, 256.8846, 256.8846, 256.8846, 256.8846, 
    256.8846, 256.8846, 256.8846, 256.8846, 256.8846, 256.8846, 256.8846, 
    256.8846, 256.8846, 256.8846, 256.8846, 256.8846, 256.8846, 256.8846, 
    256.8846, 256.8846, 256.8846, 256.8846, 256.8846, 256.8846, 256.8846, 
    256.8846, 256.8846, 256.8846, 256.8846, 256.8846, 256.8846, 256.8846, 
    256.8846, 256.8846, 256.8846, 256.8846, 256.8846, 256.8846,
  257.9225, 257.9225, 257.9225, 257.9225, 257.9225, 257.9225, 257.9225, 
    257.9225, 257.9225, 257.9225, 257.9225, 257.9225, 257.9225, 257.9225, 
    257.9225, 257.9225, 257.9225, 257.9225, 257.9225, 257.9225, 257.9225, 
    257.9225, 257.9225, 257.9225, 257.9225, 257.9225, 257.9225, 257.9225, 
    257.9225, 257.9225, 257.9225, 257.9225, 257.9225, 257.9225, 257.9225, 
    257.9225, 257.9225, 257.9225, 257.9225, 257.9225, 257.9225, 257.9225, 
    257.9225, 257.9225, 257.9225, 257.9225, 257.9225, 257.9225, 257.9225, 
    257.9225, 257.9225, 257.9225, 257.9225, 257.9225, 257.9225, 257.9225, 
    257.9225, 257.9225, 257.9225, 257.9225, 257.9225, 257.9225, 257.9225, 
    257.9225, 257.9225, 257.9225, 257.9225, 257.9225, 257.9225, 257.9225, 
    257.9225, 257.9225, 257.9225, 257.9225, 257.9225, 257.9225, 257.9225, 
    257.9225, 257.9225, 257.9225, 257.9225, 257.9225, 257.9225, 257.9225, 
    257.9225, 257.9225, 257.9225, 257.9225, 257.9225, 257.9225, 257.9225, 
    257.9225, 257.9225, 257.9225, 257.9225, 257.9225, 257.9225,
  258.9611, 258.9611, 258.9611, 258.9611, 258.9611, 258.9611, 258.9611, 
    258.9611, 258.9611, 258.9611, 258.9611, 258.9611, 258.9611, 258.9611, 
    258.9611, 258.9611, 258.9611, 258.9611, 258.9611, 258.9611, 258.9611, 
    258.9611, 258.9611, 258.9611, 258.9611, 258.9611, 258.9611, 258.9611, 
    258.9611, 258.9611, 258.9611, 258.9611, 258.9611, 258.9611, 258.9611, 
    258.9611, 258.9611, 258.9611, 258.9611, 258.9611, 258.9611, 258.9611, 
    258.9611, 258.9611, 258.9611, 258.9611, 258.9611, 258.9611, 258.9611, 
    258.9611, 258.9611, 258.9611, 258.9611, 258.9611, 258.9611, 258.9611, 
    258.9611, 258.9611, 258.9611, 258.9611, 258.9611, 258.9611, 258.9611, 
    258.9611, 258.9611, 258.9611, 258.9611, 258.9611, 258.9611, 258.9611, 
    258.9611, 258.9611, 258.9611, 258.9611, 258.9611, 258.9611, 258.9611, 
    258.9611, 258.9611, 258.9611, 258.9611, 258.9611, 258.9611, 258.9611, 
    258.9611, 258.9611, 258.9611, 258.9611, 258.9611, 258.9611, 258.9611, 
    258.9611, 258.9611, 258.9611, 258.9611, 258.9611, 258.9611,
  260, 260, 260, 260, 260, 260, 260, 260, 260, 260, 260, 260, 260, 260, 260, 
    260, 260, 260, 260, 260, 260, 260, 260, 260, 260, 260, 260, 260, 260, 
    260, 260, 260, 260, 260, 260, 260, 260, 260, 260, 260, 260, 260, 260, 
    260, 260, 260, 260, 260, 260, 260, 260, 260, 260, 260, 260, 260, 260, 
    260, 260, 260, 260, 260, 260, 260, 260, 260, 260, 260, 260, 260, 260, 
    260, 260, 260, 260, 260, 260, 260, 260, 260, 260, 260, 260, 260, 260, 
    260, 260, 260, 260, 260, 260, 260, 260, 260, 260, 260, 260,
  261.0389, 261.0389, 261.0389, 261.0389, 261.0389, 261.0389, 261.0389, 
    261.0389, 261.0389, 261.0389, 261.0389, 261.0389, 261.0389, 261.0389, 
    261.0389, 261.0389, 261.0389, 261.0389, 261.0389, 261.0389, 261.0389, 
    261.0389, 261.0389, 261.0389, 261.0389, 261.0389, 261.0389, 261.0389, 
    261.0389, 261.0389, 261.0389, 261.0389, 261.0389, 261.0389, 261.0389, 
    261.0389, 261.0389, 261.0389, 261.0389, 261.0389, 261.0389, 261.0389, 
    261.0389, 261.0389, 261.0389, 261.0389, 261.0389, 261.0389, 261.0389, 
    261.0389, 261.0389, 261.0389, 261.0389, 261.0389, 261.0389, 261.0389, 
    261.0389, 261.0389, 261.0389, 261.0389, 261.0389, 261.0389, 261.0389, 
    261.0389, 261.0389, 261.0389, 261.0389, 261.0389, 261.0389, 261.0389, 
    261.0389, 261.0389, 261.0389, 261.0389, 261.0389, 261.0389, 261.0389, 
    261.0389, 261.0389, 261.0389, 261.0389, 261.0389, 261.0389, 261.0389, 
    261.0389, 261.0389, 261.0389, 261.0389, 261.0389, 261.0389, 261.0389, 
    261.0389, 261.0389, 261.0389, 261.0389, 261.0389, 261.0389,
  262.0775, 262.0775, 262.0775, 262.0775, 262.0775, 262.0775, 262.0775, 
    262.0775, 262.0775, 262.0775, 262.0775, 262.0775, 262.0775, 262.0775, 
    262.0775, 262.0775, 262.0775, 262.0775, 262.0775, 262.0775, 262.0775, 
    262.0775, 262.0775, 262.0775, 262.0775, 262.0775, 262.0775, 262.0775, 
    262.0775, 262.0775, 262.0775, 262.0775, 262.0775, 262.0775, 262.0775, 
    262.0775, 262.0775, 262.0775, 262.0775, 262.0775, 262.0775, 262.0775, 
    262.0775, 262.0775, 262.0775, 262.0775, 262.0775, 262.0775, 262.0775, 
    262.0775, 262.0775, 262.0775, 262.0775, 262.0775, 262.0775, 262.0775, 
    262.0775, 262.0775, 262.0775, 262.0775, 262.0775, 262.0775, 262.0775, 
    262.0775, 262.0775, 262.0775, 262.0775, 262.0775, 262.0775, 262.0775, 
    262.0775, 262.0775, 262.0775, 262.0775, 262.0775, 262.0775, 262.0775, 
    262.0775, 262.0775, 262.0775, 262.0775, 262.0775, 262.0775, 262.0775, 
    262.0775, 262.0775, 262.0775, 262.0775, 262.0775, 262.0775, 262.0775, 
    262.0775, 262.0775, 262.0775, 262.0775, 262.0775, 262.0775,
  263.1154, 263.1154, 263.1154, 263.1154, 263.1154, 263.1154, 263.1154, 
    263.1154, 263.1154, 263.1154, 263.1154, 263.1154, 263.1154, 263.1154, 
    263.1154, 263.1154, 263.1154, 263.1154, 263.1154, 263.1154, 263.1154, 
    263.1154, 263.1154, 263.1154, 263.1154, 263.1154, 263.1154, 263.1154, 
    263.1154, 263.1154, 263.1154, 263.1154, 263.1154, 263.1154, 263.1154, 
    263.1154, 263.1154, 263.1154, 263.1154, 263.1154, 263.1154, 263.1154, 
    263.1154, 263.1154, 263.1154, 263.1154, 263.1154, 263.1154, 263.1154, 
    263.1154, 263.1154, 263.1154, 263.1154, 263.1154, 263.1154, 263.1154, 
    263.1154, 263.1154, 263.1154, 263.1154, 263.1154, 263.1154, 263.1154, 
    263.1154, 263.1154, 263.1154, 263.1154, 263.1154, 263.1154, 263.1154, 
    263.1154, 263.1154, 263.1154, 263.1154, 263.1154, 263.1154, 263.1154, 
    263.1154, 263.1154, 263.1154, 263.1154, 263.1154, 263.1154, 263.1154, 
    263.1154, 263.1154, 263.1154, 263.1154, 263.1154, 263.1154, 263.1154, 
    263.1154, 263.1154, 263.1154, 263.1154, 263.1154, 263.1154,
  264.1523, 264.1523, 264.1523, 264.1523, 264.1523, 264.1523, 264.1523, 
    264.1523, 264.1523, 264.1523, 264.1523, 264.1523, 264.1523, 264.1523, 
    264.1523, 264.1523, 264.1523, 264.1523, 264.1523, 264.1523, 264.1523, 
    264.1523, 264.1523, 264.1523, 264.1523, 264.1523, 264.1523, 264.1523, 
    264.1523, 264.1523, 264.1523, 264.1523, 264.1523, 264.1523, 264.1523, 
    264.1523, 264.1523, 264.1523, 264.1523, 264.1523, 264.1523, 264.1523, 
    264.1523, 264.1523, 264.1523, 264.1523, 264.1523, 264.1523, 264.1523, 
    264.1523, 264.1523, 264.1523, 264.1523, 264.1523, 264.1523, 264.1523, 
    264.1523, 264.1523, 264.1523, 264.1523, 264.1523, 264.1523, 264.1523, 
    264.1523, 264.1523, 264.1523, 264.1523, 264.1523, 264.1523, 264.1523, 
    264.1523, 264.1523, 264.1523, 264.1523, 264.1523, 264.1523, 264.1523, 
    264.1523, 264.1523, 264.1523, 264.1523, 264.1523, 264.1523, 264.1523, 
    264.1523, 264.1523, 264.1523, 264.1523, 264.1523, 264.1523, 264.1523, 
    264.1523, 264.1523, 264.1523, 264.1523, 264.1523, 264.1523,
  265.1878, 265.1878, 265.1878, 265.1878, 265.1878, 265.1878, 265.1878, 
    265.1878, 265.1878, 265.1878, 265.1878, 265.1878, 265.1878, 265.1878, 
    265.1878, 265.1878, 265.1878, 265.1878, 265.1878, 265.1878, 265.1878, 
    265.1878, 265.1878, 265.1878, 265.1878, 265.1878, 265.1878, 265.1878, 
    265.1878, 265.1878, 265.1878, 265.1878, 265.1878, 265.1878, 265.1878, 
    265.1878, 265.1878, 265.1878, 265.1878, 265.1878, 265.1878, 265.1878, 
    265.1878, 265.1878, 265.1878, 265.1878, 265.1878, 265.1878, 265.1878, 
    265.1878, 265.1878, 265.1878, 265.1878, 265.1878, 265.1878, 265.1878, 
    265.1878, 265.1878, 265.1878, 265.1878, 265.1878, 265.1878, 265.1878, 
    265.1878, 265.1878, 265.1878, 265.1878, 265.1878, 265.1878, 265.1878, 
    265.1878, 265.1878, 265.1878, 265.1878, 265.1878, 265.1878, 265.1878, 
    265.1878, 265.1878, 265.1878, 265.1878, 265.1878, 265.1878, 265.1878, 
    265.1878, 265.1878, 265.1878, 265.1878, 265.1878, 265.1878, 265.1878, 
    265.1878, 265.1878, 265.1878, 265.1878, 265.1878, 265.1878,
  266.2217, 266.2217, 266.2217, 266.2217, 266.2217, 266.2217, 266.2217, 
    266.2217, 266.2217, 266.2217, 266.2217, 266.2217, 266.2217, 266.2217, 
    266.2217, 266.2217, 266.2217, 266.2217, 266.2217, 266.2217, 266.2217, 
    266.2217, 266.2217, 266.2217, 266.2217, 266.2217, 266.2217, 266.2217, 
    266.2217, 266.2217, 266.2217, 266.2217, 266.2217, 266.2217, 266.2217, 
    266.2217, 266.2217, 266.2217, 266.2217, 266.2217, 266.2217, 266.2217, 
    266.2217, 266.2217, 266.2217, 266.2217, 266.2217, 266.2217, 266.2217, 
    266.2217, 266.2217, 266.2217, 266.2217, 266.2217, 266.2217, 266.2217, 
    266.2217, 266.2217, 266.2217, 266.2217, 266.2217, 266.2217, 266.2217, 
    266.2217, 266.2217, 266.2217, 266.2217, 266.2217, 266.2217, 266.2217, 
    266.2217, 266.2217, 266.2217, 266.2217, 266.2217, 266.2217, 266.2217, 
    266.2217, 266.2217, 266.2217, 266.2217, 266.2217, 266.2217, 266.2217, 
    266.2217, 266.2217, 266.2217, 266.2217, 266.2217, 266.2217, 266.2217, 
    266.2217, 266.2217, 266.2217, 266.2217, 266.2217, 266.2217,
  267.2535, 267.2535, 267.2535, 267.2535, 267.2535, 267.2535, 267.2535, 
    267.2535, 267.2535, 267.2535, 267.2535, 267.2535, 267.2535, 267.2535, 
    267.2535, 267.2535, 267.2535, 267.2535, 267.2535, 267.2535, 267.2535, 
    267.2535, 267.2535, 267.2535, 267.2535, 267.2535, 267.2535, 267.2535, 
    267.2535, 267.2535, 267.2535, 267.2535, 267.2535, 267.2535, 267.2535, 
    267.2535, 267.2535, 267.2535, 267.2535, 267.2535, 267.2535, 267.2535, 
    267.2535, 267.2535, 267.2535, 267.2535, 267.2535, 267.2535, 267.2535, 
    267.2535, 267.2535, 267.2535, 267.2535, 267.2535, 267.2535, 267.2535, 
    267.2535, 267.2535, 267.2535, 267.2535, 267.2535, 267.2535, 267.2535, 
    267.2535, 267.2535, 267.2535, 267.2535, 267.2535, 267.2535, 267.2535, 
    267.2535, 267.2535, 267.2535, 267.2535, 267.2535, 267.2535, 267.2535, 
    267.2535, 267.2535, 267.2535, 267.2535, 267.2535, 267.2535, 267.2535, 
    267.2535, 267.2535, 267.2535, 267.2535, 267.2535, 267.2535, 267.2535, 
    267.2535, 267.2535, 267.2535, 267.2535, 267.2535, 267.2535,
  268.283, 268.283, 268.283, 268.283, 268.283, 268.283, 268.283, 268.283, 
    268.283, 268.283, 268.283, 268.283, 268.283, 268.283, 268.283, 268.283, 
    268.283, 268.283, 268.283, 268.283, 268.283, 268.283, 268.283, 268.283, 
    268.283, 268.283, 268.283, 268.283, 268.283, 268.283, 268.283, 268.283, 
    268.283, 268.283, 268.283, 268.283, 268.283, 268.283, 268.283, 268.283, 
    268.283, 268.283, 268.283, 268.283, 268.283, 268.283, 268.283, 268.283, 
    268.283, 268.283, 268.283, 268.283, 268.283, 268.283, 268.283, 268.283, 
    268.283, 268.283, 268.283, 268.283, 268.283, 268.283, 268.283, 268.283, 
    268.283, 268.283, 268.283, 268.283, 268.283, 268.283, 268.283, 268.283, 
    268.283, 268.283, 268.283, 268.283, 268.283, 268.283, 268.283, 268.283, 
    268.283, 268.283, 268.283, 268.283, 268.283, 268.283, 268.283, 268.283, 
    268.283, 268.283, 268.283, 268.283, 268.283, 268.283, 268.283, 268.283, 
    268.283,
  269.3098, 269.3098, 269.3098, 269.3098, 269.3098, 269.3098, 269.3098, 
    269.3098, 269.3098, 269.3098, 269.3098, 269.3098, 269.3098, 269.3098, 
    269.3098, 269.3098, 269.3098, 269.3098, 269.3098, 269.3098, 269.3098, 
    269.3098, 269.3098, 269.3098, 269.3098, 269.3098, 269.3098, 269.3098, 
    269.3098, 269.3098, 269.3098, 269.3098, 269.3098, 269.3098, 269.3098, 
    269.3098, 269.3098, 269.3098, 269.3098, 269.3098, 269.3098, 269.3098, 
    269.3098, 269.3098, 269.3098, 269.3098, 269.3098, 269.3098, 269.3098, 
    269.3098, 269.3098, 269.3098, 269.3098, 269.3098, 269.3098, 269.3098, 
    269.3098, 269.3098, 269.3098, 269.3098, 269.3098, 269.3098, 269.3098, 
    269.3098, 269.3098, 269.3098, 269.3098, 269.3098, 269.3098, 269.3098, 
    269.3098, 269.3098, 269.3098, 269.3098, 269.3098, 269.3098, 269.3098, 
    269.3098, 269.3098, 269.3098, 269.3098, 269.3098, 269.3098, 269.3098, 
    269.3098, 269.3098, 269.3098, 269.3098, 269.3098, 269.3098, 269.3098, 
    269.3098, 269.3098, 269.3098, 269.3098, 269.3098, 269.3098,
  270.3337, 270.3337, 270.3337, 270.3337, 270.3337, 270.3337, 270.3337, 
    270.3337, 270.3337, 270.3337, 270.3337, 270.3337, 270.3337, 270.3337, 
    270.3337, 270.3337, 270.3337, 270.3337, 270.3337, 270.3337, 270.3337, 
    270.3337, 270.3337, 270.3337, 270.3337, 270.3337, 270.3337, 270.3337, 
    270.3337, 270.3337, 270.3337, 270.3337, 270.3337, 270.3337, 270.3337, 
    270.3337, 270.3337, 270.3337, 270.3337, 270.3337, 270.3337, 270.3337, 
    270.3337, 270.3337, 270.3337, 270.3337, 270.3337, 270.3337, 270.3337, 
    270.3337, 270.3337, 270.3337, 270.3337, 270.3337, 270.3337, 270.3337, 
    270.3337, 270.3337, 270.3337, 270.3337, 270.3337, 270.3337, 270.3337, 
    270.3337, 270.3337, 270.3337, 270.3337, 270.3337, 270.3337, 270.3337, 
    270.3337, 270.3337, 270.3337, 270.3337, 270.3337, 270.3337, 270.3337, 
    270.3337, 270.3337, 270.3337, 270.3337, 270.3337, 270.3337, 270.3337, 
    270.3337, 270.3337, 270.3337, 270.3337, 270.3337, 270.3337, 270.3337, 
    270.3337, 270.3337, 270.3337, 270.3337, 270.3337, 270.3337,
  271.3542, 271.3542, 271.3542, 271.3542, 271.3542, 271.3542, 271.3542, 
    271.3542, 271.3542, 271.3542, 271.3542, 271.3542, 271.3542, 271.3542, 
    271.3542, 271.3542, 271.3542, 271.3542, 271.3542, 271.3542, 271.3542, 
    271.3542, 271.3542, 271.3542, 271.3542, 271.3542, 271.3542, 271.3542, 
    271.3542, 271.3542, 271.3542, 271.3542, 271.3542, 271.3542, 271.3542, 
    271.3542, 271.3542, 271.3542, 271.3542, 271.3542, 271.3542, 271.3542, 
    271.3542, 271.3542, 271.3542, 271.3542, 271.3542, 271.3542, 271.3542, 
    271.3542, 271.3542, 271.3542, 271.3542, 271.3542, 271.3542, 271.3542, 
    271.3542, 271.3542, 271.3542, 271.3542, 271.3542, 271.3542, 271.3542, 
    271.3542, 271.3542, 271.3542, 271.3542, 271.3542, 271.3542, 271.3542, 
    271.3542, 271.3542, 271.3542, 271.3542, 271.3542, 271.3542, 271.3542, 
    271.3542, 271.3542, 271.3542, 271.3542, 271.3542, 271.3542, 271.3542, 
    271.3542, 271.3542, 271.3542, 271.3542, 271.3542, 271.3542, 271.3542, 
    271.3542, 271.3542, 271.3542, 271.3542, 271.3542, 271.3542,
  272.3713, 272.3713, 272.3713, 272.3713, 272.3713, 272.3713, 272.3713, 
    272.3713, 272.3713, 272.3713, 272.3713, 272.3713, 272.3713, 272.3713, 
    272.3713, 272.3713, 272.3713, 272.3713, 272.3713, 272.3713, 272.3713, 
    272.3713, 272.3713, 272.3713, 272.3713, 272.3713, 272.3713, 272.3713, 
    272.3713, 272.3713, 272.3713, 272.3713, 272.3713, 272.3713, 272.3713, 
    272.3713, 272.3713, 272.3713, 272.3713, 272.3713, 272.3713, 272.3713, 
    272.3713, 272.3713, 272.3713, 272.3713, 272.3713, 272.3713, 272.3713, 
    272.3713, 272.3713, 272.3713, 272.3713, 272.3713, 272.3713, 272.3713, 
    272.3713, 272.3713, 272.3713, 272.3713, 272.3713, 272.3713, 272.3713, 
    272.3713, 272.3713, 272.3713, 272.3713, 272.3713, 272.3713, 272.3713, 
    272.3713, 272.3713, 272.3713, 272.3713, 272.3713, 272.3713, 272.3713, 
    272.3713, 272.3713, 272.3713, 272.3713, 272.3713, 272.3713, 272.3713, 
    272.3713, 272.3713, 272.3713, 272.3713, 272.3713, 272.3713, 272.3713, 
    272.3713, 272.3713, 272.3713, 272.3713, 272.3713, 272.3713,
  273.3844, 273.3844, 273.3844, 273.3844, 273.3844, 273.3844, 273.3844, 
    273.3844, 273.3844, 273.3844, 273.3844, 273.3844, 273.3844, 273.3844, 
    273.3844, 273.3844, 273.3844, 273.3844, 273.3844, 273.3844, 273.3844, 
    273.3844, 273.3844, 273.3844, 273.3844, 273.3844, 273.3844, 273.3844, 
    273.3844, 273.3844, 273.3844, 273.3844, 273.3844, 273.3844, 273.3844, 
    273.3844, 273.3844, 273.3844, 273.3844, 273.3844, 273.3844, 273.3844, 
    273.3844, 273.3844, 273.3844, 273.3844, 273.3844, 273.3844, 273.3844, 
    273.3844, 273.3844, 273.3844, 273.3844, 273.3844, 273.3844, 273.3844, 
    273.3844, 273.3844, 273.3844, 273.3844, 273.3844, 273.3844, 273.3844, 
    273.3844, 273.3844, 273.3844, 273.3844, 273.3844, 273.3844, 273.3844, 
    273.3844, 273.3844, 273.3844, 273.3844, 273.3844, 273.3844, 273.3844, 
    273.3844, 273.3844, 273.3844, 273.3844, 273.3844, 273.3844, 273.3844, 
    273.3844, 273.3844, 273.3844, 273.3844, 273.3844, 273.3844, 273.3844, 
    273.3844, 273.3844, 273.3844, 273.3844, 273.3844, 273.3844,
  274.3935, 274.3935, 274.3935, 274.3935, 274.3935, 274.3935, 274.3935, 
    274.3935, 274.3935, 274.3935, 274.3935, 274.3935, 274.3935, 274.3935, 
    274.3935, 274.3935, 274.3935, 274.3935, 274.3935, 274.3935, 274.3935, 
    274.3935, 274.3935, 274.3935, 274.3935, 274.3935, 274.3935, 274.3935, 
    274.3935, 274.3935, 274.3935, 274.3935, 274.3935, 274.3935, 274.3935, 
    274.3935, 274.3935, 274.3935, 274.3935, 274.3935, 274.3935, 274.3935, 
    274.3935, 274.3935, 274.3935, 274.3935, 274.3935, 274.3935, 274.3935, 
    274.3935, 274.3935, 274.3935, 274.3935, 274.3935, 274.3935, 274.3935, 
    274.3935, 274.3935, 274.3935, 274.3935, 274.3935, 274.3935, 274.3935, 
    274.3935, 274.3935, 274.3935, 274.3935, 274.3935, 274.3935, 274.3935, 
    274.3935, 274.3935, 274.3935, 274.3935, 274.3935, 274.3935, 274.3935, 
    274.3935, 274.3935, 274.3935, 274.3935, 274.3935, 274.3935, 274.3935, 
    274.3935, 274.3935, 274.3935, 274.3935, 274.3935, 274.3935, 274.3935, 
    274.3935, 274.3935, 274.3935, 274.3935, 274.3935, 274.3935,
  275.3981, 275.3981, 275.3981, 275.3981, 275.3981, 275.3981, 275.3981, 
    275.3981, 275.3981, 275.3981, 275.3981, 275.3981, 275.3981, 275.3981, 
    275.3981, 275.3981, 275.3981, 275.3981, 275.3981, 275.3981, 275.3981, 
    275.3981, 275.3981, 275.3981, 275.3981, 275.3981, 275.3981, 275.3981, 
    275.3981, 275.3981, 275.3981, 275.3981, 275.3981, 275.3981, 275.3981, 
    275.3981, 275.3981, 275.3981, 275.3981, 275.3981, 275.3981, 275.3981, 
    275.3981, 275.3981, 275.3981, 275.3981, 275.3981, 275.3981, 275.3981, 
    275.3981, 275.3981, 275.3981, 275.3981, 275.3981, 275.3981, 275.3981, 
    275.3981, 275.3981, 275.3981, 275.3981, 275.3981, 275.3981, 275.3981, 
    275.3981, 275.3981, 275.3981, 275.3981, 275.3981, 275.3981, 275.3981, 
    275.3981, 275.3981, 275.3981, 275.3981, 275.3981, 275.3981, 275.3981, 
    275.3981, 275.3981, 275.3981, 275.3981, 275.3981, 275.3981, 275.3981, 
    275.3981, 275.3981, 275.3981, 275.3981, 275.3981, 275.3981, 275.3981, 
    275.3981, 275.3981, 275.3981, 275.3981, 275.3981, 275.3981,
  276.3981, 276.3981, 276.3981, 276.3981, 276.3981, 276.3981, 276.3981, 
    276.3981, 276.3981, 276.3981, 276.3981, 276.3981, 276.3981, 276.3981, 
    276.3981, 276.3981, 276.3981, 276.3981, 276.3981, 276.3981, 276.3981, 
    276.3981, 276.3981, 276.3981, 276.3981, 276.3981, 276.3981, 276.3981, 
    276.3981, 276.3981, 276.3981, 276.3981, 276.3981, 276.3981, 276.3981, 
    276.3981, 276.3981, 276.3981, 276.3981, 276.3981, 276.3981, 276.3981, 
    276.3981, 276.3981, 276.3981, 276.3981, 276.3981, 276.3981, 276.3981, 
    276.3981, 276.3981, 276.3981, 276.3981, 276.3981, 276.3981, 276.3981, 
    276.3981, 276.3981, 276.3981, 276.3981, 276.3981, 276.3981, 276.3981, 
    276.3981, 276.3981, 276.3981, 276.3981, 276.3981, 276.3981, 276.3981, 
    276.3981, 276.3981, 276.3981, 276.3981, 276.3981, 276.3981, 276.3981, 
    276.3981, 276.3981, 276.3981, 276.3981, 276.3981, 276.3981, 276.3981, 
    276.3981, 276.3981, 276.3981, 276.3981, 276.3981, 276.3981, 276.3981, 
    276.3981, 276.3981, 276.3981, 276.3981, 276.3981, 276.3981,
  277.3932, 277.3932, 277.3932, 277.3932, 277.3932, 277.3932, 277.3932, 
    277.3932, 277.3932, 277.3932, 277.3932, 277.3932, 277.3932, 277.3932, 
    277.3932, 277.3932, 277.3932, 277.3932, 277.3932, 277.3932, 277.3932, 
    277.3932, 277.3932, 277.3932, 277.3932, 277.3932, 277.3932, 277.3932, 
    277.3932, 277.3932, 277.3932, 277.3932, 277.3932, 277.3932, 277.3932, 
    277.3932, 277.3932, 277.3932, 277.3932, 277.3932, 277.3932, 277.3932, 
    277.3932, 277.3932, 277.3932, 277.3932, 277.3932, 277.3932, 277.3932, 
    277.3932, 277.3932, 277.3932, 277.3932, 277.3932, 277.3932, 277.3932, 
    277.3932, 277.3932, 277.3932, 277.3932, 277.3932, 277.3932, 277.3932, 
    277.3932, 277.3932, 277.3932, 277.3932, 277.3932, 277.3932, 277.3932, 
    277.3932, 277.3932, 277.3932, 277.3932, 277.3932, 277.3932, 277.3932, 
    277.3932, 277.3932, 277.3932, 277.3932, 277.3932, 277.3932, 277.3932, 
    277.3932, 277.3932, 277.3932, 277.3932, 277.3932, 277.3932, 277.3932, 
    277.3932, 277.3932, 277.3932, 277.3932, 277.3932, 277.3932,
  278.3832, 278.3832, 278.3832, 278.3832, 278.3832, 278.3832, 278.3832, 
    278.3832, 278.3832, 278.3832, 278.3832, 278.3832, 278.3832, 278.3832, 
    278.3832, 278.3832, 278.3832, 278.3832, 278.3832, 278.3832, 278.3832, 
    278.3832, 278.3832, 278.3832, 278.3832, 278.3832, 278.3832, 278.3832, 
    278.3832, 278.3832, 278.3832, 278.3832, 278.3832, 278.3832, 278.3832, 
    278.3832, 278.3832, 278.3832, 278.3832, 278.3832, 278.3832, 278.3832, 
    278.3832, 278.3832, 278.3832, 278.3832, 278.3832, 278.3832, 278.3832, 
    278.3832, 278.3832, 278.3832, 278.3832, 278.3832, 278.3832, 278.3832, 
    278.3832, 278.3832, 278.3832, 278.3832, 278.3832, 278.3832, 278.3832, 
    278.3832, 278.3832, 278.3832, 278.3832, 278.3832, 278.3832, 278.3832, 
    278.3832, 278.3832, 278.3832, 278.3832, 278.3832, 278.3832, 278.3832, 
    278.3832, 278.3832, 278.3832, 278.3832, 278.3832, 278.3832, 278.3832, 
    278.3832, 278.3832, 278.3832, 278.3832, 278.3832, 278.3832, 278.3832, 
    278.3832, 278.3832, 278.3832, 278.3832, 278.3832, 278.3832,
  279.3678, 279.3678, 279.3678, 279.3678, 279.3678, 279.3678, 279.3678, 
    279.3678, 279.3678, 279.3678, 279.3678, 279.3678, 279.3678, 279.3678, 
    279.3678, 279.3678, 279.3678, 279.3678, 279.3678, 279.3678, 279.3678, 
    279.3678, 279.3678, 279.3678, 279.3678, 279.3678, 279.3678, 279.3678, 
    279.3678, 279.3678, 279.3678, 279.3678, 279.3678, 279.3678, 279.3678, 
    279.3678, 279.3678, 279.3678, 279.3678, 279.3678, 279.3678, 279.3678, 
    279.3678, 279.3678, 279.3678, 279.3678, 279.3678, 279.3678, 279.3678, 
    279.3678, 279.3678, 279.3678, 279.3678, 279.3678, 279.3678, 279.3678, 
    279.3678, 279.3678, 279.3678, 279.3678, 279.3678, 279.3678, 279.3678, 
    279.3678, 279.3678, 279.3678, 279.3678, 279.3678, 279.3678, 279.3678, 
    279.3678, 279.3678, 279.3678, 279.3678, 279.3678, 279.3678, 279.3678, 
    279.3678, 279.3678, 279.3678, 279.3678, 279.3678, 279.3678, 279.3678, 
    279.3678, 279.3678, 279.3678, 279.3678, 279.3678, 279.3678, 279.3678, 
    279.3678, 279.3678, 279.3678, 279.3678, 279.3678, 279.3678,
  280.3468, 280.3468, 280.3468, 280.3468, 280.3468, 280.3468, 280.3468, 
    280.3468, 280.3468, 280.3468, 280.3468, 280.3468, 280.3468, 280.3468, 
    280.3468, 280.3468, 280.3468, 280.3468, 280.3468, 280.3468, 280.3468, 
    280.3468, 280.3468, 280.3468, 280.3468, 280.3468, 280.3468, 280.3468, 
    280.3468, 280.3468, 280.3468, 280.3468, 280.3468, 280.3468, 280.3468, 
    280.3468, 280.3468, 280.3468, 280.3468, 280.3468, 280.3468, 280.3468, 
    280.3468, 280.3468, 280.3468, 280.3468, 280.3468, 280.3468, 280.3468, 
    280.3468, 280.3468, 280.3468, 280.3468, 280.3468, 280.3468, 280.3468, 
    280.3468, 280.3468, 280.3468, 280.3468, 280.3468, 280.3468, 280.3468, 
    280.3468, 280.3468, 280.3468, 280.3468, 280.3468, 280.3468, 280.3468, 
    280.3468, 280.3468, 280.3468, 280.3468, 280.3468, 280.3468, 280.3468, 
    280.3468, 280.3468, 280.3468, 280.3468, 280.3468, 280.3468, 280.3468, 
    280.3468, 280.3468, 280.3468, 280.3468, 280.3468, 280.3468, 280.3468, 
    280.3468, 280.3468, 280.3468, 280.3468, 280.3468, 280.3468,
  281.3201, 281.3201, 281.3201, 281.3201, 281.3201, 281.3201, 281.3201, 
    281.3201, 281.3201, 281.3201, 281.3201, 281.3201, 281.3201, 281.3201, 
    281.3201, 281.3201, 281.3201, 281.3201, 281.3201, 281.3201, 281.3201, 
    281.3201, 281.3201, 281.3201, 281.3201, 281.3201, 281.3201, 281.3201, 
    281.3201, 281.3201, 281.3201, 281.3201, 281.3201, 281.3201, 281.3201, 
    281.3201, 281.3201, 281.3201, 281.3201, 281.3201, 281.3201, 281.3201, 
    281.3201, 281.3201, 281.3201, 281.3201, 281.3201, 281.3201, 281.3201, 
    281.3201, 281.3201, 281.3201, 281.3201, 281.3201, 281.3201, 281.3201, 
    281.3201, 281.3201, 281.3201, 281.3201, 281.3201, 281.3201, 281.3201, 
    281.3201, 281.3201, 281.3201, 281.3201, 281.3201, 281.3201, 281.3201, 
    281.3201, 281.3201, 281.3201, 281.3201, 281.3201, 281.3201, 281.3201, 
    281.3201, 281.3201, 281.3201, 281.3201, 281.3201, 281.3201, 281.3201, 
    281.3201, 281.3201, 281.3201, 281.3201, 281.3201, 281.3201, 281.3201, 
    281.3201, 281.3201, 281.3201, 281.3201, 281.3201, 281.3201,
  282.2874, 282.2874, 282.2874, 282.2874, 282.2874, 282.2874, 282.2874, 
    282.2874, 282.2874, 282.2874, 282.2874, 282.2874, 282.2874, 282.2874, 
    282.2874, 282.2874, 282.2874, 282.2874, 282.2874, 282.2874, 282.2874, 
    282.2874, 282.2874, 282.2874, 282.2874, 282.2874, 282.2874, 282.2874, 
    282.2874, 282.2874, 282.2874, 282.2874, 282.2874, 282.2874, 282.2874, 
    282.2874, 282.2874, 282.2874, 282.2874, 282.2874, 282.2874, 282.2874, 
    282.2874, 282.2874, 282.2874, 282.2874, 282.2874, 282.2874, 282.2874, 
    282.2874, 282.2874, 282.2874, 282.2874, 282.2874, 282.2874, 282.2874, 
    282.2874, 282.2874, 282.2874, 282.2874, 282.2874, 282.2874, 282.2874, 
    282.2874, 282.2874, 282.2874, 282.2874, 282.2874, 282.2874, 282.2874, 
    282.2874, 282.2874, 282.2874, 282.2874, 282.2874, 282.2874, 282.2874, 
    282.2874, 282.2874, 282.2874, 282.2874, 282.2874, 282.2874, 282.2874, 
    282.2874, 282.2874, 282.2874, 282.2874, 282.2874, 282.2874, 282.2874, 
    282.2874, 282.2874, 282.2874, 282.2874, 282.2874, 282.2874,
  283.2486, 283.2486, 283.2486, 283.2486, 283.2486, 283.2486, 283.2486, 
    283.2486, 283.2486, 283.2486, 283.2486, 283.2486, 283.2486, 283.2486, 
    283.2486, 283.2486, 283.2486, 283.2486, 283.2486, 283.2486, 283.2486, 
    283.2486, 283.2486, 283.2486, 283.2486, 283.2486, 283.2486, 283.2486, 
    283.2486, 283.2486, 283.2486, 283.2486, 283.2486, 283.2486, 283.2486, 
    283.2486, 283.2486, 283.2486, 283.2486, 283.2486, 283.2486, 283.2486, 
    283.2486, 283.2486, 283.2486, 283.2486, 283.2486, 283.2486, 283.2486, 
    283.2486, 283.2486, 283.2486, 283.2486, 283.2486, 283.2486, 283.2486, 
    283.2486, 283.2486, 283.2486, 283.2486, 283.2486, 283.2486, 283.2486, 
    283.2486, 283.2486, 283.2486, 283.2486, 283.2486, 283.2486, 283.2486, 
    283.2486, 283.2486, 283.2486, 283.2486, 283.2486, 283.2486, 283.2486, 
    283.2486, 283.2486, 283.2486, 283.2486, 283.2486, 283.2486, 283.2486, 
    283.2486, 283.2486, 283.2486, 283.2486, 283.2486, 283.2486, 283.2486, 
    283.2486, 283.2486, 283.2486, 283.2486, 283.2486, 283.2486,
  284.2034, 284.2034, 284.2034, 284.2034, 284.2034, 284.2034, 284.2034, 
    284.2034, 284.2034, 284.2034, 284.2034, 284.2034, 284.2034, 284.2034, 
    284.2034, 284.2034, 284.2034, 284.2034, 284.2034, 284.2034, 284.2034, 
    284.2034, 284.2034, 284.2034, 284.2034, 284.2034, 284.2034, 284.2034, 
    284.2034, 284.2034, 284.2034, 284.2034, 284.2034, 284.2034, 284.2034, 
    284.2034, 284.2034, 284.2034, 284.2034, 284.2034, 284.2034, 284.2034, 
    284.2034, 284.2034, 284.2034, 284.2034, 284.2034, 284.2034, 284.2034, 
    284.2034, 284.2034, 284.2034, 284.2034, 284.2034, 284.2034, 284.2034, 
    284.2034, 284.2034, 284.2034, 284.2034, 284.2034, 284.2034, 284.2034, 
    284.2034, 284.2034, 284.2034, 284.2034, 284.2034, 284.2034, 284.2034, 
    284.2034, 284.2034, 284.2034, 284.2034, 284.2034, 284.2034, 284.2034, 
    284.2034, 284.2034, 284.2034, 284.2034, 284.2034, 284.2034, 284.2034, 
    284.2034, 284.2034, 284.2034, 284.2034, 284.2034, 284.2034, 284.2034, 
    284.2034, 284.2034, 284.2034, 284.2034, 284.2034, 284.2034,
  285.1519, 285.1519, 285.1519, 285.1519, 285.1519, 285.1519, 285.1519, 
    285.1519, 285.1519, 285.1519, 285.1519, 285.1519, 285.1519, 285.1519, 
    285.1519, 285.1519, 285.1519, 285.1519, 285.1519, 285.1519, 285.1519, 
    285.1519, 285.1519, 285.1519, 285.1519, 285.1519, 285.1519, 285.1519, 
    285.1519, 285.1519, 285.1519, 285.1519, 285.1519, 285.1519, 285.1519, 
    285.1519, 285.1519, 285.1519, 285.1519, 285.1519, 285.1519, 285.1519, 
    285.1519, 285.1519, 285.1519, 285.1519, 285.1519, 285.1519, 285.1519, 
    285.1519, 285.1519, 285.1519, 285.1519, 285.1519, 285.1519, 285.1519, 
    285.1519, 285.1519, 285.1519, 285.1519, 285.1519, 285.1519, 285.1519, 
    285.1519, 285.1519, 285.1519, 285.1519, 285.1519, 285.1519, 285.1519, 
    285.1519, 285.1519, 285.1519, 285.1519, 285.1519, 285.1519, 285.1519, 
    285.1519, 285.1519, 285.1519, 285.1519, 285.1519, 285.1519, 285.1519, 
    285.1519, 285.1519, 285.1519, 285.1519, 285.1519, 285.1519, 285.1519, 
    285.1519, 285.1519, 285.1519, 285.1519, 285.1519, 285.1519,
  286.0937, 286.0937, 286.0937, 286.0937, 286.0937, 286.0937, 286.0937, 
    286.0937, 286.0937, 286.0937, 286.0937, 286.0937, 286.0937, 286.0937, 
    286.0937, 286.0937, 286.0937, 286.0937, 286.0937, 286.0937, 286.0937, 
    286.0937, 286.0937, 286.0937, 286.0937, 286.0937, 286.0937, 286.0937, 
    286.0937, 286.0937, 286.0937, 286.0937, 286.0937, 286.0937, 286.0937, 
    286.0937, 286.0937, 286.0937, 286.0937, 286.0937, 286.0937, 286.0937, 
    286.0937, 286.0937, 286.0937, 286.0937, 286.0937, 286.0937, 286.0937, 
    286.0937, 286.0937, 286.0937, 286.0937, 286.0937, 286.0937, 286.0937, 
    286.0937, 286.0937, 286.0937, 286.0937, 286.0937, 286.0937, 286.0937, 
    286.0937, 286.0937, 286.0937, 286.0937, 286.0937, 286.0937, 286.0937, 
    286.0937, 286.0937, 286.0937, 286.0937, 286.0937, 286.0937, 286.0937, 
    286.0937, 286.0937, 286.0937, 286.0937, 286.0937, 286.0937, 286.0937, 
    286.0937, 286.0937, 286.0937, 286.0937, 286.0937, 286.0937, 286.0937, 
    286.0937, 286.0937, 286.0937, 286.0937, 286.0937, 286.0937,
  287.0288, 287.0288, 287.0288, 287.0288, 287.0288, 287.0288, 287.0288, 
    287.0288, 287.0288, 287.0288, 287.0288, 287.0288, 287.0288, 287.0288, 
    287.0288, 287.0288, 287.0288, 287.0288, 287.0288, 287.0288, 287.0288, 
    287.0288, 287.0288, 287.0288, 287.0288, 287.0288, 287.0288, 287.0288, 
    287.0288, 287.0288, 287.0288, 287.0288, 287.0288, 287.0288, 287.0288, 
    287.0288, 287.0288, 287.0288, 287.0288, 287.0288, 287.0288, 287.0288, 
    287.0288, 287.0288, 287.0288, 287.0288, 287.0288, 287.0288, 287.0288, 
    287.0288, 287.0288, 287.0288, 287.0288, 287.0288, 287.0288, 287.0288, 
    287.0288, 287.0288, 287.0288, 287.0288, 287.0288, 287.0288, 287.0288, 
    287.0288, 287.0288, 287.0288, 287.0288, 287.0288, 287.0288, 287.0288, 
    287.0288, 287.0288, 287.0288, 287.0288, 287.0288, 287.0288, 287.0288, 
    287.0288, 287.0288, 287.0288, 287.0288, 287.0288, 287.0288, 287.0288, 
    287.0288, 287.0288, 287.0288, 287.0288, 287.0288, 287.0288, 287.0288, 
    287.0288, 287.0288, 287.0288, 287.0288, 287.0288, 287.0288,
  287.957, 287.957, 287.957, 287.957, 287.957, 287.957, 287.957, 287.957, 
    287.957, 287.957, 287.957, 287.957, 287.957, 287.957, 287.957, 287.957, 
    287.957, 287.957, 287.957, 287.957, 287.957, 287.957, 287.957, 287.957, 
    287.957, 287.957, 287.957, 287.957, 287.957, 287.957, 287.957, 287.957, 
    287.957, 287.957, 287.957, 287.957, 287.957, 287.957, 287.957, 287.957, 
    287.957, 287.957, 287.957, 287.957, 287.957, 287.957, 287.957, 287.957, 
    287.957, 287.957, 287.957, 287.957, 287.957, 287.957, 287.957, 287.957, 
    287.957, 287.957, 287.957, 287.957, 287.957, 287.957, 287.957, 287.957, 
    287.957, 287.957, 287.957, 287.957, 287.957, 287.957, 287.957, 287.957, 
    287.957, 287.957, 287.957, 287.957, 287.957, 287.957, 287.957, 287.957, 
    287.957, 287.957, 287.957, 287.957, 287.957, 287.957, 287.957, 287.957, 
    287.957, 287.957, 287.957, 287.957, 287.957, 287.957, 287.957, 287.957, 
    287.957,
  288.8784, 288.8784, 288.8784, 288.8784, 288.8784, 288.8784, 288.8784, 
    288.8784, 288.8784, 288.8784, 288.8784, 288.8784, 288.8784, 288.8784, 
    288.8784, 288.8784, 288.8784, 288.8784, 288.8784, 288.8784, 288.8784, 
    288.8784, 288.8784, 288.8784, 288.8784, 288.8784, 288.8784, 288.8784, 
    288.8784, 288.8784, 288.8784, 288.8784, 288.8784, 288.8784, 288.8784, 
    288.8784, 288.8784, 288.8784, 288.8784, 288.8784, 288.8784, 288.8784, 
    288.8784, 288.8784, 288.8784, 288.8784, 288.8784, 288.8784, 288.8784, 
    288.8784, 288.8784, 288.8784, 288.8784, 288.8784, 288.8784, 288.8784, 
    288.8784, 288.8784, 288.8784, 288.8784, 288.8784, 288.8784, 288.8784, 
    288.8784, 288.8784, 288.8784, 288.8784, 288.8784, 288.8784, 288.8784, 
    288.8784, 288.8784, 288.8784, 288.8784, 288.8784, 288.8784, 288.8784, 
    288.8784, 288.8784, 288.8784, 288.8784, 288.8784, 288.8784, 288.8784, 
    288.8784, 288.8784, 288.8784, 288.8784, 288.8784, 288.8784, 288.8784, 
    288.8784, 288.8784, 288.8784, 288.8784, 288.8784, 288.8784,
  289.7927, 289.7927, 289.7927, 289.7927, 289.7927, 289.7927, 289.7927, 
    289.7927, 289.7927, 289.7927, 289.7927, 289.7927, 289.7927, 289.7927, 
    289.7927, 289.7927, 289.7927, 289.7927, 289.7927, 289.7927, 289.7927, 
    289.7927, 289.7927, 289.7927, 289.7927, 289.7927, 289.7927, 289.7927, 
    289.7927, 289.7927, 289.7927, 289.7927, 289.7927, 289.7927, 289.7927, 
    289.7927, 289.7927, 289.7927, 289.7927, 289.7927, 289.7927, 289.7927, 
    289.7927, 289.7927, 289.7927, 289.7927, 289.7927, 289.7927, 289.7927, 
    289.7927, 289.7927, 289.7927, 289.7927, 289.7927, 289.7927, 289.7927, 
    289.7927, 289.7927, 289.7927, 289.7927, 289.7927, 289.7927, 289.7927, 
    289.7927, 289.7927, 289.7927, 289.7927, 289.7927, 289.7927, 289.7927, 
    289.7927, 289.7927, 289.7927, 289.7927, 289.7927, 289.7927, 289.7927, 
    289.7927, 289.7927, 289.7927, 289.7927, 289.7927, 289.7927, 289.7927, 
    289.7927, 289.7927, 289.7927, 289.7927, 289.7927, 289.7927, 289.7927, 
    289.7927, 289.7927, 289.7927, 289.7927, 289.7927, 289.7927,
  290.6998, 290.6998, 290.6998, 290.6998, 290.6998, 290.6998, 290.6998, 
    290.6998, 290.6998, 290.6998, 290.6998, 290.6998, 290.6998, 290.6998, 
    290.6998, 290.6998, 290.6998, 290.6998, 290.6998, 290.6998, 290.6998, 
    290.6998, 290.6998, 290.6998, 290.6998, 290.6998, 290.6998, 290.6998, 
    290.6998, 290.6998, 290.6998, 290.6998, 290.6998, 290.6998, 290.6998, 
    290.6998, 290.6998, 290.6998, 290.6998, 290.6998, 290.6998, 290.6998, 
    290.6998, 290.6998, 290.6998, 290.6998, 290.6998, 290.6998, 290.6998, 
    290.6998, 290.6998, 290.6998, 290.6998, 290.6998, 290.6998, 290.6998, 
    290.6998, 290.6998, 290.6998, 290.6998, 290.6998, 290.6998, 290.6998, 
    290.6998, 290.6998, 290.6998, 290.6998, 290.6998, 290.6998, 290.6998, 
    290.6998, 290.6998, 290.6998, 290.6998, 290.6998, 290.6998, 290.6998, 
    290.6998, 290.6998, 290.6998, 290.6998, 290.6998, 290.6998, 290.6998, 
    290.6998, 290.6998, 290.6998, 290.6998, 290.6998, 290.6998, 290.6998, 
    290.6998, 290.6998, 290.6998, 290.6998, 290.6998, 290.6998,
  291.5998, 291.5998, 291.5998, 291.5998, 291.5998, 291.5998, 291.5998, 
    291.5998, 291.5998, 291.5998, 291.5998, 291.5998, 291.5998, 291.5998, 
    291.5998, 291.5998, 291.5998, 291.5998, 291.5998, 291.5998, 291.5998, 
    291.5998, 291.5998, 291.5998, 291.5998, 291.5998, 291.5998, 291.5998, 
    291.5998, 291.5998, 291.5998, 291.5998, 291.5998, 291.5998, 291.5998, 
    291.5998, 291.5998, 291.5998, 291.5998, 291.5998, 291.5998, 291.5998, 
    291.5998, 291.5998, 291.5998, 291.5998, 291.5998, 291.5998, 291.5998, 
    291.5998, 291.5998, 291.5998, 291.5998, 291.5998, 291.5998, 291.5998, 
    291.5998, 291.5998, 291.5998, 291.5998, 291.5998, 291.5998, 291.5998, 
    291.5998, 291.5998, 291.5998, 291.5998, 291.5998, 291.5998, 291.5998, 
    291.5998, 291.5998, 291.5998, 291.5998, 291.5998, 291.5998, 291.5998, 
    291.5998, 291.5998, 291.5998, 291.5998, 291.5998, 291.5998, 291.5998, 
    291.5998, 291.5998, 291.5998, 291.5998, 291.5998, 291.5998, 291.5998, 
    291.5998, 291.5998, 291.5998, 291.5998, 291.5998, 291.5998,
  292.4925, 292.4925, 292.4925, 292.4925, 292.4925, 292.4925, 292.4925, 
    292.4925, 292.4925, 292.4925, 292.4925, 292.4925, 292.4925, 292.4925, 
    292.4925, 292.4925, 292.4925, 292.4925, 292.4925, 292.4925, 292.4925, 
    292.4925, 292.4925, 292.4925, 292.4925, 292.4925, 292.4925, 292.4925, 
    292.4925, 292.4925, 292.4925, 292.4925, 292.4925, 292.4925, 292.4925, 
    292.4925, 292.4925, 292.4925, 292.4925, 292.4925, 292.4925, 292.4925, 
    292.4925, 292.4925, 292.4925, 292.4925, 292.4925, 292.4925, 292.4925, 
    292.4925, 292.4925, 292.4925, 292.4925, 292.4925, 292.4925, 292.4925, 
    292.4925, 292.4925, 292.4925, 292.4925, 292.4925, 292.4925, 292.4925, 
    292.4925, 292.4925, 292.4925, 292.4925, 292.4925, 292.4925, 292.4925, 
    292.4925, 292.4925, 292.4925, 292.4925, 292.4925, 292.4925, 292.4925, 
    292.4925, 292.4925, 292.4925, 292.4925, 292.4925, 292.4925, 292.4925, 
    292.4925, 292.4925, 292.4925, 292.4925, 292.4925, 292.4925, 292.4925, 
    292.4925, 292.4925, 292.4925, 292.4925, 292.4925, 292.4925,
  293.3779, 293.3779, 293.3779, 293.3779, 293.3779, 293.3779, 293.3779, 
    293.3779, 293.3779, 293.3779, 293.3779, 293.3779, 293.3779, 293.3779, 
    293.3779, 293.3779, 293.3779, 293.3779, 293.3779, 293.3779, 293.3779, 
    293.3779, 293.3779, 293.3779, 293.3779, 293.3779, 293.3779, 293.3779, 
    293.3779, 293.3779, 293.3779, 293.3779, 293.3779, 293.3779, 293.3779, 
    293.3779, 293.3779, 293.3779, 293.3779, 293.3779, 293.3779, 293.3779, 
    293.3779, 293.3779, 293.3779, 293.3779, 293.3779, 293.3779, 293.3779, 
    293.3779, 293.3779, 293.3779, 293.3779, 293.3779, 293.3779, 293.3779, 
    293.3779, 293.3779, 293.3779, 293.3779, 293.3779, 293.3779, 293.3779, 
    293.3779, 293.3779, 293.3779, 293.3779, 293.3779, 293.3779, 293.3779, 
    293.3779, 293.3779, 293.3779, 293.3779, 293.3779, 293.3779, 293.3779, 
    293.3779, 293.3779, 293.3779, 293.3779, 293.3779, 293.3779, 293.3779, 
    293.3779, 293.3779, 293.3779, 293.3779, 293.3779, 293.3779, 293.3779, 
    293.3779, 293.3779, 293.3779, 293.3779, 293.3779, 293.3779,
  294.256, 294.256, 294.256, 294.256, 294.256, 294.256, 294.256, 294.256, 
    294.256, 294.256, 294.256, 294.256, 294.256, 294.256, 294.256, 294.256, 
    294.256, 294.256, 294.256, 294.256, 294.256, 294.256, 294.256, 294.256, 
    294.256, 294.256, 294.256, 294.256, 294.256, 294.256, 294.256, 294.256, 
    294.256, 294.256, 294.256, 294.256, 294.256, 294.256, 294.256, 294.256, 
    294.256, 294.256, 294.256, 294.256, 294.256, 294.256, 294.256, 294.256, 
    294.256, 294.256, 294.256, 294.256, 294.256, 294.256, 294.256, 294.256, 
    294.256, 294.256, 294.256, 294.256, 294.256, 294.256, 294.256, 294.256, 
    294.256, 294.256, 294.256, 294.256, 294.256, 294.256, 294.256, 294.256, 
    294.256, 294.256, 294.256, 294.256, 294.256, 294.256, 294.256, 294.256, 
    294.256, 294.256, 294.256, 294.256, 294.256, 294.256, 294.256, 294.256, 
    294.256, 294.256, 294.256, 294.256, 294.256, 294.256, 294.256, 294.256, 
    294.256,
  295.1267, 295.1267, 295.1267, 295.1267, 295.1267, 295.1267, 295.1267, 
    295.1267, 295.1267, 295.1267, 295.1267, 295.1267, 295.1267, 295.1267, 
    295.1267, 295.1267, 295.1267, 295.1267, 295.1267, 295.1267, 295.1267, 
    295.1267, 295.1267, 295.1267, 295.1267, 295.1267, 295.1267, 295.1267, 
    295.1267, 295.1267, 295.1267, 295.1267, 295.1267, 295.1267, 295.1267, 
    295.1267, 295.1267, 295.1267, 295.1267, 295.1267, 295.1267, 295.1267, 
    295.1267, 295.1267, 295.1267, 295.1267, 295.1267, 295.1267, 295.1267, 
    295.1267, 295.1267, 295.1267, 295.1267, 295.1267, 295.1267, 295.1267, 
    295.1267, 295.1267, 295.1267, 295.1267, 295.1267, 295.1267, 295.1267, 
    295.1267, 295.1267, 295.1267, 295.1267, 295.1267, 295.1267, 295.1267, 
    295.1267, 295.1267, 295.1267, 295.1267, 295.1267, 295.1267, 295.1267, 
    295.1267, 295.1267, 295.1267, 295.1267, 295.1267, 295.1267, 295.1267, 
    295.1267, 295.1267, 295.1267, 295.1267, 295.1267, 295.1267, 295.1267, 
    295.1267, 295.1267, 295.1267, 295.1267, 295.1267, 295.1267,
  295.99, 295.99, 295.99, 295.99, 295.99, 295.99, 295.99, 295.99, 295.99, 
    295.99, 295.99, 295.99, 295.99, 295.99, 295.99, 295.99, 295.99, 295.99, 
    295.99, 295.99, 295.99, 295.99, 295.99, 295.99, 295.99, 295.99, 295.99, 
    295.99, 295.99, 295.99, 295.99, 295.99, 295.99, 295.99, 295.99, 295.99, 
    295.99, 295.99, 295.99, 295.99, 295.99, 295.99, 295.99, 295.99, 295.99, 
    295.99, 295.99, 295.99, 295.99, 295.99, 295.99, 295.99, 295.99, 295.99, 
    295.99, 295.99, 295.99, 295.99, 295.99, 295.99, 295.99, 295.99, 295.99, 
    295.99, 295.99, 295.99, 295.99, 295.99, 295.99, 295.99, 295.99, 295.99, 
    295.99, 295.99, 295.99, 295.99, 295.99, 295.99, 295.99, 295.99, 295.99, 
    295.99, 295.99, 295.99, 295.99, 295.99, 295.99, 295.99, 295.99, 295.99, 
    295.99, 295.99, 295.99, 295.99, 295.99, 295.99, 295.99,
  296.8459, 296.8459, 296.8459, 296.8459, 296.8459, 296.8459, 296.8459, 
    296.8459, 296.8459, 296.8459, 296.8459, 296.8459, 296.8459, 296.8459, 
    296.8459, 296.8459, 296.8459, 296.8459, 296.8459, 296.8459, 296.8459, 
    296.8459, 296.8459, 296.8459, 296.8459, 296.8459, 296.8459, 296.8459, 
    296.8459, 296.8459, 296.8459, 296.8459, 296.8459, 296.8459, 296.8459, 
    296.8459, 296.8459, 296.8459, 296.8459, 296.8459, 296.8459, 296.8459, 
    296.8459, 296.8459, 296.8459, 296.8459, 296.8459, 296.8459, 296.8459, 
    296.8459, 296.8459, 296.8459, 296.8459, 296.8459, 296.8459, 296.8459, 
    296.8459, 296.8459, 296.8459, 296.8459, 296.8459, 296.8459, 296.8459, 
    296.8459, 296.8459, 296.8459, 296.8459, 296.8459, 296.8459, 296.8459, 
    296.8459, 296.8459, 296.8459, 296.8459, 296.8459, 296.8459, 296.8459, 
    296.8459, 296.8459, 296.8459, 296.8459, 296.8459, 296.8459, 296.8459, 
    296.8459, 296.8459, 296.8459, 296.8459, 296.8459, 296.8459, 296.8459, 
    296.8459, 296.8459, 296.8459, 296.8459, 296.8459, 296.8459,
  297.6943, 297.6943, 297.6943, 297.6943, 297.6943, 297.6943, 297.6943, 
    297.6943, 297.6943, 297.6943, 297.6943, 297.6943, 297.6943, 297.6943, 
    297.6943, 297.6943, 297.6943, 297.6943, 297.6943, 297.6943, 297.6943, 
    297.6943, 297.6943, 297.6943, 297.6943, 297.6943, 297.6943, 297.6943, 
    297.6943, 297.6943, 297.6943, 297.6943, 297.6943, 297.6943, 297.6943, 
    297.6943, 297.6943, 297.6943, 297.6943, 297.6943, 297.6943, 297.6943, 
    297.6943, 297.6943, 297.6943, 297.6943, 297.6943, 297.6943, 297.6943, 
    297.6943, 297.6943, 297.6943, 297.6943, 297.6943, 297.6943, 297.6943, 
    297.6943, 297.6943, 297.6943, 297.6943, 297.6943, 297.6943, 297.6943, 
    297.6943, 297.6943, 297.6943, 297.6943, 297.6943, 297.6943, 297.6943, 
    297.6943, 297.6943, 297.6943, 297.6943, 297.6943, 297.6943, 297.6943, 
    297.6943, 297.6943, 297.6943, 297.6943, 297.6943, 297.6943, 297.6943, 
    297.6943, 297.6943, 297.6943, 297.6943, 297.6943, 297.6943, 297.6943, 
    297.6943, 297.6943, 297.6943, 297.6943, 297.6943, 297.6943,
  298.5354, 298.5354, 298.5354, 298.5354, 298.5354, 298.5354, 298.5354, 
    298.5354, 298.5354, 298.5354, 298.5354, 298.5354, 298.5354, 298.5354, 
    298.5354, 298.5354, 298.5354, 298.5354, 298.5354, 298.5354, 298.5354, 
    298.5354, 298.5354, 298.5354, 298.5354, 298.5354, 298.5354, 298.5354, 
    298.5354, 298.5354, 298.5354, 298.5354, 298.5354, 298.5354, 298.5354, 
    298.5354, 298.5354, 298.5354, 298.5354, 298.5354, 298.5354, 298.5354, 
    298.5354, 298.5354, 298.5354, 298.5354, 298.5354, 298.5354, 298.5354, 
    298.5354, 298.5354, 298.5354, 298.5354, 298.5354, 298.5354, 298.5354, 
    298.5354, 298.5354, 298.5354, 298.5354, 298.5354, 298.5354, 298.5354, 
    298.5354, 298.5354, 298.5354, 298.5354, 298.5354, 298.5354, 298.5354, 
    298.5354, 298.5354, 298.5354, 298.5354, 298.5354, 298.5354, 298.5354, 
    298.5354, 298.5354, 298.5354, 298.5354, 298.5354, 298.5354, 298.5354, 
    298.5354, 298.5354, 298.5354, 298.5354, 298.5354, 298.5354, 298.5354, 
    298.5354, 298.5354, 298.5354, 298.5354, 298.5354, 298.5354,
  299.3691, 299.3691, 299.3691, 299.3691, 299.3691, 299.3691, 299.3691, 
    299.3691, 299.3691, 299.3691, 299.3691, 299.3691, 299.3691, 299.3691, 
    299.3691, 299.3691, 299.3691, 299.3691, 299.3691, 299.3691, 299.3691, 
    299.3691, 299.3691, 299.3691, 299.3691, 299.3691, 299.3691, 299.3691, 
    299.3691, 299.3691, 299.3691, 299.3691, 299.3691, 299.3691, 299.3691, 
    299.3691, 299.3691, 299.3691, 299.3691, 299.3691, 299.3691, 299.3691, 
    299.3691, 299.3691, 299.3691, 299.3691, 299.3691, 299.3691, 299.3691, 
    299.3691, 299.3691, 299.3691, 299.3691, 299.3691, 299.3691, 299.3691, 
    299.3691, 299.3691, 299.3691, 299.3691, 299.3691, 299.3691, 299.3691, 
    299.3691, 299.3691, 299.3691, 299.3691, 299.3691, 299.3691, 299.3691, 
    299.3691, 299.3691, 299.3691, 299.3691, 299.3691, 299.3691, 299.3691, 
    299.3691, 299.3691, 299.3691, 299.3691, 299.3691, 299.3691, 299.3691, 
    299.3691, 299.3691, 299.3691, 299.3691, 299.3691, 299.3691, 299.3691, 
    299.3691, 299.3691, 299.3691, 299.3691, 299.3691, 299.3691,
  300.1953, 300.1953, 300.1953, 300.1953, 300.1953, 300.1953, 300.1953, 
    300.1953, 300.1953, 300.1953, 300.1953, 300.1953, 300.1953, 300.1953, 
    300.1953, 300.1953, 300.1953, 300.1953, 300.1953, 300.1953, 300.1953, 
    300.1953, 300.1953, 300.1953, 300.1953, 300.1953, 300.1953, 300.1953, 
    300.1953, 300.1953, 300.1953, 300.1953, 300.1953, 300.1953, 300.1953, 
    300.1953, 300.1953, 300.1953, 300.1953, 300.1953, 300.1953, 300.1953, 
    300.1953, 300.1953, 300.1953, 300.1953, 300.1953, 300.1953, 300.1953, 
    300.1953, 300.1953, 300.1953, 300.1953, 300.1953, 300.1953, 300.1953, 
    300.1953, 300.1953, 300.1953, 300.1953, 300.1953, 300.1953, 300.1953, 
    300.1953, 300.1953, 300.1953, 300.1953, 300.1953, 300.1953, 300.1953, 
    300.1953, 300.1953, 300.1953, 300.1953, 300.1953, 300.1953, 300.1953, 
    300.1953, 300.1953, 300.1953, 300.1953, 300.1953, 300.1953, 300.1953, 
    300.1953, 300.1953, 300.1953, 300.1953, 300.1953, 300.1953, 300.1953, 
    300.1953, 300.1953, 300.1953, 300.1953, 300.1953, 300.1953,
  301.0143, 301.0143, 301.0143, 301.0143, 301.0143, 301.0143, 301.0143, 
    301.0143, 301.0143, 301.0143, 301.0143, 301.0143, 301.0143, 301.0143, 
    301.0143, 301.0143, 301.0143, 301.0143, 301.0143, 301.0143, 301.0143, 
    301.0143, 301.0143, 301.0143, 301.0143, 301.0143, 301.0143, 301.0143, 
    301.0143, 301.0143, 301.0143, 301.0143, 301.0143, 301.0143, 301.0143, 
    301.0143, 301.0143, 301.0143, 301.0143, 301.0143, 301.0143, 301.0143, 
    301.0143, 301.0143, 301.0143, 301.0143, 301.0143, 301.0143, 301.0143, 
    301.0143, 301.0143, 301.0143, 301.0143, 301.0143, 301.0143, 301.0143, 
    301.0143, 301.0143, 301.0143, 301.0143, 301.0143, 301.0143, 301.0143, 
    301.0143, 301.0143, 301.0143, 301.0143, 301.0143, 301.0143, 301.0143, 
    301.0143, 301.0143, 301.0143, 301.0143, 301.0143, 301.0143, 301.0143, 
    301.0143, 301.0143, 301.0143, 301.0143, 301.0143, 301.0143, 301.0143, 
    301.0143, 301.0143, 301.0143, 301.0143, 301.0143, 301.0143, 301.0143, 
    301.0143, 301.0143, 301.0143, 301.0143, 301.0143, 301.0143,
  301.8259, 301.8259, 301.8259, 301.8259, 301.8259, 301.8259, 301.8259, 
    301.8259, 301.8259, 301.8259, 301.8259, 301.8259, 301.8259, 301.8259, 
    301.8259, 301.8259, 301.8259, 301.8259, 301.8259, 301.8259, 301.8259, 
    301.8259, 301.8259, 301.8259, 301.8259, 301.8259, 301.8259, 301.8259, 
    301.8259, 301.8259, 301.8259, 301.8259, 301.8259, 301.8259, 301.8259, 
    301.8259, 301.8259, 301.8259, 301.8259, 301.8259, 301.8259, 301.8259, 
    301.8259, 301.8259, 301.8259, 301.8259, 301.8259, 301.8259, 301.8259, 
    301.8259, 301.8259, 301.8259, 301.8259, 301.8259, 301.8259, 301.8259, 
    301.8259, 301.8259, 301.8259, 301.8259, 301.8259, 301.8259, 301.8259, 
    301.8259, 301.8259, 301.8259, 301.8259, 301.8259, 301.8259, 301.8259, 
    301.8259, 301.8259, 301.8259, 301.8259, 301.8259, 301.8259, 301.8259, 
    301.8259, 301.8259, 301.8259, 301.8259, 301.8259, 301.8259, 301.8259, 
    301.8259, 301.8259, 301.8259, 301.8259, 301.8259, 301.8259, 301.8259, 
    301.8259, 301.8259, 301.8259, 301.8259, 301.8259, 301.8259,
  302.6302, 302.6302, 302.6302, 302.6302, 302.6302, 302.6302, 302.6302, 
    302.6302, 302.6302, 302.6302, 302.6302, 302.6302, 302.6302, 302.6302, 
    302.6302, 302.6302, 302.6302, 302.6302, 302.6302, 302.6302, 302.6302, 
    302.6302, 302.6302, 302.6302, 302.6302, 302.6302, 302.6302, 302.6302, 
    302.6302, 302.6302, 302.6302, 302.6302, 302.6302, 302.6302, 302.6302, 
    302.6302, 302.6302, 302.6302, 302.6302, 302.6302, 302.6302, 302.6302, 
    302.6302, 302.6302, 302.6302, 302.6302, 302.6302, 302.6302, 302.6302, 
    302.6302, 302.6302, 302.6302, 302.6302, 302.6302, 302.6302, 302.6302, 
    302.6302, 302.6302, 302.6302, 302.6302, 302.6302, 302.6302, 302.6302, 
    302.6302, 302.6302, 302.6302, 302.6302, 302.6302, 302.6302, 302.6302, 
    302.6302, 302.6302, 302.6302, 302.6302, 302.6302, 302.6302, 302.6302, 
    302.6302, 302.6302, 302.6302, 302.6302, 302.6302, 302.6302, 302.6302, 
    302.6302, 302.6302, 302.6302, 302.6302, 302.6302, 302.6302, 302.6302, 
    302.6302, 302.6302, 302.6302, 302.6302, 302.6302, 302.6302,
  303.4273, 303.4273, 303.4273, 303.4273, 303.4273, 303.4273, 303.4273, 
    303.4273, 303.4273, 303.4273, 303.4273, 303.4273, 303.4273, 303.4273, 
    303.4273, 303.4273, 303.4273, 303.4273, 303.4273, 303.4273, 303.4273, 
    303.4273, 303.4273, 303.4273, 303.4273, 303.4273, 303.4273, 303.4273, 
    303.4273, 303.4273, 303.4273, 303.4273, 303.4273, 303.4273, 303.4273, 
    303.4273, 303.4273, 303.4273, 303.4273, 303.4273, 303.4273, 303.4273, 
    303.4273, 303.4273, 303.4273, 303.4273, 303.4273, 303.4273, 303.4273, 
    303.4273, 303.4273, 303.4273, 303.4273, 303.4273, 303.4273, 303.4273, 
    303.4273, 303.4273, 303.4273, 303.4273, 303.4273, 303.4273, 303.4273, 
    303.4273, 303.4273, 303.4273, 303.4273, 303.4273, 303.4273, 303.4273, 
    303.4273, 303.4273, 303.4273, 303.4273, 303.4273, 303.4273, 303.4273, 
    303.4273, 303.4273, 303.4273, 303.4273, 303.4273, 303.4273, 303.4273, 
    303.4273, 303.4273, 303.4273, 303.4273, 303.4273, 303.4273, 303.4273, 
    303.4273, 303.4273, 303.4273, 303.4273, 303.4273, 303.4273,
  304.2172, 304.2172, 304.2172, 304.2172, 304.2172, 304.2172, 304.2172, 
    304.2172, 304.2172, 304.2172, 304.2172, 304.2172, 304.2172, 304.2172, 
    304.2172, 304.2172, 304.2172, 304.2172, 304.2172, 304.2172, 304.2172, 
    304.2172, 304.2172, 304.2172, 304.2172, 304.2172, 304.2172, 304.2172, 
    304.2172, 304.2172, 304.2172, 304.2172, 304.2172, 304.2172, 304.2172, 
    304.2172, 304.2172, 304.2172, 304.2172, 304.2172, 304.2172, 304.2172, 
    304.2172, 304.2172, 304.2172, 304.2172, 304.2172, 304.2172, 304.2172, 
    304.2172, 304.2172, 304.2172, 304.2172, 304.2172, 304.2172, 304.2172, 
    304.2172, 304.2172, 304.2172, 304.2172, 304.2172, 304.2172, 304.2172, 
    304.2172, 304.2172, 304.2172, 304.2172, 304.2172, 304.2172, 304.2172, 
    304.2172, 304.2172, 304.2172, 304.2172, 304.2172, 304.2172, 304.2172, 
    304.2172, 304.2172, 304.2172, 304.2172, 304.2172, 304.2172, 304.2172, 
    304.2172, 304.2172, 304.2172, 304.2172, 304.2172, 304.2172, 304.2172, 
    304.2172, 304.2172, 304.2172, 304.2172, 304.2172, 304.2172,
  305, 305, 305, 305, 305, 305, 305, 305, 305, 305, 305, 305, 305, 305, 305, 
    305, 305, 305, 305, 305, 305, 305, 305, 305, 305, 305, 305, 305, 305, 
    305, 305, 305, 305, 305, 305, 305, 305, 305, 305, 305, 305, 305, 305, 
    305, 305, 305, 305, 305, 305, 305, 305, 305, 305, 305, 305, 305, 305, 
    305, 305, 305, 305, 305, 305, 305, 305, 305, 305, 305, 305, 305, 305, 
    305, 305, 305, 305, 305, 305, 305, 305, 305, 305, 305, 305, 305, 305, 
    305, 305, 305, 305, 305, 305, 305, 305, 305, 305, 305, 305 ;

 grid_lat =
  35.26439, 34.52972, 33.79504, 33.06036, 32.32569, 31.59101, 30.85634, 
    30.12167, 29.38699, 28.65232, 27.91764, 27.18297, 26.44829, 25.71362, 
    24.97894, 24.24427, 23.50959, 22.77492, 22.04024, 21.30557, 20.57089, 
    19.83622, 19.10155, 18.36687, 17.63219, 16.89752, 16.16285, 15.42817, 
    14.6935, 13.95882, 13.22415, 12.48947, 11.7548, 11.02012, 10.28545, 
    9.550773, 8.816097, 8.081423, 7.346748, 6.612073, 5.877398, 5.142724, 
    4.408049, 3.673374, 2.938699, 2.204024, 1.46935, 0.7346748, 1.272222e-14, 
    -0.7346748, -1.46935, -2.204024, -2.938699, -3.673374, -4.408049, 
    -5.142724, -5.877398, -6.612073, -7.346748, -8.081423, -8.816097, 
    -9.550773, -10.28545, -11.02012, -11.7548, -12.48947, -13.22415, 
    -13.95882, -14.6935, -15.42817, -16.16285, -16.89752, -17.63219, 
    -18.36687, -19.10155, -19.83622, -20.57089, -21.30557, -22.04024, 
    -22.77492, -23.50959, -24.24427, -24.97894, -25.71362, -26.44829, 
    -27.18297, -27.91764, -28.65232, -29.38699, -30.12167, -30.85634, 
    -31.59101, -32.32569, -33.06036, -33.79504, -34.52972, -35.26439,
  35.62921, 34.89117, 34.15289, 33.41436, 32.67561, 31.93662, 31.19741, 
    30.45796, 29.7183, 28.97841, 28.23831, 27.49799, 26.75747, 26.01674, 
    25.2758, 24.53467, 23.79335, 23.05183, 22.31014, 21.56826, 20.8262, 
    20.08398, 19.34159, 18.59904, 17.85633, 17.11348, 16.37048, 15.62734, 
    14.88407, 14.14067, 13.39715, 12.65351, 11.90976, 11.16591, 10.42197, 
    9.677926, 8.933801, 8.189597, 7.445321, 6.700978, 5.956575, 5.21212, 
    4.467618, 3.723077, 2.978501, 2.233899, 1.489277, 0.744642, 0, -0.744642, 
    -1.489277, -2.233899, -2.978501, -3.723077, -4.467618, -5.21212, 
    -5.956575, -6.700978, -7.445321, -8.189597, -8.933801, -9.677926, 
    -10.42197, -11.16591, -11.90976, -12.65351, -13.39715, -14.14067, 
    -14.88407, -15.62734, -16.37048, -17.11348, -17.85633, -18.59904, 
    -19.34159, -20.08398, -20.8262, -21.56826, -22.31014, -23.05183, 
    -23.79335, -24.53467, -25.2758, -26.01674, -26.75747, -27.49799, 
    -28.23831, -28.97841, -29.7183, -30.45796, -31.19741, -31.93662, 
    -32.67561, -33.41436, -34.15289, -34.89117, -35.62921,
  35.98892, 35.24767, 34.50594, 33.76374, 33.02107, 32.27793, 31.53433, 
    30.79028, 30.04578, 29.30084, 28.55546, 27.80966, 27.06343, 26.31679, 
    25.56974, 24.82229, 24.07445, 23.32623, 22.57764, 21.82868, 21.07937, 
    20.32972, 19.57973, 18.82941, 18.07879, 17.32786, 16.57663, 15.82513, 
    15.07335, 14.32132, 13.56903, 12.81652, 12.06378, 11.31083, 10.55768, 
    9.804344, 9.050837, 8.297169, 7.543353, 6.789403, 6.035332, 5.281153, 
    4.526879, 3.772523, 3.0181, 2.263623, 1.509105, 0.7545591, 0, -0.7545591, 
    -1.509105, -2.263623, -3.0181, -3.772523, -4.526879, -5.281153, 
    -6.035332, -6.789403, -7.543353, -8.297169, -9.050837, -9.804344, 
    -10.55768, -11.31083, -12.06378, -12.81652, -13.56903, -14.32132, 
    -15.07335, -15.82513, -16.57663, -17.32786, -18.07879, -18.82941, 
    -19.57973, -20.32972, -21.07937, -21.82868, -22.57764, -23.32623, 
    -24.07445, -24.82229, -25.56974, -26.31679, -27.06343, -27.80966, 
    -28.55546, -29.30084, -30.04578, -30.79028, -31.53433, -32.27793, 
    -33.02107, -33.76374, -34.50594, -35.24767, -35.98892,
  36.34341, 35.59911, 34.8541, 34.10837, 33.36194, 32.61481, 31.86699, 
    31.11849, 30.36931, 29.61947, 28.86897, 28.11782, 27.36604, 26.61363, 
    25.86061, 25.10699, 24.35277, 23.59798, 22.84263, 22.08672, 21.33028, 
    20.57332, 19.81585, 19.05788, 18.29944, 17.54054, 16.7812, 16.02143, 
    15.26124, 14.50067, 13.73972, 12.97841, 12.21676, 11.45479, 10.69252, 
    9.929964, 9.167146, 8.404083, 7.640796, 6.877304, 6.113627, 5.349786, 
    4.5858, 3.82169, 3.057476, 2.29318, 1.528821, 0.7644209, 0, -0.7644209, 
    -1.528821, -2.29318, -3.057476, -3.82169, -4.5858, -5.349786, -6.113627, 
    -6.877304, -7.640796, -8.404083, -9.167146, -9.929964, -10.69252, 
    -11.45479, -12.21676, -12.97841, -13.73972, -14.50067, -15.26124, 
    -16.02143, -16.7812, -17.54054, -18.29944, -19.05788, -19.81585, 
    -20.57332, -21.33028, -22.08672, -22.84263, -23.59798, -24.35277, 
    -25.10699, -25.86061, -26.61363, -27.36604, -28.11782, -28.86897, 
    -29.61947, -30.36931, -31.11849, -31.86699, -32.61481, -33.36194, 
    -34.10837, -34.8541, -35.59911, -36.34341,
  36.69255, 35.94537, 35.19722, 34.44813, 33.6981, 32.94714, 32.19525, 
    31.44245, 30.68875, 29.93416, 29.17869, 28.42235, 27.66517, 26.90714, 
    26.14829, 25.38863, 24.62818, 23.86696, 23.10497, 22.34225, 21.5788, 
    20.81466, 20.04982, 19.28433, 18.51819, 17.75143, 16.98408, 16.21614, 
    15.44765, 14.67863, 13.90911, 13.1391, 12.36863, 11.59772, 10.82641, 
    10.05472, 9.282667, 8.510284, 7.737598, 6.964634, 6.19142, 5.417983, 
    4.64435, 3.870549, 3.096608, 2.322554, 1.548416, 0.7742223, 0, 
    -0.7742223, -1.548416, -2.322554, -3.096608, -3.870549, -4.64435, 
    -5.417983, -6.19142, -6.964634, -7.737598, -8.510284, -9.282667, 
    -10.05472, -10.82641, -11.59772, -12.36863, -13.1391, -13.90911, 
    -14.67863, -15.44765, -16.21614, -16.98408, -17.75143, -18.51819, 
    -19.28433, -20.04982, -20.81466, -21.5788, -22.34225, -23.10497, 
    -23.86696, -24.62818, -25.38863, -26.14829, -26.90714, -27.66517, 
    -28.42235, -29.17869, -29.93416, -30.68875, -31.44245, -32.19525, 
    -32.94714, -33.6981, -34.44813, -35.19722, -35.94537, -36.69255,
  37.03624, 36.28631, 35.53519, 34.78289, 34.02942, 33.27477, 32.51897, 
    31.76203, 31.00396, 30.24478, 29.48449, 28.72311, 27.96067, 27.19717, 
    26.43264, 25.66709, 24.90054, 24.13302, 23.36455, 22.59513, 21.82482, 
    21.05361, 20.28154, 19.50863, 18.73492, 17.96042, 17.18516, 16.40917, 
    15.63248, 14.85512, 14.07711, 13.2985, 12.5193, 11.73955, 10.95929, 
    10.17854, 9.397336, 8.615713, 7.833705, 7.051345, 6.268667, 5.485706, 
    4.702497, 3.919074, 3.135473, 2.35173, 1.56788, 0.7839577, 0, -0.7839577, 
    -1.56788, -2.35173, -3.135473, -3.919074, -4.702497, -5.485706, 
    -6.268667, -7.051345, -7.833705, -8.615713, -9.397336, -10.17854, 
    -10.95929, -11.73955, -12.5193, -13.2985, -14.07711, -14.85512, 
    -15.63248, -16.40917, -17.18516, -17.96042, -18.73492, -19.50863, 
    -20.28154, -21.05361, -21.82482, -22.59513, -23.36455, -24.13302, 
    -24.90054, -25.66709, -26.43264, -27.19717, -27.96067, -28.72311, 
    -29.48449, -30.24478, -31.00396, -31.76203, -32.51897, -33.27477, 
    -34.02942, -34.78289, -35.53519, -36.28631, -37.03624,
  37.37434, 36.62183, 35.86789, 35.11252, 34.35575, 33.59758, 32.83802, 
    32.0771, 31.31481, 30.55118, 29.78622, 29.01996, 28.25241, 27.48358, 
    26.71351, 25.94222, 25.16972, 24.39604, 23.6212, 22.84524, 22.06818, 
    21.29005, 20.51087, 19.73068, 18.9495, 18.16737, 17.38433, 16.6004, 
    15.81561, 15.03002, 14.24364, 13.45652, 12.66869, 11.88019, 11.09107, 
    10.30135, 9.511086, 8.720308, 7.929061, 7.137385, 6.345323, 5.552916, 
    4.760206, 3.967237, 3.17405, 2.38069, 1.587199, 0.7936214, 0, -0.7936214, 
    -1.587199, -2.38069, -3.17405, -3.967237, -4.760206, -5.552916, 
    -6.345323, -7.137385, -7.929061, -8.720308, -9.511086, -10.30135, 
    -11.09107, -11.88019, -12.66869, -13.45652, -14.24364, -15.03002, 
    -15.81561, -16.6004, -17.38433, -18.16737, -18.9495, -19.73068, 
    -20.51087, -21.29005, -22.06818, -22.84524, -23.6212, -24.39604, 
    -25.16972, -25.94222, -26.71351, -27.48358, -28.25241, -29.01996, 
    -29.78622, -30.55118, -31.31481, -32.0771, -32.83802, -33.59758, 
    -34.35575, -35.11252, -35.86789, -36.62183, -37.37434,
  37.70675, 36.95179, 36.19517, 35.4369, 34.67698, 33.91543, 33.15226, 
    32.3875, 31.62114, 30.85322, 30.08375, 29.31275, 28.54023, 27.76624, 
    26.99077, 26.21387, 25.43556, 24.65587, 23.87482, 23.09244, 22.30877, 
    21.52384, 20.73768, 19.95033, 19.16182, 18.37219, 17.58147, 16.78971, 
    15.99695, 15.20323, 14.40859, 13.61306, 12.81671, 12.01956, 11.22167, 
    10.42309, 9.623848, 8.824006, 8.023608, 7.222704, 6.421341, 5.619571, 
    4.817443, 4.015007, 3.212315, 2.409416, 1.606363, 0.8032075, 0, 
    -0.8032075, -1.606363, -2.409416, -3.212315, -4.015007, -4.817443, 
    -5.619571, -6.421341, -7.222704, -8.023608, -8.824006, -9.623848, 
    -10.42309, -11.22167, -12.01956, -12.81671, -13.61306, -14.40859, 
    -15.20323, -15.99695, -16.78971, -17.58147, -18.37219, -19.16182, 
    -19.95033, -20.73768, -21.52384, -22.30877, -23.09244, -23.87482, 
    -24.65587, -25.43556, -26.21387, -26.99077, -27.76624, -28.54023, 
    -29.31275, -30.08375, -30.85322, -31.62114, -32.3875, -33.15226, 
    -33.91543, -34.67698, -35.4369, -36.19517, -36.95179, -37.70675,
  38.03334, 37.27608, 36.51693, 35.75588, 34.99296, 34.22818, 33.46156, 
    32.6931, 31.92283, 31.15076, 30.37692, 29.60133, 28.82401, 28.04498, 
    27.26427, 26.48191, 25.69794, 24.91236, 24.12524, 23.33659, 22.54645, 
    21.75485, 20.96184, 20.16746, 19.37174, 18.57473, 17.77647, 16.97701, 
    16.17639, 15.37465, 14.57185, 13.76804, 12.96326, 12.15757, 11.35102, 
    10.54366, 9.735553, 8.926742, 8.117288, 7.307246, 6.496675, 5.68563, 
    4.874171, 4.062356, 3.250242, 2.437891, 1.62536, 0.8127099, 0, 
    -0.8127099, -1.62536, -2.437891, -3.250242, -4.062356, -4.874171, 
    -5.68563, -6.496675, -7.307246, -8.117288, -8.926742, -9.735553, 
    -10.54366, -11.35102, -12.15757, -12.96326, -13.76804, -14.57185, 
    -15.37465, -16.17639, -16.97701, -17.77647, -18.57473, -19.37174, 
    -20.16746, -20.96184, -21.75485, -22.54645, -23.33659, -24.12524, 
    -24.91236, -25.69794, -26.48191, -27.26427, -28.04498, -28.82401, 
    -29.60133, -30.37692, -31.15076, -31.92283, -32.6931, -33.46156, 
    -34.22818, -34.99296, -35.75588, -36.51693, -37.27608, -38.03334,
  38.354, 37.59457, 36.83301, 36.06934, 35.30357, 34.5357, 33.76576, 
    32.99376, 32.21972, 31.44366, 30.6656, 29.88556, 29.10357, 28.31966, 
    27.53386, 26.74619, 25.95669, 25.16539, 24.37232, 23.57754, 22.78106, 
    21.98295, 21.18322, 20.38194, 19.57915, 18.77489, 17.96921, 17.16216, 
    16.3538, 15.54417, 14.73334, 13.92135, 13.10826, 12.29414, 11.47903, 
    10.66301, 9.846126, 9.028447, 8.210036, 7.390956, 6.571271, 5.751048, 
    4.930352, 4.10925, 3.287808, 2.466094, 1.644176, 0.8221223, 0, 
    -0.8221223, -1.644176, -2.466094, -3.287808, -4.10925, -4.930352, 
    -5.751048, -6.571271, -7.390956, -8.210036, -9.028447, -9.846126, 
    -10.66301, -11.47903, -12.29414, -13.10826, -13.92135, -14.73334, 
    -15.54417, -16.3538, -17.16216, -17.96921, -18.77489, -19.57915, 
    -20.38194, -21.18322, -21.98295, -22.78106, -23.57754, -24.37232, 
    -25.16539, -25.95669, -26.74619, -27.53386, -28.31966, -29.10357, 
    -29.88556, -30.6656, -31.44366, -32.21972, -32.99376, -33.76576, 
    -34.5357, -35.30357, -36.06934, -36.83301, -37.59457, -38.354,
  38.66859, 37.90713, 37.14331, 36.37715, 35.60866, 34.83784, 34.06473, 
    33.28933, 32.51167, 31.73176, 30.94962, 30.16529, 29.37879, 28.59014, 
    27.79938, 27.00655, 26.21167, 25.41478, 24.61593, 23.81515, 23.01249, 
    22.20798, 21.40168, 20.59364, 19.7839, 18.97252, 18.15956, 17.34505, 
    16.52908, 15.71168, 14.89293, 14.07288, 13.2516, 12.42916, 11.60561, 
    10.78103, 9.955491, 9.129053, 8.30179, 7.473776, 6.645081, 5.815781, 
    4.985948, 4.155657, 3.324986, 2.494007, 1.662799, 0.8314381, 0, 
    -0.8314381, -1.662799, -2.494007, -3.324986, -4.155657, -4.985948, 
    -5.815781, -6.645081, -7.473776, -8.30179, -9.129053, -9.955491, 
    -10.78103, -11.60561, -12.42916, -13.2516, -14.07288, -14.89293, 
    -15.71168, -16.52908, -17.34505, -18.15956, -18.97252, -19.7839, 
    -20.59364, -21.40168, -22.20798, -23.01249, -23.81515, -24.61593, 
    -25.41478, -26.21167, -27.00655, -27.79938, -28.59014, -29.37879, 
    -30.16529, -30.94962, -31.73176, -32.51167, -33.28933, -34.06473, 
    -34.83784, -35.60866, -36.37715, -37.14331, -37.90713, -38.66859,
  38.977, 38.21363, 37.44768, 36.67916, 35.90809, 35.13448, 34.35833, 
    33.57967, 32.79853, 32.01491, 31.22885, 30.44036, 29.64949, 28.85626, 
    28.0607, 27.26284, 26.46273, 25.6604, 24.85591, 24.04927, 23.24056, 
    22.42981, 21.61708, 20.80241, 19.98587, 19.16751, 18.34738, 17.52556, 
    16.7021, 15.87706, 15.05052, 14.22254, 13.39319, 12.56255, 11.73068, 
    10.89766, 10.06357, 9.228487, 8.392486, 7.555646, 6.718051, 5.87978, 
    5.040917, 4.201545, 3.361748, 2.52161, 1.681216, 0.8406506, 0, 
    -0.8406506, -1.681216, -2.52161, -3.361748, -4.201545, -5.040917, 
    -5.87978, -6.718051, -7.555646, -8.392486, -9.228487, -10.06357, 
    -10.89766, -11.73068, -12.56255, -13.39319, -14.22254, -15.05052, 
    -15.87706, -16.7021, -17.52556, -18.34738, -19.16751, -19.98587, 
    -20.80241, -21.61708, -22.42981, -23.24056, -24.04927, -24.85591, 
    -25.6604, -26.46273, -27.26284, -28.0607, -28.85626, -29.64949, 
    -30.44036, -31.22885, -32.01491, -32.79853, -33.57967, -34.35833, 
    -35.13448, -35.90809, -36.67916, -37.44768, -38.21363, -38.977,
  39.27911, 38.51395, 37.746, 36.97525, 36.20173, 35.42545, 34.64641, 
    33.86464, 33.08015, 32.29297, 31.50312, 30.71063, 29.91554, 29.11786, 
    28.31764, 27.51491, 26.70972, 25.9021, 25.0921, 24.27976, 23.46515, 
    22.6483, 21.82927, 21.00812, 20.18491, 19.35971, 18.53256, 17.70355, 
    16.87274, 16.0402, 15.20599, 14.37021, 13.53292, 12.6942, 11.85414, 
    11.0128, 10.17029, 9.326677, 8.482054, 7.636507, 6.790126, 5.943, 
    5.095221, 4.246879, 3.398068, 2.548881, 1.699411, 0.8497528, 0, 
    -0.8497528, -1.699411, -2.548881, -3.398068, -4.246879, -5.095221, 
    -5.943, -6.790126, -7.636507, -8.482054, -9.326677, -10.17029, -11.0128, 
    -11.85414, -12.6942, -13.53292, -14.37021, -15.20599, -16.0402, 
    -16.87274, -17.70355, -18.53256, -19.35971, -20.18491, -21.00812, 
    -21.82927, -22.6483, -23.46515, -24.27976, -25.0921, -25.9021, -26.70972, 
    -27.51491, -28.31764, -29.11786, -29.91554, -30.71063, -31.50312, 
    -32.29297, -33.08015, -33.86464, -34.64641, -35.42545, -36.20173, 
    -36.97525, -37.746, -38.51395, -39.27911,
  39.57478, 38.80796, 38.03813, 37.26529, 36.48944, 35.71062, 34.92882, 
    34.14407, 33.35638, 32.56578, 31.77229, 30.97594, 30.17676, 29.37479, 
    28.57006, 27.76261, 26.95247, 26.13971, 25.32435, 24.50646, 23.68609, 
    22.86328, 22.03811, 21.21062, 20.38089, 19.54898, 18.71496, 17.8789, 
    17.04088, 16.20097, 15.35924, 14.51579, 13.67069, 12.82403, 11.97589, 
    11.12637, 10.27556, 9.423547, 8.570426, 7.716295, 6.86125, 6.00539, 
    5.148814, 4.291623, 3.433917, 2.575799, 1.717372, 0.8587376, 0, 
    -0.8587376, -1.717372, -2.575799, -3.433917, -4.291623, -5.148814, 
    -6.00539, -6.86125, -7.716295, -8.570426, -9.423547, -10.27556, 
    -11.12637, -11.97589, -12.82403, -13.67069, -14.51579, -15.35924, 
    -16.20097, -17.04088, -17.8789, -18.71496, -19.54898, -20.38089, 
    -21.21062, -22.03811, -22.86328, -23.68609, -24.50646, -25.32435, 
    -26.13971, -26.95247, -27.76261, -28.57006, -29.37479, -30.17676, 
    -30.97594, -31.77229, -32.56578, -33.35638, -34.14407, -34.92882, 
    -35.71062, -36.48944, -37.26529, -38.03813, -38.80796, -39.57478,
  39.8639, 39.09554, 38.32394, 37.54912, 36.77109, 35.98985, 35.20542, 
    34.41782, 33.62707, 32.83318, 32.03619, 31.23613, 30.43301, 29.62689, 
    28.81779, 28.00576, 27.19084, 26.37307, 25.55252, 24.72922, 23.90323, 
    23.07462, 22.24345, 21.40977, 20.57367, 19.7352, 18.89445, 18.05148, 
    17.20639, 16.35925, 15.51014, 14.65916, 13.80638, 12.95192, 12.09585, 
    11.23828, 10.3793, 9.519018, 8.657532, 7.794946, 6.931367, 6.066901, 
    5.201655, 4.335741, 3.469266, 2.602343, 1.735083, 0.8675976, 0, 
    -0.8675976, -1.735083, -2.602343, -3.469266, -4.335741, -5.201655, 
    -6.066901, -6.931367, -7.794946, -8.657532, -9.519018, -10.3793, 
    -11.23828, -12.09585, -12.95192, -13.80638, -14.65916, -15.51014, 
    -16.35925, -17.20639, -18.05148, -18.89445, -19.7352, -20.57367, 
    -21.40977, -22.24345, -23.07462, -23.90323, -24.72922, -25.55252, 
    -26.37307, -27.19084, -28.00576, -28.81779, -29.62689, -30.43301, 
    -31.23613, -32.03619, -32.83318, -33.62707, -34.41782, -35.20542, 
    -35.98985, -36.77109, -37.54912, -38.32394, -39.09554, -39.8639,
  40.14635, 39.37654, 38.6033, 37.82662, 37.04652, 36.26299, 35.47607, 
    34.68575, 33.89207, 33.09504, 32.29469, 31.49104, 30.68413, 29.874, 
    29.06068, 28.24422, 27.42466, 26.60204, 25.77643, 24.94787, 24.11643, 
    23.28216, 22.44514, 21.60542, 20.76309, 19.91821, 19.07088, 18.22116, 
    17.36914, 16.51492, 15.65857, 14.8002, 13.9399, 13.07777, 12.21391, 
    11.34843, 10.48143, 9.613013, 8.743299, 7.872395, 7.000417, 6.12748, 
    5.253699, 4.379195, 3.504085, 2.628489, 1.752529, 0.8763254, 0, 
    -0.8763254, -1.752529, -2.628489, -3.504085, -4.379195, -5.253699, 
    -6.12748, -7.000417, -7.872395, -8.743299, -9.613013, -10.48143, 
    -11.34843, -12.21391, -13.07777, -13.9399, -14.8002, -15.65857, 
    -16.51492, -17.36914, -18.22116, -19.07088, -19.91821, -20.76309, 
    -21.60542, -22.44514, -23.28216, -24.11643, -24.94787, -25.77643, 
    -26.60204, -27.42466, -28.24422, -29.06068, -29.874, -30.68413, 
    -31.49104, -32.29469, -33.09504, -33.89207, -34.68575, -35.47607, 
    -36.26299, -37.04652, -37.82662, -38.6033, -39.37654, -40.14635,
  40.42199, 39.65086, 38.87608, 38.09766, 37.3156, 36.52991, 35.74061, 
    34.94771, 34.15122, 33.35118, 32.5476, 31.74052, 30.92996, 30.11596, 
    29.29857, 28.47782, 27.65377, 26.82645, 25.99593, 25.16227, 24.32551, 
    23.48574, 22.64302, 21.79742, 20.94901, 20.09789, 19.24412, 18.38779, 
    17.52901, 16.66785, 15.80442, 14.93881, 14.07113, 13.20149, 12.32998, 
    11.45673, 10.58185, 9.705451, 8.827652, 7.948575, 7.068341, 6.187074, 
    5.304901, 4.421948, 3.538343, 2.654216, 1.769696, 0.8849133, 0, 
    -0.8849133, -1.769696, -2.654216, -3.538343, -4.421948, -5.304901, 
    -6.187074, -7.068341, -7.948575, -8.827652, -9.705451, -10.58185, 
    -11.45673, -12.32998, -13.20149, -14.07113, -14.93881, -15.80442, 
    -16.66785, -17.52901, -18.38779, -19.24412, -20.09789, -20.94901, 
    -21.79742, -22.64302, -23.48574, -24.32551, -25.16227, -25.99593, 
    -26.82645, -27.65377, -28.47782, -29.29857, -30.11596, -30.92996, 
    -31.74052, -32.5476, -33.35118, -34.15122, -34.94771, -35.74061, 
    -36.52991, -37.3156, -38.09766, -38.87608, -39.65086, -40.42199,
  40.69072, 39.91835, 39.14214, 38.36209, 37.57819, 36.79046, 35.9989, 
    35.20354, 34.40438, 33.60146, 32.79479, 31.98441, 31.17034, 30.35262, 
    29.5313, 28.70641, 27.87801, 27.04614, 26.21087, 25.37224, 24.53034, 
    23.68522, 22.83695, 21.98561, 21.13129, 20.27407, 19.41402, 18.55125, 
    17.68585, 16.81791, 15.94755, 15.07486, 14.19996, 13.32295, 12.44396, 
    11.5631, 10.68048, 9.79625, 8.910519, 8.023417, 7.135077, 6.245632, 
    5.355214, 4.463961, 3.57201, 2.679499, 1.786567, 0.8933536, 0, 
    -0.8933536, -1.786567, -2.679499, -3.57201, -4.463961, -5.355214, 
    -6.245632, -7.135077, -8.023417, -8.910519, -9.79625, -10.68048, 
    -11.5631, -12.44396, -13.32295, -14.19996, -15.07486, -15.94755, 
    -16.81791, -17.68585, -18.55125, -19.41402, -20.27407, -21.13129, 
    -21.98561, -22.83695, -23.68522, -24.53034, -25.37224, -26.21087, 
    -27.04614, -27.87801, -28.70641, -29.5313, -30.35262, -31.17034, 
    -31.98441, -32.79479, -33.60146, -34.40438, -35.20354, -35.9989, 
    -36.79046, -37.57819, -38.36209, -39.14214, -39.91835, -40.69072,
  40.9524, 40.1789, 39.40136, 38.61978, 37.83415, 37.04449, 36.2508, 
    35.45309, 34.6514, 33.84572, 33.03609, 32.22254, 31.4051, 30.5838, 
    29.75869, 28.92981, 28.09721, 27.26094, 26.42107, 25.57764, 24.73074, 
    23.88042, 23.02677, 22.16986, 21.30978, 20.44661, 19.58045, 18.71139, 
    17.83953, 16.96498, 16.08784, 15.20823, 14.32627, 13.44206, 12.55573, 
    11.66742, 10.77724, 9.885328, 8.99182, 8.096853, 7.200565, 6.303097, 
    5.404592, 4.505196, 3.605054, 2.704315, 1.803126, 0.9016382, 0, 
    -0.9016382, -1.803126, -2.704315, -3.605054, -4.505196, -5.404592, 
    -6.303097, -7.200565, -8.096853, -8.99182, -9.885328, -10.77724, 
    -11.66742, -12.55573, -13.44206, -14.32627, -15.20823, -16.08784, 
    -16.96498, -17.83953, -18.71139, -19.58045, -20.44661, -21.30978, 
    -22.16986, -23.02677, -23.88042, -24.73074, -25.57764, -26.42107, 
    -27.26094, -28.09721, -28.92981, -29.75869, -30.5838, -31.4051, 
    -32.22254, -33.03609, -33.84572, -34.6514, -35.45309, -36.2508, 
    -37.04449, -37.83415, -38.61978, -39.40136, -40.1789, -40.9524,
  41.20691, 40.43238, 39.6536, 38.87059, 38.08334, 37.29186, 36.49615, 
    35.69623, 34.89211, 34.08381, 33.27135, 32.45477, 31.63409, 30.80936, 
    29.9806, 29.14787, 28.31122, 27.47071, 26.62638, 25.77831, 24.92656, 
    24.0712, 23.21232, 22.35, 21.48432, 20.61537, 19.74325, 18.86807, 
    17.98992, 17.10892, 16.22518, 15.33881, 14.44994, 13.5587, 12.66521, 
    11.7696, 10.87202, 9.972599, 9.071482, 8.168813, 7.26474, 6.359414, 
    5.452987, 4.545611, 3.637443, 2.72864, 1.819359, 0.9097592, 0, 
    -0.9097592, -1.819359, -2.72864, -3.637443, -4.545611, -5.452987, 
    -6.359414, -7.26474, -8.168813, -9.071482, -9.972599, -10.87202, 
    -11.7696, -12.66521, -13.5587, -14.44994, -15.33881, -16.22518, 
    -17.10892, -17.98992, -18.86807, -19.74325, -20.61537, -21.48432, -22.35, 
    -23.21232, -24.0712, -24.92656, -25.77831, -26.62638, -27.47071, 
    -28.31122, -29.14787, -29.9806, -30.80936, -31.63409, -32.45477, 
    -33.27135, -34.08381, -34.89211, -35.69623, -36.49615, -37.29186, 
    -38.08334, -38.87059, -39.6536, -40.43238, -41.20691,
  41.45414, 40.67865, 39.89874, 39.1144, 38.32563, 37.53244, 36.73482, 
    35.9328, 35.12637, 34.31557, 33.50042, 32.68093, 31.85715, 31.02912, 
    30.19686, 29.36043, 28.51988, 27.67526, 26.82663, 25.97407, 25.11763, 
    24.2574, 23.39345, 22.52588, 21.65476, 20.7802, 19.9023, 19.02115, 
    18.13688, 17.2496, 16.35942, 15.46647, 14.57087, 13.67276, 12.77227, 
    11.86955, 10.96474, 10.05798, 9.149424, 8.239225, 7.327541, 6.414529, 
    5.50035, 4.585167, 3.669145, 2.752449, 1.835248, 0.9177083, 0, 
    -0.9177083, -1.835248, -2.752449, -3.669145, -4.585167, -5.50035, 
    -6.414529, -7.327541, -8.239225, -9.149424, -10.05798, -10.96474, 
    -11.86955, -12.77227, -13.67276, -14.57087, -15.46647, -16.35942, 
    -17.2496, -18.13688, -19.02115, -19.9023, -20.7802, -21.65476, -22.52588, 
    -23.39345, -24.2574, -25.11763, -25.97407, -26.82663, -27.67526, 
    -28.51988, -29.36043, -30.19686, -31.02912, -31.85715, -32.68093, 
    -33.50042, -34.31557, -35.12637, -35.9328, -36.73482, -37.53244, 
    -38.32563, -39.1144, -39.89874, -40.67865, -41.45414,
  41.69396, 40.9176, 40.13664, 39.35107, 38.56088, 37.76608, 36.96666, 
    36.16264, 35.35404, 34.54086, 33.72313, 32.90088, 32.07413, 31.24292, 
    30.4073, 29.56732, 28.72301, 27.87444, 27.02167, 26.16477, 25.3038, 
    24.43885, 23.57, 22.69734, 21.82095, 20.94095, 20.05743, 19.1705, 
    18.28028, 17.38689, 16.49044, 15.59108, 14.68893, 13.78413, 12.87683, 
    11.96717, 11.0553, 10.14138, 9.225567, 8.308019, 7.388902, 6.468383, 
    5.546633, 4.623823, 3.700126, 2.775718, 1.850776, 0.9254774, 0, 
    -0.9254774, -1.850776, -2.775718, -3.700126, -4.623823, -5.546633, 
    -6.468383, -7.388902, -8.308019, -9.225567, -10.14138, -11.0553, 
    -11.96717, -12.87683, -13.78413, -14.68893, -15.59108, -16.49044, 
    -17.38689, -18.28028, -19.1705, -20.05743, -20.94095, -21.82095, 
    -22.69734, -23.57, -24.43885, -25.3038, -26.16477, -27.02167, -27.87444, 
    -28.72301, -29.56732, -30.4073, -31.24292, -32.07413, -32.90088, 
    -33.72313, -34.54086, -35.35404, -36.16264, -36.96666, -37.76608, 
    -38.56088, -39.35107, -40.13664, -40.9176, -41.69396,
  41.92625, 41.14911, 40.36718, 39.58046, 38.78895, 37.99264, 37.19153, 
    36.38563, 35.57495, 34.75951, 33.93933, 33.11443, 32.28485, 31.45062, 
    30.61178, 29.76838, 28.92046, 28.06809, 27.21133, 26.35024, 25.48491, 
    24.6154, 23.74181, 22.86423, 21.98275, 21.09747, 20.20851, 19.31597, 
    18.41997, 17.52065, 16.61812, 15.71253, 14.804, 13.8927, 12.97877, 
    12.06235, 11.14361, 10.22272, 9.299832, 8.375121, 7.448759, 6.520922, 
    5.591787, 4.661538, 3.730354, 2.798423, 1.865928, 0.9330581, 0, 
    -0.9330581, -1.865928, -2.798423, -3.730354, -4.661538, -5.591787, 
    -6.520922, -7.448759, -8.375121, -9.299832, -10.22272, -11.14361, 
    -12.06235, -12.97877, -13.8927, -14.804, -15.71253, -16.61812, -17.52065, 
    -18.41997, -19.31597, -20.20851, -21.09747, -21.98275, -22.86423, 
    -23.74181, -24.6154, -25.48491, -26.35024, -27.21133, -28.06809, 
    -28.92046, -29.76838, -30.61178, -31.45062, -32.28485, -33.11443, 
    -33.93933, -34.75951, -35.57495, -36.38563, -37.19153, -37.99264, 
    -38.78895, -39.58046, -40.36718, -41.14911, -41.92625,
  42.15091, 41.37305, 40.59023, 39.80246, 39.00971, 38.21198, 37.40928, 
    36.6016, 35.78897, 34.97139, 34.14888, 33.32146, 32.48917, 31.65205, 
    30.81012, 29.96344, 29.11207, 28.25605, 27.39545, 26.53034, 25.6608, 
    24.7869, 23.90874, 23.0264, 22.13999, 21.24961, 20.35538, 19.45741, 
    18.55582, 17.65075, 16.74232, 15.83068, 14.91598, 13.99836, 13.07798, 
    12.155, 11.22959, 10.30191, 9.372141, 8.44046, 7.507047, 6.572086, 
    5.635764, 4.69827, 3.759796, 2.820537, 1.880687, 0.9404421, 0, 
    -0.9404421, -1.880687, -2.820537, -3.759796, -4.69827, -5.635764, 
    -6.572086, -7.507047, -8.44046, -9.372141, -10.30191, -11.22959, -12.155, 
    -13.07798, -13.99836, -14.91598, -15.83068, -16.74232, -17.65075, 
    -18.55582, -19.45741, -20.35538, -21.24961, -22.13999, -23.0264, 
    -23.90874, -24.7869, -25.6608, -26.53034, -27.39545, -28.25605, 
    -29.11207, -29.96344, -30.81012, -31.65205, -32.48917, -33.32146, 
    -34.14888, -34.97139, -35.78897, -36.6016, -37.40928, -38.21198, 
    -39.00971, -39.80246, -40.59023, -41.37305, -42.15091,
  42.36781, 41.5893, 40.80568, 40.01692, 39.22302, 38.42397, 37.61977, 
    36.81043, 35.99594, 35.17633, 34.35161, 33.5218, 32.68693, 31.84704, 
    31.00217, 30.15236, 29.29767, 28.43815, 27.57387, 26.70489, 25.8313, 
    24.95318, 24.07061, 23.18369, 22.29253, 21.39723, 20.49791, 19.59469, 
    18.68769, 17.77705, 16.86292, 15.94542, 15.02473, 14.10098, 13.17436, 
    12.24501, 11.31312, 10.37886, 9.442413, 8.503963, 7.563702, 6.621819, 
    5.678512, 4.733978, 3.788419, 2.842036, 1.895035, 0.947621, 0, -0.947621, 
    -1.895035, -2.842036, -3.788419, -4.733978, -5.678512, -6.621819, 
    -7.563702, -8.503963, -9.442413, -10.37886, -11.31312, -12.24501, 
    -13.17436, -14.10098, -15.02473, -15.94542, -16.86292, -17.77705, 
    -18.68769, -19.59469, -20.49791, -21.39723, -22.29253, -23.18369, 
    -24.07061, -24.95318, -25.8313, -26.70489, -27.57387, -28.43815, 
    -29.29767, -30.15236, -31.00217, -31.84704, -32.68693, -33.5218, 
    -34.35161, -35.17633, -35.99594, -36.81043, -37.61977, -38.42397, 
    -39.22302, -40.01692, -40.80568, -41.5893, -42.36781,
  42.57683, 41.79774, 41.01338, 40.22372, 39.42876, 38.62848, 37.82288, 
    37.01196, 36.19573, 35.3742, 34.54738, 33.7153, 32.87798, 32.03546, 
    31.18778, 30.33498, 29.47712, 28.61425, 27.74643, 26.87375, 25.99627, 
    25.11408, 24.22728, 23.33596, 22.44022, 21.54018, 20.63595, 19.72766, 
    18.81544, 17.89944, 16.97978, 16.05663, 15.13014, 14.20047, 13.2678, 
    12.33229, 11.39412, 10.45349, 9.510569, 8.565559, 7.618658, 6.670065, 
    5.719984, 4.768622, 3.816189, 2.862896, 1.908957, 0.9545865, 0, 
    -0.9545865, -1.908957, -2.862896, -3.816189, -4.768622, -5.719984, 
    -6.670065, -7.618658, -8.565559, -9.510569, -10.45349, -11.39412, 
    -12.33229, -13.2678, -14.20047, -15.13014, -16.05663, -16.97978, 
    -17.89944, -18.81544, -19.72766, -20.63595, -21.54018, -22.44022, 
    -23.33596, -24.22728, -25.11408, -25.99627, -26.87375, -27.74643, 
    -28.61425, -29.47712, -30.33498, -31.18778, -32.03546, -32.87798, 
    -33.7153, -34.54738, -35.3742, -36.19573, -37.01196, -37.82288, 
    -38.62848, -39.42876, -40.22372, -41.01338, -41.79774, -42.57683,
  42.77788, 41.99827, 41.21324, 40.42275, 39.6268, 38.82537, 38.01846, 
    37.20607, 36.38819, 35.56485, 34.73605, 33.90181, 33.06216, 32.21714, 
    31.36679, 30.51114, 29.65025, 28.78417, 27.91298, 27.03675, 26.15555, 
    25.26947, 24.3786, 23.48304, 22.5829, 21.6783, 20.76936, 19.85619, 
    18.93895, 18.01776, 17.09279, 16.16418, 15.2321, 14.29671, 13.3582, 
    12.41673, 11.47251, 10.52571, 9.576528, 8.625175, 7.671851, 6.716765, 
    5.760129, 4.802159, 3.843073, 2.883091, 1.922435, 0.9613302, 0, 
    -0.9613302, -1.922435, -2.883091, -3.843073, -4.802159, -5.760129, 
    -6.716765, -7.671851, -8.625175, -9.576528, -10.52571, -11.47251, 
    -12.41673, -13.3582, -14.29671, -15.2321, -16.16418, -17.09279, 
    -18.01776, -18.93895, -19.85619, -20.76936, -21.6783, -22.5829, 
    -23.48304, -24.3786, -25.26947, -26.15555, -27.03675, -27.91298, 
    -28.78417, -29.65025, -30.51114, -31.36679, -32.21714, -33.06216, 
    -33.90181, -34.73605, -35.56485, -36.38819, -37.20607, -38.01846, 
    -38.82537, -39.6268, -40.42275, -41.21324, -41.99827, -42.77788,
  42.97084, 42.19077, 41.40512, 40.61388, 39.81702, 39.01452, 38.20639, 
    37.39261, 36.57319, 35.74813, 34.91746, 34.08119, 33.23934, 32.39194, 
    31.53904, 30.68068, 29.8169, 28.94778, 28.07337, 27.19374, 26.30898, 
    25.41917, 24.52441, 23.6248, 22.72045, 21.81147, 20.89799, 19.98014, 
    19.05806, 18.1319, 17.20181, 16.26795, 15.33048, 14.38959, 13.44545, 
    12.49824, 11.54817, 10.59543, 9.640213, 8.682739, 7.723217, 6.761864, 
    5.7989, 4.834549, 3.869038, 2.902596, 1.935454, 0.9678438, 0, -0.9678438, 
    -1.935454, -2.902596, -3.869038, -4.834549, -5.7989, -6.761864, 
    -7.723217, -8.682739, -9.640213, -10.59543, -11.54817, -12.49824, 
    -13.44545, -14.38959, -15.33048, -16.26795, -17.20181, -18.1319, 
    -19.05806, -19.98014, -20.89799, -21.81147, -22.72045, -23.6248, 
    -24.52441, -25.41917, -26.30898, -27.19374, -28.07337, -28.94778, 
    -29.8169, -30.68068, -31.53904, -32.39194, -33.23934, -34.08119, 
    -34.91746, -35.74813, -36.57319, -37.39261, -38.20639, -39.01452, 
    -39.81702, -40.61388, -41.40512, -42.19077, -42.97084,
  43.1556, 42.37512, 41.58892, 40.79699, 39.99928, 39.1958, 38.38652, 
    37.57145, 36.75058, 35.92393, 35.09149, 34.25329, 33.40936, 32.55971, 
    31.7044, 30.84346, 29.97694, 29.10491, 28.22743, 27.34457, 26.45642, 
    25.56305, 24.66457, 23.76108, 22.85269, 21.93953, 21.02171, 20.09937, 
    19.17266, 18.24172, 17.30672, 16.36782, 15.42518, 14.479, 13.52945, 
    12.57673, 11.62103, 10.66257, 9.701547, 8.738181, 7.772693, 6.805305, 
    5.836247, 4.865752, 3.894052, 2.921387, 1.947996, 0.9741191, 0, 
    -0.9741191, -1.947996, -2.921387, -3.894052, -4.865752, -5.836247, 
    -6.805305, -7.772693, -8.738181, -9.701547, -10.66257, -11.62103, 
    -12.57673, -13.52945, -14.479, -15.42518, -16.36782, -17.30672, 
    -18.24172, -19.17266, -20.09937, -21.02171, -21.93953, -22.85269, 
    -23.76108, -24.66457, -25.56305, -26.45642, -27.34457, -28.22743, 
    -29.10491, -29.97694, -30.84346, -31.7044, -32.55971, -33.40936, 
    -34.25329, -35.09149, -35.92393, -36.75058, -37.57145, -38.38652, 
    -39.1958, -39.99928, -40.79699, -41.58892, -42.37512, -43.1556,
  43.33206, 42.55122, 41.76453, 40.97196, 40.17348, 39.36908, 38.55875, 
    37.74247, 36.92025, 36.09208, 35.25799, 34.41798, 33.57207, 32.7203, 
    31.86271, 30.99933, 30.13022, 29.25543, 28.37503, 27.4891, 26.59771, 
    25.70096, 24.79893, 23.89175, 22.97951, 22.06234, 21.14038, 20.21375, 
    19.28261, 18.34711, 17.4074, 16.46367, 15.51608, 14.56483, 13.61009, 
    12.65208, 11.691, 10.72705, 9.760451, 8.791431, 7.820215, 6.847034, 
    5.872125, 4.895727, 3.918083, 2.93944, 1.960045, 0.9801481, 0, 
    -0.9801481, -1.960045, -2.93944, -3.918083, -4.895727, -5.872125, 
    -6.847034, -7.820215, -8.791431, -9.760451, -10.72705, -11.691, 
    -12.65208, -13.61009, -14.56483, -15.51608, -16.46367, -17.4074, 
    -18.34711, -19.28261, -20.21375, -21.14038, -22.06234, -22.97951, 
    -23.89175, -24.79893, -25.70096, -26.59771, -27.4891, -28.37503, 
    -29.25543, -30.13022, -30.99933, -31.86271, -32.7203, -33.57207, 
    -34.41798, -35.25799, -36.09208, -36.92025, -37.74247, -38.55875, 
    -39.36908, -40.17348, -40.97196, -41.76453, -42.55122, -43.33206,
  43.50012, 42.71897, 41.93184, 41.13869, 40.3395, 39.53426, 38.72294, 
    37.90554, 37.08205, 36.25248, 35.41682, 34.57511, 33.72735, 32.87358, 
    32.01384, 31.14815, 30.27658, 29.39919, 28.51603, 27.62718, 26.73272, 
    25.83275, 24.92736, 24.01665, 23.10075, 22.17978, 21.25386, 20.32315, 
    19.38778, 18.44792, 17.50373, 16.55539, 15.60307, 14.64697, 13.68729, 
    12.72422, 11.75798, 10.78878, 9.816853, 8.842422, 7.865723, 6.886996, 
    5.906484, 4.924435, 3.941099, 2.956731, 1.971586, 0.9859229, 0, 
    -0.9859229, -1.971586, -2.956731, -3.941099, -4.924435, -5.906484, 
    -6.886996, -7.865723, -8.842422, -9.816853, -10.78878, -11.75798, 
    -12.72422, -13.68729, -14.64697, -15.60307, -16.55539, -17.50373, 
    -18.44792, -19.38778, -20.32315, -21.25386, -22.17978, -23.10075, 
    -24.01665, -24.92736, -25.83275, -26.73272, -27.62718, -28.51603, 
    -29.39919, -30.27658, -31.14815, -32.01384, -32.87358, -33.72735, 
    -34.57511, -35.41682, -36.25248, -37.08205, -37.90554, -38.72294, 
    -39.53426, -40.3395, -41.13869, -41.93184, -42.71897, -43.50012,
  43.65969, 42.87827, 42.09073, 41.29707, 40.49723, 39.69121, 38.87898, 
    38.06054, 37.23587, 36.40498, 35.56787, 34.72456, 33.87507, 33.01942, 
    32.15764, 31.28979, 30.4159, 29.53604, 28.65027, 27.75867, 26.86131, 
    25.95829, 25.0497, 24.13567, 23.21629, 22.2917, 21.36204, 20.42744, 
    19.48806, 18.54405, 17.5956, 16.64287, 15.68605, 14.72534, 13.76093, 
    12.79304, 11.82189, 10.84769, 9.870676, 8.891085, 7.909157, 6.925138, 
    5.939281, 4.951838, 3.963069, 2.973237, 1.982603, 0.9914355, 0, 
    -0.9914355, -1.982603, -2.973237, -3.963069, -4.951838, -5.939281, 
    -6.925138, -7.909157, -8.891085, -9.870676, -10.84769, -11.82189, 
    -12.79304, -13.76093, -14.72534, -15.68605, -16.64287, -17.5956, 
    -18.54405, -19.48806, -20.42744, -21.36204, -22.2917, -23.21629, 
    -24.13567, -25.0497, -25.95829, -26.86131, -27.75867, -28.65027, 
    -29.53604, -30.4159, -31.28979, -32.15764, -33.01942, -33.87507, 
    -34.72456, -35.56787, -36.40498, -37.23587, -38.06054, -38.87898, 
    -39.69121, -40.49723, -41.29707, -42.09073, -42.87827, -43.65969,
  43.81068, 43.02901, 42.24112, 41.44698, 40.64656, 39.83982, 39.02676, 
    38.20735, 37.38158, 36.54947, 35.71101, 34.8662, 34.01508, 33.15767, 
    32.29399, 31.4241, 30.54803, 29.66586, 28.77763, 27.88343, 26.98333, 
    26.07744, 25.16584, 24.24865, 23.32599, 22.39799, 21.46477, 20.5265, 
    19.58331, 18.63538, 17.68288, 16.72599, 15.7649, 14.79981, 13.83093, 
    12.85847, 11.88264, 10.90369, 9.92185, 8.937356, 7.950458, 6.96141, 
    5.970469, 4.977899, 3.983964, 2.988935, 1.993082, 0.9966785, 0, 
    -0.9966785, -1.993082, -2.988935, -3.983964, -4.977899, -5.970469, 
    -6.96141, -7.950458, -8.937356, -9.92185, -10.90369, -11.88264, 
    -12.85847, -13.83093, -14.79981, -15.7649, -16.72599, -17.68288, 
    -18.63538, -19.58331, -20.5265, -21.46477, -22.39799, -23.32599, 
    -24.24865, -25.16584, -26.07744, -26.98333, -27.88343, -28.77763, 
    -29.66586, -30.54803, -31.4241, -32.29399, -33.15767, -34.01508, 
    -34.8662, -35.71101, -36.54947, -37.38158, -38.20735, -39.02676, 
    -39.83982, -40.64656, -41.44698, -42.24112, -43.02901, -43.81068,
  43.95298, 43.17111, 42.38291, 41.58834, 40.78738, 39.97999, 39.16616, 
    38.34586, 37.51908, 36.68583, 35.8461, 34.99992, 34.14728, 33.28822, 
    32.42276, 31.55096, 30.67286, 29.78851, 28.89797, 28.00133, 27.09867, 
    26.19007, 25.27564, 24.35549, 23.42973, 22.49851, 21.56195, 20.6202, 
    19.67343, 18.7218, 17.76548, 16.80466, 15.83954, 14.87031, 13.89719, 
    12.9204, 11.94017, 10.95672, 9.970306, 8.981172, 7.989569, 6.995759, 
    6.000007, 5.002581, 4.003754, 3.003803, 2.003006, 1.001644, 0, -1.001644, 
    -2.003006, -3.003803, -4.003754, -5.002581, -6.000007, -6.995759, 
    -7.989569, -8.981172, -9.970306, -10.95672, -11.94017, -12.9204, 
    -13.89719, -14.87031, -15.83954, -16.80466, -17.76548, -18.7218, 
    -19.67343, -20.6202, -21.56195, -22.49851, -23.42973, -24.35549, 
    -25.27564, -26.19007, -27.09867, -28.00133, -28.89797, -29.78851, 
    -30.67286, -31.55096, -32.42276, -33.28822, -34.14728, -34.99992, 
    -35.8461, -36.68583, -37.51908, -38.34586, -39.16616, -39.97999, 
    -40.78738, -41.58834, -42.38291, -43.17111, -43.95298,
  44.08652, 43.30448, 42.516, 41.72106, 40.91961, 40.11162, 39.29708, 
    38.47596, 37.64825, 36.81395, 35.97306, 35.12558, 34.27153, 33.41094, 
    32.54383, 31.67025, 30.79025, 29.90387, 29.01118, 28.11226, 27.20719, 
    26.29606, 25.37897, 24.45604, 23.52739, 22.59314, 21.65344, 20.70844, 
    19.7583, 18.80319, 17.84328, 16.87877, 15.90985, 14.93673, 13.95963, 
    12.97877, 11.99438, 11.0067, 10.01598, 9.02247, 8.026436, 7.02814, 
    6.027852, 5.025849, 4.022411, 3.017821, 2.012363, 1.006326, 0, -1.006326, 
    -2.012363, -3.017821, -4.022411, -5.025849, -6.027852, -7.02814, 
    -8.026436, -9.02247, -10.01598, -11.0067, -11.99438, -12.97877, 
    -13.95963, -14.93673, -15.90985, -16.87877, -17.84328, -18.80319, 
    -19.7583, -20.70844, -21.65344, -22.59314, -23.52739, -24.45604, 
    -25.37897, -26.29606, -27.20719, -28.11226, -29.01118, -29.90387, 
    -30.79025, -31.67025, -32.54383, -33.41094, -34.27153, -35.12558, 
    -35.97306, -36.81395, -37.64825, -38.47596, -39.29708, -40.11162, 
    -40.91961, -41.72106, -42.516, -43.30448, -44.08652,
  44.21122, 43.42903, 42.64032, 41.84503, 41.04314, 40.23461, 39.41943, 
    38.59755, 37.76899, 36.93372, 36.09175, 35.24308, 34.38773, 33.52573, 
    32.65709, 31.78186, 30.90008, 30.01182, 29.11712, 28.21608, 27.30877, 
    26.39529, 25.47573, 24.55021, 23.61885, 22.68178, 21.73915, 20.79111, 
    19.83782, 18.87945, 17.91618, 16.94822, 15.97575, 14.99899, 14.01815, 
    13.03348, 12.0452, 11.05355, 10.0588, 9.061195, 8.061007, 7.058504, 
    6.053965, 5.047671, 4.039908, 3.030967, 2.021138, 1.010717, 0, -1.010717, 
    -2.021138, -3.030967, -4.039908, -5.047671, -6.053965, -7.058504, 
    -8.061007, -9.061195, -10.0588, -11.05355, -12.0452, -13.03348, 
    -14.01815, -14.99899, -15.97575, -16.94822, -17.91618, -18.87945, 
    -19.83782, -20.79111, -21.73915, -22.68178, -23.61885, -24.55021, 
    -25.47573, -26.39529, -27.30877, -28.21608, -29.11712, -30.01182, 
    -30.90008, -31.78186, -32.65709, -33.52573, -34.38773, -35.24308, 
    -36.09175, -36.93372, -37.76899, -38.59755, -39.41943, -40.23461, 
    -41.04314, -41.84503, -42.64032, -43.42903, -44.21122,
  44.32701, 43.54469, 42.75576, 41.96017, 41.15789, 40.34887, 39.5331, 
    38.71054, 37.8812, 37.04504, 36.20208, 35.35233, 34.49578, 33.63246, 
    32.76241, 31.88566, 31.00225, 30.11224, 29.2157, 28.3127, 27.40331, 
    26.48764, 25.56579, 24.63787, 23.704, 22.76431, 21.81896, 20.8681, 
    19.91188, 18.95048, 17.9841, 17.01292, 16.03714, 15.05699, 14.07269, 
    13.08447, 12.09256, 11.09722, 10.09871, 9.097291, 8.09323, 7.086808, 
    6.078306, 5.068013, 4.05622, 3.043222, 2.029319, 1.014811, 0, -1.014811, 
    -2.029319, -3.043222, -4.05622, -5.068013, -6.078306, -7.086808, 
    -8.09323, -9.097291, -10.09871, -11.09722, -12.09256, -13.08447, 
    -14.07269, -15.05699, -16.03714, -17.01292, -17.9841, -18.95048, 
    -19.91188, -20.8681, -21.81896, -22.76431, -23.704, -24.63787, -25.56579, 
    -26.48764, -27.40331, -28.3127, -29.2157, -30.11224, -31.00225, 
    -31.88566, -32.76241, -33.63246, -34.49578, -35.35233, -36.20208, 
    -37.04504, -37.8812, -38.71054, -39.5331, -40.34887, -41.15789, 
    -41.96017, -42.75576, -43.54469, -44.32701,
  44.4338, 43.65138, 42.86227, 42.06641, 41.26377, 40.45432, 39.63801, 
    38.81484, 37.98478, 37.14782, 36.30396, 35.45321, 34.59556, 33.73105, 
    32.85971, 31.98156, 31.09665, 30.20505, 29.3068, 28.40199, 27.4907, 
    26.57302, 25.64905, 24.71892, 23.78273, 22.84064, 21.89278, 20.9393, 
    19.98038, 19.0162, 18.04693, 17.07278, 16.09396, 15.11067, 14.12316, 
    13.13165, 12.1364, 11.13764, 10.13566, 9.130703, 8.123061, 7.113011, 
    6.100842, 5.086846, 4.071321, 3.054569, 2.036894, 1.018601, 0, -1.018601, 
    -2.036894, -3.054569, -4.071321, -5.086846, -6.100842, -7.113011, 
    -8.123061, -9.130703, -10.13566, -11.13764, -12.1364, -13.13165, 
    -14.12316, -15.11067, -16.09396, -17.07278, -18.04693, -19.0162, 
    -19.98038, -20.9393, -21.89278, -22.84064, -23.78273, -24.71892, 
    -25.64905, -26.57302, -27.4907, -28.40199, -29.3068, -30.20505, 
    -31.09665, -31.98156, -32.85971, -33.73105, -34.59556, -35.45321, 
    -36.30396, -37.14782, -37.98478, -38.81484, -39.63801, -40.45432, 
    -41.26377, -42.06641, -42.86227, -43.65138, -44.4338,
  44.53154, 43.74903, 42.95976, 42.16367, 41.36071, 40.55087, 39.73409, 
    38.91036, 38.07965, 37.24197, 36.39729, 35.54563, 34.68699, 33.8214, 
    32.94887, 32.06945, 31.18319, 30.29012, 29.39032, 28.48387, 27.57083, 
    26.65132, 25.72542, 24.79326, 23.85496, 22.91066, 21.9605, 21.00464, 
    20.04325, 19.0765, 18.1046, 17.12773, 16.1461, 15.15995, 14.16949, 
    13.17497, 12.17664, 11.17476, 10.16958, 9.161384, 8.150454, 7.137073, 
    6.121536, 5.104141, 4.08519, 3.06499, 2.04385, 1.022082, 0, -1.022082, 
    -2.04385, -3.06499, -4.08519, -5.104141, -6.121536, -7.137073, -8.150454, 
    -9.161384, -10.16958, -11.17476, -12.17664, -13.17497, -14.16949, 
    -15.15995, -16.1461, -17.12773, -18.1046, -19.0765, -20.04325, -21.00464, 
    -21.9605, -22.91066, -23.85496, -24.79326, -25.72542, -26.65132, 
    -27.57083, -28.48387, -29.39032, -30.29012, -31.18319, -32.06945, 
    -32.94887, -33.8214, -34.68699, -35.54563, -36.39729, -37.24197, 
    -38.07965, -38.91036, -39.73409, -40.55087, -41.36071, -42.16367, 
    -42.95976, -43.74903, -44.53154,
  44.62016, 43.83758, 43.04817, 42.25187, 41.44865, 40.63845, 39.82125, 
    38.99702, 38.16574, 37.3274, 36.48199, 35.62952, 34.76999, 33.90341, 
    33.02983, 32.14926, 31.26176, 30.36738, 29.46618, 28.55823, 27.64362, 
    26.72244, 25.7948, 24.86081, 23.92059, 22.97429, 22.02205, 21.06402, 
    20.10039, 19.13132, 18.15702, 17.17768, 16.19351, 15.20475, 14.21162, 
    13.21437, 12.21324, 11.2085, 10.20043, 9.189286, 8.175366, 7.158958, 
    6.140359, 5.119872, 4.097805, 3.074468, 2.050177, 1.025248, 0, -1.025248, 
    -2.050177, -3.074468, -4.097805, -5.119872, -6.140359, -7.158958, 
    -8.175366, -9.189286, -10.20043, -11.2085, -12.21324, -13.21437, 
    -14.21162, -15.20475, -16.19351, -17.17768, -18.15702, -19.13132, 
    -20.10039, -21.06402, -22.02205, -22.97429, -23.92059, -24.86081, 
    -25.7948, -26.72244, -27.64362, -28.55823, -29.46618, -30.36738, 
    -31.26176, -32.14926, -33.02983, -33.90341, -34.76999, -35.62952, 
    -36.48199, -37.3274, -38.16574, -38.99702, -39.82125, -40.63845, 
    -41.44865, -42.25187, -43.04817, -43.83758, -44.62016,
  44.6996, 43.91697, 43.12745, 42.33097, 41.5275, 40.717, 39.89942, 39.07475, 
    38.24297, 37.40405, 36.55799, 35.70479, 34.84446, 33.97701, 33.10248, 
    32.22089, 31.33229, 30.43673, 29.53428, 28.625, 27.70898, 26.78632, 
    25.85711, 24.92148, 23.97954, 23.03145, 22.07734, 21.11737, 20.15172, 
    19.18058, 18.20412, 17.22256, 16.23612, 15.24501, 14.24948, 13.24977, 
    12.24614, 11.23884, 10.22816, 9.21437, 8.197762, 7.178632, 6.157281, 
    5.134015, 4.109146, 3.08299, 2.055866, 1.028095, 0, -1.028095, -2.055866, 
    -3.08299, -4.109146, -5.134015, -6.157281, -7.178632, -8.197762, 
    -9.21437, -10.22816, -11.23884, -12.24614, -13.24977, -14.24948, 
    -15.24501, -16.23612, -17.22256, -18.20412, -19.18058, -20.15172, 
    -21.11737, -22.07734, -23.03145, -23.97954, -24.92148, -25.85711, 
    -26.78632, -27.70898, -28.625, -29.53428, -30.43673, -31.33229, 
    -32.22089, -33.10248, -33.97701, -34.84446, -35.70479, -36.55799, 
    -37.40405, -38.24297, -39.07475, -39.89942, -40.717, -41.5275, -42.33097, 
    -43.12745, -43.91697, -44.6996,
  44.76982, 43.98714, 43.19752, 42.40089, 41.59722, 40.78645, 39.96855, 
    39.1435, 38.31126, 37.47184, 36.62521, 35.77137, 34.91034, 34.04213, 
    33.16676, 32.28428, 31.39471, 30.49811, 29.59455, 28.6841, 27.76684, 
    26.84286, 25.91227, 24.97519, 24.03174, 23.08206, 22.1263, 21.16462, 
    20.19719, 19.2242, 18.24584, 17.26232, 16.27386, 15.28068, 14.28303, 
    13.28114, 12.27528, 11.26572, 10.25273, 9.236594, 8.217607, 7.196066, 
    6.172276, 5.146547, 4.119196, 3.090542, 2.060907, 1.030618, 0, -1.030618, 
    -2.060907, -3.090542, -4.119196, -5.146547, -6.172276, -7.196066, 
    -8.217607, -9.236594, -10.25273, -11.26572, -12.27528, -13.28114, 
    -14.28303, -15.28068, -16.27386, -17.26232, -18.24584, -19.2242, 
    -20.19719, -21.16462, -22.1263, -23.08206, -24.03174, -24.97519, 
    -25.91227, -26.84286, -27.76684, -28.6841, -29.59455, -30.49811, 
    -31.39471, -32.28428, -33.16676, -34.04213, -34.91034, -35.77137, 
    -36.62521, -37.47184, -38.31126, -39.1435, -39.96855, -40.78645, 
    -41.59722, -42.40089, -43.19752, -43.98714, -44.76982,
  44.83077, 44.04806, 43.25835, 42.4616, 41.65775, 40.84675, 40.02857, 
    39.20319, 38.37057, 37.53071, 36.68359, 35.8292, 34.96757, 34.0987, 
    33.22261, 32.33934, 31.44894, 30.55145, 29.64693, 28.73546, 27.81712, 
    26.892, 25.96022, 25.02188, 24.07711, 23.12605, 22.16886, 21.20569, 
    20.23672, 19.26213, 18.28212, 17.2969, 16.30668, 15.3117, 14.3122, 
    13.30842, 12.30063, 11.2891, 10.2741, 9.255927, 8.23487, 7.211231, 
    6.18532, 5.15745, 4.127939, 3.097111, 2.065293, 1.032812, 0, -1.032812, 
    -2.065293, -3.097111, -4.127939, -5.15745, -6.18532, -7.211231, -8.23487, 
    -9.255927, -10.2741, -11.2891, -12.30063, -13.30842, -14.3122, -15.3117, 
    -16.30668, -17.2969, -18.28212, -19.26213, -20.23672, -21.20569, 
    -22.16886, -23.12605, -24.07711, -25.02188, -25.96022, -26.892, 
    -27.81712, -28.73546, -29.64693, -30.55145, -31.44894, -32.33934, 
    -33.22261, -34.0987, -34.96757, -35.8292, -36.68359, -37.53071, 
    -38.37057, -39.20319, -40.02857, -40.84675, -41.65775, -42.4616, 
    -43.25835, -44.04806, -44.83077,
  44.88241, 44.09967, 43.3099, 42.51304, 41.70904, 40.89785, 40.07944, 
    39.25378, 38.42085, 37.58062, 36.73308, 35.87823, 35.01609, 34.14666, 
    33.26997, 32.38604, 31.49493, 30.59668, 29.69135, 28.77902, 27.85977, 
    26.93369, 26.00089, 25.06149, 24.1156, 23.16338, 22.20498, 21.24054, 
    20.27026, 19.29432, 18.31291, 17.32624, 16.33454, 15.33803, 14.33696, 
    13.33158, 12.32215, 11.30894, 10.29224, 9.272337, 8.249522, 7.224104, 
    6.196393, 5.166705, 4.135361, 3.102689, 2.069016, 1.034675, 0, -1.034675, 
    -2.069016, -3.102689, -4.135361, -5.166705, -6.196393, -7.224104, 
    -8.249522, -9.272337, -10.29224, -11.30894, -12.32215, -13.33158, 
    -14.33696, -15.33803, -16.33454, -17.32624, -18.31291, -19.29432, 
    -20.27026, -21.24054, -22.20498, -23.16338, -24.1156, -25.06149, 
    -26.00089, -26.93369, -27.85977, -28.77902, -29.69135, -30.59668, 
    -31.49493, -32.38604, -33.26997, -34.14666, -35.01609, -35.87823, 
    -36.73308, -37.58062, -38.42085, -39.25378, -40.07944, -40.89785, 
    -41.70904, -42.51304, -43.3099, -44.09967, -44.88241,
  44.9247, 44.14195, 43.35213, 42.55518, 41.75106, 40.93972, 40.12112, 
    39.29524, 38.46204, 37.62151, 36.77364, 35.91842, 35.05586, 34.18597, 
    33.30878, 32.42432, 31.53263, 30.63375, 29.72776, 28.81473, 27.89473, 
    26.96786, 26.03424, 25.09396, 24.14717, 23.19399, 22.23459, 21.26912, 
    20.29777, 19.32071, 18.33815, 17.3503, 16.35738, 15.35962, 14.35726, 
    13.35057, 12.3398, 11.32522, 10.30712, 9.285798, 8.261543, 7.234665, 
    6.205477, 5.174297, 4.14145, 3.107264, 2.07207, 1.036204, 0, -1.036204, 
    -2.07207, -3.107264, -4.14145, -5.174297, -6.205477, -7.234665, 
    -8.261543, -9.285798, -10.30712, -11.32522, -12.3398, -13.35057, 
    -14.35726, -15.35962, -16.35738, -17.3503, -18.33815, -19.32071, 
    -20.29777, -21.26912, -22.23459, -23.19399, -24.14717, -25.09396, 
    -26.03424, -26.96786, -27.89473, -28.81473, -29.72776, -30.63375, 
    -31.53263, -32.42432, -33.30878, -34.18597, -35.05586, -35.91842, 
    -36.77364, -37.62151, -38.46204, -39.29524, -40.12112, -40.93972, 
    -41.75106, -42.55518, -43.35213, -44.14195, -44.9247,
  44.95763, 44.17486, 43.385, 42.58799, 41.78378, 40.97232, 40.15358, 
    39.32752, 38.49412, 37.65335, 36.80522, 35.94971, 35.08683, 34.21658, 
    33.33901, 32.45413, 31.56199, 30.66263, 29.75613, 28.84255, 27.92197, 
    26.99449, 26.06021, 25.11926, 24.17175, 23.21784, 22.25766, 21.29139, 
    20.3192, 19.34128, 18.35783, 17.36906, 16.37519, 15.37645, 14.37309, 
    13.36537, 12.35355, 11.33791, 10.31872, 9.29629, 8.270913, 7.242897, 
    6.212557, 5.180215, 4.146196, 3.11083, 2.074451, 1.037395, 0, -1.037395, 
    -2.074451, -3.11083, -4.146196, -5.180215, -6.212557, -7.242897, 
    -8.270913, -9.29629, -10.31872, -11.33791, -12.35355, -13.36537, 
    -14.37309, -15.37645, -16.37519, -17.36906, -18.35783, -19.34128, 
    -20.3192, -21.29139, -22.25766, -23.21784, -24.17175, -25.11926, 
    -26.06021, -26.99449, -27.92197, -28.84255, -29.75613, -30.66263, 
    -31.56199, -32.45413, -33.33901, -34.21658, -35.08683, -35.94971, 
    -36.80522, -37.65335, -38.49412, -39.32752, -40.15358, -40.97232, 
    -41.78378, -42.58799, -43.385, -44.17486, -44.95763,
  44.98116, 44.19839, 43.4085, 42.61144, 41.80717, 40.99562, 40.17678, 
    39.3506, 38.51705, 37.67612, 36.8278, 35.97208, 35.10897, 34.23848, 
    33.36062, 32.47544, 31.58298, 30.68328, 29.77641, 28.86244, 27.94145, 
    27.01353, 26.0788, 25.13736, 24.18934, 23.2349, 22.27417, 21.30732, 
    20.33454, 19.356, 18.3719, 17.38247, 16.38792, 15.38849, 14.38441, 
    13.37596, 12.36339, 11.34698, 10.32702, 9.303797, 8.277617, 7.248786, 
    6.217623, 5.184449, 4.149592, 3.113382, 2.076154, 1.038247, 0, -1.038247, 
    -2.076154, -3.113382, -4.149592, -5.184449, -6.217623, -7.248786, 
    -8.277617, -9.303797, -10.32702, -11.34698, -12.36339, -13.37596, 
    -14.38441, -15.38849, -16.38792, -17.38247, -18.3719, -19.356, -20.33454, 
    -21.30732, -22.27417, -23.2349, -24.18934, -25.13736, -26.0788, 
    -27.01353, -27.94145, -28.86244, -29.77641, -30.68328, -31.58298, 
    -32.47544, -33.36062, -34.23848, -35.10897, -35.97208, -36.8278, 
    -37.67612, -38.51705, -39.3506, -40.17678, -40.99562, -41.80717, 
    -42.61144, -43.4085, -44.19839, -44.98116,
  44.99529, 44.21251, 43.4226, 42.62552, 41.82121, 41.00961, 40.1907, 
    39.36445, 38.53082, 37.68979, 36.84136, 35.98551, 35.12226, 34.25162, 
    33.3736, 32.48825, 31.59559, 30.69568, 29.78859, 28.87439, 27.95315, 
    27.02497, 26.08995, 25.14822, 24.19991, 23.24514, 22.28408, 21.31689, 
    20.34374, 19.36483, 18.38036, 17.39053, 16.39557, 15.39572, 14.39121, 
    13.38232, 12.3693, 11.35243, 10.332, 9.308306, 8.281642, 7.252323, 
    6.220666, 5.186993, 4.151631, 3.114914, 2.077178, 1.038759, 0, -1.038759, 
    -2.077178, -3.114914, -4.151631, -5.186993, -6.220666, -7.252323, 
    -8.281642, -9.308306, -10.332, -11.35243, -12.3693, -13.38232, -14.39121, 
    -15.39572, -16.39557, -17.39053, -18.38036, -19.36483, -20.34374, 
    -21.31689, -22.28408, -23.24514, -24.19991, -25.14822, -26.08995, 
    -27.02497, -27.95315, -28.87439, -29.78859, -30.69568, -31.59559, 
    -32.48825, -33.3736, -34.25162, -35.12226, -35.98551, -36.84136, 
    -37.68979, -38.53082, -39.36445, -40.1907, -41.00961, -41.82121, 
    -42.62552, -43.4226, -44.21251, -44.99529,
  45, 44.21722, 43.42731, 42.63021, 41.82589, 41.01428, 40.19535, 39.36907, 
    38.53541, 37.69435, 36.84588, 35.98999, 35.12669, 34.256, 33.37793, 
    32.49251, 31.59979, 30.69982, 29.79265, 28.87837, 27.95705, 27.02878, 
    26.09367, 25.15185, 24.20343, 23.24856, 22.28739, 21.32008, 20.34682, 
    19.36778, 18.38318, 17.39322, 16.39812, 15.39813, 14.39348, 13.38444, 
    12.37127, 11.35425, 10.33367, 9.30981, 8.282985, 7.253503, 6.221681, 
    5.187841, 4.152311, 3.115426, 2.077519, 1.03893, 0, -1.03893, -2.077519, 
    -3.115426, -4.152311, -5.187841, -6.221681, -7.253503, -8.282985, 
    -9.30981, -10.33367, -11.35425, -12.37127, -13.38444, -14.39348, 
    -15.39813, -16.39812, -17.39322, -18.38318, -19.36778, -20.34682, 
    -21.32008, -22.28739, -23.24856, -24.20343, -25.15185, -26.09367, 
    -27.02878, -27.95705, -28.87837, -29.79265, -30.69982, -31.59979, 
    -32.49251, -33.37793, -34.256, -35.12669, -35.98999, -36.84588, 
    -37.69435, -38.53541, -39.36907, -40.19535, -41.01428, -41.82589, 
    -42.63021, -43.42731, -44.21722, -45,
  44.99529, 44.21251, 43.4226, 42.62552, 41.82121, 41.00961, 40.1907, 
    39.36445, 38.53082, 37.68979, 36.84136, 35.98551, 35.12226, 34.25162, 
    33.3736, 32.48825, 31.59559, 30.69568, 29.78859, 28.87439, 27.95315, 
    27.02497, 26.08995, 25.14822, 24.19991, 23.24514, 22.28408, 21.31689, 
    20.34374, 19.36483, 18.38036, 17.39053, 16.39557, 15.39572, 14.39121, 
    13.38232, 12.3693, 11.35243, 10.332, 9.308306, 8.281642, 7.252323, 
    6.220666, 5.186993, 4.151631, 3.114914, 2.077178, 1.038759, 0, -1.038759, 
    -2.077178, -3.114914, -4.151631, -5.186993, -6.220666, -7.252323, 
    -8.281642, -9.308306, -10.332, -11.35243, -12.3693, -13.38232, -14.39121, 
    -15.39572, -16.39557, -17.39053, -18.38036, -19.36483, -20.34374, 
    -21.31689, -22.28408, -23.24514, -24.19991, -25.14822, -26.08995, 
    -27.02497, -27.95315, -28.87439, -29.78859, -30.69568, -31.59559, 
    -32.48825, -33.3736, -34.25162, -35.12226, -35.98551, -36.84136, 
    -37.68979, -38.53082, -39.36445, -40.1907, -41.00961, -41.82121, 
    -42.62552, -43.4226, -44.21251, -44.99529,
  44.98116, 44.19839, 43.4085, 42.61144, 41.80717, 40.99562, 40.17678, 
    39.3506, 38.51705, 37.67612, 36.8278, 35.97208, 35.10897, 34.23848, 
    33.36062, 32.47544, 31.58298, 30.68328, 29.77641, 28.86244, 27.94145, 
    27.01353, 26.0788, 25.13736, 24.18934, 23.2349, 22.27417, 21.30732, 
    20.33454, 19.356, 18.3719, 17.38247, 16.38792, 15.38849, 14.38441, 
    13.37596, 12.36339, 11.34698, 10.32702, 9.303797, 8.277617, 7.248786, 
    6.217623, 5.184449, 4.149592, 3.113382, 2.076154, 1.038247, 0, -1.038247, 
    -2.076154, -3.113382, -4.149592, -5.184449, -6.217623, -7.248786, 
    -8.277617, -9.303797, -10.32702, -11.34698, -12.36339, -13.37596, 
    -14.38441, -15.38849, -16.38792, -17.38247, -18.3719, -19.356, -20.33454, 
    -21.30732, -22.27417, -23.2349, -24.18934, -25.13736, -26.0788, 
    -27.01353, -27.94145, -28.86244, -29.77641, -30.68328, -31.58298, 
    -32.47544, -33.36062, -34.23848, -35.10897, -35.97208, -36.8278, 
    -37.67612, -38.51705, -39.3506, -40.17678, -40.99562, -41.80717, 
    -42.61144, -43.4085, -44.19839, -44.98116,
  44.95763, 44.17486, 43.385, 42.58799, 41.78378, 40.97232, 40.15358, 
    39.32752, 38.49412, 37.65335, 36.80522, 35.94971, 35.08683, 34.21658, 
    33.33901, 32.45413, 31.56199, 30.66263, 29.75613, 28.84255, 27.92197, 
    26.99449, 26.06021, 25.11926, 24.17175, 23.21784, 22.25766, 21.29139, 
    20.3192, 19.34128, 18.35783, 17.36906, 16.37519, 15.37645, 14.37309, 
    13.36537, 12.35355, 11.33791, 10.31872, 9.29629, 8.270913, 7.242897, 
    6.212557, 5.180215, 4.146196, 3.11083, 2.074451, 1.037395, 0, -1.037395, 
    -2.074451, -3.11083, -4.146196, -5.180215, -6.212557, -7.242897, 
    -8.270913, -9.29629, -10.31872, -11.33791, -12.35355, -13.36537, 
    -14.37309, -15.37645, -16.37519, -17.36906, -18.35783, -19.34128, 
    -20.3192, -21.29139, -22.25766, -23.21784, -24.17175, -25.11926, 
    -26.06021, -26.99449, -27.92197, -28.84255, -29.75613, -30.66263, 
    -31.56199, -32.45413, -33.33901, -34.21658, -35.08683, -35.94971, 
    -36.80522, -37.65335, -38.49412, -39.32752, -40.15358, -40.97232, 
    -41.78378, -42.58799, -43.385, -44.17486, -44.95763,
  44.9247, 44.14195, 43.35213, 42.55518, 41.75106, 40.93972, 40.12112, 
    39.29524, 38.46204, 37.62151, 36.77364, 35.91842, 35.05586, 34.18597, 
    33.30878, 32.42432, 31.53263, 30.63375, 29.72776, 28.81473, 27.89473, 
    26.96786, 26.03424, 25.09396, 24.14717, 23.19399, 22.23459, 21.26912, 
    20.29777, 19.32071, 18.33815, 17.3503, 16.35738, 15.35962, 14.35726, 
    13.35057, 12.3398, 11.32522, 10.30712, 9.285798, 8.261543, 7.234665, 
    6.205477, 5.174297, 4.14145, 3.107264, 2.07207, 1.036204, 0, -1.036204, 
    -2.07207, -3.107264, -4.14145, -5.174297, -6.205477, -7.234665, 
    -8.261543, -9.285798, -10.30712, -11.32522, -12.3398, -13.35057, 
    -14.35726, -15.35962, -16.35738, -17.3503, -18.33815, -19.32071, 
    -20.29777, -21.26912, -22.23459, -23.19399, -24.14717, -25.09396, 
    -26.03424, -26.96786, -27.89473, -28.81473, -29.72776, -30.63375, 
    -31.53263, -32.42432, -33.30878, -34.18597, -35.05586, -35.91842, 
    -36.77364, -37.62151, -38.46204, -39.29524, -40.12112, -40.93972, 
    -41.75106, -42.55518, -43.35213, -44.14195, -44.9247,
  44.88241, 44.09967, 43.3099, 42.51304, 41.70904, 40.89785, 40.07944, 
    39.25378, 38.42085, 37.58062, 36.73308, 35.87823, 35.01609, 34.14666, 
    33.26997, 32.38604, 31.49493, 30.59668, 29.69135, 28.77902, 27.85977, 
    26.93369, 26.00089, 25.06149, 24.1156, 23.16338, 22.20498, 21.24054, 
    20.27026, 19.29432, 18.31291, 17.32624, 16.33454, 15.33803, 14.33696, 
    13.33158, 12.32215, 11.30894, 10.29224, 9.272337, 8.249522, 7.224104, 
    6.196393, 5.166705, 4.135361, 3.102689, 2.069016, 1.034675, 0, -1.034675, 
    -2.069016, -3.102689, -4.135361, -5.166705, -6.196393, -7.224104, 
    -8.249522, -9.272337, -10.29224, -11.30894, -12.32215, -13.33158, 
    -14.33696, -15.33803, -16.33454, -17.32624, -18.31291, -19.29432, 
    -20.27026, -21.24054, -22.20498, -23.16338, -24.1156, -25.06149, 
    -26.00089, -26.93369, -27.85977, -28.77902, -29.69135, -30.59668, 
    -31.49493, -32.38604, -33.26997, -34.14666, -35.01609, -35.87823, 
    -36.73308, -37.58062, -38.42085, -39.25378, -40.07944, -40.89785, 
    -41.70904, -42.51304, -43.3099, -44.09967, -44.88241,
  44.83077, 44.04806, 43.25835, 42.4616, 41.65775, 40.84675, 40.02857, 
    39.20319, 38.37057, 37.53071, 36.68359, 35.8292, 34.96757, 34.0987, 
    33.22261, 32.33934, 31.44894, 30.55145, 29.64693, 28.73546, 27.81712, 
    26.892, 25.96022, 25.02188, 24.07711, 23.12605, 22.16886, 21.20569, 
    20.23672, 19.26213, 18.28212, 17.2969, 16.30668, 15.3117, 14.3122, 
    13.30842, 12.30063, 11.2891, 10.2741, 9.255927, 8.23487, 7.211231, 
    6.18532, 5.15745, 4.127939, 3.097111, 2.065293, 1.032812, 0, -1.032812, 
    -2.065293, -3.097111, -4.127939, -5.15745, -6.18532, -7.211231, -8.23487, 
    -9.255927, -10.2741, -11.2891, -12.30063, -13.30842, -14.3122, -15.3117, 
    -16.30668, -17.2969, -18.28212, -19.26213, -20.23672, -21.20569, 
    -22.16886, -23.12605, -24.07711, -25.02188, -25.96022, -26.892, 
    -27.81712, -28.73546, -29.64693, -30.55145, -31.44894, -32.33934, 
    -33.22261, -34.0987, -34.96757, -35.8292, -36.68359, -37.53071, 
    -38.37057, -39.20319, -40.02857, -40.84675, -41.65775, -42.4616, 
    -43.25835, -44.04806, -44.83077,
  44.76982, 43.98714, 43.19752, 42.40089, 41.59722, 40.78645, 39.96855, 
    39.1435, 38.31126, 37.47184, 36.62521, 35.77137, 34.91034, 34.04213, 
    33.16676, 32.28428, 31.39471, 30.49811, 29.59455, 28.6841, 27.76684, 
    26.84286, 25.91227, 24.97519, 24.03174, 23.08206, 22.1263, 21.16462, 
    20.19719, 19.2242, 18.24584, 17.26232, 16.27386, 15.28068, 14.28303, 
    13.28114, 12.27528, 11.26572, 10.25273, 9.236594, 8.217607, 7.196066, 
    6.172276, 5.146547, 4.119196, 3.090542, 2.060907, 1.030618, 0, -1.030618, 
    -2.060907, -3.090542, -4.119196, -5.146547, -6.172276, -7.196066, 
    -8.217607, -9.236594, -10.25273, -11.26572, -12.27528, -13.28114, 
    -14.28303, -15.28068, -16.27386, -17.26232, -18.24584, -19.2242, 
    -20.19719, -21.16462, -22.1263, -23.08206, -24.03174, -24.97519, 
    -25.91227, -26.84286, -27.76684, -28.6841, -29.59455, -30.49811, 
    -31.39471, -32.28428, -33.16676, -34.04213, -34.91034, -35.77137, 
    -36.62521, -37.47184, -38.31126, -39.1435, -39.96855, -40.78645, 
    -41.59722, -42.40089, -43.19752, -43.98714, -44.76982,
  44.6996, 43.91697, 43.12745, 42.33097, 41.5275, 40.717, 39.89942, 39.07475, 
    38.24297, 37.40405, 36.55799, 35.70479, 34.84446, 33.97701, 33.10248, 
    32.22089, 31.33229, 30.43673, 29.53428, 28.625, 27.70898, 26.78632, 
    25.85711, 24.92148, 23.97954, 23.03145, 22.07734, 21.11737, 20.15172, 
    19.18058, 18.20412, 17.22256, 16.23612, 15.24501, 14.24948, 13.24977, 
    12.24614, 11.23884, 10.22816, 9.21437, 8.197762, 7.178632, 6.157281, 
    5.134015, 4.109146, 3.08299, 2.055866, 1.028095, 0, -1.028095, -2.055866, 
    -3.08299, -4.109146, -5.134015, -6.157281, -7.178632, -8.197762, 
    -9.21437, -10.22816, -11.23884, -12.24614, -13.24977, -14.24948, 
    -15.24501, -16.23612, -17.22256, -18.20412, -19.18058, -20.15172, 
    -21.11737, -22.07734, -23.03145, -23.97954, -24.92148, -25.85711, 
    -26.78632, -27.70898, -28.625, -29.53428, -30.43673, -31.33229, 
    -32.22089, -33.10248, -33.97701, -34.84446, -35.70479, -36.55799, 
    -37.40405, -38.24297, -39.07475, -39.89942, -40.717, -41.5275, -42.33097, 
    -43.12745, -43.91697, -44.6996,
  44.62016, 43.83758, 43.04817, 42.25187, 41.44865, 40.63845, 39.82125, 
    38.99702, 38.16574, 37.3274, 36.48199, 35.62952, 34.76999, 33.90341, 
    33.02983, 32.14926, 31.26176, 30.36738, 29.46618, 28.55823, 27.64362, 
    26.72244, 25.7948, 24.86081, 23.92059, 22.97429, 22.02205, 21.06402, 
    20.10039, 19.13132, 18.15702, 17.17768, 16.19351, 15.20475, 14.21162, 
    13.21437, 12.21324, 11.2085, 10.20043, 9.189286, 8.175366, 7.158958, 
    6.140359, 5.119872, 4.097805, 3.074468, 2.050177, 1.025248, 0, -1.025248, 
    -2.050177, -3.074468, -4.097805, -5.119872, -6.140359, -7.158958, 
    -8.175366, -9.189286, -10.20043, -11.2085, -12.21324, -13.21437, 
    -14.21162, -15.20475, -16.19351, -17.17768, -18.15702, -19.13132, 
    -20.10039, -21.06402, -22.02205, -22.97429, -23.92059, -24.86081, 
    -25.7948, -26.72244, -27.64362, -28.55823, -29.46618, -30.36738, 
    -31.26176, -32.14926, -33.02983, -33.90341, -34.76999, -35.62952, 
    -36.48199, -37.3274, -38.16574, -38.99702, -39.82125, -40.63845, 
    -41.44865, -42.25187, -43.04817, -43.83758, -44.62016,
  44.53154, 43.74903, 42.95976, 42.16367, 41.36071, 40.55087, 39.73409, 
    38.91036, 38.07965, 37.24197, 36.39729, 35.54563, 34.68699, 33.8214, 
    32.94887, 32.06945, 31.18319, 30.29012, 29.39032, 28.48387, 27.57083, 
    26.65132, 25.72542, 24.79326, 23.85496, 22.91066, 21.9605, 21.00464, 
    20.04325, 19.0765, 18.1046, 17.12773, 16.1461, 15.15995, 14.16949, 
    13.17497, 12.17664, 11.17476, 10.16958, 9.161384, 8.150454, 7.137073, 
    6.121536, 5.104141, 4.08519, 3.06499, 2.04385, 1.022082, 0, -1.022082, 
    -2.04385, -3.06499, -4.08519, -5.104141, -6.121536, -7.137073, -8.150454, 
    -9.161384, -10.16958, -11.17476, -12.17664, -13.17497, -14.16949, 
    -15.15995, -16.1461, -17.12773, -18.1046, -19.0765, -20.04325, -21.00464, 
    -21.9605, -22.91066, -23.85496, -24.79326, -25.72542, -26.65132, 
    -27.57083, -28.48387, -29.39032, -30.29012, -31.18319, -32.06945, 
    -32.94887, -33.8214, -34.68699, -35.54563, -36.39729, -37.24197, 
    -38.07965, -38.91036, -39.73409, -40.55087, -41.36071, -42.16367, 
    -42.95976, -43.74903, -44.53154,
  44.4338, 43.65138, 42.86227, 42.06641, 41.26377, 40.45432, 39.63801, 
    38.81484, 37.98478, 37.14782, 36.30396, 35.45321, 34.59556, 33.73105, 
    32.85971, 31.98156, 31.09665, 30.20505, 29.3068, 28.40199, 27.4907, 
    26.57302, 25.64905, 24.71892, 23.78273, 22.84064, 21.89278, 20.9393, 
    19.98038, 19.0162, 18.04693, 17.07278, 16.09396, 15.11067, 14.12316, 
    13.13165, 12.1364, 11.13764, 10.13566, 9.130703, 8.123061, 7.113011, 
    6.100842, 5.086846, 4.071321, 3.054569, 2.036894, 1.018601, 0, -1.018601, 
    -2.036894, -3.054569, -4.071321, -5.086846, -6.100842, -7.113011, 
    -8.123061, -9.130703, -10.13566, -11.13764, -12.1364, -13.13165, 
    -14.12316, -15.11067, -16.09396, -17.07278, -18.04693, -19.0162, 
    -19.98038, -20.9393, -21.89278, -22.84064, -23.78273, -24.71892, 
    -25.64905, -26.57302, -27.4907, -28.40199, -29.3068, -30.20505, 
    -31.09665, -31.98156, -32.85971, -33.73105, -34.59556, -35.45321, 
    -36.30396, -37.14782, -37.98478, -38.81484, -39.63801, -40.45432, 
    -41.26377, -42.06641, -42.86227, -43.65138, -44.4338,
  44.32701, 43.54469, 42.75576, 41.96017, 41.15789, 40.34887, 39.5331, 
    38.71054, 37.8812, 37.04504, 36.20208, 35.35233, 34.49578, 33.63246, 
    32.76241, 31.88566, 31.00225, 30.11224, 29.2157, 28.3127, 27.40331, 
    26.48764, 25.56579, 24.63787, 23.704, 22.76431, 21.81896, 20.8681, 
    19.91188, 18.95048, 17.9841, 17.01292, 16.03714, 15.05699, 14.07269, 
    13.08447, 12.09256, 11.09722, 10.09871, 9.097291, 8.09323, 7.086808, 
    6.078306, 5.068013, 4.05622, 3.043222, 2.029319, 1.014811, 0, -1.014811, 
    -2.029319, -3.043222, -4.05622, -5.068013, -6.078306, -7.086808, 
    -8.09323, -9.097291, -10.09871, -11.09722, -12.09256, -13.08447, 
    -14.07269, -15.05699, -16.03714, -17.01292, -17.9841, -18.95048, 
    -19.91188, -20.8681, -21.81896, -22.76431, -23.704, -24.63787, -25.56579, 
    -26.48764, -27.40331, -28.3127, -29.2157, -30.11224, -31.00225, 
    -31.88566, -32.76241, -33.63246, -34.49578, -35.35233, -36.20208, 
    -37.04504, -37.8812, -38.71054, -39.5331, -40.34887, -41.15789, 
    -41.96017, -42.75576, -43.54469, -44.32701,
  44.21122, 43.42903, 42.64032, 41.84503, 41.04314, 40.23461, 39.41943, 
    38.59755, 37.76899, 36.93372, 36.09175, 35.24308, 34.38773, 33.52573, 
    32.65709, 31.78186, 30.90008, 30.01182, 29.11712, 28.21608, 27.30877, 
    26.39529, 25.47573, 24.55021, 23.61885, 22.68178, 21.73915, 20.79111, 
    19.83782, 18.87945, 17.91618, 16.94822, 15.97575, 14.99899, 14.01815, 
    13.03348, 12.0452, 11.05355, 10.0588, 9.061195, 8.061007, 7.058504, 
    6.053965, 5.047671, 4.039908, 3.030967, 2.021138, 1.010717, 0, -1.010717, 
    -2.021138, -3.030967, -4.039908, -5.047671, -6.053965, -7.058504, 
    -8.061007, -9.061195, -10.0588, -11.05355, -12.0452, -13.03348, 
    -14.01815, -14.99899, -15.97575, -16.94822, -17.91618, -18.87945, 
    -19.83782, -20.79111, -21.73915, -22.68178, -23.61885, -24.55021, 
    -25.47573, -26.39529, -27.30877, -28.21608, -29.11712, -30.01182, 
    -30.90008, -31.78186, -32.65709, -33.52573, -34.38773, -35.24308, 
    -36.09175, -36.93372, -37.76899, -38.59755, -39.41943, -40.23461, 
    -41.04314, -41.84503, -42.64032, -43.42903, -44.21122,
  44.08652, 43.30448, 42.516, 41.72106, 40.91961, 40.11162, 39.29708, 
    38.47596, 37.64825, 36.81395, 35.97306, 35.12558, 34.27153, 33.41094, 
    32.54383, 31.67025, 30.79025, 29.90387, 29.01118, 28.11226, 27.20719, 
    26.29606, 25.37897, 24.45604, 23.52739, 22.59314, 21.65344, 20.70844, 
    19.7583, 18.80319, 17.84328, 16.87877, 15.90985, 14.93673, 13.95963, 
    12.97877, 11.99438, 11.0067, 10.01598, 9.02247, 8.026436, 7.02814, 
    6.027852, 5.025849, 4.022411, 3.017821, 2.012363, 1.006326, 0, -1.006326, 
    -2.012363, -3.017821, -4.022411, -5.025849, -6.027852, -7.02814, 
    -8.026436, -9.02247, -10.01598, -11.0067, -11.99438, -12.97877, 
    -13.95963, -14.93673, -15.90985, -16.87877, -17.84328, -18.80319, 
    -19.7583, -20.70844, -21.65344, -22.59314, -23.52739, -24.45604, 
    -25.37897, -26.29606, -27.20719, -28.11226, -29.01118, -29.90387, 
    -30.79025, -31.67025, -32.54383, -33.41094, -34.27153, -35.12558, 
    -35.97306, -36.81395, -37.64825, -38.47596, -39.29708, -40.11162, 
    -40.91961, -41.72106, -42.516, -43.30448, -44.08652,
  43.95298, 43.17111, 42.38291, 41.58834, 40.78738, 39.97999, 39.16616, 
    38.34586, 37.51908, 36.68583, 35.8461, 34.99992, 34.14728, 33.28822, 
    32.42276, 31.55096, 30.67286, 29.78851, 28.89797, 28.00133, 27.09867, 
    26.19007, 25.27564, 24.35549, 23.42973, 22.49851, 21.56195, 20.6202, 
    19.67343, 18.7218, 17.76548, 16.80466, 15.83954, 14.87031, 13.89719, 
    12.9204, 11.94017, 10.95672, 9.970306, 8.981172, 7.989569, 6.995759, 
    6.000007, 5.002581, 4.003754, 3.003803, 2.003006, 1.001644, 0, -1.001644, 
    -2.003006, -3.003803, -4.003754, -5.002581, -6.000007, -6.995759, 
    -7.989569, -8.981172, -9.970306, -10.95672, -11.94017, -12.9204, 
    -13.89719, -14.87031, -15.83954, -16.80466, -17.76548, -18.7218, 
    -19.67343, -20.6202, -21.56195, -22.49851, -23.42973, -24.35549, 
    -25.27564, -26.19007, -27.09867, -28.00133, -28.89797, -29.78851, 
    -30.67286, -31.55096, -32.42276, -33.28822, -34.14728, -34.99992, 
    -35.8461, -36.68583, -37.51908, -38.34586, -39.16616, -39.97999, 
    -40.78738, -41.58834, -42.38291, -43.17111, -43.95298,
  43.81068, 43.02901, 42.24112, 41.44698, 40.64656, 39.83982, 39.02676, 
    38.20735, 37.38158, 36.54947, 35.71101, 34.8662, 34.01508, 33.15767, 
    32.29399, 31.4241, 30.54803, 29.66586, 28.77763, 27.88343, 26.98333, 
    26.07744, 25.16584, 24.24865, 23.32599, 22.39799, 21.46477, 20.5265, 
    19.58331, 18.63538, 17.68288, 16.72599, 15.7649, 14.79981, 13.83093, 
    12.85847, 11.88264, 10.90369, 9.92185, 8.937356, 7.950458, 6.96141, 
    5.970469, 4.977899, 3.983964, 2.988935, 1.993082, 0.9966785, 0, 
    -0.9966785, -1.993082, -2.988935, -3.983964, -4.977899, -5.970469, 
    -6.96141, -7.950458, -8.937356, -9.92185, -10.90369, -11.88264, 
    -12.85847, -13.83093, -14.79981, -15.7649, -16.72599, -17.68288, 
    -18.63538, -19.58331, -20.5265, -21.46477, -22.39799, -23.32599, 
    -24.24865, -25.16584, -26.07744, -26.98333, -27.88343, -28.77763, 
    -29.66586, -30.54803, -31.4241, -32.29399, -33.15767, -34.01508, 
    -34.8662, -35.71101, -36.54947, -37.38158, -38.20735, -39.02676, 
    -39.83982, -40.64656, -41.44698, -42.24112, -43.02901, -43.81068,
  43.65969, 42.87827, 42.09073, 41.29707, 40.49723, 39.69121, 38.87898, 
    38.06054, 37.23587, 36.40498, 35.56787, 34.72456, 33.87507, 33.01942, 
    32.15764, 31.28979, 30.4159, 29.53604, 28.65027, 27.75867, 26.86131, 
    25.95829, 25.0497, 24.13567, 23.21629, 22.2917, 21.36204, 20.42744, 
    19.48806, 18.54405, 17.5956, 16.64287, 15.68605, 14.72534, 13.76093, 
    12.79304, 11.82189, 10.84769, 9.870676, 8.891085, 7.909157, 6.925138, 
    5.939281, 4.951838, 3.963069, 2.973237, 1.982603, 0.9914355, 0, 
    -0.9914355, -1.982603, -2.973237, -3.963069, -4.951838, -5.939281, 
    -6.925138, -7.909157, -8.891085, -9.870676, -10.84769, -11.82189, 
    -12.79304, -13.76093, -14.72534, -15.68605, -16.64287, -17.5956, 
    -18.54405, -19.48806, -20.42744, -21.36204, -22.2917, -23.21629, 
    -24.13567, -25.0497, -25.95829, -26.86131, -27.75867, -28.65027, 
    -29.53604, -30.4159, -31.28979, -32.15764, -33.01942, -33.87507, 
    -34.72456, -35.56787, -36.40498, -37.23587, -38.06054, -38.87898, 
    -39.69121, -40.49723, -41.29707, -42.09073, -42.87827, -43.65969,
  43.50012, 42.71897, 41.93184, 41.13869, 40.3395, 39.53426, 38.72294, 
    37.90554, 37.08205, 36.25248, 35.41682, 34.57511, 33.72735, 32.87358, 
    32.01384, 31.14815, 30.27658, 29.39919, 28.51603, 27.62718, 26.73272, 
    25.83275, 24.92736, 24.01665, 23.10075, 22.17978, 21.25386, 20.32315, 
    19.38778, 18.44792, 17.50373, 16.55539, 15.60307, 14.64697, 13.68729, 
    12.72422, 11.75798, 10.78878, 9.816853, 8.842422, 7.865723, 6.886996, 
    5.906484, 4.924435, 3.941099, 2.956731, 1.971586, 0.9859229, 0, 
    -0.9859229, -1.971586, -2.956731, -3.941099, -4.924435, -5.906484, 
    -6.886996, -7.865723, -8.842422, -9.816853, -10.78878, -11.75798, 
    -12.72422, -13.68729, -14.64697, -15.60307, -16.55539, -17.50373, 
    -18.44792, -19.38778, -20.32315, -21.25386, -22.17978, -23.10075, 
    -24.01665, -24.92736, -25.83275, -26.73272, -27.62718, -28.51603, 
    -29.39919, -30.27658, -31.14815, -32.01384, -32.87358, -33.72735, 
    -34.57511, -35.41682, -36.25248, -37.08205, -37.90554, -38.72294, 
    -39.53426, -40.3395, -41.13869, -41.93184, -42.71897, -43.50012,
  43.33206, 42.55122, 41.76453, 40.97196, 40.17348, 39.36908, 38.55875, 
    37.74247, 36.92025, 36.09208, 35.25799, 34.41798, 33.57207, 32.7203, 
    31.86271, 30.99933, 30.13022, 29.25543, 28.37503, 27.4891, 26.59771, 
    25.70096, 24.79893, 23.89175, 22.97951, 22.06234, 21.14038, 20.21375, 
    19.28261, 18.34711, 17.4074, 16.46367, 15.51608, 14.56483, 13.61009, 
    12.65208, 11.691, 10.72705, 9.760451, 8.791431, 7.820215, 6.847034, 
    5.872125, 4.895727, 3.918083, 2.93944, 1.960045, 0.9801481, 0, 
    -0.9801481, -1.960045, -2.93944, -3.918083, -4.895727, -5.872125, 
    -6.847034, -7.820215, -8.791431, -9.760451, -10.72705, -11.691, 
    -12.65208, -13.61009, -14.56483, -15.51608, -16.46367, -17.4074, 
    -18.34711, -19.28261, -20.21375, -21.14038, -22.06234, -22.97951, 
    -23.89175, -24.79893, -25.70096, -26.59771, -27.4891, -28.37503, 
    -29.25543, -30.13022, -30.99933, -31.86271, -32.7203, -33.57207, 
    -34.41798, -35.25799, -36.09208, -36.92025, -37.74247, -38.55875, 
    -39.36908, -40.17348, -40.97196, -41.76453, -42.55122, -43.33206,
  43.1556, 42.37512, 41.58892, 40.79699, 39.99928, 39.1958, 38.38652, 
    37.57145, 36.75058, 35.92393, 35.09149, 34.25329, 33.40936, 32.55971, 
    31.7044, 30.84346, 29.97694, 29.10491, 28.22743, 27.34457, 26.45642, 
    25.56305, 24.66457, 23.76108, 22.85269, 21.93953, 21.02171, 20.09937, 
    19.17266, 18.24172, 17.30672, 16.36782, 15.42518, 14.479, 13.52945, 
    12.57673, 11.62103, 10.66257, 9.701547, 8.738181, 7.772693, 6.805305, 
    5.836247, 4.865752, 3.894052, 2.921387, 1.947996, 0.9741191, 0, 
    -0.9741191, -1.947996, -2.921387, -3.894052, -4.865752, -5.836247, 
    -6.805305, -7.772693, -8.738181, -9.701547, -10.66257, -11.62103, 
    -12.57673, -13.52945, -14.479, -15.42518, -16.36782, -17.30672, 
    -18.24172, -19.17266, -20.09937, -21.02171, -21.93953, -22.85269, 
    -23.76108, -24.66457, -25.56305, -26.45642, -27.34457, -28.22743, 
    -29.10491, -29.97694, -30.84346, -31.7044, -32.55971, -33.40936, 
    -34.25329, -35.09149, -35.92393, -36.75058, -37.57145, -38.38652, 
    -39.1958, -39.99928, -40.79699, -41.58892, -42.37512, -43.1556,
  42.97084, 42.19077, 41.40512, 40.61388, 39.81702, 39.01452, 38.20639, 
    37.39261, 36.57319, 35.74813, 34.91746, 34.08119, 33.23934, 32.39194, 
    31.53904, 30.68068, 29.8169, 28.94778, 28.07337, 27.19374, 26.30898, 
    25.41917, 24.52441, 23.6248, 22.72045, 21.81147, 20.89799, 19.98014, 
    19.05806, 18.1319, 17.20181, 16.26795, 15.33048, 14.38959, 13.44545, 
    12.49824, 11.54817, 10.59543, 9.640213, 8.682739, 7.723217, 6.761864, 
    5.7989, 4.834549, 3.869038, 2.902596, 1.935454, 0.9678438, 0, -0.9678438, 
    -1.935454, -2.902596, -3.869038, -4.834549, -5.7989, -6.761864, 
    -7.723217, -8.682739, -9.640213, -10.59543, -11.54817, -12.49824, 
    -13.44545, -14.38959, -15.33048, -16.26795, -17.20181, -18.1319, 
    -19.05806, -19.98014, -20.89799, -21.81147, -22.72045, -23.6248, 
    -24.52441, -25.41917, -26.30898, -27.19374, -28.07337, -28.94778, 
    -29.8169, -30.68068, -31.53904, -32.39194, -33.23934, -34.08119, 
    -34.91746, -35.74813, -36.57319, -37.39261, -38.20639, -39.01452, 
    -39.81702, -40.61388, -41.40512, -42.19077, -42.97084,
  42.77788, 41.99827, 41.21324, 40.42275, 39.6268, 38.82537, 38.01846, 
    37.20607, 36.38819, 35.56485, 34.73605, 33.90181, 33.06216, 32.21714, 
    31.36679, 30.51114, 29.65025, 28.78417, 27.91298, 27.03675, 26.15555, 
    25.26947, 24.3786, 23.48304, 22.5829, 21.6783, 20.76936, 19.85619, 
    18.93895, 18.01776, 17.09279, 16.16418, 15.2321, 14.29671, 13.3582, 
    12.41673, 11.47251, 10.52571, 9.576528, 8.625175, 7.671851, 6.716765, 
    5.760129, 4.802159, 3.843073, 2.883091, 1.922435, 0.9613302, 0, 
    -0.9613302, -1.922435, -2.883091, -3.843073, -4.802159, -5.760129, 
    -6.716765, -7.671851, -8.625175, -9.576528, -10.52571, -11.47251, 
    -12.41673, -13.3582, -14.29671, -15.2321, -16.16418, -17.09279, 
    -18.01776, -18.93895, -19.85619, -20.76936, -21.6783, -22.5829, 
    -23.48304, -24.3786, -25.26947, -26.15555, -27.03675, -27.91298, 
    -28.78417, -29.65025, -30.51114, -31.36679, -32.21714, -33.06216, 
    -33.90181, -34.73605, -35.56485, -36.38819, -37.20607, -38.01846, 
    -38.82537, -39.6268, -40.42275, -41.21324, -41.99827, -42.77788,
  42.57683, 41.79774, 41.01338, 40.22372, 39.42876, 38.62848, 37.82288, 
    37.01196, 36.19573, 35.3742, 34.54738, 33.7153, 32.87798, 32.03546, 
    31.18778, 30.33498, 29.47712, 28.61425, 27.74643, 26.87375, 25.99627, 
    25.11408, 24.22728, 23.33596, 22.44022, 21.54018, 20.63595, 19.72766, 
    18.81544, 17.89944, 16.97978, 16.05663, 15.13014, 14.20047, 13.2678, 
    12.33229, 11.39412, 10.45349, 9.510569, 8.565559, 7.618658, 6.670065, 
    5.719984, 4.768622, 3.816189, 2.862896, 1.908957, 0.9545865, 0, 
    -0.9545865, -1.908957, -2.862896, -3.816189, -4.768622, -5.719984, 
    -6.670065, -7.618658, -8.565559, -9.510569, -10.45349, -11.39412, 
    -12.33229, -13.2678, -14.20047, -15.13014, -16.05663, -16.97978, 
    -17.89944, -18.81544, -19.72766, -20.63595, -21.54018, -22.44022, 
    -23.33596, -24.22728, -25.11408, -25.99627, -26.87375, -27.74643, 
    -28.61425, -29.47712, -30.33498, -31.18778, -32.03546, -32.87798, 
    -33.7153, -34.54738, -35.3742, -36.19573, -37.01196, -37.82288, 
    -38.62848, -39.42876, -40.22372, -41.01338, -41.79774, -42.57683,
  42.36781, 41.5893, 40.80568, 40.01692, 39.22302, 38.42397, 37.61977, 
    36.81043, 35.99594, 35.17633, 34.35161, 33.5218, 32.68693, 31.84704, 
    31.00217, 30.15236, 29.29767, 28.43815, 27.57387, 26.70489, 25.8313, 
    24.95318, 24.07061, 23.18369, 22.29253, 21.39723, 20.49791, 19.59469, 
    18.68769, 17.77705, 16.86292, 15.94542, 15.02473, 14.10098, 13.17436, 
    12.24501, 11.31312, 10.37886, 9.442413, 8.503963, 7.563702, 6.621819, 
    5.678512, 4.733978, 3.788419, 2.842036, 1.895035, 0.947621, 0, -0.947621, 
    -1.895035, -2.842036, -3.788419, -4.733978, -5.678512, -6.621819, 
    -7.563702, -8.503963, -9.442413, -10.37886, -11.31312, -12.24501, 
    -13.17436, -14.10098, -15.02473, -15.94542, -16.86292, -17.77705, 
    -18.68769, -19.59469, -20.49791, -21.39723, -22.29253, -23.18369, 
    -24.07061, -24.95318, -25.8313, -26.70489, -27.57387, -28.43815, 
    -29.29767, -30.15236, -31.00217, -31.84704, -32.68693, -33.5218, 
    -34.35161, -35.17633, -35.99594, -36.81043, -37.61977, -38.42397, 
    -39.22302, -40.01692, -40.80568, -41.5893, -42.36781,
  42.15091, 41.37305, 40.59023, 39.80246, 39.00971, 38.21198, 37.40928, 
    36.6016, 35.78897, 34.97139, 34.14888, 33.32146, 32.48917, 31.65205, 
    30.81012, 29.96344, 29.11207, 28.25605, 27.39545, 26.53034, 25.6608, 
    24.7869, 23.90874, 23.0264, 22.13999, 21.24961, 20.35538, 19.45741, 
    18.55582, 17.65075, 16.74232, 15.83068, 14.91598, 13.99836, 13.07798, 
    12.155, 11.22959, 10.30191, 9.372141, 8.44046, 7.507047, 6.572086, 
    5.635764, 4.69827, 3.759796, 2.820537, 1.880687, 0.9404421, 0, 
    -0.9404421, -1.880687, -2.820537, -3.759796, -4.69827, -5.635764, 
    -6.572086, -7.507047, -8.44046, -9.372141, -10.30191, -11.22959, -12.155, 
    -13.07798, -13.99836, -14.91598, -15.83068, -16.74232, -17.65075, 
    -18.55582, -19.45741, -20.35538, -21.24961, -22.13999, -23.0264, 
    -23.90874, -24.7869, -25.6608, -26.53034, -27.39545, -28.25605, 
    -29.11207, -29.96344, -30.81012, -31.65205, -32.48917, -33.32146, 
    -34.14888, -34.97139, -35.78897, -36.6016, -37.40928, -38.21198, 
    -39.00971, -39.80246, -40.59023, -41.37305, -42.15091,
  41.92625, 41.14911, 40.36718, 39.58046, 38.78895, 37.99264, 37.19153, 
    36.38563, 35.57495, 34.75951, 33.93933, 33.11443, 32.28485, 31.45062, 
    30.61178, 29.76838, 28.92046, 28.06809, 27.21133, 26.35024, 25.48491, 
    24.6154, 23.74181, 22.86423, 21.98275, 21.09747, 20.20851, 19.31597, 
    18.41997, 17.52065, 16.61812, 15.71253, 14.804, 13.8927, 12.97877, 
    12.06235, 11.14361, 10.22272, 9.299832, 8.375121, 7.448759, 6.520922, 
    5.591787, 4.661538, 3.730354, 2.798423, 1.865928, 0.9330581, 0, 
    -0.9330581, -1.865928, -2.798423, -3.730354, -4.661538, -5.591787, 
    -6.520922, -7.448759, -8.375121, -9.299832, -10.22272, -11.14361, 
    -12.06235, -12.97877, -13.8927, -14.804, -15.71253, -16.61812, -17.52065, 
    -18.41997, -19.31597, -20.20851, -21.09747, -21.98275, -22.86423, 
    -23.74181, -24.6154, -25.48491, -26.35024, -27.21133, -28.06809, 
    -28.92046, -29.76838, -30.61178, -31.45062, -32.28485, -33.11443, 
    -33.93933, -34.75951, -35.57495, -36.38563, -37.19153, -37.99264, 
    -38.78895, -39.58046, -40.36718, -41.14911, -41.92625,
  41.69396, 40.9176, 40.13664, 39.35107, 38.56088, 37.76608, 36.96666, 
    36.16264, 35.35404, 34.54086, 33.72313, 32.90088, 32.07413, 31.24292, 
    30.4073, 29.56732, 28.72301, 27.87444, 27.02167, 26.16477, 25.3038, 
    24.43885, 23.57, 22.69734, 21.82095, 20.94095, 20.05743, 19.1705, 
    18.28028, 17.38689, 16.49044, 15.59108, 14.68893, 13.78413, 12.87683, 
    11.96717, 11.0553, 10.14138, 9.225567, 8.308019, 7.388902, 6.468383, 
    5.546633, 4.623823, 3.700126, 2.775718, 1.850776, 0.9254774, 0, 
    -0.9254774, -1.850776, -2.775718, -3.700126, -4.623823, -5.546633, 
    -6.468383, -7.388902, -8.308019, -9.225567, -10.14138, -11.0553, 
    -11.96717, -12.87683, -13.78413, -14.68893, -15.59108, -16.49044, 
    -17.38689, -18.28028, -19.1705, -20.05743, -20.94095, -21.82095, 
    -22.69734, -23.57, -24.43885, -25.3038, -26.16477, -27.02167, -27.87444, 
    -28.72301, -29.56732, -30.4073, -31.24292, -32.07413, -32.90088, 
    -33.72313, -34.54086, -35.35404, -36.16264, -36.96666, -37.76608, 
    -38.56088, -39.35107, -40.13664, -40.9176, -41.69396,
  41.45414, 40.67865, 39.89874, 39.1144, 38.32563, 37.53244, 36.73482, 
    35.9328, 35.12637, 34.31557, 33.50042, 32.68093, 31.85715, 31.02912, 
    30.19686, 29.36043, 28.51988, 27.67526, 26.82663, 25.97407, 25.11763, 
    24.2574, 23.39345, 22.52588, 21.65476, 20.7802, 19.9023, 19.02115, 
    18.13688, 17.2496, 16.35942, 15.46647, 14.57087, 13.67276, 12.77227, 
    11.86955, 10.96474, 10.05798, 9.149424, 8.239225, 7.327541, 6.414529, 
    5.50035, 4.585167, 3.669145, 2.752449, 1.835248, 0.9177083, 0, 
    -0.9177083, -1.835248, -2.752449, -3.669145, -4.585167, -5.50035, 
    -6.414529, -7.327541, -8.239225, -9.149424, -10.05798, -10.96474, 
    -11.86955, -12.77227, -13.67276, -14.57087, -15.46647, -16.35942, 
    -17.2496, -18.13688, -19.02115, -19.9023, -20.7802, -21.65476, -22.52588, 
    -23.39345, -24.2574, -25.11763, -25.97407, -26.82663, -27.67526, 
    -28.51988, -29.36043, -30.19686, -31.02912, -31.85715, -32.68093, 
    -33.50042, -34.31557, -35.12637, -35.9328, -36.73482, -37.53244, 
    -38.32563, -39.1144, -39.89874, -40.67865, -41.45414,
  41.20691, 40.43238, 39.6536, 38.87059, 38.08334, 37.29186, 36.49615, 
    35.69623, 34.89211, 34.08381, 33.27135, 32.45477, 31.63409, 30.80936, 
    29.9806, 29.14787, 28.31122, 27.47071, 26.62638, 25.77831, 24.92656, 
    24.0712, 23.21232, 22.35, 21.48432, 20.61537, 19.74325, 18.86807, 
    17.98992, 17.10892, 16.22518, 15.33881, 14.44994, 13.5587, 12.66521, 
    11.7696, 10.87202, 9.972599, 9.071482, 8.168813, 7.26474, 6.359414, 
    5.452987, 4.545611, 3.637443, 2.72864, 1.819359, 0.9097592, 0, 
    -0.9097592, -1.819359, -2.72864, -3.637443, -4.545611, -5.452987, 
    -6.359414, -7.26474, -8.168813, -9.071482, -9.972599, -10.87202, 
    -11.7696, -12.66521, -13.5587, -14.44994, -15.33881, -16.22518, 
    -17.10892, -17.98992, -18.86807, -19.74325, -20.61537, -21.48432, -22.35, 
    -23.21232, -24.0712, -24.92656, -25.77831, -26.62638, -27.47071, 
    -28.31122, -29.14787, -29.9806, -30.80936, -31.63409, -32.45477, 
    -33.27135, -34.08381, -34.89211, -35.69623, -36.49615, -37.29186, 
    -38.08334, -38.87059, -39.6536, -40.43238, -41.20691,
  40.9524, 40.1789, 39.40136, 38.61978, 37.83415, 37.04449, 36.2508, 
    35.45309, 34.6514, 33.84572, 33.03609, 32.22254, 31.4051, 30.5838, 
    29.75869, 28.92981, 28.09721, 27.26094, 26.42107, 25.57764, 24.73074, 
    23.88042, 23.02677, 22.16986, 21.30978, 20.44661, 19.58045, 18.71139, 
    17.83953, 16.96498, 16.08784, 15.20823, 14.32627, 13.44206, 12.55573, 
    11.66742, 10.77724, 9.885328, 8.99182, 8.096853, 7.200565, 6.303097, 
    5.404592, 4.505196, 3.605054, 2.704315, 1.803126, 0.9016382, 0, 
    -0.9016382, -1.803126, -2.704315, -3.605054, -4.505196, -5.404592, 
    -6.303097, -7.200565, -8.096853, -8.99182, -9.885328, -10.77724, 
    -11.66742, -12.55573, -13.44206, -14.32627, -15.20823, -16.08784, 
    -16.96498, -17.83953, -18.71139, -19.58045, -20.44661, -21.30978, 
    -22.16986, -23.02677, -23.88042, -24.73074, -25.57764, -26.42107, 
    -27.26094, -28.09721, -28.92981, -29.75869, -30.5838, -31.4051, 
    -32.22254, -33.03609, -33.84572, -34.6514, -35.45309, -36.2508, 
    -37.04449, -37.83415, -38.61978, -39.40136, -40.1789, -40.9524,
  40.69072, 39.91835, 39.14214, 38.36209, 37.57819, 36.79046, 35.9989, 
    35.20354, 34.40438, 33.60146, 32.79479, 31.98441, 31.17034, 30.35262, 
    29.5313, 28.70641, 27.87801, 27.04614, 26.21087, 25.37224, 24.53034, 
    23.68522, 22.83695, 21.98561, 21.13129, 20.27407, 19.41402, 18.55125, 
    17.68585, 16.81791, 15.94755, 15.07486, 14.19996, 13.32295, 12.44396, 
    11.5631, 10.68048, 9.79625, 8.910519, 8.023417, 7.135077, 6.245632, 
    5.355214, 4.463961, 3.57201, 2.679499, 1.786567, 0.8933536, 0, 
    -0.8933536, -1.786567, -2.679499, -3.57201, -4.463961, -5.355214, 
    -6.245632, -7.135077, -8.023417, -8.910519, -9.79625, -10.68048, 
    -11.5631, -12.44396, -13.32295, -14.19996, -15.07486, -15.94755, 
    -16.81791, -17.68585, -18.55125, -19.41402, -20.27407, -21.13129, 
    -21.98561, -22.83695, -23.68522, -24.53034, -25.37224, -26.21087, 
    -27.04614, -27.87801, -28.70641, -29.5313, -30.35262, -31.17034, 
    -31.98441, -32.79479, -33.60146, -34.40438, -35.20354, -35.9989, 
    -36.79046, -37.57819, -38.36209, -39.14214, -39.91835, -40.69072,
  40.42199, 39.65086, 38.87608, 38.09766, 37.3156, 36.52991, 35.74061, 
    34.94771, 34.15122, 33.35118, 32.5476, 31.74052, 30.92996, 30.11596, 
    29.29857, 28.47782, 27.65377, 26.82645, 25.99593, 25.16227, 24.32551, 
    23.48574, 22.64302, 21.79742, 20.94901, 20.09789, 19.24412, 18.38779, 
    17.52901, 16.66785, 15.80442, 14.93881, 14.07113, 13.20149, 12.32998, 
    11.45673, 10.58185, 9.705451, 8.827652, 7.948575, 7.068341, 6.187074, 
    5.304901, 4.421948, 3.538343, 2.654216, 1.769696, 0.8849133, 0, 
    -0.8849133, -1.769696, -2.654216, -3.538343, -4.421948, -5.304901, 
    -6.187074, -7.068341, -7.948575, -8.827652, -9.705451, -10.58185, 
    -11.45673, -12.32998, -13.20149, -14.07113, -14.93881, -15.80442, 
    -16.66785, -17.52901, -18.38779, -19.24412, -20.09789, -20.94901, 
    -21.79742, -22.64302, -23.48574, -24.32551, -25.16227, -25.99593, 
    -26.82645, -27.65377, -28.47782, -29.29857, -30.11596, -30.92996, 
    -31.74052, -32.5476, -33.35118, -34.15122, -34.94771, -35.74061, 
    -36.52991, -37.3156, -38.09766, -38.87608, -39.65086, -40.42199,
  40.14635, 39.37654, 38.6033, 37.82662, 37.04652, 36.26299, 35.47607, 
    34.68575, 33.89207, 33.09504, 32.29469, 31.49104, 30.68413, 29.874, 
    29.06068, 28.24422, 27.42466, 26.60204, 25.77643, 24.94787, 24.11643, 
    23.28216, 22.44514, 21.60542, 20.76309, 19.91821, 19.07088, 18.22116, 
    17.36914, 16.51492, 15.65857, 14.8002, 13.9399, 13.07777, 12.21391, 
    11.34843, 10.48143, 9.613013, 8.743299, 7.872395, 7.000417, 6.12748, 
    5.253699, 4.379195, 3.504085, 2.628489, 1.752529, 0.8763254, 0, 
    -0.8763254, -1.752529, -2.628489, -3.504085, -4.379195, -5.253699, 
    -6.12748, -7.000417, -7.872395, -8.743299, -9.613013, -10.48143, 
    -11.34843, -12.21391, -13.07777, -13.9399, -14.8002, -15.65857, 
    -16.51492, -17.36914, -18.22116, -19.07088, -19.91821, -20.76309, 
    -21.60542, -22.44514, -23.28216, -24.11643, -24.94787, -25.77643, 
    -26.60204, -27.42466, -28.24422, -29.06068, -29.874, -30.68413, 
    -31.49104, -32.29469, -33.09504, -33.89207, -34.68575, -35.47607, 
    -36.26299, -37.04652, -37.82662, -38.6033, -39.37654, -40.14635,
  39.8639, 39.09554, 38.32394, 37.54912, 36.77109, 35.98985, 35.20542, 
    34.41782, 33.62707, 32.83318, 32.03619, 31.23613, 30.43301, 29.62689, 
    28.81779, 28.00576, 27.19084, 26.37307, 25.55252, 24.72922, 23.90323, 
    23.07462, 22.24345, 21.40977, 20.57367, 19.7352, 18.89445, 18.05148, 
    17.20639, 16.35925, 15.51014, 14.65916, 13.80638, 12.95192, 12.09585, 
    11.23828, 10.3793, 9.519018, 8.657532, 7.794946, 6.931367, 6.066901, 
    5.201655, 4.335741, 3.469266, 2.602343, 1.735083, 0.8675976, 0, 
    -0.8675976, -1.735083, -2.602343, -3.469266, -4.335741, -5.201655, 
    -6.066901, -6.931367, -7.794946, -8.657532, -9.519018, -10.3793, 
    -11.23828, -12.09585, -12.95192, -13.80638, -14.65916, -15.51014, 
    -16.35925, -17.20639, -18.05148, -18.89445, -19.7352, -20.57367, 
    -21.40977, -22.24345, -23.07462, -23.90323, -24.72922, -25.55252, 
    -26.37307, -27.19084, -28.00576, -28.81779, -29.62689, -30.43301, 
    -31.23613, -32.03619, -32.83318, -33.62707, -34.41782, -35.20542, 
    -35.98985, -36.77109, -37.54912, -38.32394, -39.09554, -39.8639,
  39.57478, 38.80796, 38.03813, 37.26529, 36.48944, 35.71062, 34.92882, 
    34.14407, 33.35638, 32.56578, 31.77229, 30.97594, 30.17676, 29.37479, 
    28.57006, 27.76261, 26.95247, 26.13971, 25.32435, 24.50646, 23.68609, 
    22.86328, 22.03811, 21.21062, 20.38089, 19.54898, 18.71496, 17.8789, 
    17.04088, 16.20097, 15.35924, 14.51579, 13.67069, 12.82403, 11.97589, 
    11.12637, 10.27556, 9.423547, 8.570426, 7.716295, 6.86125, 6.00539, 
    5.148814, 4.291623, 3.433917, 2.575799, 1.717372, 0.8587376, 0, 
    -0.8587376, -1.717372, -2.575799, -3.433917, -4.291623, -5.148814, 
    -6.00539, -6.86125, -7.716295, -8.570426, -9.423547, -10.27556, 
    -11.12637, -11.97589, -12.82403, -13.67069, -14.51579, -15.35924, 
    -16.20097, -17.04088, -17.8789, -18.71496, -19.54898, -20.38089, 
    -21.21062, -22.03811, -22.86328, -23.68609, -24.50646, -25.32435, 
    -26.13971, -26.95247, -27.76261, -28.57006, -29.37479, -30.17676, 
    -30.97594, -31.77229, -32.56578, -33.35638, -34.14407, -34.92882, 
    -35.71062, -36.48944, -37.26529, -38.03813, -38.80796, -39.57478,
  39.27911, 38.51395, 37.746, 36.97525, 36.20173, 35.42545, 34.64641, 
    33.86464, 33.08015, 32.29297, 31.50312, 30.71063, 29.91554, 29.11786, 
    28.31764, 27.51491, 26.70972, 25.9021, 25.0921, 24.27976, 23.46515, 
    22.6483, 21.82927, 21.00812, 20.18491, 19.35971, 18.53256, 17.70355, 
    16.87274, 16.0402, 15.20599, 14.37021, 13.53292, 12.6942, 11.85414, 
    11.0128, 10.17029, 9.326677, 8.482054, 7.636507, 6.790126, 5.943, 
    5.095221, 4.246879, 3.398068, 2.548881, 1.699411, 0.8497528, 0, 
    -0.8497528, -1.699411, -2.548881, -3.398068, -4.246879, -5.095221, 
    -5.943, -6.790126, -7.636507, -8.482054, -9.326677, -10.17029, -11.0128, 
    -11.85414, -12.6942, -13.53292, -14.37021, -15.20599, -16.0402, 
    -16.87274, -17.70355, -18.53256, -19.35971, -20.18491, -21.00812, 
    -21.82927, -22.6483, -23.46515, -24.27976, -25.0921, -25.9021, -26.70972, 
    -27.51491, -28.31764, -29.11786, -29.91554, -30.71063, -31.50312, 
    -32.29297, -33.08015, -33.86464, -34.64641, -35.42545, -36.20173, 
    -36.97525, -37.746, -38.51395, -39.27911,
  38.977, 38.21363, 37.44768, 36.67916, 35.90809, 35.13448, 34.35833, 
    33.57967, 32.79853, 32.01491, 31.22885, 30.44036, 29.64949, 28.85626, 
    28.0607, 27.26284, 26.46273, 25.6604, 24.85591, 24.04927, 23.24056, 
    22.42981, 21.61708, 20.80241, 19.98587, 19.16751, 18.34738, 17.52556, 
    16.7021, 15.87706, 15.05052, 14.22254, 13.39319, 12.56255, 11.73068, 
    10.89766, 10.06357, 9.228487, 8.392486, 7.555646, 6.718051, 5.87978, 
    5.040917, 4.201545, 3.361748, 2.52161, 1.681216, 0.8406506, 0, 
    -0.8406506, -1.681216, -2.52161, -3.361748, -4.201545, -5.040917, 
    -5.87978, -6.718051, -7.555646, -8.392486, -9.228487, -10.06357, 
    -10.89766, -11.73068, -12.56255, -13.39319, -14.22254, -15.05052, 
    -15.87706, -16.7021, -17.52556, -18.34738, -19.16751, -19.98587, 
    -20.80241, -21.61708, -22.42981, -23.24056, -24.04927, -24.85591, 
    -25.6604, -26.46273, -27.26284, -28.0607, -28.85626, -29.64949, 
    -30.44036, -31.22885, -32.01491, -32.79853, -33.57967, -34.35833, 
    -35.13448, -35.90809, -36.67916, -37.44768, -38.21363, -38.977,
  38.66859, 37.90713, 37.14331, 36.37715, 35.60866, 34.83784, 34.06473, 
    33.28933, 32.51167, 31.73176, 30.94962, 30.16529, 29.37879, 28.59014, 
    27.79938, 27.00655, 26.21167, 25.41478, 24.61593, 23.81515, 23.01249, 
    22.20798, 21.40168, 20.59364, 19.7839, 18.97252, 18.15956, 17.34505, 
    16.52908, 15.71168, 14.89293, 14.07288, 13.2516, 12.42916, 11.60561, 
    10.78103, 9.955491, 9.129053, 8.30179, 7.473776, 6.645081, 5.815781, 
    4.985948, 4.155657, 3.324986, 2.494007, 1.662799, 0.8314381, 0, 
    -0.8314381, -1.662799, -2.494007, -3.324986, -4.155657, -4.985948, 
    -5.815781, -6.645081, -7.473776, -8.30179, -9.129053, -9.955491, 
    -10.78103, -11.60561, -12.42916, -13.2516, -14.07288, -14.89293, 
    -15.71168, -16.52908, -17.34505, -18.15956, -18.97252, -19.7839, 
    -20.59364, -21.40168, -22.20798, -23.01249, -23.81515, -24.61593, 
    -25.41478, -26.21167, -27.00655, -27.79938, -28.59014, -29.37879, 
    -30.16529, -30.94962, -31.73176, -32.51167, -33.28933, -34.06473, 
    -34.83784, -35.60866, -36.37715, -37.14331, -37.90713, -38.66859,
  38.354, 37.59457, 36.83301, 36.06934, 35.30357, 34.5357, 33.76576, 
    32.99376, 32.21972, 31.44366, 30.6656, 29.88556, 29.10357, 28.31966, 
    27.53386, 26.74619, 25.95669, 25.16539, 24.37232, 23.57754, 22.78106, 
    21.98295, 21.18322, 20.38194, 19.57915, 18.77489, 17.96921, 17.16216, 
    16.3538, 15.54417, 14.73334, 13.92135, 13.10826, 12.29414, 11.47903, 
    10.66301, 9.846126, 9.028447, 8.210036, 7.390956, 6.571271, 5.751048, 
    4.930352, 4.10925, 3.287808, 2.466094, 1.644176, 0.8221223, 0, 
    -0.8221223, -1.644176, -2.466094, -3.287808, -4.10925, -4.930352, 
    -5.751048, -6.571271, -7.390956, -8.210036, -9.028447, -9.846126, 
    -10.66301, -11.47903, -12.29414, -13.10826, -13.92135, -14.73334, 
    -15.54417, -16.3538, -17.16216, -17.96921, -18.77489, -19.57915, 
    -20.38194, -21.18322, -21.98295, -22.78106, -23.57754, -24.37232, 
    -25.16539, -25.95669, -26.74619, -27.53386, -28.31966, -29.10357, 
    -29.88556, -30.6656, -31.44366, -32.21972, -32.99376, -33.76576, 
    -34.5357, -35.30357, -36.06934, -36.83301, -37.59457, -38.354,
  38.03334, 37.27608, 36.51693, 35.75588, 34.99296, 34.22818, 33.46156, 
    32.6931, 31.92283, 31.15076, 30.37692, 29.60133, 28.82401, 28.04498, 
    27.26427, 26.48191, 25.69794, 24.91236, 24.12524, 23.33659, 22.54645, 
    21.75485, 20.96184, 20.16746, 19.37174, 18.57473, 17.77647, 16.97701, 
    16.17639, 15.37465, 14.57185, 13.76804, 12.96326, 12.15757, 11.35102, 
    10.54366, 9.735553, 8.926742, 8.117288, 7.307246, 6.496675, 5.68563, 
    4.874171, 4.062356, 3.250242, 2.437891, 1.62536, 0.8127099, 0, 
    -0.8127099, -1.62536, -2.437891, -3.250242, -4.062356, -4.874171, 
    -5.68563, -6.496675, -7.307246, -8.117288, -8.926742, -9.735553, 
    -10.54366, -11.35102, -12.15757, -12.96326, -13.76804, -14.57185, 
    -15.37465, -16.17639, -16.97701, -17.77647, -18.57473, -19.37174, 
    -20.16746, -20.96184, -21.75485, -22.54645, -23.33659, -24.12524, 
    -24.91236, -25.69794, -26.48191, -27.26427, -28.04498, -28.82401, 
    -29.60133, -30.37692, -31.15076, -31.92283, -32.6931, -33.46156, 
    -34.22818, -34.99296, -35.75588, -36.51693, -37.27608, -38.03334,
  37.70675, 36.95179, 36.19517, 35.4369, 34.67698, 33.91543, 33.15226, 
    32.3875, 31.62114, 30.85322, 30.08375, 29.31275, 28.54023, 27.76624, 
    26.99077, 26.21387, 25.43556, 24.65587, 23.87482, 23.09244, 22.30877, 
    21.52384, 20.73768, 19.95033, 19.16182, 18.37219, 17.58147, 16.78971, 
    15.99695, 15.20323, 14.40859, 13.61306, 12.81671, 12.01956, 11.22167, 
    10.42309, 9.623848, 8.824006, 8.023608, 7.222704, 6.421341, 5.619571, 
    4.817443, 4.015007, 3.212315, 2.409416, 1.606363, 0.8032075, 0, 
    -0.8032075, -1.606363, -2.409416, -3.212315, -4.015007, -4.817443, 
    -5.619571, -6.421341, -7.222704, -8.023608, -8.824006, -9.623848, 
    -10.42309, -11.22167, -12.01956, -12.81671, -13.61306, -14.40859, 
    -15.20323, -15.99695, -16.78971, -17.58147, -18.37219, -19.16182, 
    -19.95033, -20.73768, -21.52384, -22.30877, -23.09244, -23.87482, 
    -24.65587, -25.43556, -26.21387, -26.99077, -27.76624, -28.54023, 
    -29.31275, -30.08375, -30.85322, -31.62114, -32.3875, -33.15226, 
    -33.91543, -34.67698, -35.4369, -36.19517, -36.95179, -37.70675,
  37.37434, 36.62183, 35.86789, 35.11252, 34.35575, 33.59758, 32.83802, 
    32.0771, 31.31481, 30.55118, 29.78622, 29.01996, 28.25241, 27.48358, 
    26.71351, 25.94222, 25.16972, 24.39604, 23.6212, 22.84524, 22.06818, 
    21.29005, 20.51087, 19.73068, 18.9495, 18.16737, 17.38433, 16.6004, 
    15.81561, 15.03002, 14.24364, 13.45652, 12.66869, 11.88019, 11.09107, 
    10.30135, 9.511086, 8.720308, 7.929061, 7.137385, 6.345323, 5.552916, 
    4.760206, 3.967237, 3.17405, 2.38069, 1.587199, 0.7936214, 0, -0.7936214, 
    -1.587199, -2.38069, -3.17405, -3.967237, -4.760206, -5.552916, 
    -6.345323, -7.137385, -7.929061, -8.720308, -9.511086, -10.30135, 
    -11.09107, -11.88019, -12.66869, -13.45652, -14.24364, -15.03002, 
    -15.81561, -16.6004, -17.38433, -18.16737, -18.9495, -19.73068, 
    -20.51087, -21.29005, -22.06818, -22.84524, -23.6212, -24.39604, 
    -25.16972, -25.94222, -26.71351, -27.48358, -28.25241, -29.01996, 
    -29.78622, -30.55118, -31.31481, -32.0771, -32.83802, -33.59758, 
    -34.35575, -35.11252, -35.86789, -36.62183, -37.37434,
  37.03624, 36.28631, 35.53519, 34.78289, 34.02942, 33.27477, 32.51897, 
    31.76203, 31.00396, 30.24478, 29.48449, 28.72311, 27.96067, 27.19717, 
    26.43264, 25.66709, 24.90054, 24.13302, 23.36455, 22.59513, 21.82482, 
    21.05361, 20.28154, 19.50863, 18.73492, 17.96042, 17.18516, 16.40917, 
    15.63248, 14.85512, 14.07711, 13.2985, 12.5193, 11.73955, 10.95929, 
    10.17854, 9.397336, 8.615713, 7.833705, 7.051345, 6.268667, 5.485706, 
    4.702497, 3.919074, 3.135473, 2.35173, 1.56788, 0.7839577, 0, -0.7839577, 
    -1.56788, -2.35173, -3.135473, -3.919074, -4.702497, -5.485706, 
    -6.268667, -7.051345, -7.833705, -8.615713, -9.397336, -10.17854, 
    -10.95929, -11.73955, -12.5193, -13.2985, -14.07711, -14.85512, 
    -15.63248, -16.40917, -17.18516, -17.96042, -18.73492, -19.50863, 
    -20.28154, -21.05361, -21.82482, -22.59513, -23.36455, -24.13302, 
    -24.90054, -25.66709, -26.43264, -27.19717, -27.96067, -28.72311, 
    -29.48449, -30.24478, -31.00396, -31.76203, -32.51897, -33.27477, 
    -34.02942, -34.78289, -35.53519, -36.28631, -37.03624,
  36.69255, 35.94537, 35.19722, 34.44813, 33.6981, 32.94714, 32.19525, 
    31.44245, 30.68875, 29.93416, 29.17869, 28.42235, 27.66517, 26.90714, 
    26.14829, 25.38863, 24.62818, 23.86696, 23.10497, 22.34225, 21.5788, 
    20.81466, 20.04982, 19.28433, 18.51819, 17.75143, 16.98408, 16.21614, 
    15.44765, 14.67863, 13.90911, 13.1391, 12.36863, 11.59772, 10.82641, 
    10.05472, 9.282667, 8.510284, 7.737598, 6.964634, 6.19142, 5.417983, 
    4.64435, 3.870549, 3.096608, 2.322554, 1.548416, 0.7742223, 0, 
    -0.7742223, -1.548416, -2.322554, -3.096608, -3.870549, -4.64435, 
    -5.417983, -6.19142, -6.964634, -7.737598, -8.510284, -9.282667, 
    -10.05472, -10.82641, -11.59772, -12.36863, -13.1391, -13.90911, 
    -14.67863, -15.44765, -16.21614, -16.98408, -17.75143, -18.51819, 
    -19.28433, -20.04982, -20.81466, -21.5788, -22.34225, -23.10497, 
    -23.86696, -24.62818, -25.38863, -26.14829, -26.90714, -27.66517, 
    -28.42235, -29.17869, -29.93416, -30.68875, -31.44245, -32.19525, 
    -32.94714, -33.6981, -34.44813, -35.19722, -35.94537, -36.69255,
  36.34341, 35.59911, 34.8541, 34.10837, 33.36194, 32.61481, 31.86699, 
    31.11849, 30.36931, 29.61947, 28.86897, 28.11782, 27.36604, 26.61363, 
    25.86061, 25.10699, 24.35277, 23.59798, 22.84263, 22.08672, 21.33028, 
    20.57332, 19.81585, 19.05788, 18.29944, 17.54054, 16.7812, 16.02143, 
    15.26124, 14.50067, 13.73972, 12.97841, 12.21676, 11.45479, 10.69252, 
    9.929964, 9.167146, 8.404083, 7.640796, 6.877304, 6.113627, 5.349786, 
    4.5858, 3.82169, 3.057476, 2.29318, 1.528821, 0.7644209, 0, -0.7644209, 
    -1.528821, -2.29318, -3.057476, -3.82169, -4.5858, -5.349786, -6.113627, 
    -6.877304, -7.640796, -8.404083, -9.167146, -9.929964, -10.69252, 
    -11.45479, -12.21676, -12.97841, -13.73972, -14.50067, -15.26124, 
    -16.02143, -16.7812, -17.54054, -18.29944, -19.05788, -19.81585, 
    -20.57332, -21.33028, -22.08672, -22.84263, -23.59798, -24.35277, 
    -25.10699, -25.86061, -26.61363, -27.36604, -28.11782, -28.86897, 
    -29.61947, -30.36931, -31.11849, -31.86699, -32.61481, -33.36194, 
    -34.10837, -34.8541, -35.59911, -36.34341,
  35.98892, 35.24767, 34.50594, 33.76374, 33.02107, 32.27793, 31.53433, 
    30.79028, 30.04578, 29.30084, 28.55546, 27.80966, 27.06343, 26.31679, 
    25.56974, 24.82229, 24.07445, 23.32623, 22.57764, 21.82868, 21.07937, 
    20.32972, 19.57973, 18.82941, 18.07879, 17.32786, 16.57663, 15.82513, 
    15.07335, 14.32132, 13.56903, 12.81652, 12.06378, 11.31083, 10.55768, 
    9.804344, 9.050837, 8.297169, 7.543353, 6.789403, 6.035332, 5.281153, 
    4.526879, 3.772523, 3.0181, 2.263623, 1.509105, 0.7545591, 0, -0.7545591, 
    -1.509105, -2.263623, -3.0181, -3.772523, -4.526879, -5.281153, 
    -6.035332, -6.789403, -7.543353, -8.297169, -9.050837, -9.804344, 
    -10.55768, -11.31083, -12.06378, -12.81652, -13.56903, -14.32132, 
    -15.07335, -15.82513, -16.57663, -17.32786, -18.07879, -18.82941, 
    -19.57973, -20.32972, -21.07937, -21.82868, -22.57764, -23.32623, 
    -24.07445, -24.82229, -25.56974, -26.31679, -27.06343, -27.80966, 
    -28.55546, -29.30084, -30.04578, -30.79028, -31.53433, -32.27793, 
    -33.02107, -33.76374, -34.50594, -35.24767, -35.98892,
  35.62921, 34.89117, 34.15289, 33.41436, 32.67561, 31.93662, 31.19741, 
    30.45796, 29.7183, 28.97841, 28.23831, 27.49799, 26.75747, 26.01674, 
    25.2758, 24.53467, 23.79335, 23.05183, 22.31014, 21.56826, 20.8262, 
    20.08398, 19.34159, 18.59904, 17.85633, 17.11348, 16.37048, 15.62734, 
    14.88407, 14.14067, 13.39715, 12.65351, 11.90976, 11.16591, 10.42197, 
    9.677926, 8.933801, 8.189597, 7.445321, 6.700978, 5.956575, 5.21212, 
    4.467618, 3.723077, 2.978501, 2.233899, 1.489277, 0.744642, 0, -0.744642, 
    -1.489277, -2.233899, -2.978501, -3.723077, -4.467618, -5.21212, 
    -5.956575, -6.700978, -7.445321, -8.189597, -8.933801, -9.677926, 
    -10.42197, -11.16591, -11.90976, -12.65351, -13.39715, -14.14067, 
    -14.88407, -15.62734, -16.37048, -17.11348, -17.85633, -18.59904, 
    -19.34159, -20.08398, -20.8262, -21.56826, -22.31014, -23.05183, 
    -23.79335, -24.53467, -25.2758, -26.01674, -26.75747, -27.49799, 
    -28.23831, -28.97841, -29.7183, -30.45796, -31.19741, -31.93662, 
    -32.67561, -33.41436, -34.15289, -34.89117, -35.62921,
  35.26439, 34.52972, 33.79504, 33.06036, 32.32569, 31.59101, 30.85634, 
    30.12167, 29.38699, 28.65232, 27.91764, 27.18297, 26.44829, 25.71362, 
    24.97894, 24.24427, 23.50959, 22.77492, 22.04024, 21.30557, 20.57089, 
    19.83622, 19.10155, 18.36687, 17.63219, 16.89752, 16.16285, 15.42817, 
    14.6935, 13.95882, 13.22415, 12.48947, 11.7548, 11.02012, 10.28545, 
    9.550773, 8.816097, 8.081423, 7.346748, 6.612073, 5.877398, 5.142724, 
    4.408049, 3.673374, 2.938699, 2.204024, 1.46935, 0.7346748, 0, 
    -0.7346748, -1.46935, -2.204024, -2.938699, -3.673374, -4.408049, 
    -5.142724, -5.877398, -6.612073, -7.346748, -8.081423, -8.816097, 
    -9.550773, -10.28545, -11.02012, -11.7548, -12.48947, -13.22415, 
    -13.95882, -14.6935, -15.42817, -16.16285, -16.89752, -17.63219, 
    -18.36687, -19.10155, -19.83622, -20.57089, -21.30557, -22.04024, 
    -22.77492, -23.50959, -24.24427, -24.97894, -25.71362, -26.44829, 
    -27.18297, -27.91764, -28.65232, -29.38699, -30.12167, -30.85634, 
    -31.59101, -32.32569, -33.06036, -33.79504, -34.52972, -35.26439 ;

 grid_lont =
  215.3905, 215.3905, 215.3906, 215.3906, 215.3906, 215.3907, 215.3907, 
    215.3907, 215.3908, 215.3908, 215.3908, 215.3909, 215.3909, 215.3909, 
    215.3909, 215.391, 215.391, 215.391, 215.391, 215.3911, 215.3911, 
    215.3911, 215.3911, 215.3911, 215.3912, 215.3912, 215.3912, 215.3912, 
    215.3912, 215.3913, 215.3913, 215.3913, 215.3913, 215.3913, 215.3913, 
    215.3913, 215.3913, 215.3913, 215.3914, 215.3914, 215.3914, 215.3914, 
    215.3914, 215.3914, 215.3914, 215.3914, 215.3914, 215.3914, 215.3914, 
    215.3914, 215.3914, 215.3914, 215.3914, 215.3914, 215.3914, 215.3914, 
    215.3914, 215.3914, 215.3913, 215.3913, 215.3913, 215.3913, 215.3913, 
    215.3913, 215.3913, 215.3913, 215.3913, 215.3912, 215.3912, 215.3912, 
    215.3912, 215.3912, 215.3911, 215.3911, 215.3911, 215.3911, 215.3911, 
    215.391, 215.391, 215.391, 215.391, 215.3909, 215.3909, 215.3909, 
    215.3909, 215.3908, 215.3908, 215.3908, 215.3907, 215.3907, 215.3907, 
    215.3906, 215.3906, 215.3906, 215.3905, 215.3905,
  216.1769, 216.1769, 216.1769, 216.177, 216.177, 216.177, 216.177, 216.1771, 
    216.1771, 216.1771, 216.1772, 216.1772, 216.1772, 216.1772, 216.1773, 
    216.1773, 216.1773, 216.1774, 216.1774, 216.1774, 216.1774, 216.1774, 
    216.1775, 216.1775, 216.1775, 216.1775, 216.1775, 216.1776, 216.1776, 
    216.1776, 216.1776, 216.1776, 216.1776, 216.1776, 216.1777, 216.1777, 
    216.1777, 216.1777, 216.1777, 216.1777, 216.1777, 216.1777, 216.1777, 
    216.1777, 216.1777, 216.1777, 216.1777, 216.1777, 216.1777, 216.1777, 
    216.1777, 216.1777, 216.1777, 216.1777, 216.1777, 216.1777, 216.1777, 
    216.1777, 216.1777, 216.1777, 216.1777, 216.1777, 216.1776, 216.1776, 
    216.1776, 216.1776, 216.1776, 216.1776, 216.1776, 216.1775, 216.1775, 
    216.1775, 216.1775, 216.1775, 216.1774, 216.1774, 216.1774, 216.1774, 
    216.1774, 216.1773, 216.1773, 216.1773, 216.1772, 216.1772, 216.1772, 
    216.1772, 216.1771, 216.1771, 216.1771, 216.177, 216.177, 216.177, 
    216.177, 216.1769, 216.1769, 216.1769,
  216.9704, 216.9704, 216.9704, 216.9704, 216.9705, 216.9705, 216.9705, 
    216.9706, 216.9706, 216.9706, 216.9707, 216.9707, 216.9707, 216.9707, 
    216.9708, 216.9708, 216.9708, 216.9708, 216.9709, 216.9709, 216.9709, 
    216.9709, 216.971, 216.971, 216.971, 216.971, 216.971, 216.9711, 
    216.9711, 216.9711, 216.9711, 216.9711, 216.9711, 216.9711, 216.9712, 
    216.9712, 216.9712, 216.9712, 216.9712, 216.9712, 216.9712, 216.9712, 
    216.9712, 216.9712, 216.9712, 216.9712, 216.9712, 216.9712, 216.9712, 
    216.9712, 216.9712, 216.9712, 216.9712, 216.9712, 216.9712, 216.9712, 
    216.9712, 216.9712, 216.9712, 216.9712, 216.9712, 216.9712, 216.9711, 
    216.9711, 216.9711, 216.9711, 216.9711, 216.9711, 216.9711, 216.971, 
    216.971, 216.971, 216.971, 216.971, 216.9709, 216.9709, 216.9709, 
    216.9709, 216.9708, 216.9708, 216.9708, 216.9708, 216.9707, 216.9707, 
    216.9707, 216.9707, 216.9706, 216.9706, 216.9706, 216.9705, 216.9705, 
    216.9705, 216.9704, 216.9704, 216.9704, 216.9704,
  217.7711, 217.7711, 217.7711, 217.7711, 217.7712, 217.7712, 217.7712, 
    217.7713, 217.7713, 217.7713, 217.7714, 217.7714, 217.7714, 217.7714, 
    217.7715, 217.7715, 217.7715, 217.7715, 217.7716, 217.7716, 217.7716, 
    217.7716, 217.7717, 217.7717, 217.7717, 217.7717, 217.7717, 217.7718, 
    217.7718, 217.7718, 217.7718, 217.7718, 217.7718, 217.7719, 217.7719, 
    217.7719, 217.7719, 217.7719, 217.7719, 217.7719, 217.7719, 217.7719, 
    217.7719, 217.7719, 217.7719, 217.7719, 217.7719, 217.772, 217.772, 
    217.7719, 217.7719, 217.7719, 217.7719, 217.7719, 217.7719, 217.7719, 
    217.7719, 217.7719, 217.7719, 217.7719, 217.7719, 217.7719, 217.7719, 
    217.7718, 217.7718, 217.7718, 217.7718, 217.7718, 217.7718, 217.7717, 
    217.7717, 217.7717, 217.7717, 217.7717, 217.7716, 217.7716, 217.7716, 
    217.7716, 217.7715, 217.7715, 217.7715, 217.7715, 217.7714, 217.7714, 
    217.7714, 217.7714, 217.7713, 217.7713, 217.7713, 217.7712, 217.7712, 
    217.7712, 217.7711, 217.7711, 217.7711, 217.7711,
  218.579, 218.5791, 218.5791, 218.5791, 218.5791, 218.5792, 218.5792, 
    218.5792, 218.5793, 218.5793, 218.5793, 218.5793, 218.5794, 218.5794, 
    218.5794, 218.5795, 218.5795, 218.5795, 218.5795, 218.5796, 218.5796, 
    218.5796, 218.5796, 218.5797, 218.5797, 218.5797, 218.5797, 218.5797, 
    218.5797, 218.5798, 218.5798, 218.5798, 218.5798, 218.5798, 218.5798, 
    218.5798, 218.5798, 218.5799, 218.5799, 218.5799, 218.5799, 218.5799, 
    218.5799, 218.5799, 218.5799, 218.5799, 218.5799, 218.5799, 218.5799, 
    218.5799, 218.5799, 218.5799, 218.5799, 218.5799, 218.5799, 218.5799, 
    218.5799, 218.5799, 218.5799, 218.5798, 218.5798, 218.5798, 218.5798, 
    218.5798, 218.5798, 218.5798, 218.5798, 218.5797, 218.5797, 218.5797, 
    218.5797, 218.5797, 218.5797, 218.5796, 218.5796, 218.5796, 218.5796, 
    218.5795, 218.5795, 218.5795, 218.5795, 218.5794, 218.5794, 218.5794, 
    218.5793, 218.5793, 218.5793, 218.5793, 218.5792, 218.5792, 218.5792, 
    218.5791, 218.5791, 218.5791, 218.5791, 218.579,
  219.3943, 219.3943, 219.3943, 219.3944, 219.3944, 219.3944, 219.3945, 
    219.3945, 219.3945, 219.3946, 219.3946, 219.3946, 219.3946, 219.3947, 
    219.3947, 219.3947, 219.3947, 219.3948, 219.3948, 219.3948, 219.3949, 
    219.3949, 219.3949, 219.3949, 219.3949, 219.395, 219.395, 219.395, 
    219.395, 219.395, 219.3951, 219.3951, 219.3951, 219.3951, 219.3951, 
    219.3951, 219.3951, 219.3951, 219.3951, 219.3952, 219.3952, 219.3952, 
    219.3952, 219.3952, 219.3952, 219.3952, 219.3952, 219.3952, 219.3952, 
    219.3952, 219.3952, 219.3952, 219.3952, 219.3952, 219.3952, 219.3952, 
    219.3952, 219.3951, 219.3951, 219.3951, 219.3951, 219.3951, 219.3951, 
    219.3951, 219.3951, 219.3951, 219.395, 219.395, 219.395, 219.395, 
    219.395, 219.3949, 219.3949, 219.3949, 219.3949, 219.3949, 219.3948, 
    219.3948, 219.3948, 219.3947, 219.3947, 219.3947, 219.3947, 219.3946, 
    219.3946, 219.3946, 219.3946, 219.3945, 219.3945, 219.3945, 219.3944, 
    219.3944, 219.3944, 219.3943, 219.3943, 219.3943,
  220.2169, 220.2169, 220.2169, 220.217, 220.217, 220.217, 220.2171, 
    220.2171, 220.2171, 220.2172, 220.2172, 220.2172, 220.2172, 220.2173, 
    220.2173, 220.2173, 220.2173, 220.2174, 220.2174, 220.2174, 220.2175, 
    220.2175, 220.2175, 220.2175, 220.2175, 220.2176, 220.2176, 220.2176, 
    220.2176, 220.2176, 220.2177, 220.2177, 220.2177, 220.2177, 220.2177, 
    220.2177, 220.2177, 220.2177, 220.2177, 220.2178, 220.2178, 220.2178, 
    220.2178, 220.2178, 220.2178, 220.2178, 220.2178, 220.2178, 220.2178, 
    220.2178, 220.2178, 220.2178, 220.2178, 220.2178, 220.2178, 220.2178, 
    220.2178, 220.2177, 220.2177, 220.2177, 220.2177, 220.2177, 220.2177, 
    220.2177, 220.2177, 220.2177, 220.2176, 220.2176, 220.2176, 220.2176, 
    220.2176, 220.2175, 220.2175, 220.2175, 220.2175, 220.2175, 220.2174, 
    220.2174, 220.2174, 220.2173, 220.2173, 220.2173, 220.2173, 220.2172, 
    220.2172, 220.2172, 220.2172, 220.2171, 220.2171, 220.2171, 220.217, 
    220.217, 220.217, 220.2169, 220.2169, 220.2169,
  221.0469, 221.0469, 221.0469, 221.047, 221.047, 221.047, 221.047, 221.0471, 
    221.0471, 221.0471, 221.0471, 221.0472, 221.0472, 221.0472, 221.0473, 
    221.0473, 221.0473, 221.0473, 221.0474, 221.0474, 221.0474, 221.0474, 
    221.0475, 221.0475, 221.0475, 221.0475, 221.0475, 221.0476, 221.0476, 
    221.0476, 221.0476, 221.0476, 221.0477, 221.0477, 221.0477, 221.0477, 
    221.0477, 221.0477, 221.0477, 221.0477, 221.0477, 221.0477, 221.0477, 
    221.0477, 221.0478, 221.0478, 221.0478, 221.0478, 221.0478, 221.0478, 
    221.0478, 221.0478, 221.0477, 221.0477, 221.0477, 221.0477, 221.0477, 
    221.0477, 221.0477, 221.0477, 221.0477, 221.0477, 221.0477, 221.0477, 
    221.0476, 221.0476, 221.0476, 221.0476, 221.0476, 221.0475, 221.0475, 
    221.0475, 221.0475, 221.0475, 221.0474, 221.0474, 221.0474, 221.0474, 
    221.0473, 221.0473, 221.0473, 221.0473, 221.0472, 221.0472, 221.0472, 
    221.0471, 221.0471, 221.0471, 221.0471, 221.047, 221.047, 221.047, 
    221.047, 221.0469, 221.0469, 221.0469,
  221.8842, 221.8842, 221.8843, 221.8843, 221.8843, 221.8844, 221.8844, 
    221.8844, 221.8845, 221.8845, 221.8845, 221.8845, 221.8846, 221.8846, 
    221.8846, 221.8846, 221.8847, 221.8847, 221.8847, 221.8848, 221.8848, 
    221.8848, 221.8848, 221.8848, 221.8849, 221.8849, 221.8849, 221.8849, 
    221.8849, 221.885, 221.885, 221.885, 221.885, 221.885, 221.885, 221.885, 
    221.8851, 221.8851, 221.8851, 221.8851, 221.8851, 221.8851, 221.8851, 
    221.8851, 221.8851, 221.8851, 221.8851, 221.8851, 221.8851, 221.8851, 
    221.8851, 221.8851, 221.8851, 221.8851, 221.8851, 221.8851, 221.8851, 
    221.8851, 221.8851, 221.8851, 221.885, 221.885, 221.885, 221.885, 
    221.885, 221.885, 221.885, 221.8849, 221.8849, 221.8849, 221.8849, 
    221.8849, 221.8848, 221.8848, 221.8848, 221.8848, 221.8848, 221.8847, 
    221.8847, 221.8847, 221.8846, 221.8846, 221.8846, 221.8846, 221.8845, 
    221.8845, 221.8845, 221.8845, 221.8844, 221.8844, 221.8844, 221.8843, 
    221.8843, 221.8843, 221.8842, 221.8842,
  222.729, 222.729, 222.729, 222.7291, 222.7291, 222.7291, 222.7292, 
    222.7292, 222.7292, 222.7292, 222.7293, 222.7293, 222.7293, 222.7294, 
    222.7294, 222.7294, 222.7294, 222.7295, 222.7295, 222.7295, 222.7295, 
    222.7296, 222.7296, 222.7296, 222.7296, 222.7296, 222.7297, 222.7297, 
    222.7297, 222.7297, 222.7297, 222.7298, 222.7298, 222.7298, 222.7298, 
    222.7298, 222.7298, 222.7298, 222.7298, 222.7299, 222.7299, 222.7299, 
    222.7299, 222.7299, 222.7299, 222.7299, 222.7299, 222.7299, 222.7299, 
    222.7299, 222.7299, 222.7299, 222.7299, 222.7299, 222.7299, 222.7299, 
    222.7299, 222.7298, 222.7298, 222.7298, 222.7298, 222.7298, 222.7298, 
    222.7298, 222.7298, 222.7297, 222.7297, 222.7297, 222.7297, 222.7297, 
    222.7296, 222.7296, 222.7296, 222.7296, 222.7296, 222.7295, 222.7295, 
    222.7295, 222.7295, 222.7294, 222.7294, 222.7294, 222.7294, 222.7293, 
    222.7293, 222.7293, 222.7292, 222.7292, 222.7292, 222.7292, 222.7291, 
    222.7291, 222.7291, 222.729, 222.729, 222.729,
  223.5812, 223.5812, 223.5812, 223.5813, 223.5813, 223.5813, 223.5813, 
    223.5814, 223.5814, 223.5814, 223.5815, 223.5815, 223.5815, 223.5815, 
    223.5816, 223.5816, 223.5816, 223.5816, 223.5817, 223.5817, 223.5817, 
    223.5817, 223.5818, 223.5818, 223.5818, 223.5818, 223.5818, 223.5819, 
    223.5819, 223.5819, 223.5819, 223.5819, 223.582, 223.582, 223.582, 
    223.582, 223.582, 223.582, 223.582, 223.582, 223.582, 223.582, 223.582, 
    223.5821, 223.5821, 223.5821, 223.5821, 223.5821, 223.5821, 223.5821, 
    223.5821, 223.5821, 223.5821, 223.582, 223.582, 223.582, 223.582, 
    223.582, 223.582, 223.582, 223.582, 223.582, 223.582, 223.582, 223.5819, 
    223.5819, 223.5819, 223.5819, 223.5819, 223.5818, 223.5818, 223.5818, 
    223.5818, 223.5818, 223.5817, 223.5817, 223.5817, 223.5817, 223.5816, 
    223.5816, 223.5816, 223.5816, 223.5815, 223.5815, 223.5815, 223.5815, 
    223.5814, 223.5814, 223.5814, 223.5813, 223.5813, 223.5813, 223.5813, 
    223.5812, 223.5812, 223.5812,
  224.4408, 224.4408, 224.4408, 224.4408, 224.4409, 224.4409, 224.4409, 
    224.4409, 224.441, 224.441, 224.441, 224.4411, 224.4411, 224.4411, 
    224.4411, 224.4412, 224.4412, 224.4412, 224.4413, 224.4413, 224.4413, 
    224.4413, 224.4413, 224.4414, 224.4414, 224.4414, 224.4414, 224.4415, 
    224.4415, 224.4415, 224.4415, 224.4415, 224.4415, 224.4416, 224.4416, 
    224.4416, 224.4416, 224.4416, 224.4416, 224.4416, 224.4416, 224.4416, 
    224.4416, 224.4417, 224.4417, 224.4417, 224.4417, 224.4417, 224.4417, 
    224.4417, 224.4417, 224.4417, 224.4417, 224.4416, 224.4416, 224.4416, 
    224.4416, 224.4416, 224.4416, 224.4416, 224.4416, 224.4416, 224.4416, 
    224.4415, 224.4415, 224.4415, 224.4415, 224.4415, 224.4415, 224.4414, 
    224.4414, 224.4414, 224.4414, 224.4413, 224.4413, 224.4413, 224.4413, 
    224.4413, 224.4412, 224.4412, 224.4412, 224.4411, 224.4411, 224.4411, 
    224.4411, 224.441, 224.441, 224.441, 224.4409, 224.4409, 224.4409, 
    224.4409, 224.4408, 224.4408, 224.4408, 224.4408,
  225.3077, 225.3078, 225.3078, 225.3078, 225.3079, 225.3079, 225.3079, 
    225.308, 225.308, 225.308, 225.308, 225.3081, 225.3081, 225.3081, 
    225.3082, 225.3082, 225.3082, 225.3082, 225.3082, 225.3083, 225.3083, 
    225.3083, 225.3083, 225.3084, 225.3084, 225.3084, 225.3084, 225.3084, 
    225.3085, 225.3085, 225.3085, 225.3085, 225.3085, 225.3085, 225.3086, 
    225.3086, 225.3086, 225.3086, 225.3086, 225.3086, 225.3086, 225.3086, 
    225.3086, 225.3086, 225.3086, 225.3087, 225.3087, 225.3087, 225.3087, 
    225.3087, 225.3087, 225.3086, 225.3086, 225.3086, 225.3086, 225.3086, 
    225.3086, 225.3086, 225.3086, 225.3086, 225.3086, 225.3086, 225.3085, 
    225.3085, 225.3085, 225.3085, 225.3085, 225.3085, 225.3084, 225.3084, 
    225.3084, 225.3084, 225.3084, 225.3083, 225.3083, 225.3083, 225.3083, 
    225.3082, 225.3082, 225.3082, 225.3082, 225.3082, 225.3081, 225.3081, 
    225.3081, 225.308, 225.308, 225.308, 225.308, 225.3079, 225.3079, 
    225.3079, 225.3078, 225.3078, 225.3078, 225.3077,
  226.1821, 226.1822, 226.1822, 226.1822, 226.1823, 226.1823, 226.1823, 
    226.1823, 226.1824, 226.1824, 226.1824, 226.1824, 226.1825, 226.1825, 
    226.1825, 226.1826, 226.1826, 226.1826, 226.1826, 226.1827, 226.1827, 
    226.1827, 226.1827, 226.1828, 226.1828, 226.1828, 226.1828, 226.1828, 
    226.1828, 226.1829, 226.1829, 226.1829, 226.1829, 226.1829, 226.1829, 
    226.183, 226.183, 226.183, 226.183, 226.183, 226.183, 226.183, 226.183, 
    226.183, 226.183, 226.183, 226.183, 226.183, 226.183, 226.183, 226.183, 
    226.183, 226.183, 226.183, 226.183, 226.183, 226.183, 226.183, 226.183, 
    226.183, 226.183, 226.1829, 226.1829, 226.1829, 226.1829, 226.1829, 
    226.1829, 226.1828, 226.1828, 226.1828, 226.1828, 226.1828, 226.1828, 
    226.1827, 226.1827, 226.1827, 226.1827, 226.1826, 226.1826, 226.1826, 
    226.1826, 226.1825, 226.1825, 226.1825, 226.1824, 226.1824, 226.1824, 
    226.1824, 226.1823, 226.1823, 226.1823, 226.1823, 226.1822, 226.1822, 
    226.1822, 226.1821,
  227.0639, 227.0639, 227.0639, 227.064, 227.064, 227.064, 227.0641, 
    227.0641, 227.0641, 227.0641, 227.0642, 227.0642, 227.0642, 227.0642, 
    227.0643, 227.0643, 227.0643, 227.0643, 227.0644, 227.0644, 227.0644, 
    227.0645, 227.0645, 227.0645, 227.0645, 227.0645, 227.0646, 227.0646, 
    227.0646, 227.0646, 227.0646, 227.0646, 227.0647, 227.0647, 227.0647, 
    227.0647, 227.0647, 227.0647, 227.0647, 227.0647, 227.0647, 227.0648, 
    227.0648, 227.0648, 227.0648, 227.0648, 227.0648, 227.0648, 227.0648, 
    227.0648, 227.0648, 227.0648, 227.0648, 227.0648, 227.0648, 227.0647, 
    227.0647, 227.0647, 227.0647, 227.0647, 227.0647, 227.0647, 227.0647, 
    227.0647, 227.0646, 227.0646, 227.0646, 227.0646, 227.0646, 227.0646, 
    227.0645, 227.0645, 227.0645, 227.0645, 227.0645, 227.0644, 227.0644, 
    227.0644, 227.0643, 227.0643, 227.0643, 227.0643, 227.0642, 227.0642, 
    227.0642, 227.0642, 227.0641, 227.0641, 227.0641, 227.0641, 227.064, 
    227.064, 227.064, 227.0639, 227.0639, 227.0639,
  227.953, 227.953, 227.953, 227.953, 227.9531, 227.9531, 227.9531, 227.9532, 
    227.9532, 227.9532, 227.9532, 227.9533, 227.9533, 227.9533, 227.9533, 
    227.9534, 227.9534, 227.9534, 227.9534, 227.9535, 227.9535, 227.9535, 
    227.9535, 227.9536, 227.9536, 227.9536, 227.9536, 227.9536, 227.9537, 
    227.9537, 227.9537, 227.9537, 227.9537, 227.9537, 227.9538, 227.9538, 
    227.9538, 227.9538, 227.9538, 227.9538, 227.9538, 227.9538, 227.9538, 
    227.9538, 227.9538, 227.9538, 227.9538, 227.9538, 227.9538, 227.9538, 
    227.9538, 227.9538, 227.9538, 227.9538, 227.9538, 227.9538, 227.9538, 
    227.9538, 227.9538, 227.9538, 227.9538, 227.9538, 227.9537, 227.9537, 
    227.9537, 227.9537, 227.9537, 227.9537, 227.9536, 227.9536, 227.9536, 
    227.9536, 227.9536, 227.9535, 227.9535, 227.9535, 227.9535, 227.9534, 
    227.9534, 227.9534, 227.9534, 227.9533, 227.9533, 227.9533, 227.9533, 
    227.9532, 227.9532, 227.9532, 227.9532, 227.9531, 227.9531, 227.9531, 
    227.953, 227.953, 227.953, 227.953,
  228.8493, 228.8493, 228.8494, 228.8494, 228.8494, 228.8494, 228.8495, 
    228.8495, 228.8495, 228.8496, 228.8496, 228.8496, 228.8496, 228.8497, 
    228.8497, 228.8497, 228.8497, 228.8498, 228.8498, 228.8498, 228.8498, 
    228.8499, 228.8499, 228.8499, 228.8499, 228.8499, 228.85, 228.85, 228.85, 
    228.85, 228.85, 228.8501, 228.8501, 228.8501, 228.8501, 228.8501, 
    228.8501, 228.8501, 228.8501, 228.8502, 228.8502, 228.8502, 228.8502, 
    228.8502, 228.8502, 228.8502, 228.8502, 228.8502, 228.8502, 228.8502, 
    228.8502, 228.8502, 228.8502, 228.8502, 228.8502, 228.8502, 228.8502, 
    228.8501, 228.8501, 228.8501, 228.8501, 228.8501, 228.8501, 228.8501, 
    228.8501, 228.85, 228.85, 228.85, 228.85, 228.85, 228.8499, 228.8499, 
    228.8499, 228.8499, 228.8499, 228.8498, 228.8498, 228.8498, 228.8498, 
    228.8497, 228.8497, 228.8497, 228.8497, 228.8496, 228.8496, 228.8496, 
    228.8496, 228.8495, 228.8495, 228.8495, 228.8494, 228.8494, 228.8494, 
    228.8494, 228.8493, 228.8493,
  229.7529, 229.7529, 229.7529, 229.753, 229.753, 229.753, 229.7531, 
    229.7531, 229.7531, 229.7531, 229.7532, 229.7532, 229.7532, 229.7532, 
    229.7533, 229.7533, 229.7533, 229.7533, 229.7534, 229.7534, 229.7534, 
    229.7534, 229.7534, 229.7535, 229.7535, 229.7535, 229.7535, 229.7536, 
    229.7536, 229.7536, 229.7536, 229.7536, 229.7536, 229.7537, 229.7537, 
    229.7537, 229.7537, 229.7537, 229.7537, 229.7537, 229.7537, 229.7537, 
    229.7538, 229.7538, 229.7538, 229.7538, 229.7538, 229.7538, 229.7538, 
    229.7538, 229.7538, 229.7538, 229.7538, 229.7538, 229.7537, 229.7537, 
    229.7537, 229.7537, 229.7537, 229.7537, 229.7537, 229.7537, 229.7537, 
    229.7536, 229.7536, 229.7536, 229.7536, 229.7536, 229.7536, 229.7535, 
    229.7535, 229.7535, 229.7535, 229.7534, 229.7534, 229.7534, 229.7534, 
    229.7534, 229.7533, 229.7533, 229.7533, 229.7533, 229.7532, 229.7532, 
    229.7532, 229.7532, 229.7531, 229.7531, 229.7531, 229.7531, 229.753, 
    229.753, 229.753, 229.7529, 229.7529, 229.7529,
  230.6636, 230.6637, 230.6637, 230.6637, 230.6637, 230.6638, 230.6638, 
    230.6638, 230.6638, 230.6639, 230.6639, 230.6639, 230.6639, 230.664, 
    230.664, 230.664, 230.664, 230.6641, 230.6641, 230.6641, 230.6641, 
    230.6642, 230.6642, 230.6642, 230.6642, 230.6642, 230.6643, 230.6643, 
    230.6643, 230.6643, 230.6643, 230.6644, 230.6644, 230.6644, 230.6644, 
    230.6644, 230.6644, 230.6644, 230.6644, 230.6644, 230.6645, 230.6645, 
    230.6645, 230.6645, 230.6645, 230.6645, 230.6645, 230.6645, 230.6645, 
    230.6645, 230.6645, 230.6645, 230.6645, 230.6645, 230.6645, 230.6645, 
    230.6644, 230.6644, 230.6644, 230.6644, 230.6644, 230.6644, 230.6644, 
    230.6644, 230.6644, 230.6643, 230.6643, 230.6643, 230.6643, 230.6643, 
    230.6642, 230.6642, 230.6642, 230.6642, 230.6642, 230.6641, 230.6641, 
    230.6641, 230.6641, 230.664, 230.664, 230.664, 230.664, 230.6639, 
    230.6639, 230.6639, 230.6639, 230.6638, 230.6638, 230.6638, 230.6638, 
    230.6637, 230.6637, 230.6637, 230.6637, 230.6636,
  231.5814, 231.5815, 231.5815, 231.5815, 231.5815, 231.5816, 231.5816, 
    231.5816, 231.5816, 231.5817, 231.5817, 231.5817, 231.5818, 231.5818, 
    231.5818, 231.5818, 231.5818, 231.5819, 231.5819, 231.5819, 231.5819, 
    231.582, 231.582, 231.582, 231.582, 231.582, 231.5821, 231.5821, 
    231.5821, 231.5821, 231.5821, 231.5822, 231.5822, 231.5822, 231.5822, 
    231.5822, 231.5822, 231.5822, 231.5822, 231.5823, 231.5823, 231.5823, 
    231.5823, 231.5823, 231.5823, 231.5823, 231.5823, 231.5823, 231.5823, 
    231.5823, 231.5823, 231.5823, 231.5823, 231.5823, 231.5823, 231.5823, 
    231.5823, 231.5822, 231.5822, 231.5822, 231.5822, 231.5822, 231.5822, 
    231.5822, 231.5822, 231.5821, 231.5821, 231.5821, 231.5821, 231.5821, 
    231.582, 231.582, 231.582, 231.582, 231.582, 231.5819, 231.5819, 
    231.5819, 231.5819, 231.5818, 231.5818, 231.5818, 231.5818, 231.5818, 
    231.5817, 231.5817, 231.5817, 231.5816, 231.5816, 231.5816, 231.5816, 
    231.5815, 231.5815, 231.5815, 231.5815, 231.5814,
  232.5062, 232.5063, 232.5063, 232.5063, 232.5063, 232.5064, 232.5064, 
    232.5064, 232.5065, 232.5065, 232.5065, 232.5065, 232.5065, 232.5066, 
    232.5066, 232.5066, 232.5067, 232.5067, 232.5067, 232.5067, 232.5067, 
    232.5068, 232.5068, 232.5068, 232.5068, 232.5069, 232.5069, 232.5069, 
    232.5069, 232.5069, 232.5069, 232.507, 232.507, 232.507, 232.507, 
    232.507, 232.507, 232.507, 232.507, 232.507, 232.5071, 232.5071, 
    232.5071, 232.5071, 232.5071, 232.5071, 232.5071, 232.5071, 232.5071, 
    232.5071, 232.5071, 232.5071, 232.5071, 232.5071, 232.5071, 232.5071, 
    232.507, 232.507, 232.507, 232.507, 232.507, 232.507, 232.507, 232.507, 
    232.507, 232.5069, 232.5069, 232.5069, 232.5069, 232.5069, 232.5069, 
    232.5068, 232.5068, 232.5068, 232.5068, 232.5067, 232.5067, 232.5067, 
    232.5067, 232.5067, 232.5066, 232.5066, 232.5066, 232.5065, 232.5065, 
    232.5065, 232.5065, 232.5065, 232.5064, 232.5064, 232.5064, 232.5063, 
    232.5063, 232.5063, 232.5063, 232.5062,
  233.4379, 233.438, 233.438, 233.438, 233.438, 233.4381, 233.4381, 233.4381, 
    233.4381, 233.4382, 233.4382, 233.4382, 233.4382, 233.4383, 233.4383, 
    233.4383, 233.4383, 233.4384, 233.4384, 233.4384, 233.4384, 233.4385, 
    233.4385, 233.4385, 233.4385, 233.4385, 233.4386, 233.4386, 233.4386, 
    233.4386, 233.4386, 233.4386, 233.4387, 233.4387, 233.4387, 233.4387, 
    233.4387, 233.4387, 233.4387, 233.4387, 233.4388, 233.4388, 233.4388, 
    233.4388, 233.4388, 233.4388, 233.4388, 233.4388, 233.4388, 233.4388, 
    233.4388, 233.4388, 233.4388, 233.4388, 233.4388, 233.4388, 233.4387, 
    233.4387, 233.4387, 233.4387, 233.4387, 233.4387, 233.4387, 233.4387, 
    233.4386, 233.4386, 233.4386, 233.4386, 233.4386, 233.4386, 233.4385, 
    233.4385, 233.4385, 233.4385, 233.4385, 233.4384, 233.4384, 233.4384, 
    233.4384, 233.4383, 233.4383, 233.4383, 233.4383, 233.4382, 233.4382, 
    233.4382, 233.4382, 233.4381, 233.4381, 233.4381, 233.4381, 233.438, 
    233.438, 233.438, 233.438, 233.4379,
  234.3764, 234.3764, 234.3765, 234.3765, 234.3765, 234.3765, 234.3766, 
    234.3766, 234.3766, 234.3766, 234.3767, 234.3767, 234.3767, 234.3767, 
    234.3768, 234.3768, 234.3768, 234.3768, 234.3769, 234.3769, 234.3769, 
    234.3769, 234.377, 234.377, 234.377, 234.377, 234.377, 234.377, 234.3771, 
    234.3771, 234.3771, 234.3771, 234.3771, 234.3771, 234.3772, 234.3772, 
    234.3772, 234.3772, 234.3772, 234.3772, 234.3772, 234.3772, 234.3772, 
    234.3772, 234.3772, 234.3772, 234.3772, 234.3772, 234.3772, 234.3772, 
    234.3772, 234.3772, 234.3772, 234.3772, 234.3772, 234.3772, 234.3772, 
    234.3772, 234.3772, 234.3772, 234.3772, 234.3772, 234.3771, 234.3771, 
    234.3771, 234.3771, 234.3771, 234.3771, 234.377, 234.377, 234.377, 
    234.377, 234.377, 234.377, 234.3769, 234.3769, 234.3769, 234.3769, 
    234.3768, 234.3768, 234.3768, 234.3768, 234.3767, 234.3767, 234.3767, 
    234.3767, 234.3766, 234.3766, 234.3766, 234.3766, 234.3765, 234.3765, 
    234.3765, 234.3765, 234.3764, 234.3764,
  235.3216, 235.3216, 235.3216, 235.3216, 235.3217, 235.3217, 235.3217, 
    235.3217, 235.3217, 235.3218, 235.3218, 235.3218, 235.3219, 235.3219, 
    235.3219, 235.3219, 235.3219, 235.322, 235.322, 235.322, 235.322, 
    235.3221, 235.3221, 235.3221, 235.3221, 235.3221, 235.3222, 235.3222, 
    235.3222, 235.3222, 235.3222, 235.3222, 235.3223, 235.3223, 235.3223, 
    235.3223, 235.3223, 235.3223, 235.3223, 235.3223, 235.3223, 235.3223, 
    235.3223, 235.3224, 235.3224, 235.3224, 235.3224, 235.3224, 235.3224, 
    235.3224, 235.3224, 235.3224, 235.3224, 235.3223, 235.3223, 235.3223, 
    235.3223, 235.3223, 235.3223, 235.3223, 235.3223, 235.3223, 235.3223, 
    235.3223, 235.3222, 235.3222, 235.3222, 235.3222, 235.3222, 235.3222, 
    235.3221, 235.3221, 235.3221, 235.3221, 235.3221, 235.322, 235.322, 
    235.322, 235.322, 235.3219, 235.3219, 235.3219, 235.3219, 235.3219, 
    235.3218, 235.3218, 235.3218, 235.3217, 235.3217, 235.3217, 235.3217, 
    235.3217, 235.3216, 235.3216, 235.3216, 235.3216,
  236.2732, 236.2732, 236.2733, 236.2733, 236.2733, 236.2733, 236.2734, 
    236.2734, 236.2734, 236.2734, 236.2735, 236.2735, 236.2735, 236.2735, 
    236.2736, 236.2736, 236.2736, 236.2736, 236.2736, 236.2737, 236.2737, 
    236.2737, 236.2737, 236.2737, 236.2738, 236.2738, 236.2738, 236.2738, 
    236.2738, 236.2738, 236.2739, 236.2739, 236.2739, 236.2739, 236.2739, 
    236.2739, 236.2739, 236.274, 236.274, 236.274, 236.274, 236.274, 236.274, 
    236.274, 236.274, 236.274, 236.274, 236.274, 236.274, 236.274, 236.274, 
    236.274, 236.274, 236.274, 236.274, 236.274, 236.274, 236.274, 236.274, 
    236.2739, 236.2739, 236.2739, 236.2739, 236.2739, 236.2739, 236.2739, 
    236.2738, 236.2738, 236.2738, 236.2738, 236.2738, 236.2738, 236.2737, 
    236.2737, 236.2737, 236.2737, 236.2737, 236.2736, 236.2736, 236.2736, 
    236.2736, 236.2736, 236.2735, 236.2735, 236.2735, 236.2735, 236.2734, 
    236.2734, 236.2734, 236.2734, 236.2733, 236.2733, 236.2733, 236.2733, 
    236.2732, 236.2732,
  237.2313, 237.2313, 237.2313, 237.2313, 237.2314, 237.2314, 237.2314, 
    237.2314, 237.2314, 237.2315, 237.2315, 237.2315, 237.2315, 237.2316, 
    237.2316, 237.2316, 237.2316, 237.2316, 237.2317, 237.2317, 237.2317, 
    237.2317, 237.2318, 237.2318, 237.2318, 237.2318, 237.2318, 237.2318, 
    237.2319, 237.2319, 237.2319, 237.2319, 237.2319, 237.2319, 237.2319, 
    237.232, 237.232, 237.232, 237.232, 237.232, 237.232, 237.232, 237.232, 
    237.232, 237.232, 237.232, 237.232, 237.232, 237.232, 237.232, 237.232, 
    237.232, 237.232, 237.232, 237.232, 237.232, 237.232, 237.232, 237.232, 
    237.232, 237.232, 237.2319, 237.2319, 237.2319, 237.2319, 237.2319, 
    237.2319, 237.2319, 237.2318, 237.2318, 237.2318, 237.2318, 237.2318, 
    237.2318, 237.2317, 237.2317, 237.2317, 237.2317, 237.2316, 237.2316, 
    237.2316, 237.2316, 237.2316, 237.2315, 237.2315, 237.2315, 237.2315, 
    237.2314, 237.2314, 237.2314, 237.2314, 237.2314, 237.2313, 237.2313, 
    237.2313, 237.2313,
  238.1955, 238.1955, 238.1956, 238.1956, 238.1956, 238.1956, 238.1957, 
    238.1957, 238.1957, 238.1957, 238.1957, 238.1958, 238.1958, 238.1958, 
    238.1958, 238.1959, 238.1959, 238.1959, 238.1959, 238.1959, 238.196, 
    238.196, 238.196, 238.196, 238.196, 238.196, 238.1961, 238.1961, 
    238.1961, 238.1961, 238.1961, 238.1962, 238.1962, 238.1962, 238.1962, 
    238.1962, 238.1962, 238.1962, 238.1962, 238.1962, 238.1962, 238.1962, 
    238.1963, 238.1963, 238.1963, 238.1963, 238.1963, 238.1963, 238.1963, 
    238.1963, 238.1963, 238.1963, 238.1963, 238.1963, 238.1962, 238.1962, 
    238.1962, 238.1962, 238.1962, 238.1962, 238.1962, 238.1962, 238.1962, 
    238.1962, 238.1962, 238.1961, 238.1961, 238.1961, 238.1961, 238.1961, 
    238.196, 238.196, 238.196, 238.196, 238.196, 238.196, 238.1959, 238.1959, 
    238.1959, 238.1959, 238.1959, 238.1958, 238.1958, 238.1958, 238.1958, 
    238.1957, 238.1957, 238.1957, 238.1957, 238.1957, 238.1956, 238.1956, 
    238.1956, 238.1956, 238.1955, 238.1955,
  239.1658, 239.1658, 239.1659, 239.1659, 239.1659, 239.1659, 239.166, 
    239.166, 239.166, 239.166, 239.166, 239.1661, 239.1661, 239.1661, 
    239.1661, 239.1662, 239.1662, 239.1662, 239.1662, 239.1662, 239.1662, 
    239.1663, 239.1663, 239.1663, 239.1663, 239.1663, 239.1664, 239.1664, 
    239.1664, 239.1664, 239.1664, 239.1664, 239.1664, 239.1665, 239.1665, 
    239.1665, 239.1665, 239.1665, 239.1665, 239.1665, 239.1665, 239.1665, 
    239.1665, 239.1665, 239.1665, 239.1665, 239.1665, 239.1665, 239.1665, 
    239.1665, 239.1665, 239.1665, 239.1665, 239.1665, 239.1665, 239.1665, 
    239.1665, 239.1665, 239.1665, 239.1665, 239.1665, 239.1665, 239.1665, 
    239.1664, 239.1664, 239.1664, 239.1664, 239.1664, 239.1664, 239.1664, 
    239.1663, 239.1663, 239.1663, 239.1663, 239.1663, 239.1662, 239.1662, 
    239.1662, 239.1662, 239.1662, 239.1662, 239.1661, 239.1661, 239.1661, 
    239.1661, 239.166, 239.166, 239.166, 239.166, 239.166, 239.1659, 
    239.1659, 239.1659, 239.1659, 239.1658, 239.1658,
  240.142, 240.142, 240.142, 240.1421, 240.1421, 240.1421, 240.1421, 
    240.1422, 240.1422, 240.1422, 240.1422, 240.1422, 240.1423, 240.1423, 
    240.1423, 240.1423, 240.1423, 240.1423, 240.1424, 240.1424, 240.1424, 
    240.1424, 240.1424, 240.1425, 240.1425, 240.1425, 240.1425, 240.1425, 
    240.1425, 240.1426, 240.1426, 240.1426, 240.1426, 240.1426, 240.1426, 
    240.1426, 240.1426, 240.1427, 240.1427, 240.1427, 240.1427, 240.1427, 
    240.1427, 240.1427, 240.1427, 240.1427, 240.1427, 240.1427, 240.1427, 
    240.1427, 240.1427, 240.1427, 240.1427, 240.1427, 240.1427, 240.1427, 
    240.1427, 240.1427, 240.1427, 240.1426, 240.1426, 240.1426, 240.1426, 
    240.1426, 240.1426, 240.1426, 240.1426, 240.1425, 240.1425, 240.1425, 
    240.1425, 240.1425, 240.1425, 240.1424, 240.1424, 240.1424, 240.1424, 
    240.1424, 240.1423, 240.1423, 240.1423, 240.1423, 240.1423, 240.1423, 
    240.1422, 240.1422, 240.1422, 240.1422, 240.1422, 240.1421, 240.1421, 
    240.1421, 240.1421, 240.142, 240.142, 240.142,
  241.1239, 241.1239, 241.1239, 241.1239, 241.1239, 241.1239, 241.124, 
    241.124, 241.124, 241.124, 241.1241, 241.1241, 241.1241, 241.1241, 
    241.1241, 241.1241, 241.1242, 241.1242, 241.1242, 241.1242, 241.1242, 
    241.1243, 241.1243, 241.1243, 241.1243, 241.1243, 241.1243, 241.1244, 
    241.1244, 241.1244, 241.1244, 241.1244, 241.1244, 241.1244, 241.1245, 
    241.1245, 241.1245, 241.1245, 241.1245, 241.1245, 241.1245, 241.1245, 
    241.1245, 241.1245, 241.1245, 241.1245, 241.1245, 241.1245, 241.1245, 
    241.1245, 241.1245, 241.1245, 241.1245, 241.1245, 241.1245, 241.1245, 
    241.1245, 241.1245, 241.1245, 241.1245, 241.1245, 241.1245, 241.1244, 
    241.1244, 241.1244, 241.1244, 241.1244, 241.1244, 241.1244, 241.1243, 
    241.1243, 241.1243, 241.1243, 241.1243, 241.1243, 241.1242, 241.1242, 
    241.1242, 241.1242, 241.1242, 241.1241, 241.1241, 241.1241, 241.1241, 
    241.1241, 241.1241, 241.124, 241.124, 241.124, 241.124, 241.1239, 
    241.1239, 241.1239, 241.1239, 241.1239, 241.1239,
  242.1112, 242.1112, 242.1112, 242.1112, 242.1112, 242.1113, 242.1113, 
    242.1113, 242.1113, 242.1113, 242.1113, 242.1114, 242.1114, 242.1114, 
    242.1114, 242.1115, 242.1115, 242.1115, 242.1115, 242.1115, 242.1115, 
    242.1116, 242.1116, 242.1116, 242.1116, 242.1116, 242.1116, 242.1116, 
    242.1117, 242.1117, 242.1117, 242.1117, 242.1117, 242.1117, 242.1117, 
    242.1117, 242.1118, 242.1118, 242.1118, 242.1118, 242.1118, 242.1118, 
    242.1118, 242.1118, 242.1118, 242.1118, 242.1118, 242.1118, 242.1118, 
    242.1118, 242.1118, 242.1118, 242.1118, 242.1118, 242.1118, 242.1118, 
    242.1118, 242.1118, 242.1118, 242.1118, 242.1117, 242.1117, 242.1117, 
    242.1117, 242.1117, 242.1117, 242.1117, 242.1117, 242.1116, 242.1116, 
    242.1116, 242.1116, 242.1116, 242.1116, 242.1116, 242.1115, 242.1115, 
    242.1115, 242.1115, 242.1115, 242.1115, 242.1114, 242.1114, 242.1114, 
    242.1114, 242.1113, 242.1113, 242.1113, 242.1113, 242.1113, 242.1113, 
    242.1112, 242.1112, 242.1112, 242.1112, 242.1112,
  243.1037, 243.1037, 243.1037, 243.1038, 243.1038, 243.1038, 243.1038, 
    243.1038, 243.1039, 243.1039, 243.1039, 243.1039, 243.1039, 243.1039, 
    243.104, 243.104, 243.104, 243.104, 243.104, 243.104, 243.1041, 243.1041, 
    243.1041, 243.1041, 243.1041, 243.1042, 243.1042, 243.1042, 243.1042, 
    243.1042, 243.1042, 243.1042, 243.1042, 243.1042, 243.1043, 243.1043, 
    243.1043, 243.1043, 243.1043, 243.1043, 243.1043, 243.1043, 243.1043, 
    243.1043, 243.1043, 243.1043, 243.1043, 243.1043, 243.1043, 243.1043, 
    243.1043, 243.1043, 243.1043, 243.1043, 243.1043, 243.1043, 243.1043, 
    243.1043, 243.1043, 243.1043, 243.1043, 243.1043, 243.1042, 243.1042, 
    243.1042, 243.1042, 243.1042, 243.1042, 243.1042, 243.1042, 243.1042, 
    243.1041, 243.1041, 243.1041, 243.1041, 243.1041, 243.104, 243.104, 
    243.104, 243.104, 243.104, 243.104, 243.1039, 243.1039, 243.1039, 
    243.1039, 243.1039, 243.1039, 243.1038, 243.1038, 243.1038, 243.1038, 
    243.1038, 243.1037, 243.1037, 243.1037,
  244.1013, 244.1013, 244.1013, 244.1013, 244.1013, 244.1014, 244.1014, 
    244.1014, 244.1014, 244.1014, 244.1015, 244.1015, 244.1015, 244.1015, 
    244.1015, 244.1015, 244.1016, 244.1016, 244.1016, 244.1016, 244.1016, 
    244.1016, 244.1017, 244.1017, 244.1017, 244.1017, 244.1017, 244.1017, 
    244.1017, 244.1018, 244.1018, 244.1018, 244.1018, 244.1018, 244.1018, 
    244.1018, 244.1018, 244.1018, 244.1018, 244.1019, 244.1019, 244.1019, 
    244.1019, 244.1019, 244.1019, 244.1019, 244.1019, 244.1019, 244.1019, 
    244.1019, 244.1019, 244.1019, 244.1019, 244.1019, 244.1019, 244.1019, 
    244.1019, 244.1018, 244.1018, 244.1018, 244.1018, 244.1018, 244.1018, 
    244.1018, 244.1018, 244.1018, 244.1018, 244.1017, 244.1017, 244.1017, 
    244.1017, 244.1017, 244.1017, 244.1017, 244.1016, 244.1016, 244.1016, 
    244.1016, 244.1016, 244.1016, 244.1015, 244.1015, 244.1015, 244.1015, 
    244.1015, 244.1015, 244.1014, 244.1014, 244.1014, 244.1014, 244.1014, 
    244.1013, 244.1013, 244.1013, 244.1013, 244.1013,
  245.1036, 245.1037, 245.1037, 245.1037, 245.1037, 245.1037, 245.1037, 
    245.1037, 245.1038, 245.1038, 245.1038, 245.1038, 245.1038, 245.1039, 
    245.1039, 245.1039, 245.1039, 245.1039, 245.1039, 245.1039, 245.104, 
    245.104, 245.104, 245.104, 245.104, 245.104, 245.104, 245.104, 245.1041, 
    245.1041, 245.1041, 245.1041, 245.1041, 245.1041, 245.1041, 245.1041, 
    245.1041, 245.1042, 245.1042, 245.1042, 245.1042, 245.1042, 245.1042, 
    245.1042, 245.1042, 245.1042, 245.1042, 245.1042, 245.1042, 245.1042, 
    245.1042, 245.1042, 245.1042, 245.1042, 245.1042, 245.1042, 245.1042, 
    245.1042, 245.1042, 245.1041, 245.1041, 245.1041, 245.1041, 245.1041, 
    245.1041, 245.1041, 245.1041, 245.1041, 245.104, 245.104, 245.104, 
    245.104, 245.104, 245.104, 245.104, 245.104, 245.1039, 245.1039, 
    245.1039, 245.1039, 245.1039, 245.1039, 245.1039, 245.1038, 245.1038, 
    245.1038, 245.1038, 245.1038, 245.1037, 245.1037, 245.1037, 245.1037, 
    245.1037, 245.1037, 245.1037, 245.1036,
  246.1105, 246.1105, 246.1105, 246.1106, 246.1106, 246.1106, 246.1106, 
    246.1106, 246.1106, 246.1107, 246.1107, 246.1107, 246.1107, 246.1107, 
    246.1107, 246.1107, 246.1108, 246.1108, 246.1108, 246.1108, 246.1108, 
    246.1108, 246.1108, 246.1109, 246.1109, 246.1109, 246.1109, 246.1109, 
    246.1109, 246.1109, 246.1109, 246.1109, 246.111, 246.111, 246.111, 
    246.111, 246.111, 246.111, 246.111, 246.111, 246.111, 246.111, 246.111, 
    246.111, 246.111, 246.111, 246.111, 246.111, 246.111, 246.111, 246.111, 
    246.111, 246.111, 246.111, 246.111, 246.111, 246.111, 246.111, 246.111, 
    246.111, 246.111, 246.111, 246.111, 246.111, 246.1109, 246.1109, 
    246.1109, 246.1109, 246.1109, 246.1109, 246.1109, 246.1109, 246.1109, 
    246.1108, 246.1108, 246.1108, 246.1108, 246.1108, 246.1108, 246.1108, 
    246.1107, 246.1107, 246.1107, 246.1107, 246.1107, 246.1107, 246.1107, 
    246.1106, 246.1106, 246.1106, 246.1106, 246.1106, 246.1106, 246.1105, 
    246.1105, 246.1105,
  247.1217, 247.1217, 247.1217, 247.1217, 247.1217, 247.1217, 247.1217, 
    247.1217, 247.1218, 247.1218, 247.1218, 247.1218, 247.1218, 247.1218, 
    247.1219, 247.1219, 247.1219, 247.1219, 247.1219, 247.1219, 247.1219, 
    247.1219, 247.122, 247.122, 247.122, 247.122, 247.122, 247.122, 247.122, 
    247.122, 247.1221, 247.1221, 247.1221, 247.1221, 247.1221, 247.1221, 
    247.1221, 247.1221, 247.1221, 247.1221, 247.1221, 247.1221, 247.1221, 
    247.1221, 247.1221, 247.1221, 247.1221, 247.1221, 247.1221, 247.1221, 
    247.1221, 247.1221, 247.1221, 247.1221, 247.1221, 247.1221, 247.1221, 
    247.1221, 247.1221, 247.1221, 247.1221, 247.1221, 247.1221, 247.1221, 
    247.1221, 247.1221, 247.122, 247.122, 247.122, 247.122, 247.122, 247.122, 
    247.122, 247.122, 247.1219, 247.1219, 247.1219, 247.1219, 247.1219, 
    247.1219, 247.1219, 247.1219, 247.1218, 247.1218, 247.1218, 247.1218, 
    247.1218, 247.1218, 247.1217, 247.1217, 247.1217, 247.1217, 247.1217, 
    247.1217, 247.1217, 247.1217,
  248.1368, 248.1368, 248.1368, 248.1368, 248.1368, 248.1368, 248.1369, 
    248.1369, 248.1369, 248.1369, 248.1369, 248.1369, 248.1369, 248.1369, 
    248.137, 248.137, 248.137, 248.137, 248.137, 248.137, 248.137, 248.1371, 
    248.1371, 248.1371, 248.1371, 248.1371, 248.1371, 248.1371, 248.1371, 
    248.1371, 248.1371, 248.1372, 248.1372, 248.1372, 248.1372, 248.1372, 
    248.1372, 248.1372, 248.1372, 248.1372, 248.1372, 248.1372, 248.1372, 
    248.1372, 248.1372, 248.1372, 248.1372, 248.1372, 248.1372, 248.1372, 
    248.1372, 248.1372, 248.1372, 248.1372, 248.1372, 248.1372, 248.1372, 
    248.1372, 248.1372, 248.1372, 248.1372, 248.1372, 248.1372, 248.1372, 
    248.1372, 248.1371, 248.1371, 248.1371, 248.1371, 248.1371, 248.1371, 
    248.1371, 248.1371, 248.1371, 248.1371, 248.137, 248.137, 248.137, 
    248.137, 248.137, 248.137, 248.137, 248.1369, 248.1369, 248.1369, 
    248.1369, 248.1369, 248.1369, 248.1369, 248.1369, 248.1368, 248.1368, 
    248.1368, 248.1368, 248.1368, 248.1368,
  249.1556, 249.1556, 249.1556, 249.1557, 249.1557, 249.1557, 249.1557, 
    249.1557, 249.1557, 249.1557, 249.1557, 249.1557, 249.1558, 249.1558, 
    249.1558, 249.1558, 249.1558, 249.1558, 249.1558, 249.1559, 249.1559, 
    249.1559, 249.1559, 249.1559, 249.1559, 249.1559, 249.1559, 249.1559, 
    249.1559, 249.156, 249.156, 249.156, 249.156, 249.156, 249.156, 249.156, 
    249.156, 249.156, 249.156, 249.156, 249.156, 249.156, 249.156, 249.156, 
    249.156, 249.156, 249.156, 249.156, 249.156, 249.156, 249.156, 249.156, 
    249.156, 249.156, 249.156, 249.156, 249.156, 249.156, 249.156, 249.156, 
    249.156, 249.156, 249.156, 249.156, 249.156, 249.156, 249.156, 249.1559, 
    249.1559, 249.1559, 249.1559, 249.1559, 249.1559, 249.1559, 249.1559, 
    249.1559, 249.1559, 249.1558, 249.1558, 249.1558, 249.1558, 249.1558, 
    249.1558, 249.1558, 249.1557, 249.1557, 249.1557, 249.1557, 249.1557, 
    249.1557, 249.1557, 249.1557, 249.1557, 249.1556, 249.1556, 249.1556,
  250.1779, 250.1779, 250.1779, 250.1779, 250.1779, 250.1779, 250.1779, 
    250.1779, 250.178, 250.178, 250.178, 250.178, 250.178, 250.178, 250.178, 
    250.178, 250.1781, 250.1781, 250.1781, 250.1781, 250.1781, 250.1781, 
    250.1781, 250.1781, 250.1781, 250.1781, 250.1782, 250.1782, 250.1782, 
    250.1782, 250.1782, 250.1782, 250.1782, 250.1782, 250.1782, 250.1782, 
    250.1782, 250.1782, 250.1782, 250.1782, 250.1783, 250.1783, 250.1783, 
    250.1783, 250.1783, 250.1783, 250.1783, 250.1783, 250.1783, 250.1783, 
    250.1783, 250.1783, 250.1783, 250.1783, 250.1783, 250.1783, 250.1782, 
    250.1782, 250.1782, 250.1782, 250.1782, 250.1782, 250.1782, 250.1782, 
    250.1782, 250.1782, 250.1782, 250.1782, 250.1782, 250.1782, 250.1781, 
    250.1781, 250.1781, 250.1781, 250.1781, 250.1781, 250.1781, 250.1781, 
    250.1781, 250.1781, 250.178, 250.178, 250.178, 250.178, 250.178, 250.178, 
    250.178, 250.178, 250.1779, 250.1779, 250.1779, 250.1779, 250.1779, 
    250.1779, 250.1779, 250.1779,
  251.2033, 251.2033, 251.2033, 251.2033, 251.2033, 251.2033, 251.2033, 
    251.2033, 251.2033, 251.2033, 251.2034, 251.2034, 251.2034, 251.2034, 
    251.2034, 251.2034, 251.2034, 251.2034, 251.2034, 251.2034, 251.2035, 
    251.2035, 251.2035, 251.2035, 251.2035, 251.2035, 251.2035, 251.2035, 
    251.2035, 251.2035, 251.2035, 251.2035, 251.2036, 251.2036, 251.2036, 
    251.2036, 251.2036, 251.2036, 251.2036, 251.2036, 251.2036, 251.2036, 
    251.2036, 251.2036, 251.2036, 251.2036, 251.2036, 251.2036, 251.2036, 
    251.2036, 251.2036, 251.2036, 251.2036, 251.2036, 251.2036, 251.2036, 
    251.2036, 251.2036, 251.2036, 251.2036, 251.2036, 251.2036, 251.2036, 
    251.2036, 251.2035, 251.2035, 251.2035, 251.2035, 251.2035, 251.2035, 
    251.2035, 251.2035, 251.2035, 251.2035, 251.2035, 251.2035, 251.2034, 
    251.2034, 251.2034, 251.2034, 251.2034, 251.2034, 251.2034, 251.2034, 
    251.2034, 251.2034, 251.2033, 251.2033, 251.2033, 251.2033, 251.2033, 
    251.2033, 251.2033, 251.2033, 251.2033, 251.2033,
  252.2314, 252.2315, 252.2315, 252.2315, 252.2315, 252.2315, 252.2315, 
    252.2315, 252.2315, 252.2315, 252.2315, 252.2316, 252.2316, 252.2316, 
    252.2316, 252.2316, 252.2316, 252.2316, 252.2316, 252.2316, 252.2316, 
    252.2316, 252.2316, 252.2316, 252.2317, 252.2317, 252.2317, 252.2317, 
    252.2317, 252.2317, 252.2317, 252.2317, 252.2317, 252.2317, 252.2317, 
    252.2317, 252.2317, 252.2317, 252.2317, 252.2317, 252.2318, 252.2318, 
    252.2318, 252.2318, 252.2318, 252.2318, 252.2318, 252.2318, 252.2318, 
    252.2318, 252.2318, 252.2318, 252.2318, 252.2318, 252.2318, 252.2318, 
    252.2317, 252.2317, 252.2317, 252.2317, 252.2317, 252.2317, 252.2317, 
    252.2317, 252.2317, 252.2317, 252.2317, 252.2317, 252.2317, 252.2317, 
    252.2317, 252.2317, 252.2316, 252.2316, 252.2316, 252.2316, 252.2316, 
    252.2316, 252.2316, 252.2316, 252.2316, 252.2316, 252.2316, 252.2316, 
    252.2316, 252.2315, 252.2315, 252.2315, 252.2315, 252.2315, 252.2315, 
    252.2315, 252.2315, 252.2315, 252.2315, 252.2314,
  253.2621, 253.2621, 253.2622, 253.2622, 253.2622, 253.2622, 253.2622, 
    253.2622, 253.2622, 253.2622, 253.2622, 253.2622, 253.2622, 253.2622, 
    253.2623, 253.2623, 253.2623, 253.2623, 253.2623, 253.2623, 253.2623, 
    253.2623, 253.2623, 253.2623, 253.2623, 253.2623, 253.2623, 253.2623, 
    253.2623, 253.2623, 253.2624, 253.2624, 253.2624, 253.2624, 253.2624, 
    253.2624, 253.2624, 253.2624, 253.2624, 253.2624, 253.2624, 253.2624, 
    253.2624, 253.2624, 253.2624, 253.2624, 253.2624, 253.2624, 253.2624, 
    253.2624, 253.2624, 253.2624, 253.2624, 253.2624, 253.2624, 253.2624, 
    253.2624, 253.2624, 253.2624, 253.2624, 253.2624, 253.2624, 253.2624, 
    253.2624, 253.2624, 253.2624, 253.2623, 253.2623, 253.2623, 253.2623, 
    253.2623, 253.2623, 253.2623, 253.2623, 253.2623, 253.2623, 253.2623, 
    253.2623, 253.2623, 253.2623, 253.2623, 253.2623, 253.2622, 253.2622, 
    253.2622, 253.2622, 253.2622, 253.2622, 253.2622, 253.2622, 253.2622, 
    253.2622, 253.2622, 253.2622, 253.2621, 253.2621,
  254.295, 254.295, 254.295, 254.295, 254.295, 254.295, 254.295, 254.2951, 
    254.2951, 254.2951, 254.2951, 254.2951, 254.2951, 254.2951, 254.2951, 
    254.2951, 254.2951, 254.2951, 254.2951, 254.2951, 254.2951, 254.2952, 
    254.2952, 254.2952, 254.2952, 254.2952, 254.2952, 254.2952, 254.2952, 
    254.2952, 254.2952, 254.2952, 254.2952, 254.2952, 254.2952, 254.2952, 
    254.2952, 254.2952, 254.2952, 254.2952, 254.2952, 254.2952, 254.2952, 
    254.2952, 254.2952, 254.2952, 254.2952, 254.2952, 254.2952, 254.2952, 
    254.2952, 254.2952, 254.2952, 254.2952, 254.2952, 254.2952, 254.2952, 
    254.2952, 254.2952, 254.2952, 254.2952, 254.2952, 254.2952, 254.2952, 
    254.2952, 254.2952, 254.2952, 254.2952, 254.2952, 254.2952, 254.2952, 
    254.2952, 254.2952, 254.2952, 254.2952, 254.2951, 254.2951, 254.2951, 
    254.2951, 254.2951, 254.2951, 254.2951, 254.2951, 254.2951, 254.2951, 
    254.2951, 254.2951, 254.2951, 254.2951, 254.295, 254.295, 254.295, 
    254.295, 254.295, 254.295, 254.295,
  255.3297, 255.3297, 255.3297, 255.3298, 255.3298, 255.3298, 255.3298, 
    255.3298, 255.3298, 255.3298, 255.3298, 255.3298, 255.3298, 255.3298, 
    255.3298, 255.3298, 255.3298, 255.3298, 255.3298, 255.3298, 255.3298, 
    255.3298, 255.3298, 255.3299, 255.3299, 255.3299, 255.3299, 255.3299, 
    255.3299, 255.3299, 255.3299, 255.3299, 255.3299, 255.3299, 255.3299, 
    255.3299, 255.3299, 255.3299, 255.3299, 255.3299, 255.3299, 255.3299, 
    255.3299, 255.3299, 255.3299, 255.3299, 255.3299, 255.3299, 255.3299, 
    255.3299, 255.3299, 255.3299, 255.3299, 255.3299, 255.3299, 255.3299, 
    255.3299, 255.3299, 255.3299, 255.3299, 255.3299, 255.3299, 255.3299, 
    255.3299, 255.3299, 255.3299, 255.3299, 255.3299, 255.3299, 255.3299, 
    255.3299, 255.3299, 255.3299, 255.3298, 255.3298, 255.3298, 255.3298, 
    255.3298, 255.3298, 255.3298, 255.3298, 255.3298, 255.3298, 255.3298, 
    255.3298, 255.3298, 255.3298, 255.3298, 255.3298, 255.3298, 255.3298, 
    255.3298, 255.3298, 255.3297, 255.3297, 255.3297,
  256.366, 256.366, 256.366, 256.366, 256.366, 256.366, 256.366, 256.366, 
    256.366, 256.366, 256.366, 256.366, 256.366, 256.366, 256.3661, 256.3661, 
    256.3661, 256.3661, 256.3661, 256.3661, 256.3661, 256.3661, 256.3661, 
    256.3661, 256.3661, 256.3661, 256.3661, 256.3661, 256.3661, 256.3661, 
    256.3661, 256.3661, 256.3661, 256.3661, 256.3661, 256.3661, 256.3661, 
    256.3661, 256.3661, 256.3661, 256.3661, 256.3661, 256.3661, 256.3661, 
    256.3661, 256.3661, 256.3661, 256.3661, 256.3661, 256.3661, 256.3661, 
    256.3661, 256.3661, 256.3661, 256.3661, 256.3661, 256.3661, 256.3661, 
    256.3661, 256.3661, 256.3661, 256.3661, 256.3661, 256.3661, 256.3661, 
    256.3661, 256.3661, 256.3661, 256.3661, 256.3661, 256.3661, 256.3661, 
    256.3661, 256.3661, 256.3661, 256.3661, 256.3661, 256.3661, 256.3661, 
    256.3661, 256.3661, 256.3661, 256.366, 256.366, 256.366, 256.366, 
    256.366, 256.366, 256.366, 256.366, 256.366, 256.366, 256.366, 256.366, 
    256.366, 256.366,
  257.4034, 257.4034, 257.4034, 257.4034, 257.4034, 257.4034, 257.4034, 
    257.4034, 257.4034, 257.4034, 257.4034, 257.4034, 257.4035, 257.4035, 
    257.4035, 257.4035, 257.4035, 257.4035, 257.4035, 257.4035, 257.4035, 
    257.4035, 257.4035, 257.4035, 257.4035, 257.4035, 257.4035, 257.4035, 
    257.4035, 257.4035, 257.4035, 257.4035, 257.4035, 257.4035, 257.4035, 
    257.4035, 257.4035, 257.4035, 257.4035, 257.4035, 257.4035, 257.4035, 
    257.4035, 257.4035, 257.4035, 257.4035, 257.4035, 257.4035, 257.4035, 
    257.4035, 257.4035, 257.4035, 257.4035, 257.4035, 257.4035, 257.4035, 
    257.4035, 257.4035, 257.4035, 257.4035, 257.4035, 257.4035, 257.4035, 
    257.4035, 257.4035, 257.4035, 257.4035, 257.4035, 257.4035, 257.4035, 
    257.4035, 257.4035, 257.4035, 257.4035, 257.4035, 257.4035, 257.4035, 
    257.4035, 257.4035, 257.4035, 257.4035, 257.4035, 257.4035, 257.4035, 
    257.4034, 257.4034, 257.4034, 257.4034, 257.4034, 257.4034, 257.4034, 
    257.4034, 257.4034, 257.4034, 257.4034, 257.4034,
  258.4417, 258.4417, 258.4417, 258.4417, 258.4417, 258.4417, 258.4417, 
    258.4417, 258.4417, 258.4417, 258.4417, 258.4417, 258.4417, 258.4417, 
    258.4417, 258.4417, 258.4417, 258.4417, 258.4417, 258.4417, 258.4417, 
    258.4417, 258.4417, 258.4417, 258.4417, 258.4417, 258.4418, 258.4418, 
    258.4418, 258.4418, 258.4418, 258.4418, 258.4418, 258.4418, 258.4418, 
    258.4418, 258.4418, 258.4418, 258.4418, 258.4418, 258.4418, 258.4418, 
    258.4418, 258.4418, 258.4418, 258.4418, 258.4418, 258.4418, 258.4418, 
    258.4418, 258.4418, 258.4418, 258.4418, 258.4418, 258.4418, 258.4418, 
    258.4418, 258.4418, 258.4418, 258.4418, 258.4418, 258.4418, 258.4418, 
    258.4418, 258.4418, 258.4418, 258.4418, 258.4418, 258.4418, 258.4418, 
    258.4417, 258.4417, 258.4417, 258.4417, 258.4417, 258.4417, 258.4417, 
    258.4417, 258.4417, 258.4417, 258.4417, 258.4417, 258.4417, 258.4417, 
    258.4417, 258.4417, 258.4417, 258.4417, 258.4417, 258.4417, 258.4417, 
    258.4417, 258.4417, 258.4417, 258.4417, 258.4417,
  259.4805, 259.4805, 259.4805, 259.4805, 259.4805, 259.4805, 259.4805, 
    259.4805, 259.4805, 259.4805, 259.4805, 259.4805, 259.4805, 259.4805, 
    259.4805, 259.4805, 259.4805, 259.4805, 259.4805, 259.4805, 259.4805, 
    259.4805, 259.4805, 259.4805, 259.4805, 259.4805, 259.4805, 259.4805, 
    259.4805, 259.4805, 259.4805, 259.4805, 259.4805, 259.4805, 259.4805, 
    259.4805, 259.4805, 259.4805, 259.4805, 259.4805, 259.4805, 259.4805, 
    259.4805, 259.4805, 259.4805, 259.4805, 259.4805, 259.4805, 259.4805, 
    259.4805, 259.4805, 259.4805, 259.4805, 259.4805, 259.4805, 259.4805, 
    259.4805, 259.4805, 259.4805, 259.4805, 259.4805, 259.4805, 259.4805, 
    259.4805, 259.4805, 259.4805, 259.4805, 259.4805, 259.4805, 259.4805, 
    259.4805, 259.4805, 259.4805, 259.4805, 259.4805, 259.4805, 259.4805, 
    259.4805, 259.4805, 259.4805, 259.4805, 259.4805, 259.4805, 259.4805, 
    259.4805, 259.4805, 259.4805, 259.4805, 259.4805, 259.4805, 259.4805, 
    259.4805, 259.4805, 259.4805, 259.4805, 259.4805,
  260.5195, 260.5195, 260.5195, 260.5195, 260.5195, 260.5195, 260.5195, 
    260.5195, 260.5195, 260.5195, 260.5195, 260.5195, 260.5195, 260.5195, 
    260.5195, 260.5195, 260.5195, 260.5195, 260.5195, 260.5195, 260.5195, 
    260.5195, 260.5195, 260.5195, 260.5195, 260.5195, 260.5195, 260.5195, 
    260.5195, 260.5195, 260.5195, 260.5195, 260.5195, 260.5195, 260.5195, 
    260.5195, 260.5195, 260.5195, 260.5195, 260.5195, 260.5195, 260.5195, 
    260.5195, 260.5195, 260.5195, 260.5195, 260.5195, 260.5195, 260.5195, 
    260.5195, 260.5195, 260.5195, 260.5195, 260.5195, 260.5195, 260.5195, 
    260.5195, 260.5195, 260.5195, 260.5195, 260.5195, 260.5195, 260.5195, 
    260.5195, 260.5195, 260.5195, 260.5195, 260.5195, 260.5195, 260.5195, 
    260.5195, 260.5195, 260.5195, 260.5195, 260.5195, 260.5195, 260.5195, 
    260.5195, 260.5195, 260.5195, 260.5195, 260.5195, 260.5195, 260.5195, 
    260.5195, 260.5195, 260.5195, 260.5195, 260.5195, 260.5195, 260.5195, 
    260.5195, 260.5195, 260.5195, 260.5195, 260.5195,
  261.5583, 261.5583, 261.5583, 261.5583, 261.5583, 261.5583, 261.5583, 
    261.5583, 261.5583, 261.5583, 261.5583, 261.5583, 261.5583, 261.5583, 
    261.5583, 261.5583, 261.5583, 261.5583, 261.5583, 261.5583, 261.5583, 
    261.5583, 261.5583, 261.5583, 261.5583, 261.5583, 261.5582, 261.5582, 
    261.5582, 261.5582, 261.5582, 261.5582, 261.5582, 261.5582, 261.5582, 
    261.5582, 261.5582, 261.5582, 261.5582, 261.5582, 261.5582, 261.5582, 
    261.5582, 261.5582, 261.5582, 261.5582, 261.5582, 261.5582, 261.5582, 
    261.5582, 261.5582, 261.5582, 261.5582, 261.5582, 261.5582, 261.5582, 
    261.5582, 261.5582, 261.5582, 261.5582, 261.5582, 261.5582, 261.5582, 
    261.5582, 261.5582, 261.5582, 261.5582, 261.5582, 261.5582, 261.5582, 
    261.5583, 261.5583, 261.5583, 261.5583, 261.5583, 261.5583, 261.5583, 
    261.5583, 261.5583, 261.5583, 261.5583, 261.5583, 261.5583, 261.5583, 
    261.5583, 261.5583, 261.5583, 261.5583, 261.5583, 261.5583, 261.5583, 
    261.5583, 261.5583, 261.5583, 261.5583, 261.5583,
  262.5966, 262.5966, 262.5966, 262.5966, 262.5966, 262.5966, 262.5966, 
    262.5966, 262.5966, 262.5966, 262.5966, 262.5966, 262.5965, 262.5965, 
    262.5965, 262.5965, 262.5965, 262.5965, 262.5965, 262.5965, 262.5965, 
    262.5965, 262.5965, 262.5965, 262.5965, 262.5965, 262.5965, 262.5965, 
    262.5965, 262.5965, 262.5965, 262.5965, 262.5965, 262.5965, 262.5965, 
    262.5965, 262.5965, 262.5965, 262.5965, 262.5965, 262.5965, 262.5965, 
    262.5965, 262.5965, 262.5965, 262.5965, 262.5965, 262.5965, 262.5965, 
    262.5965, 262.5965, 262.5965, 262.5965, 262.5965, 262.5965, 262.5965, 
    262.5965, 262.5965, 262.5965, 262.5965, 262.5965, 262.5965, 262.5965, 
    262.5965, 262.5965, 262.5965, 262.5965, 262.5965, 262.5965, 262.5965, 
    262.5965, 262.5965, 262.5965, 262.5965, 262.5965, 262.5965, 262.5965, 
    262.5965, 262.5965, 262.5965, 262.5965, 262.5965, 262.5965, 262.5965, 
    262.5966, 262.5966, 262.5966, 262.5966, 262.5966, 262.5966, 262.5966, 
    262.5966, 262.5966, 262.5966, 262.5966, 262.5966,
  263.634, 263.634, 263.634, 263.634, 263.634, 263.634, 263.634, 263.634, 
    263.634, 263.634, 263.634, 263.634, 263.634, 263.634, 263.6339, 263.6339, 
    263.6339, 263.6339, 263.6339, 263.6339, 263.6339, 263.6339, 263.6339, 
    263.6339, 263.6339, 263.6339, 263.6339, 263.6339, 263.6339, 263.6339, 
    263.6339, 263.6339, 263.6339, 263.6339, 263.6339, 263.6339, 263.6339, 
    263.6339, 263.6339, 263.6339, 263.6339, 263.6339, 263.6339, 263.6339, 
    263.6339, 263.6339, 263.6339, 263.6339, 263.6339, 263.6339, 263.6339, 
    263.6339, 263.6339, 263.6339, 263.6339, 263.6339, 263.6339, 263.6339, 
    263.6339, 263.6339, 263.6339, 263.6339, 263.6339, 263.6339, 263.6339, 
    263.6339, 263.6339, 263.6339, 263.6339, 263.6339, 263.6339, 263.6339, 
    263.6339, 263.6339, 263.6339, 263.6339, 263.6339, 263.6339, 263.6339, 
    263.6339, 263.6339, 263.6339, 263.634, 263.634, 263.634, 263.634, 
    263.634, 263.634, 263.634, 263.634, 263.634, 263.634, 263.634, 263.634, 
    263.634, 263.634,
  264.6703, 264.6703, 264.6703, 264.6703, 264.6703, 264.6702, 264.6702, 
    264.6702, 264.6702, 264.6702, 264.6702, 264.6702, 264.6702, 264.6702, 
    264.6702, 264.6702, 264.6702, 264.6702, 264.6702, 264.6702, 264.6702, 
    264.6702, 264.6701, 264.6701, 264.6701, 264.6701, 264.6701, 264.6701, 
    264.6701, 264.6701, 264.6701, 264.6701, 264.6701, 264.6701, 264.6701, 
    264.6701, 264.6701, 264.6701, 264.6701, 264.6701, 264.6701, 264.6701, 
    264.6701, 264.6701, 264.6701, 264.6701, 264.6701, 264.6701, 264.6701, 
    264.6701, 264.6701, 264.6701, 264.6701, 264.6701, 264.6701, 264.6701, 
    264.6701, 264.6701, 264.6701, 264.6701, 264.6701, 264.6701, 264.6701, 
    264.6701, 264.6701, 264.6701, 264.6701, 264.6701, 264.6701, 264.6701, 
    264.6701, 264.6701, 264.6701, 264.6701, 264.6702, 264.6702, 264.6702, 
    264.6702, 264.6702, 264.6702, 264.6702, 264.6702, 264.6702, 264.6702, 
    264.6702, 264.6702, 264.6702, 264.6702, 264.6702, 264.6702, 264.6702, 
    264.6703, 264.6703, 264.6703, 264.6703, 264.6703,
  265.705, 265.705, 265.705, 265.705, 265.705, 265.705, 265.705, 265.705, 
    265.7049, 265.7049, 265.7049, 265.7049, 265.7049, 265.7049, 265.7049, 
    265.7049, 265.7049, 265.7049, 265.7049, 265.7049, 265.7049, 265.7049, 
    265.7048, 265.7048, 265.7048, 265.7048, 265.7048, 265.7048, 265.7048, 
    265.7048, 265.7048, 265.7048, 265.7048, 265.7048, 265.7048, 265.7048, 
    265.7048, 265.7048, 265.7048, 265.7048, 265.7048, 265.7048, 265.7048, 
    265.7048, 265.7048, 265.7048, 265.7048, 265.7048, 265.7048, 265.7048, 
    265.7048, 265.7048, 265.7048, 265.7048, 265.7048, 265.7048, 265.7048, 
    265.7048, 265.7048, 265.7048, 265.7048, 265.7048, 265.7048, 265.7048, 
    265.7048, 265.7048, 265.7048, 265.7048, 265.7048, 265.7048, 265.7048, 
    265.7048, 265.7048, 265.7048, 265.7049, 265.7049, 265.7049, 265.7049, 
    265.7049, 265.7049, 265.7049, 265.7049, 265.7049, 265.7049, 265.7049, 
    265.7049, 265.7049, 265.7049, 265.705, 265.705, 265.705, 265.705, 
    265.705, 265.705, 265.705, 265.705,
  266.7379, 266.7379, 266.7379, 266.7378, 266.7378, 266.7378, 266.7378, 
    266.7378, 266.7378, 266.7378, 266.7378, 266.7378, 266.7378, 266.7378, 
    266.7378, 266.7377, 266.7377, 266.7377, 266.7377, 266.7377, 266.7377, 
    266.7377, 266.7377, 266.7377, 266.7377, 266.7377, 266.7377, 266.7377, 
    266.7376, 266.7376, 266.7376, 266.7376, 266.7376, 266.7376, 266.7376, 
    266.7376, 266.7376, 266.7376, 266.7376, 266.7376, 266.7376, 266.7376, 
    266.7376, 266.7376, 266.7376, 266.7376, 266.7376, 266.7376, 266.7376, 
    266.7376, 266.7376, 266.7376, 266.7376, 266.7376, 266.7376, 266.7376, 
    266.7376, 266.7376, 266.7376, 266.7376, 266.7376, 266.7376, 266.7376, 
    266.7376, 266.7376, 266.7376, 266.7376, 266.7376, 266.7377, 266.7377, 
    266.7377, 266.7377, 266.7377, 266.7377, 266.7377, 266.7377, 266.7377, 
    266.7377, 266.7377, 266.7377, 266.7377, 266.7378, 266.7378, 266.7378, 
    266.7378, 266.7378, 266.7378, 266.7378, 266.7378, 266.7378, 266.7378, 
    266.7378, 266.7378, 266.7379, 266.7379, 266.7379,
  267.7686, 267.7686, 267.7685, 267.7685, 267.7685, 267.7685, 267.7685, 
    267.7685, 267.7685, 267.7685, 267.7685, 267.7685, 267.7684, 267.7684, 
    267.7684, 267.7684, 267.7684, 267.7684, 267.7684, 267.7684, 267.7684, 
    267.7684, 267.7684, 267.7683, 267.7683, 267.7683, 267.7683, 267.7683, 
    267.7683, 267.7683, 267.7683, 267.7683, 267.7683, 267.7683, 267.7683, 
    267.7683, 267.7683, 267.7683, 267.7682, 267.7682, 267.7682, 267.7682, 
    267.7682, 267.7682, 267.7682, 267.7682, 267.7682, 267.7682, 267.7682, 
    267.7682, 267.7682, 267.7682, 267.7682, 267.7682, 267.7682, 267.7682, 
    267.7682, 267.7682, 267.7683, 267.7683, 267.7683, 267.7683, 267.7683, 
    267.7683, 267.7683, 267.7683, 267.7683, 267.7683, 267.7683, 267.7683, 
    267.7683, 267.7683, 267.7683, 267.7684, 267.7684, 267.7684, 267.7684, 
    267.7684, 267.7684, 267.7684, 267.7684, 267.7684, 267.7684, 267.7684, 
    267.7685, 267.7685, 267.7685, 267.7685, 267.7685, 267.7685, 267.7685, 
    267.7685, 267.7685, 267.7685, 267.7686, 267.7686,
  268.7968, 268.7967, 268.7967, 268.7967, 268.7967, 268.7967, 268.7967, 
    268.7967, 268.7967, 268.7967, 268.7966, 268.7966, 268.7966, 268.7966, 
    268.7966, 268.7966, 268.7966, 268.7966, 268.7966, 268.7966, 268.7965, 
    268.7965, 268.7965, 268.7965, 268.7965, 268.7965, 268.7965, 268.7965, 
    268.7965, 268.7965, 268.7965, 268.7964, 268.7964, 268.7964, 268.7964, 
    268.7964, 268.7964, 268.7964, 268.7964, 268.7964, 268.7964, 268.7964, 
    268.7964, 268.7964, 268.7964, 268.7964, 268.7964, 268.7964, 268.7964, 
    268.7964, 268.7964, 268.7964, 268.7964, 268.7964, 268.7964, 268.7964, 
    268.7964, 268.7964, 268.7964, 268.7964, 268.7964, 268.7964, 268.7964, 
    268.7964, 268.7964, 268.7965, 268.7965, 268.7965, 268.7965, 268.7965, 
    268.7965, 268.7965, 268.7965, 268.7965, 268.7965, 268.7965, 268.7966, 
    268.7966, 268.7966, 268.7966, 268.7966, 268.7966, 268.7966, 268.7966, 
    268.7966, 268.7966, 268.7967, 268.7967, 268.7967, 268.7967, 268.7967, 
    268.7967, 268.7967, 268.7967, 268.7967, 268.7968,
  269.8221, 269.8221, 269.8221, 269.8221, 269.8221, 269.8221, 269.8221, 
    269.8221, 269.822, 269.822, 269.822, 269.822, 269.822, 269.822, 269.822, 
    269.822, 269.8219, 269.8219, 269.8219, 269.8219, 269.8219, 269.8219, 
    269.8219, 269.8219, 269.8219, 269.8218, 269.8218, 269.8218, 269.8218, 
    269.8218, 269.8218, 269.8218, 269.8218, 269.8218, 269.8218, 269.8218, 
    269.8218, 269.8218, 269.8217, 269.8217, 269.8217, 269.8217, 269.8217, 
    269.8217, 269.8217, 269.8217, 269.8217, 269.8217, 269.8217, 269.8217, 
    269.8217, 269.8217, 269.8217, 269.8217, 269.8217, 269.8217, 269.8217, 
    269.8217, 269.8218, 269.8218, 269.8218, 269.8218, 269.8218, 269.8218, 
    269.8218, 269.8218, 269.8218, 269.8218, 269.8218, 269.8218, 269.8218, 
    269.8219, 269.8219, 269.8219, 269.8219, 269.8219, 269.8219, 269.8219, 
    269.8219, 269.8219, 269.822, 269.822, 269.822, 269.822, 269.822, 269.822, 
    269.822, 269.822, 269.8221, 269.8221, 269.8221, 269.8221, 269.8221, 
    269.8221, 269.8221, 269.8221,
  270.8444, 270.8444, 270.8444, 270.8443, 270.8443, 270.8443, 270.8443, 
    270.8443, 270.8443, 270.8443, 270.8443, 270.8442, 270.8442, 270.8442, 
    270.8442, 270.8442, 270.8442, 270.8442, 270.8442, 270.8441, 270.8441, 
    270.8441, 270.8441, 270.8441, 270.8441, 270.8441, 270.8441, 270.8441, 
    270.8441, 270.8441, 270.844, 270.844, 270.844, 270.844, 270.844, 270.844, 
    270.844, 270.844, 270.844, 270.844, 270.844, 270.844, 270.844, 270.844, 
    270.844, 270.844, 270.844, 270.844, 270.844, 270.844, 270.844, 270.844, 
    270.844, 270.844, 270.844, 270.844, 270.844, 270.844, 270.844, 270.844, 
    270.844, 270.844, 270.844, 270.844, 270.844, 270.844, 270.8441, 270.8441, 
    270.8441, 270.8441, 270.8441, 270.8441, 270.8441, 270.8441, 270.8441, 
    270.8441, 270.8441, 270.8442, 270.8442, 270.8442, 270.8442, 270.8442, 
    270.8442, 270.8442, 270.8442, 270.8443, 270.8443, 270.8443, 270.8443, 
    270.8443, 270.8443, 270.8443, 270.8443, 270.8444, 270.8444, 270.8444,
  271.8632, 271.8632, 271.8632, 271.8632, 271.8632, 271.8632, 271.8631, 
    271.8631, 271.8631, 271.8631, 271.8631, 271.8631, 271.8631, 271.863, 
    271.863, 271.863, 271.863, 271.863, 271.863, 271.863, 271.8629, 271.8629, 
    271.8629, 271.8629, 271.8629, 271.8629, 271.8629, 271.8629, 271.8629, 
    271.8629, 271.8629, 271.8629, 271.8628, 271.8628, 271.8628, 271.8628, 
    271.8628, 271.8628, 271.8628, 271.8628, 271.8628, 271.8628, 271.8628, 
    271.8628, 271.8628, 271.8628, 271.8628, 271.8628, 271.8628, 271.8628, 
    271.8628, 271.8628, 271.8628, 271.8628, 271.8628, 271.8628, 271.8628, 
    271.8628, 271.8628, 271.8628, 271.8628, 271.8628, 271.8628, 271.8628, 
    271.8629, 271.8629, 271.8629, 271.8629, 271.8629, 271.8629, 271.8629, 
    271.8629, 271.8629, 271.8629, 271.8629, 271.8629, 271.863, 271.863, 
    271.863, 271.863, 271.863, 271.863, 271.863, 271.8631, 271.8631, 
    271.8631, 271.8631, 271.8631, 271.8631, 271.8631, 271.8632, 271.8632, 
    271.8632, 271.8632, 271.8632, 271.8632,
  272.8784, 272.8783, 272.8783, 272.8783, 272.8783, 272.8783, 272.8783, 
    272.8782, 272.8782, 272.8782, 272.8782, 272.8782, 272.8782, 272.8782, 
    272.8781, 272.8781, 272.8781, 272.8781, 272.8781, 272.8781, 272.8781, 
    272.8781, 272.8781, 272.878, 272.878, 272.878, 272.878, 272.878, 272.878, 
    272.878, 272.878, 272.8779, 272.8779, 272.8779, 272.8779, 272.8779, 
    272.8779, 272.8779, 272.8779, 272.8779, 272.8779, 272.8779, 272.8779, 
    272.8779, 272.8779, 272.8779, 272.8779, 272.8779, 272.8779, 272.8779, 
    272.8779, 272.8779, 272.8779, 272.8779, 272.8779, 272.8779, 272.8779, 
    272.8779, 272.8779, 272.8779, 272.8779, 272.8779, 272.8779, 272.8779, 
    272.8779, 272.878, 272.878, 272.878, 272.878, 272.878, 272.878, 272.878, 
    272.878, 272.8781, 272.8781, 272.8781, 272.8781, 272.8781, 272.8781, 
    272.8781, 272.8781, 272.8781, 272.8782, 272.8782, 272.8782, 272.8782, 
    272.8782, 272.8782, 272.8782, 272.8783, 272.8783, 272.8783, 272.8783, 
    272.8783, 272.8783, 272.8784,
  273.8895, 273.8895, 273.8895, 273.8894, 273.8894, 273.8894, 273.8894, 
    273.8894, 273.8894, 273.8893, 273.8893, 273.8893, 273.8893, 273.8893, 
    273.8893, 273.8893, 273.8893, 273.8892, 273.8892, 273.8892, 273.8892, 
    273.8892, 273.8892, 273.8891, 273.8891, 273.8891, 273.8891, 273.8891, 
    273.8891, 273.8891, 273.8891, 273.889, 273.889, 273.889, 273.889, 
    273.889, 273.889, 273.889, 273.889, 273.889, 273.889, 273.889, 273.889, 
    273.889, 273.889, 273.889, 273.889, 273.889, 273.889, 273.889, 273.889, 
    273.889, 273.889, 273.889, 273.889, 273.889, 273.889, 273.889, 273.889, 
    273.889, 273.889, 273.889, 273.889, 273.889, 273.889, 273.8891, 273.8891, 
    273.8891, 273.8891, 273.8891, 273.8891, 273.8891, 273.8891, 273.8892, 
    273.8892, 273.8892, 273.8892, 273.8892, 273.8892, 273.8893, 273.8893, 
    273.8893, 273.8893, 273.8893, 273.8893, 273.8893, 273.8893, 273.8894, 
    273.8894, 273.8894, 273.8894, 273.8894, 273.8894, 273.8895, 273.8895, 
    273.8895,
  274.8964, 274.8963, 274.8963, 274.8963, 274.8963, 274.8963, 274.8963, 
    274.8962, 274.8962, 274.8962, 274.8962, 274.8962, 274.8962, 274.8961, 
    274.8961, 274.8961, 274.8961, 274.8961, 274.8961, 274.8961, 274.896, 
    274.896, 274.896, 274.896, 274.896, 274.896, 274.896, 274.8959, 274.8959, 
    274.8959, 274.8959, 274.8959, 274.8959, 274.8959, 274.8959, 274.8959, 
    274.8958, 274.8958, 274.8958, 274.8958, 274.8958, 274.8958, 274.8958, 
    274.8958, 274.8958, 274.8958, 274.8958, 274.8958, 274.8958, 274.8958, 
    274.8958, 274.8958, 274.8958, 274.8958, 274.8958, 274.8958, 274.8958, 
    274.8958, 274.8958, 274.8958, 274.8959, 274.8959, 274.8959, 274.8959, 
    274.8959, 274.8959, 274.8959, 274.8959, 274.8959, 274.896, 274.896, 
    274.896, 274.896, 274.896, 274.896, 274.896, 274.8961, 274.8961, 
    274.8961, 274.8961, 274.8961, 274.8961, 274.8961, 274.8962, 274.8962, 
    274.8962, 274.8962, 274.8962, 274.8962, 274.8963, 274.8963, 274.8963, 
    274.8963, 274.8963, 274.8963, 274.8964,
  275.8987, 275.8987, 275.8987, 275.8987, 275.8987, 275.8986, 275.8986, 
    275.8986, 275.8986, 275.8986, 275.8985, 275.8985, 275.8985, 275.8985, 
    275.8985, 275.8985, 275.8984, 275.8984, 275.8984, 275.8984, 275.8984, 
    275.8983, 275.8983, 275.8983, 275.8983, 275.8983, 275.8983, 275.8983, 
    275.8983, 275.8983, 275.8982, 275.8982, 275.8982, 275.8982, 275.8982, 
    275.8982, 275.8982, 275.8982, 275.8982, 275.8982, 275.8981, 275.8981, 
    275.8981, 275.8981, 275.8981, 275.8981, 275.8981, 275.8981, 275.8981, 
    275.8981, 275.8981, 275.8981, 275.8981, 275.8981, 275.8981, 275.8981, 
    275.8982, 275.8982, 275.8982, 275.8982, 275.8982, 275.8982, 275.8982, 
    275.8982, 275.8982, 275.8982, 275.8983, 275.8983, 275.8983, 275.8983, 
    275.8983, 275.8983, 275.8983, 275.8983, 275.8983, 275.8984, 275.8984, 
    275.8984, 275.8984, 275.8984, 275.8985, 275.8985, 275.8985, 275.8985, 
    275.8985, 275.8985, 275.8986, 275.8986, 275.8986, 275.8986, 275.8986, 
    275.8987, 275.8987, 275.8987, 275.8987, 275.8987,
  276.8963, 276.8963, 276.8962, 276.8962, 276.8962, 276.8962, 276.8962, 
    276.8961, 276.8961, 276.8961, 276.8961, 276.8961, 276.8961, 276.8961, 
    276.896, 276.896, 276.896, 276.896, 276.896, 276.8959, 276.8959, 
    276.8959, 276.8959, 276.8959, 276.8959, 276.8958, 276.8958, 276.8958, 
    276.8958, 276.8958, 276.8958, 276.8958, 276.8958, 276.8958, 276.8958, 
    276.8957, 276.8957, 276.8957, 276.8957, 276.8957, 276.8957, 276.8957, 
    276.8957, 276.8957, 276.8957, 276.8957, 276.8957, 276.8957, 276.8957, 
    276.8957, 276.8957, 276.8957, 276.8957, 276.8957, 276.8957, 276.8957, 
    276.8957, 276.8957, 276.8957, 276.8957, 276.8957, 276.8958, 276.8958, 
    276.8958, 276.8958, 276.8958, 276.8958, 276.8958, 276.8958, 276.8958, 
    276.8958, 276.8959, 276.8959, 276.8959, 276.8959, 276.8959, 276.8959, 
    276.896, 276.896, 276.896, 276.896, 276.896, 276.8961, 276.8961, 
    276.8961, 276.8961, 276.8961, 276.8961, 276.8961, 276.8962, 276.8962, 
    276.8962, 276.8962, 276.8962, 276.8963, 276.8963,
  277.8889, 277.8888, 277.8888, 277.8888, 277.8888, 277.8887, 277.8887, 
    277.8887, 277.8887, 277.8887, 277.8886, 277.8886, 277.8886, 277.8886, 
    277.8886, 277.8885, 277.8885, 277.8885, 277.8885, 277.8885, 277.8885, 
    277.8885, 277.8884, 277.8884, 277.8884, 277.8884, 277.8884, 277.8884, 
    277.8883, 277.8883, 277.8883, 277.8883, 277.8883, 277.8883, 277.8883, 
    277.8882, 277.8882, 277.8882, 277.8882, 277.8882, 277.8882, 277.8882, 
    277.8882, 277.8882, 277.8882, 277.8882, 277.8882, 277.8882, 277.8882, 
    277.8882, 277.8882, 277.8882, 277.8882, 277.8882, 277.8882, 277.8882, 
    277.8882, 277.8882, 277.8882, 277.8882, 277.8882, 277.8883, 277.8883, 
    277.8883, 277.8883, 277.8883, 277.8883, 277.8883, 277.8884, 277.8884, 
    277.8884, 277.8884, 277.8884, 277.8884, 277.8885, 277.8885, 277.8885, 
    277.8885, 277.8885, 277.8885, 277.8885, 277.8886, 277.8886, 277.8886, 
    277.8886, 277.8886, 277.8887, 277.8887, 277.8887, 277.8887, 277.8887, 
    277.8888, 277.8888, 277.8888, 277.8888, 277.8889,
  278.8762, 278.8761, 278.8761, 278.8761, 278.8761, 278.876, 278.876, 
    278.876, 278.876, 278.876, 278.8759, 278.8759, 278.8759, 278.8759, 
    278.8759, 278.8759, 278.8758, 278.8758, 278.8758, 278.8758, 278.8758, 
    278.8757, 278.8757, 278.8757, 278.8757, 278.8757, 278.8757, 278.8756, 
    278.8756, 278.8756, 278.8756, 278.8756, 278.8756, 278.8756, 278.8755, 
    278.8755, 278.8755, 278.8755, 278.8755, 278.8755, 278.8755, 278.8755, 
    278.8755, 278.8755, 278.8755, 278.8755, 278.8755, 278.8755, 278.8755, 
    278.8755, 278.8755, 278.8755, 278.8755, 278.8755, 278.8755, 278.8755, 
    278.8755, 278.8755, 278.8755, 278.8755, 278.8755, 278.8755, 278.8756, 
    278.8756, 278.8756, 278.8756, 278.8756, 278.8756, 278.8756, 278.8757, 
    278.8757, 278.8757, 278.8757, 278.8757, 278.8757, 278.8758, 278.8758, 
    278.8758, 278.8758, 278.8758, 278.8759, 278.8759, 278.8759, 278.8759, 
    278.8759, 278.8759, 278.876, 278.876, 278.876, 278.876, 278.876, 
    278.8761, 278.8761, 278.8761, 278.8761, 278.8762,
  279.858, 279.858, 279.8579, 279.8579, 279.8579, 279.8579, 279.8579, 
    279.8578, 279.8578, 279.8578, 279.8578, 279.8578, 279.8578, 279.8577, 
    279.8577, 279.8577, 279.8577, 279.8576, 279.8576, 279.8576, 279.8576, 
    279.8576, 279.8575, 279.8575, 279.8575, 279.8575, 279.8575, 279.8575, 
    279.8575, 279.8575, 279.8574, 279.8574, 279.8574, 279.8574, 279.8574, 
    279.8574, 279.8574, 279.8573, 279.8573, 279.8573, 279.8573, 279.8573, 
    279.8573, 279.8573, 279.8573, 279.8573, 279.8573, 279.8573, 279.8573, 
    279.8573, 279.8573, 279.8573, 279.8573, 279.8573, 279.8573, 279.8573, 
    279.8573, 279.8573, 279.8573, 279.8574, 279.8574, 279.8574, 279.8574, 
    279.8574, 279.8574, 279.8574, 279.8575, 279.8575, 279.8575, 279.8575, 
    279.8575, 279.8575, 279.8575, 279.8575, 279.8576, 279.8576, 279.8576, 
    279.8576, 279.8576, 279.8577, 279.8577, 279.8577, 279.8577, 279.8578, 
    279.8578, 279.8578, 279.8578, 279.8578, 279.8578, 279.8579, 279.8579, 
    279.8579, 279.8579, 279.8579, 279.858, 279.858,
  280.8342, 280.8341, 280.8341, 280.8341, 280.8341, 280.8341, 280.834, 
    280.834, 280.834, 280.834, 280.834, 280.8339, 280.8339, 280.8339, 
    280.8339, 280.8339, 280.8338, 280.8338, 280.8338, 280.8338, 280.8337, 
    280.8337, 280.8337, 280.8337, 280.8337, 280.8336, 280.8336, 280.8336, 
    280.8336, 280.8336, 280.8336, 280.8336, 280.8336, 280.8335, 280.8335, 
    280.8335, 280.8335, 280.8335, 280.8335, 280.8335, 280.8335, 280.8335, 
    280.8335, 280.8335, 280.8335, 280.8335, 280.8334, 280.8334, 280.8334, 
    280.8334, 280.8335, 280.8335, 280.8335, 280.8335, 280.8335, 280.8335, 
    280.8335, 280.8335, 280.8335, 280.8335, 280.8335, 280.8335, 280.8335, 
    280.8336, 280.8336, 280.8336, 280.8336, 280.8336, 280.8336, 280.8336, 
    280.8336, 280.8337, 280.8337, 280.8337, 280.8337, 280.8337, 280.8338, 
    280.8338, 280.8338, 280.8338, 280.8339, 280.8339, 280.8339, 280.8339, 
    280.8339, 280.834, 280.834, 280.834, 280.834, 280.834, 280.8341, 
    280.8341, 280.8341, 280.8341, 280.8341, 280.8342,
  281.8045, 281.8044, 281.8044, 281.8044, 281.8044, 281.8044, 281.8044, 
    281.8043, 281.8043, 281.8043, 281.8043, 281.8042, 281.8042, 281.8042, 
    281.8042, 281.8041, 281.8041, 281.8041, 281.8041, 281.8041, 281.804, 
    281.804, 281.804, 281.804, 281.804, 281.804, 281.8039, 281.8039, 
    281.8039, 281.8039, 281.8039, 281.8039, 281.8038, 281.8038, 281.8038, 
    281.8038, 281.8038, 281.8038, 281.8038, 281.8038, 281.8038, 281.8037, 
    281.8037, 281.8037, 281.8037, 281.8037, 281.8037, 281.8037, 281.8037, 
    281.8037, 281.8037, 281.8037, 281.8037, 281.8037, 281.8037, 281.8038, 
    281.8038, 281.8038, 281.8038, 281.8038, 281.8038, 281.8038, 281.8038, 
    281.8038, 281.8039, 281.8039, 281.8039, 281.8039, 281.8039, 281.8039, 
    281.804, 281.804, 281.804, 281.804, 281.804, 281.804, 281.8041, 281.8041, 
    281.8041, 281.8041, 281.8041, 281.8042, 281.8042, 281.8042, 281.8042, 
    281.8043, 281.8043, 281.8043, 281.8043, 281.8044, 281.8044, 281.8044, 
    281.8044, 281.8044, 281.8044, 281.8045,
  282.7687, 282.7687, 282.7687, 282.7687, 282.7686, 282.7686, 282.7686, 
    282.7686, 282.7686, 282.7685, 282.7685, 282.7685, 282.7685, 282.7684, 
    282.7684, 282.7684, 282.7684, 282.7683, 282.7683, 282.7683, 282.7683, 
    282.7683, 282.7682, 282.7682, 282.7682, 282.7682, 282.7682, 282.7682, 
    282.7681, 282.7681, 282.7681, 282.7681, 282.7681, 282.7681, 282.7681, 
    282.768, 282.768, 282.768, 282.768, 282.768, 282.768, 282.768, 282.768, 
    282.768, 282.768, 282.768, 282.768, 282.768, 282.768, 282.768, 282.768, 
    282.768, 282.768, 282.768, 282.768, 282.768, 282.768, 282.768, 282.768, 
    282.768, 282.768, 282.7681, 282.7681, 282.7681, 282.7681, 282.7681, 
    282.7681, 282.7681, 282.7682, 282.7682, 282.7682, 282.7682, 282.7682, 
    282.7682, 282.7683, 282.7683, 282.7683, 282.7683, 282.7683, 282.7684, 
    282.7684, 282.7684, 282.7684, 282.7685, 282.7685, 282.7685, 282.7685, 
    282.7686, 282.7686, 282.7686, 282.7686, 282.7686, 282.7687, 282.7687, 
    282.7687, 282.7687,
  283.7268, 283.7267, 283.7267, 283.7267, 283.7267, 283.7267, 283.7266, 
    283.7266, 283.7266, 283.7266, 283.7265, 283.7265, 283.7265, 283.7265, 
    283.7264, 283.7264, 283.7264, 283.7264, 283.7263, 283.7263, 283.7263, 
    283.7263, 283.7263, 283.7263, 283.7262, 283.7262, 283.7262, 283.7262, 
    283.7262, 283.7261, 283.7261, 283.7261, 283.7261, 283.7261, 283.7261, 
    283.7261, 283.726, 283.726, 283.726, 283.726, 283.726, 283.726, 283.726, 
    283.726, 283.726, 283.726, 283.726, 283.726, 283.726, 283.726, 283.726, 
    283.726, 283.726, 283.726, 283.726, 283.726, 283.726, 283.726, 283.726, 
    283.726, 283.7261, 283.7261, 283.7261, 283.7261, 283.7261, 283.7261, 
    283.7261, 283.7262, 283.7262, 283.7262, 283.7262, 283.7262, 283.7263, 
    283.7263, 283.7263, 283.7263, 283.7263, 283.7263, 283.7264, 283.7264, 
    283.7264, 283.7264, 283.7265, 283.7265, 283.7265, 283.7265, 283.7266, 
    283.7266, 283.7266, 283.7266, 283.7267, 283.7267, 283.7267, 283.7267, 
    283.7267, 283.7268,
  284.6784, 284.6784, 284.6784, 284.6784, 284.6783, 284.6783, 284.6783, 
    284.6783, 284.6783, 284.6782, 284.6782, 284.6782, 284.6782, 284.6781, 
    284.6781, 284.6781, 284.6781, 284.678, 284.678, 284.678, 284.678, 
    284.6779, 284.6779, 284.6779, 284.6779, 284.6779, 284.6779, 284.6778, 
    284.6778, 284.6778, 284.6778, 284.6778, 284.6778, 284.6777, 284.6777, 
    284.6777, 284.6777, 284.6777, 284.6777, 284.6777, 284.6777, 284.6777, 
    284.6776, 284.6776, 284.6776, 284.6776, 284.6776, 284.6776, 284.6776, 
    284.6776, 284.6776, 284.6776, 284.6776, 284.6776, 284.6777, 284.6777, 
    284.6777, 284.6777, 284.6777, 284.6777, 284.6777, 284.6777, 284.6777, 
    284.6778, 284.6778, 284.6778, 284.6778, 284.6778, 284.6778, 284.6779, 
    284.6779, 284.6779, 284.6779, 284.6779, 284.6779, 284.678, 284.678, 
    284.678, 284.678, 284.6781, 284.6781, 284.6781, 284.6781, 284.6782, 
    284.6782, 284.6782, 284.6782, 284.6783, 284.6783, 284.6783, 284.6783, 
    284.6783, 284.6784, 284.6784, 284.6784, 284.6784,
  285.6236, 285.6236, 285.6235, 285.6235, 285.6235, 285.6234, 285.6234, 
    285.6234, 285.6234, 285.6234, 285.6233, 285.6233, 285.6233, 285.6233, 
    285.6232, 285.6232, 285.6232, 285.6232, 285.6231, 285.6231, 285.6231, 
    285.6231, 285.623, 285.623, 285.623, 285.623, 285.623, 285.623, 285.6229, 
    285.6229, 285.6229, 285.6229, 285.6229, 285.6229, 285.6229, 285.6228, 
    285.6228, 285.6228, 285.6228, 285.6228, 285.6228, 285.6228, 285.6228, 
    285.6228, 285.6228, 285.6228, 285.6228, 285.6228, 285.6228, 285.6228, 
    285.6228, 285.6228, 285.6228, 285.6228, 285.6228, 285.6228, 285.6228, 
    285.6228, 285.6228, 285.6228, 285.6228, 285.6229, 285.6229, 285.6229, 
    285.6229, 285.6229, 285.6229, 285.6229, 285.623, 285.623, 285.623, 
    285.623, 285.623, 285.623, 285.6231, 285.6231, 285.6231, 285.6231, 
    285.6232, 285.6232, 285.6232, 285.6232, 285.6233, 285.6233, 285.6233, 
    285.6233, 285.6234, 285.6234, 285.6234, 285.6234, 285.6234, 285.6235, 
    285.6235, 285.6235, 285.6236, 285.6236,
  286.5621, 286.562, 286.562, 286.562, 286.562, 286.5619, 286.5619, 286.5619, 
    286.5619, 286.5618, 286.5618, 286.5618, 286.5618, 286.5617, 286.5617, 
    286.5617, 286.5616, 286.5616, 286.5616, 286.5616, 286.5616, 286.5616, 
    286.5615, 286.5615, 286.5615, 286.5615, 286.5614, 286.5614, 286.5614, 
    286.5614, 286.5614, 286.5614, 286.5613, 286.5613, 286.5613, 286.5613, 
    286.5613, 286.5613, 286.5613, 286.5612, 286.5612, 286.5612, 286.5612, 
    286.5612, 286.5612, 286.5612, 286.5612, 286.5612, 286.5612, 286.5612, 
    286.5612, 286.5612, 286.5612, 286.5612, 286.5612, 286.5612, 286.5612, 
    286.5613, 286.5613, 286.5613, 286.5613, 286.5613, 286.5613, 286.5613, 
    286.5614, 286.5614, 286.5614, 286.5614, 286.5614, 286.5614, 286.5615, 
    286.5615, 286.5615, 286.5615, 286.5616, 286.5616, 286.5616, 286.5616, 
    286.5616, 286.5616, 286.5617, 286.5617, 286.5617, 286.5618, 286.5618, 
    286.5618, 286.5618, 286.5619, 286.5619, 286.5619, 286.5619, 286.562, 
    286.562, 286.562, 286.562, 286.5621,
  287.4938, 287.4937, 287.4937, 287.4937, 287.4937, 287.4936, 287.4936, 
    287.4936, 287.4936, 287.4935, 287.4935, 287.4935, 287.4934, 287.4934, 
    287.4934, 287.4934, 287.4933, 287.4933, 287.4933, 287.4933, 287.4933, 
    287.4932, 287.4932, 287.4932, 287.4932, 287.4932, 287.4931, 287.4931, 
    287.4931, 287.4931, 287.4931, 287.493, 287.493, 287.493, 287.493, 
    287.493, 287.493, 287.493, 287.493, 287.493, 287.493, 287.4929, 287.4929, 
    287.4929, 287.4929, 287.4929, 287.4929, 287.4929, 287.4929, 287.4929, 
    287.4929, 287.4929, 287.4929, 287.4929, 287.4929, 287.493, 287.493, 
    287.493, 287.493, 287.493, 287.493, 287.493, 287.493, 287.493, 287.493, 
    287.4931, 287.4931, 287.4931, 287.4931, 287.4931, 287.4932, 287.4932, 
    287.4932, 287.4932, 287.4932, 287.4933, 287.4933, 287.4933, 287.4933, 
    287.4933, 287.4934, 287.4934, 287.4934, 287.4934, 287.4935, 287.4935, 
    287.4935, 287.4936, 287.4936, 287.4936, 287.4936, 287.4937, 287.4937, 
    287.4937, 287.4937, 287.4938,
  288.4186, 288.4185, 288.4185, 288.4185, 288.4185, 288.4184, 288.4184, 
    288.4184, 288.4184, 288.4183, 288.4183, 288.4183, 288.4182, 288.4182, 
    288.4182, 288.4182, 288.4182, 288.4181, 288.4181, 288.4181, 288.4181, 
    288.418, 288.418, 288.418, 288.418, 288.4179, 288.4179, 288.4179, 
    288.4179, 288.4179, 288.4178, 288.4178, 288.4178, 288.4178, 288.4178, 
    288.4178, 288.4178, 288.4178, 288.4178, 288.4178, 288.4177, 288.4177, 
    288.4177, 288.4177, 288.4177, 288.4177, 288.4177, 288.4177, 288.4177, 
    288.4177, 288.4177, 288.4177, 288.4177, 288.4177, 288.4177, 288.4177, 
    288.4178, 288.4178, 288.4178, 288.4178, 288.4178, 288.4178, 288.4178, 
    288.4178, 288.4178, 288.4178, 288.4179, 288.4179, 288.4179, 288.4179, 
    288.4179, 288.418, 288.418, 288.418, 288.418, 288.4181, 288.4181, 
    288.4181, 288.4181, 288.4182, 288.4182, 288.4182, 288.4182, 288.4182, 
    288.4183, 288.4183, 288.4183, 288.4184, 288.4184, 288.4184, 288.4184, 
    288.4185, 288.4185, 288.4185, 288.4185, 288.4186,
  289.3364, 289.3364, 289.3363, 289.3363, 289.3363, 289.3362, 289.3362, 
    289.3362, 289.3362, 289.3362, 289.3361, 289.3361, 289.3361, 289.336, 
    289.336, 289.336, 289.336, 289.3359, 289.3359, 289.3359, 289.3359, 
    289.3358, 289.3358, 289.3358, 289.3358, 289.3358, 289.3357, 289.3357, 
    289.3357, 289.3357, 289.3357, 289.3356, 289.3356, 289.3356, 289.3356, 
    289.3356, 289.3356, 289.3356, 289.3356, 289.3355, 289.3355, 289.3355, 
    289.3355, 289.3355, 289.3355, 289.3355, 289.3355, 289.3355, 289.3355, 
    289.3355, 289.3355, 289.3355, 289.3355, 289.3355, 289.3355, 289.3355, 
    289.3355, 289.3356, 289.3356, 289.3356, 289.3356, 289.3356, 289.3356, 
    289.3356, 289.3356, 289.3357, 289.3357, 289.3357, 289.3357, 289.3357, 
    289.3358, 289.3358, 289.3358, 289.3358, 289.3358, 289.3359, 289.3359, 
    289.3359, 289.3359, 289.336, 289.336, 289.336, 289.336, 289.3361, 
    289.3361, 289.3361, 289.3362, 289.3362, 289.3362, 289.3362, 289.3362, 
    289.3363, 289.3363, 289.3363, 289.3364, 289.3364,
  290.2471, 290.2471, 290.2471, 290.247, 290.247, 290.247, 290.2469, 
    290.2469, 290.2469, 290.2469, 290.2469, 290.2468, 290.2468, 290.2468, 
    290.2467, 290.2467, 290.2467, 290.2467, 290.2466, 290.2466, 290.2466, 
    290.2466, 290.2466, 290.2465, 290.2465, 290.2465, 290.2465, 290.2464, 
    290.2464, 290.2464, 290.2464, 290.2464, 290.2464, 290.2463, 290.2463, 
    290.2463, 290.2463, 290.2463, 290.2463, 290.2463, 290.2463, 290.2462, 
    290.2462, 290.2462, 290.2462, 290.2462, 290.2462, 290.2462, 290.2462, 
    290.2462, 290.2462, 290.2462, 290.2462, 290.2462, 290.2462, 290.2463, 
    290.2463, 290.2463, 290.2463, 290.2463, 290.2463, 290.2463, 290.2463, 
    290.2464, 290.2464, 290.2464, 290.2464, 290.2464, 290.2464, 290.2465, 
    290.2465, 290.2465, 290.2465, 290.2466, 290.2466, 290.2466, 290.2466, 
    290.2466, 290.2467, 290.2467, 290.2467, 290.2467, 290.2468, 290.2468, 
    290.2468, 290.2469, 290.2469, 290.2469, 290.2469, 290.2469, 290.247, 
    290.247, 290.247, 290.2471, 290.2471, 290.2471,
  291.1507, 291.1507, 291.1506, 291.1506, 291.1506, 291.1505, 291.1505, 
    291.1505, 291.1505, 291.1505, 291.1504, 291.1504, 291.1504, 291.1503, 
    291.1503, 291.1503, 291.1503, 291.1502, 291.1502, 291.1502, 291.1501, 
    291.1501, 291.1501, 291.1501, 291.1501, 291.1501, 291.15, 291.15, 291.15, 
    291.15, 291.15, 291.1499, 291.1499, 291.1499, 291.1499, 291.1499, 
    291.1499, 291.1499, 291.1498, 291.1498, 291.1498, 291.1498, 291.1498, 
    291.1498, 291.1498, 291.1498, 291.1498, 291.1498, 291.1498, 291.1498, 
    291.1498, 291.1498, 291.1498, 291.1498, 291.1498, 291.1498, 291.1498, 
    291.1498, 291.1499, 291.1499, 291.1499, 291.1499, 291.1499, 291.1499, 
    291.1499, 291.15, 291.15, 291.15, 291.15, 291.15, 291.1501, 291.1501, 
    291.1501, 291.1501, 291.1501, 291.1501, 291.1502, 291.1502, 291.1502, 
    291.1503, 291.1503, 291.1503, 291.1503, 291.1504, 291.1504, 291.1504, 
    291.1505, 291.1505, 291.1505, 291.1505, 291.1505, 291.1506, 291.1506, 
    291.1506, 291.1507, 291.1507,
  292.0471, 292.047, 292.047, 292.047, 292.0469, 292.0469, 292.0469, 
    292.0468, 292.0468, 292.0468, 292.0468, 292.0468, 292.0467, 292.0467, 
    292.0467, 292.0466, 292.0466, 292.0466, 292.0466, 292.0465, 292.0465, 
    292.0465, 292.0464, 292.0464, 292.0464, 292.0464, 292.0464, 292.0464, 
    292.0463, 292.0463, 292.0463, 292.0463, 292.0463, 292.0463, 292.0462, 
    292.0462, 292.0462, 292.0462, 292.0462, 292.0462, 292.0462, 292.0462, 
    292.0462, 292.0462, 292.0462, 292.0461, 292.0461, 292.0461, 292.0461, 
    292.0461, 292.0461, 292.0462, 292.0462, 292.0462, 292.0462, 292.0462, 
    292.0462, 292.0462, 292.0462, 292.0462, 292.0462, 292.0462, 292.0463, 
    292.0463, 292.0463, 292.0463, 292.0463, 292.0463, 292.0464, 292.0464, 
    292.0464, 292.0464, 292.0464, 292.0464, 292.0465, 292.0465, 292.0465, 
    292.0466, 292.0466, 292.0466, 292.0466, 292.0467, 292.0467, 292.0467, 
    292.0468, 292.0468, 292.0468, 292.0468, 292.0468, 292.0469, 292.0469, 
    292.0469, 292.047, 292.047, 292.047, 292.0471,
  292.9361, 292.9361, 292.9361, 292.936, 292.936, 292.936, 292.9359, 
    292.9359, 292.9359, 292.9359, 292.9358, 292.9358, 292.9358, 292.9358, 
    292.9357, 292.9357, 292.9357, 292.9356, 292.9356, 292.9356, 292.9356, 
    292.9355, 292.9355, 292.9355, 292.9355, 292.9355, 292.9355, 292.9354, 
    292.9354, 292.9354, 292.9354, 292.9354, 292.9353, 292.9353, 292.9353, 
    292.9353, 292.9353, 292.9353, 292.9353, 292.9353, 292.9352, 292.9352, 
    292.9352, 292.9352, 292.9352, 292.9352, 292.9352, 292.9352, 292.9352, 
    292.9352, 292.9352, 292.9352, 292.9352, 292.9352, 292.9352, 292.9352, 
    292.9353, 292.9353, 292.9353, 292.9353, 292.9353, 292.9353, 292.9353, 
    292.9353, 292.9354, 292.9354, 292.9354, 292.9354, 292.9354, 292.9355, 
    292.9355, 292.9355, 292.9355, 292.9355, 292.9355, 292.9356, 292.9356, 
    292.9356, 292.9356, 292.9357, 292.9357, 292.9357, 292.9358, 292.9358, 
    292.9358, 292.9358, 292.9359, 292.9359, 292.9359, 292.9359, 292.936, 
    292.936, 292.936, 292.9361, 292.9361, 292.9361,
  293.8179, 293.8178, 293.8178, 293.8178, 293.8177, 293.8177, 293.8177, 
    293.8177, 293.8176, 293.8176, 293.8176, 293.8176, 293.8175, 293.8175, 
    293.8175, 293.8174, 293.8174, 293.8174, 293.8174, 293.8174, 293.8173, 
    293.8173, 293.8173, 293.8173, 293.8172, 293.8172, 293.8172, 293.8172, 
    293.8171, 293.8171, 293.8171, 293.8171, 293.8171, 293.8171, 293.817, 
    293.817, 293.817, 293.817, 293.817, 293.817, 293.817, 293.817, 293.817, 
    293.817, 293.817, 293.817, 293.817, 293.817, 293.817, 293.817, 293.817, 
    293.817, 293.817, 293.817, 293.817, 293.817, 293.817, 293.817, 293.817, 
    293.817, 293.817, 293.817, 293.8171, 293.8171, 293.8171, 293.8171, 
    293.8171, 293.8171, 293.8172, 293.8172, 293.8172, 293.8172, 293.8173, 
    293.8173, 293.8173, 293.8173, 293.8174, 293.8174, 293.8174, 293.8174, 
    293.8174, 293.8175, 293.8175, 293.8175, 293.8176, 293.8176, 293.8176, 
    293.8176, 293.8177, 293.8177, 293.8177, 293.8177, 293.8178, 293.8178, 
    293.8178, 293.8179,
  294.6923, 294.6922, 294.6922, 294.6922, 294.6921, 294.6921, 294.6921, 
    294.692, 294.692, 294.692, 294.692, 294.6919, 294.6919, 294.6919, 
    294.6919, 294.6918, 294.6918, 294.6918, 294.6917, 294.6917, 294.6917, 
    294.6917, 294.6917, 294.6916, 294.6916, 294.6916, 294.6916, 294.6916, 
    294.6915, 294.6915, 294.6915, 294.6915, 294.6915, 294.6914, 294.6914, 
    294.6914, 294.6914, 294.6914, 294.6914, 294.6914, 294.6914, 294.6914, 
    294.6914, 294.6913, 294.6913, 294.6913, 294.6913, 294.6913, 294.6913, 
    294.6913, 294.6913, 294.6913, 294.6913, 294.6914, 294.6914, 294.6914, 
    294.6914, 294.6914, 294.6914, 294.6914, 294.6914, 294.6914, 294.6914, 
    294.6915, 294.6915, 294.6915, 294.6915, 294.6915, 294.6916, 294.6916, 
    294.6916, 294.6916, 294.6916, 294.6917, 294.6917, 294.6917, 294.6917, 
    294.6917, 294.6918, 294.6918, 294.6918, 294.6919, 294.6919, 294.6919, 
    294.6919, 294.692, 294.692, 294.692, 294.692, 294.6921, 294.6921, 
    294.6921, 294.6922, 294.6922, 294.6922, 294.6923,
  295.5593, 295.5592, 295.5592, 295.5592, 295.5591, 295.5591, 295.5591, 
    295.5591, 295.559, 295.559, 295.559, 295.5589, 295.5589, 295.5589, 
    295.5588, 295.5588, 295.5588, 295.5588, 295.5587, 295.5587, 295.5587, 
    295.5587, 295.5587, 295.5586, 295.5586, 295.5586, 295.5586, 295.5585, 
    295.5585, 295.5585, 295.5585, 295.5585, 295.5585, 295.5584, 295.5584, 
    295.5584, 295.5584, 295.5584, 295.5584, 295.5584, 295.5584, 295.5583, 
    295.5583, 295.5583, 295.5583, 295.5583, 295.5583, 295.5583, 295.5583, 
    295.5583, 295.5583, 295.5583, 295.5583, 295.5583, 295.5583, 295.5584, 
    295.5584, 295.5584, 295.5584, 295.5584, 295.5584, 295.5584, 295.5584, 
    295.5585, 295.5585, 295.5585, 295.5585, 295.5585, 295.5585, 295.5586, 
    295.5586, 295.5586, 295.5586, 295.5587, 295.5587, 295.5587, 295.5587, 
    295.5587, 295.5588, 295.5588, 295.5588, 295.5588, 295.5589, 295.5589, 
    295.5589, 295.559, 295.559, 295.559, 295.5591, 295.5591, 295.5591, 
    295.5591, 295.5592, 295.5592, 295.5592, 295.5593,
  296.4189, 296.4188, 296.4188, 296.4188, 296.4187, 296.4187, 296.4187, 
    296.4186, 296.4186, 296.4186, 296.4185, 296.4185, 296.4185, 296.4185, 
    296.4184, 296.4184, 296.4184, 296.4184, 296.4183, 296.4183, 296.4183, 
    296.4183, 296.4182, 296.4182, 296.4182, 296.4182, 296.4182, 296.4181, 
    296.4181, 296.4181, 296.4181, 296.4181, 296.4181, 296.418, 296.418, 
    296.418, 296.418, 296.418, 296.418, 296.418, 296.418, 296.418, 296.4179, 
    296.4179, 296.4179, 296.4179, 296.4179, 296.4179, 296.4179, 296.4179, 
    296.4179, 296.4179, 296.4179, 296.4179, 296.418, 296.418, 296.418, 
    296.418, 296.418, 296.418, 296.418, 296.418, 296.418, 296.4181, 296.4181, 
    296.4181, 296.4181, 296.4181, 296.4181, 296.4182, 296.4182, 296.4182, 
    296.4182, 296.4182, 296.4183, 296.4183, 296.4183, 296.4183, 296.4184, 
    296.4184, 296.4184, 296.4184, 296.4185, 296.4185, 296.4185, 296.4185, 
    296.4186, 296.4186, 296.4186, 296.4187, 296.4187, 296.4187, 296.4188, 
    296.4188, 296.4188, 296.4189,
  297.271, 297.271, 297.271, 297.2709, 297.2709, 297.2709, 297.2708, 
    297.2708, 297.2708, 297.2708, 297.2707, 297.2707, 297.2707, 297.2706, 
    297.2706, 297.2706, 297.2706, 297.2705, 297.2705, 297.2705, 297.2705, 
    297.2704, 297.2704, 297.2704, 297.2704, 297.2704, 297.2703, 297.2703, 
    297.2703, 297.2703, 297.2703, 297.2702, 297.2702, 297.2702, 297.2702, 
    297.2702, 297.2702, 297.2702, 297.2702, 297.2701, 297.2701, 297.2701, 
    297.2701, 297.2701, 297.2701, 297.2701, 297.2701, 297.2701, 297.2701, 
    297.2701, 297.2701, 297.2701, 297.2701, 297.2701, 297.2701, 297.2701, 
    297.2701, 297.2702, 297.2702, 297.2702, 297.2702, 297.2702, 297.2702, 
    297.2702, 297.2702, 297.2703, 297.2703, 297.2703, 297.2703, 297.2703, 
    297.2704, 297.2704, 297.2704, 297.2704, 297.2704, 297.2705, 297.2705, 
    297.2705, 297.2705, 297.2706, 297.2706, 297.2706, 297.2706, 297.2707, 
    297.2707, 297.2707, 297.2708, 297.2708, 297.2708, 297.2708, 297.2709, 
    297.2709, 297.2709, 297.271, 297.271, 297.271,
  298.1158, 298.1158, 298.1157, 298.1157, 298.1157, 298.1156, 298.1156, 
    298.1156, 298.1155, 298.1155, 298.1155, 298.1154, 298.1154, 298.1154, 
    298.1154, 298.1154, 298.1153, 298.1153, 298.1153, 298.1153, 298.1152, 
    298.1152, 298.1152, 298.1151, 298.1151, 298.1151, 298.1151, 298.1151, 
    298.1151, 298.1151, 298.115, 298.115, 298.115, 298.115, 298.115, 298.115, 
    298.1149, 298.1149, 298.1149, 298.1149, 298.1149, 298.1149, 298.1149, 
    298.1149, 298.1149, 298.1149, 298.1149, 298.1149, 298.1149, 298.1149, 
    298.1149, 298.1149, 298.1149, 298.1149, 298.1149, 298.1149, 298.1149, 
    298.1149, 298.1149, 298.1149, 298.115, 298.115, 298.115, 298.115, 
    298.115, 298.115, 298.1151, 298.1151, 298.1151, 298.1151, 298.1151, 
    298.1151, 298.1151, 298.1152, 298.1152, 298.1152, 298.1153, 298.1153, 
    298.1153, 298.1153, 298.1154, 298.1154, 298.1154, 298.1154, 298.1154, 
    298.1155, 298.1155, 298.1155, 298.1156, 298.1156, 298.1156, 298.1157, 
    298.1157, 298.1157, 298.1158, 298.1158,
  298.9532, 298.9531, 298.9531, 298.9531, 298.953, 298.953, 298.953, 
    298.9529, 298.9529, 298.9529, 298.9529, 298.9528, 298.9528, 298.9528, 
    298.9527, 298.9527, 298.9527, 298.9527, 298.9526, 298.9526, 298.9526, 
    298.9525, 298.9525, 298.9525, 298.9525, 298.9525, 298.9525, 298.9524, 
    298.9524, 298.9524, 298.9524, 298.9524, 298.9524, 298.9523, 298.9523, 
    298.9523, 298.9523, 298.9523, 298.9523, 298.9523, 298.9523, 298.9523, 
    298.9522, 298.9522, 298.9522, 298.9522, 298.9522, 298.9522, 298.9522, 
    298.9522, 298.9522, 298.9522, 298.9522, 298.9522, 298.9523, 298.9523, 
    298.9523, 298.9523, 298.9523, 298.9523, 298.9523, 298.9523, 298.9523, 
    298.9524, 298.9524, 298.9524, 298.9524, 298.9524, 298.9524, 298.9525, 
    298.9525, 298.9525, 298.9525, 298.9525, 298.9525, 298.9526, 298.9526, 
    298.9526, 298.9527, 298.9527, 298.9527, 298.9527, 298.9528, 298.9528, 
    298.9528, 298.9529, 298.9529, 298.9529, 298.9529, 298.953, 298.953, 
    298.953, 298.9531, 298.9531, 298.9531, 298.9532,
  299.7831, 299.7831, 299.7831, 299.783, 299.783, 299.783, 299.7829, 
    299.7829, 299.7829, 299.7828, 299.7828, 299.7828, 299.7827, 299.7827, 
    299.7827, 299.7827, 299.7827, 299.7826, 299.7826, 299.7826, 299.7826, 
    299.7825, 299.7825, 299.7825, 299.7825, 299.7824, 299.7824, 299.7824, 
    299.7824, 299.7824, 299.7823, 299.7823, 299.7823, 299.7823, 299.7823, 
    299.7823, 299.7823, 299.7823, 299.7823, 299.7823, 299.7822, 299.7822, 
    299.7822, 299.7822, 299.7822, 299.7822, 299.7822, 299.7822, 299.7822, 
    299.7822, 299.7822, 299.7822, 299.7822, 299.7822, 299.7822, 299.7822, 
    299.7823, 299.7823, 299.7823, 299.7823, 299.7823, 299.7823, 299.7823, 
    299.7823, 299.7823, 299.7823, 299.7824, 299.7824, 299.7824, 299.7824, 
    299.7824, 299.7825, 299.7825, 299.7825, 299.7825, 299.7826, 299.7826, 
    299.7826, 299.7826, 299.7827, 299.7827, 299.7827, 299.7827, 299.7827, 
    299.7828, 299.7828, 299.7828, 299.7829, 299.7829, 299.7829, 299.783, 
    299.783, 299.783, 299.7831, 299.7831, 299.7831,
  300.6057, 300.6057, 300.6057, 300.6056, 300.6056, 300.6056, 300.6055, 
    300.6055, 300.6055, 300.6054, 300.6054, 300.6054, 300.6053, 300.6053, 
    300.6053, 300.6053, 300.6053, 300.6052, 300.6052, 300.6052, 300.6052, 
    300.6051, 300.6051, 300.6051, 300.6051, 300.605, 300.605, 300.605, 
    300.605, 300.605, 300.6049, 300.6049, 300.6049, 300.6049, 300.6049, 
    300.6049, 300.6049, 300.6049, 300.6049, 300.6049, 300.6048, 300.6048, 
    300.6048, 300.6048, 300.6048, 300.6048, 300.6048, 300.6048, 300.6048, 
    300.6048, 300.6048, 300.6048, 300.6048, 300.6048, 300.6048, 300.6048, 
    300.6049, 300.6049, 300.6049, 300.6049, 300.6049, 300.6049, 300.6049, 
    300.6049, 300.6049, 300.6049, 300.605, 300.605, 300.605, 300.605, 
    300.605, 300.6051, 300.6051, 300.6051, 300.6051, 300.6052, 300.6052, 
    300.6052, 300.6052, 300.6053, 300.6053, 300.6053, 300.6053, 300.6053, 
    300.6054, 300.6054, 300.6054, 300.6055, 300.6055, 300.6055, 300.6056, 
    300.6056, 300.6056, 300.6057, 300.6057, 300.6057,
  301.421, 301.421, 301.4209, 301.4209, 301.4209, 301.4208, 301.4208, 
    301.4208, 301.4207, 301.4207, 301.4207, 301.4207, 301.4206, 301.4206, 
    301.4206, 301.4205, 301.4205, 301.4205, 301.4205, 301.4204, 301.4204, 
    301.4204, 301.4204, 301.4203, 301.4203, 301.4203, 301.4203, 301.4203, 
    301.4203, 301.4202, 301.4202, 301.4202, 301.4202, 301.4202, 301.4202, 
    301.4202, 301.4201, 301.4201, 301.4201, 301.4201, 301.4201, 301.4201, 
    301.4201, 301.4201, 301.4201, 301.4201, 301.4201, 301.4201, 301.4201, 
    301.4201, 301.4201, 301.4201, 301.4201, 301.4201, 301.4201, 301.4201, 
    301.4201, 301.4201, 301.4201, 301.4201, 301.4202, 301.4202, 301.4202, 
    301.4202, 301.4202, 301.4202, 301.4202, 301.4203, 301.4203, 301.4203, 
    301.4203, 301.4203, 301.4203, 301.4204, 301.4204, 301.4204, 301.4204, 
    301.4205, 301.4205, 301.4205, 301.4205, 301.4206, 301.4206, 301.4206, 
    301.4207, 301.4207, 301.4207, 301.4207, 301.4208, 301.4208, 301.4208, 
    301.4209, 301.4209, 301.4209, 301.421, 301.421,
  302.2289, 302.2289, 302.2289, 302.2289, 302.2288, 302.2288, 302.2288, 
    302.2287, 302.2287, 302.2287, 302.2286, 302.2286, 302.2286, 302.2285, 
    302.2285, 302.2285, 302.2285, 302.2285, 302.2284, 302.2284, 302.2284, 
    302.2284, 302.2283, 302.2283, 302.2283, 302.2283, 302.2283, 302.2282, 
    302.2282, 302.2282, 302.2282, 302.2282, 302.2281, 302.2281, 302.2281, 
    302.2281, 302.2281, 302.2281, 302.2281, 302.2281, 302.2281, 302.2281, 
    302.2281, 302.2281, 302.2281, 302.2281, 302.2281, 302.2281, 302.2281, 
    302.2281, 302.2281, 302.2281, 302.2281, 302.2281, 302.2281, 302.2281, 
    302.2281, 302.2281, 302.2281, 302.2281, 302.2281, 302.2281, 302.2281, 
    302.2281, 302.2282, 302.2282, 302.2282, 302.2282, 302.2282, 302.2283, 
    302.2283, 302.2283, 302.2283, 302.2283, 302.2284, 302.2284, 302.2284, 
    302.2284, 302.2285, 302.2285, 302.2285, 302.2285, 302.2285, 302.2286, 
    302.2286, 302.2286, 302.2287, 302.2287, 302.2287, 302.2288, 302.2288, 
    302.2288, 302.2289, 302.2289, 302.2289, 302.2289,
  303.0296, 303.0296, 303.0296, 303.0295, 303.0295, 303.0295, 303.0294, 
    303.0294, 303.0294, 303.0294, 303.0294, 303.0293, 303.0293, 303.0293, 
    303.0292, 303.0292, 303.0292, 303.0291, 303.0291, 303.0291, 303.0291, 
    303.0291, 303.0291, 303.029, 303.029, 303.029, 303.029, 303.029, 
    303.0289, 303.0289, 303.0289, 303.0289, 303.0289, 303.0289, 303.0288, 
    303.0288, 303.0288, 303.0288, 303.0288, 303.0288, 303.0288, 303.0288, 
    303.0288, 303.0288, 303.0288, 303.0288, 303.0287, 303.0287, 303.0287, 
    303.0287, 303.0288, 303.0288, 303.0288, 303.0288, 303.0288, 303.0288, 
    303.0288, 303.0288, 303.0288, 303.0288, 303.0288, 303.0288, 303.0289, 
    303.0289, 303.0289, 303.0289, 303.0289, 303.0289, 303.029, 303.029, 
    303.029, 303.029, 303.029, 303.0291, 303.0291, 303.0291, 303.0291, 
    303.0291, 303.0291, 303.0292, 303.0292, 303.0292, 303.0293, 303.0293, 
    303.0293, 303.0294, 303.0294, 303.0294, 303.0294, 303.0294, 303.0295, 
    303.0295, 303.0295, 303.0296, 303.0296, 303.0296,
  303.8232, 303.8231, 303.8231, 303.8231, 303.823, 303.823, 303.823, 
    303.8229, 303.8229, 303.8229, 303.8228, 303.8228, 303.8228, 303.8228, 
    303.8227, 303.8227, 303.8227, 303.8227, 303.8226, 303.8226, 303.8226, 
    303.8226, 303.8225, 303.8225, 303.8225, 303.8225, 303.8224, 303.8224, 
    303.8224, 303.8224, 303.8224, 303.8224, 303.8224, 303.8224, 303.8224, 
    303.8223, 303.8223, 303.8223, 303.8223, 303.8223, 303.8223, 303.8223, 
    303.8223, 303.8223, 303.8223, 303.8223, 303.8223, 303.8223, 303.8223, 
    303.8223, 303.8223, 303.8223, 303.8223, 303.8223, 303.8223, 303.8223, 
    303.8223, 303.8223, 303.8223, 303.8223, 303.8223, 303.8224, 303.8224, 
    303.8224, 303.8224, 303.8224, 303.8224, 303.8224, 303.8224, 303.8224, 
    303.8225, 303.8225, 303.8225, 303.8225, 303.8226, 303.8226, 303.8226, 
    303.8226, 303.8227, 303.8227, 303.8227, 303.8227, 303.8228, 303.8228, 
    303.8228, 303.8228, 303.8229, 303.8229, 303.8229, 303.823, 303.823, 
    303.823, 303.8231, 303.8231, 303.8231, 303.8232,
  304.6095, 304.6094, 304.6094, 304.6094, 304.6093, 304.6093, 304.6093, 
    304.6093, 304.6092, 304.6092, 304.6092, 304.6092, 304.6091, 304.6091, 
    304.6091, 304.609, 304.609, 304.609, 304.609, 304.6089, 304.6089, 
    304.6089, 304.6089, 304.6089, 304.6089, 304.6088, 304.6088, 304.6088, 
    304.6088, 304.6088, 304.6087, 304.6087, 304.6087, 304.6087, 304.6087, 
    304.6087, 304.6087, 304.6086, 304.6086, 304.6086, 304.6086, 304.6086, 
    304.6086, 304.6086, 304.6086, 304.6086, 304.6086, 304.6086, 304.6086, 
    304.6086, 304.6086, 304.6086, 304.6086, 304.6086, 304.6086, 304.6086, 
    304.6086, 304.6086, 304.6086, 304.6087, 304.6087, 304.6087, 304.6087, 
    304.6087, 304.6087, 304.6087, 304.6088, 304.6088, 304.6088, 304.6088, 
    304.6088, 304.6089, 304.6089, 304.6089, 304.6089, 304.6089, 304.6089, 
    304.609, 304.609, 304.609, 304.609, 304.6091, 304.6091, 304.6091, 
    304.6092, 304.6092, 304.6092, 304.6092, 304.6093, 304.6093, 304.6093, 
    304.6093, 304.6094, 304.6094, 304.6094, 304.6095 ;

 grid_latt =
  35.07925, 34.34282, 33.60628, 32.86962, 32.13284, 31.39594, 30.65893, 
    29.92181, 29.18457, 28.44723, 27.70978, 26.97222, 26.23456, 25.4968, 
    24.75893, 24.02097, 23.28291, 22.54476, 21.80651, 21.06818, 20.32976, 
    19.59126, 18.85267, 18.114, 17.37526, 16.63645, 15.89756, 15.15861, 
    14.41959, 13.6805, 12.94136, 12.20216, 11.46291, 10.72361, 9.984256, 
    9.244861, 8.505425, 7.765951, 7.026442, 6.286901, 5.547333, 4.807739, 
    4.068124, 3.32849, 2.588841, 1.849181, 1.109512, 0.3698378, -0.3698378, 
    -1.109512, -1.849181, -2.588841, -3.32849, -4.068124, -4.807739, 
    -5.547333, -6.286901, -7.026442, -7.765951, -8.505425, -9.244861, 
    -9.984256, -10.72361, -11.46291, -12.20216, -12.94136, -13.6805, 
    -14.41959, -15.15861, -15.89756, -16.63645, -17.37526, -18.114, 
    -18.85267, -19.59126, -20.32976, -21.06818, -21.80651, -22.54476, 
    -23.28291, -24.02097, -24.75893, -25.4968, -26.23456, -26.97222, 
    -27.70978, -28.44723, -29.18457, -29.92181, -30.65893, -31.39594, 
    -32.13284, -32.86962, -33.60628, -34.34282, -35.07925,
  35.43988, 34.70005, 33.95987, 33.21932, 32.47842, 31.73718, 30.9956, 
    30.25368, 29.51142, 28.76883, 28.02592, 27.28269, 26.53915, 25.7953, 
    25.05115, 24.3067, 23.56197, 22.81695, 22.07165, 21.32609, 20.58027, 
    19.83419, 19.08786, 18.3413, 17.59451, 16.84749, 16.10026, 15.35282, 
    14.60518, 13.85736, 13.10935, 12.36118, 11.61284, 10.86435, 10.11571, 
    9.366945, 8.618052, 7.869044, 7.119931, 6.370722, 5.621428, 4.872057, 
    4.122622, 3.37313, 2.623593, 1.87402, 1.124422, 0.3748092, -0.3748092, 
    -1.124422, -1.87402, -2.623593, -3.37313, -4.122622, -4.872057, 
    -5.621428, -6.370722, -7.119931, -7.869044, -8.618052, -9.366945, 
    -10.11571, -10.86435, -11.61284, -12.36118, -13.10935, -13.85736, 
    -14.60518, -15.35282, -16.10026, -16.84749, -17.59451, -18.3413, 
    -19.08786, -19.83419, -20.58027, -21.32609, -22.07165, -22.81695, 
    -23.56197, -24.3067, -25.05115, -25.7953, -26.53915, -27.28269, 
    -28.02592, -28.76883, -29.51142, -30.25368, -30.9956, -31.73718, 
    -32.47842, -33.21932, -33.95987, -34.70005, -35.43988,
  35.79544, 35.05236, 34.30869, 33.56442, 32.81957, 32.07414, 31.32814, 
    30.58158, 29.83445, 29.08677, 28.33856, 27.58981, 26.84053, 26.09074, 
    25.34044, 24.58965, 23.83837, 23.08662, 22.33441, 21.58174, 20.82863, 
    20.0751, 19.32115, 18.5668, 17.81206, 17.05695, 16.30147, 15.54564, 
    14.78949, 14.03301, 13.27623, 12.51916, 11.76182, 11.00421, 10.24637, 
    9.488298, 8.730017, 7.971541, 7.212887, 6.454072, 5.695111, 4.936023, 
    4.176824, 3.41753, 2.658159, 1.898728, 1.139254, 0.3797542, -0.3797542, 
    -1.139254, -1.898728, -2.658159, -3.41753, -4.176824, -4.936023, 
    -5.695111, -6.454072, -7.212887, -7.971541, -8.730017, -9.488298, 
    -10.24637, -11.00421, -11.76182, -12.51916, -13.27623, -14.03301, 
    -14.78949, -15.54564, -16.30147, -17.05695, -17.81206, -18.5668, 
    -19.32115, -20.0751, -20.82863, -21.58174, -22.33441, -23.08662, 
    -23.83837, -24.58965, -25.34044, -26.09074, -26.84053, -27.58981, 
    -28.33856, -29.08677, -29.83445, -30.58158, -31.32814, -32.07414, 
    -32.81957, -33.56442, -34.30869, -35.05236, -35.79544,
  36.14578, 35.39962, 34.65261, 33.90479, 33.15614, 32.40669, 31.65643, 
    30.90537, 30.15354, 29.40093, 28.64755, 27.89343, 27.13857, 26.38298, 
    25.62668, 24.86968, 24.112, 23.35365, 22.59464, 21.835, 21.07474, 
    20.31387, 19.55242, 18.79039, 18.02782, 17.26471, 16.50109, 15.73699, 
    14.9724, 14.20737, 13.4419, 12.67602, 11.90976, 11.14313, 10.37615, 
    9.608856, 8.84126, 8.073387, 7.305261, 6.536906, 5.768345, 4.999602, 
    4.230701, 3.461666, 2.692521, 1.92329, 1.153999, 0.3846703, -0.3846703, 
    -1.153999, -1.92329, -2.692521, -3.461666, -4.230701, -4.999602, 
    -5.768345, -6.536906, -7.305261, -8.073387, -8.84126, -9.608856, 
    -10.37615, -11.14313, -11.90976, -12.67602, -13.4419, -14.20737, 
    -14.9724, -15.73699, -16.50109, -17.26471, -18.02782, -18.79039, 
    -19.55242, -20.31387, -21.07474, -21.835, -22.59464, -23.35365, -24.112, 
    -24.86968, -25.62668, -26.38298, -27.13857, -27.89343, -28.64755, 
    -29.40093, -30.15354, -30.90537, -31.65643, -32.40669, -33.15614, 
    -33.90479, -34.65261, -35.39962, -36.14578,
  36.4908, 35.7417, 34.99154, 34.2403, 33.48802, 32.73469, 31.98032, 
    31.22494, 30.46854, 29.71115, 28.95277, 28.19342, 27.43312, 26.67189, 
    25.90973, 25.14667, 24.38272, 23.6179, 22.85224, 22.08575, 21.31846, 
    20.55038, 19.78154, 19.01196, 18.24167, 17.47068, 16.69903, 15.92674, 
    15.15383, 14.38034, 13.60628, 12.83169, 12.05659, 11.28102, 10.505, 
    9.728554, 8.951721, 8.174527, 7.397004, 6.619181, 5.84109, 5.06276, 
    4.284225, 3.505514, 2.72666, 1.947694, 1.168648, 0.3895547, -0.3895547, 
    -1.168648, -1.947694, -2.72666, -3.505514, -4.284225, -5.06276, -5.84109, 
    -6.619181, -7.397004, -8.174527, -8.951721, -9.728554, -10.505, 
    -11.28102, -12.05659, -12.83169, -13.60628, -14.38034, -15.15383, 
    -15.92674, -16.69903, -17.47068, -18.24167, -19.01196, -19.78154, 
    -20.55038, -21.31846, -22.08575, -22.85224, -23.6179, -24.38272, 
    -25.14667, -25.90973, -26.67189, -27.43312, -28.19342, -28.95277, 
    -29.71115, -30.46854, -31.22494, -31.98032, -32.73469, -33.48802, 
    -34.2403, -34.99154, -35.7417, -36.4908,
  36.83038, 36.0785, 35.32531, 34.57083, 33.81506, 33.05801, 32.29969, 
    31.54013, 30.77932, 30.0173, 29.25407, 28.48965, 27.72406, 26.95732, 
    26.18944, 25.42046, 24.65038, 23.87924, 23.10706, 22.33386, 21.55966, 
    20.7845, 20.0084, 19.23139, 18.45349, 17.67474, 16.89517, 16.11481, 
    15.33368, 14.55183, 13.76928, 12.98607, 12.20224, 11.41781, 10.63283, 
    9.847324, 9.061338, 8.274905, 7.488063, 6.70085, 5.913303, 5.125462, 
    4.337364, 3.549049, 2.760556, 1.971925, 1.183195, 0.3944048, -0.3944048, 
    -1.183195, -1.971925, -2.760556, -3.549049, -4.337364, -5.125462, 
    -5.913303, -6.70085, -7.488063, -8.274905, -9.061338, -9.847324, 
    -10.63283, -11.41781, -12.20224, -12.98607, -13.76928, -14.55183, 
    -15.33368, -16.11481, -16.89517, -17.67474, -18.45349, -19.23139, 
    -20.0084, -20.7845, -21.55966, -22.33386, -23.10706, -23.87924, 
    -24.65038, -25.42046, -26.18944, -26.95732, -27.72406, -28.48965, 
    -29.25407, -30.0173, -30.77932, -31.54013, -32.29969, -33.05801, 
    -33.81506, -34.57083, -35.32531, -36.0785, -36.83038,
  37.1644, 36.40988, 35.65382, 34.89624, 34.13713, 33.37651, 32.6144, 
    31.8508, 31.08575, 30.31924, 29.55131, 28.78197, 28.01123, 27.23913, 
    26.46569, 25.69092, 24.91487, 24.13754, 23.35897, 22.57919, 21.79822, 
    21.01611, 20.23287, 19.44855, 18.66317, 17.87678, 17.0894, 16.30107, 
    15.51184, 14.72173, 13.9308, 13.13908, 12.3466, 11.55342, 10.75957, 
    9.965097, 9.170046, 8.37446, 7.578384, 6.781863, 5.984942, 5.187668, 
    4.390087, 3.592245, 2.79419, 1.995969, 1.197629, 0.3992176, -0.3992176, 
    -1.197629, -1.995969, -2.79419, -3.592245, -4.390087, -5.187668, 
    -5.984942, -6.781863, -7.578384, -8.37446, -9.170046, -9.965097, 
    -10.75957, -11.55342, -12.3466, -13.13908, -13.9308, -14.72173, 
    -15.51184, -16.30107, -17.0894, -17.87678, -18.66317, -19.44855, 
    -20.23287, -21.01611, -21.79822, -22.57919, -23.35897, -24.13754, 
    -24.91487, -25.69092, -26.46569, -27.23913, -28.01123, -28.78197, 
    -29.55131, -30.31924, -31.08575, -31.8508, -32.6144, -33.37651, 
    -34.13713, -34.89624, -35.65382, -36.40988, -37.1644,
  37.49273, 36.73572, 35.97694, 35.2164, 34.4541, 33.69006, 32.9243, 
    32.15683, 31.38766, 30.61683, 29.84434, 29.07022, 28.29449, 27.51719, 
    26.73832, 25.95792, 25.17602, 24.39264, 23.60783, 22.8216, 22.034, 
    21.24507, 20.45482, 19.66332, 18.87058, 18.07666, 17.2816, 16.48543, 
    15.6882, 14.88996, 14.09074, 13.29061, 12.4896, 11.68776, 10.88514, 
    10.0818, 9.277779, 8.473132, 7.667912, 6.862171, 6.055964, 5.249342, 
    4.442361, 3.635076, 2.827541, 2.019811, 1.211942, 0.40399, -0.40399, 
    -1.211942, -2.019811, -2.827541, -3.635076, -4.442361, -5.249342, 
    -6.055964, -6.862171, -7.667912, -8.473132, -9.277779, -10.0818, 
    -10.88514, -11.68776, -12.4896, -13.29061, -14.09074, -14.88996, 
    -15.6882, -16.48543, -17.2816, -18.07666, -18.87058, -19.66332, 
    -20.45482, -21.24507, -22.034, -22.8216, -23.60783, -24.39264, -25.17602, 
    -25.95792, -26.73832, -27.51719, -28.29449, -29.07022, -29.84434, 
    -30.61683, -31.38766, -32.15683, -32.9243, -33.69006, -34.4541, -35.2164, 
    -35.97694, -36.73572, -37.49273,
  37.81525, 37.05589, 36.29453, 35.53117, 34.76583, 33.99852, 33.22925, 
    32.45805, 31.68493, 30.90992, 30.13302, 29.35428, 28.5737, 27.79133, 
    27.00718, 26.22129, 25.43369, 24.64441, 23.85349, 23.06096, 22.26687, 
    21.47124, 20.67413, 19.87557, 19.07561, 18.27429, 17.47165, 16.66776, 
    15.86266, 15.05639, 14.24901, 13.44058, 12.63114, 11.82075, 11.00947, 
    10.19736, 9.384465, 8.570855, 7.756588, 6.941722, 6.12632, 5.310442, 
    4.494153, 3.677513, 2.860586, 2.043435, 1.226125, 0.4087191, -0.4087191, 
    -1.226125, -2.043435, -2.860586, -3.677513, -4.494153, -5.310442, 
    -6.12632, -6.941722, -7.756588, -8.570855, -9.384465, -10.19736, 
    -11.00947, -11.82075, -12.63114, -13.44058, -14.24901, -15.05639, 
    -15.86266, -16.66776, -17.47165, -18.27429, -19.07561, -19.87557, 
    -20.67413, -21.47124, -22.26687, -23.06096, -23.85349, -24.64441, 
    -25.43369, -26.22129, -27.00718, -27.79133, -28.5737, -29.35428, 
    -30.13302, -30.90992, -31.68493, -32.45805, -33.22925, -33.99852, 
    -34.76583, -35.53117, -36.29453, -37.05589, -37.81525,
  38.13184, 37.37026, 36.60646, 35.84042, 35.07218, 34.30174, 33.52912, 
    32.75434, 31.97741, 31.19835, 30.4172, 29.63398, 28.84871, 28.06141, 
    27.27213, 26.4809, 25.68774, 24.89271, 24.09582, 23.29713, 22.49667, 
    21.6945, 20.89065, 20.08517, 19.2781, 18.46952, 17.65945, 16.84796, 
    16.0351, 15.22093, 14.4055, 13.58888, 12.77113, 11.9523, 11.13247, 
    10.31169, 9.490034, 8.667565, 7.844352, 7.020462, 6.195964, 5.370928, 
    4.545426, 3.719527, 2.893303, 2.066826, 1.240168, 0.4134014, -0.4134014, 
    -1.240168, -2.066826, -2.893303, -3.719527, -4.545426, -5.370928, 
    -6.195964, -7.020462, -7.844352, -8.667565, -9.490034, -10.31169, 
    -11.13247, -11.9523, -12.77113, -13.58888, -14.4055, -15.22093, -16.0351, 
    -16.84796, -17.65945, -18.46952, -19.2781, -20.08517, -20.89065, 
    -21.6945, -22.49667, -23.29713, -24.09582, -24.89271, -25.68774, 
    -26.4809, -27.27213, -28.06141, -28.84871, -29.63398, -30.4172, 
    -31.19835, -31.97741, -32.75434, -33.52912, -34.30174, -35.07218, 
    -35.84042, -36.60646, -37.37026, -38.13184,
  38.44237, 37.67871, 36.91259, 36.14403, 35.37302, 34.59959, 33.82376, 
    33.04553, 32.26494, 31.482, 30.69673, 29.90917, 29.11935, 28.32729, 
    27.53302, 26.73659, 25.93803, 25.13737, 24.33467, 23.52995, 22.72328, 
    21.91469, 21.10424, 20.29198, 19.47795, 18.66223, 17.84485, 17.02589, 
    16.20541, 15.38346, 14.56011, 13.73542, 12.90947, 12.08233, 11.25405, 
    10.42472, 9.594414, 8.763195, 7.931143, 7.098334, 6.264847, 5.430757, 
    4.596145, 3.761089, 2.925669, 2.089966, 1.254061, 0.4180338, -0.4180338, 
    -1.254061, -2.089966, -2.925669, -3.761089, -4.596145, -5.430757, 
    -6.264847, -7.098334, -7.931143, -8.763195, -9.594414, -10.42472, 
    -11.25405, -12.08233, -12.90947, -13.73542, -14.56011, -15.38346, 
    -16.20541, -17.02589, -17.84485, -18.66223, -19.47795, -20.29198, 
    -21.10424, -21.91469, -22.72328, -23.52995, -24.33467, -25.13737, 
    -25.93803, -26.73659, -27.53302, -28.32729, -29.11935, -29.90917, 
    -30.69673, -31.482, -32.26494, -33.04553, -33.82376, -34.59959, 
    -35.37302, -36.14403, -36.91259, -37.67871, -38.44237,
  38.74672, 37.9811, 37.21281, 36.44184, 35.66821, 34.89193, 34.11302, 
    33.33149, 32.54737, 31.76069, 30.97146, 30.17971, 29.38548, 28.5888, 
    27.78969, 26.98821, 26.18438, 25.37826, 24.56988, 23.75929, 22.94654, 
    22.13168, 21.31477, 20.49586, 19.67501, 18.85229, 18.02774, 17.20144, 
    16.37346, 15.54386, 14.71272, 13.88009, 13.04607, 12.21073, 11.37413, 
    10.53637, 9.697527, 8.857674, 8.016898, 7.175284, 6.332918, 5.489884, 
    4.646272, 3.802168, 2.957661, 2.112839, 1.267794, 0.4226128, -0.4226128, 
    -1.267794, -2.112839, -2.957661, -3.802168, -4.646272, -5.489884, 
    -6.332918, -7.175284, -8.016898, -8.857674, -9.697527, -10.53637, 
    -11.37413, -12.21073, -13.04607, -13.88009, -14.71272, -15.54386, 
    -16.37346, -17.20144, -18.02774, -18.85229, -19.67501, -20.49586, 
    -21.31477, -22.13168, -22.94654, -23.75929, -24.56988, -25.37826, 
    -26.18438, -26.98821, -27.78969, -28.5888, -29.38548, -30.17971, 
    -30.97146, -31.76069, -32.54737, -33.33149, -34.11302, -34.89193, 
    -35.66821, -36.44184, -37.21281, -37.9811, -38.74672,
  39.04476, 38.27731, 37.50697, 36.73372, 35.9576, 35.1786, 34.39675, 
    33.61207, 32.82457, 32.03428, 31.24123, 30.44544, 29.64695, 28.84579, 
    28.04199, 27.2356, 26.42666, 25.61521, 24.8013, 23.98498, 23.1663, 
    22.34532, 21.52209, 20.69669, 19.86915, 19.03956, 18.20799, 17.37449, 
    16.53915, 15.70203, 14.86322, 14.02279, 13.18083, 12.33741, 11.49262, 
    10.64656, 9.799295, 8.95093, 8.101551, 7.251252, 6.400125, 5.548265, 
    4.695769, 3.842732, 2.989253, 2.135427, 1.281355, 0.4271349, -0.4271349, 
    -1.281355, -2.135427, -2.989253, -3.842732, -4.695769, -5.548265, 
    -6.400125, -7.251252, -8.101551, -8.95093, -9.799295, -10.64656, 
    -11.49262, -12.33741, -13.18083, -14.02279, -14.86322, -15.70203, 
    -16.53915, -17.37449, -18.20799, -19.03956, -19.86915, -20.69669, 
    -21.52209, -22.34532, -23.1663, -23.98498, -24.8013, -25.61521, 
    -26.42666, -27.2356, -28.04199, -28.84579, -29.64695, -30.44544, 
    -31.24123, -32.03428, -32.82457, -33.61207, -34.39675, -35.1786, 
    -35.9576, -36.73372, -37.50697, -38.27731, -39.04476,
  39.33637, 38.56721, 37.79493, 37.01954, 36.24105, 35.45947, 34.67482, 
    33.88711, 33.09637, 32.30262, 31.50589, 30.7062, 29.90359, 29.0981, 
    28.28975, 27.47861, 26.6647, 25.84807, 25.02878, 24.20688, 23.38242, 
    22.55546, 21.72607, 20.8943, 20.06023, 19.22392, 18.38545, 17.5449, 
    16.70233, 15.85784, 15.0115, 14.1634, 13.31363, 12.46228, 11.60943, 
    10.75519, 9.899641, 9.042892, 8.185037, 7.326178, 6.466415, 5.605854, 
    4.744597, 3.88275, 3.02042, 2.157712, 1.294735, 0.4315965, -0.4315965, 
    -1.294735, -2.157712, -3.02042, -3.88275, -4.744597, -5.605854, 
    -6.466415, -7.326178, -8.185037, -9.042892, -9.899641, -10.75519, 
    -11.60943, -12.46228, -13.31363, -14.1634, -15.0115, -15.85784, 
    -16.70233, -17.5449, -18.38545, -19.22392, -20.06023, -20.8943, 
    -21.72607, -22.55546, -23.38242, -24.20688, -25.02878, -25.84807, 
    -26.6647, -27.47861, -28.28975, -29.0981, -29.90359, -30.7062, -31.50589, 
    -32.30262, -33.09637, -33.88711, -34.67482, -35.45947, -36.24105, 
    -37.01954, -37.79493, -38.56721, -39.33637,
  39.62142, 38.85067, 38.07658, 37.29916, 36.51843, 35.73439, 34.94707, 
    34.15647, 33.36263, 32.56555, 31.76528, 30.96183, 30.15525, 29.34557, 
    28.53283, 27.71707, 26.89834, 26.07669, 25.25217, 24.42483, 23.59474, 
    22.76195, 21.92654, 21.08856, 20.2481, 19.40522, 18.56001, 17.71254, 
    16.8629, 16.01117, 15.15745, 14.30182, 13.44438, 12.58523, 11.72446, 
    10.86218, 9.998483, 9.133484, 8.267286, 7.4, 6.531734, 5.662601, 
    4.792715, 3.922188, 3.051136, 2.179676, 1.307923, 0.4359938, -0.4359938, 
    -1.307923, -2.179676, -3.051136, -3.922188, -4.792715, -5.662601, 
    -6.531734, -7.4, -8.267286, -9.133484, -9.998483, -10.86218, -11.72446, 
    -12.58523, -13.44438, -14.30182, -15.15745, -16.01117, -16.8629, 
    -17.71254, -18.56001, -19.40522, -20.2481, -21.08856, -21.92654, 
    -22.76195, -23.59474, -24.42483, -25.25217, -26.07669, -26.89834, 
    -27.71707, -28.53283, -29.34557, -30.15525, -30.96183, -31.76528, 
    -32.56555, -33.36263, -34.15647, -34.94707, -35.73439, -36.51843, 
    -37.29916, -38.07658, -38.85067, -39.62142,
  39.89979, 39.12755, 38.35176, 37.57244, 36.78959, 36.00322, 35.21335, 
    34.42, 33.62318, 32.82292, 32.01924, 31.21218, 30.40177, 29.58805, 
    28.77106, 27.95084, 27.12744, 26.30091, 25.4713, 24.63868, 23.8031, 
    22.96464, 22.12335, 21.27932, 20.43262, 19.58332, 18.73152, 17.87728, 
    17.02072, 16.1619, 15.30094, 14.43793, 13.57297, 12.70616, 11.83762, 
    10.96744, 10.09574, 9.222629, 8.34823, 7.472656, 6.596026, 5.718461, 
    4.840082, 3.961012, 3.081377, 2.201299, 1.320906, 0.4403231, -0.4403231, 
    -1.320906, -2.201299, -3.081377, -3.961012, -4.840082, -5.718461, 
    -6.596026, -7.472656, -8.34823, -9.222629, -10.09574, -10.96744, 
    -11.83762, -12.70616, -13.57297, -14.43793, -15.30094, -16.1619, 
    -17.02072, -17.87728, -18.73152, -19.58332, -20.43262, -21.27932, 
    -22.12335, -22.96464, -23.8031, -24.63868, -25.4713, -26.30091, 
    -27.12744, -27.95084, -28.77106, -29.58805, -30.40177, -31.21218, 
    -32.01924, -32.82292, -33.62318, -34.42, -35.21335, -36.00322, -36.78959, 
    -37.57244, -38.35176, -39.12755, -39.89979,
  40.17135, 39.39772, 38.62035, 37.83924, 37.05439, 36.26581, 35.47353, 
    34.67754, 33.87788, 33.07457, 32.26763, 31.45709, 30.643, 29.82537, 
    29.00427, 28.17974, 27.35181, 26.52055, 25.68602, 24.84826, 24.00736, 
    23.16337, 22.31637, 21.46644, 20.61365, 19.75808, 18.89984, 18.03899, 
    17.17565, 16.30991, 15.44186, 14.57162, 13.69929, 12.82498, 11.9488, 
    11.07087, 10.19132, 9.31025, 8.427797, 7.544083, 6.659235, 5.773382, 
    4.886656, 3.999188, 3.111113, 2.222563, 1.333673, 0.4445804, -0.4445804, 
    -1.333673, -2.222563, -3.111113, -3.999188, -4.886656, -5.773382, 
    -6.659235, -7.544083, -8.427797, -9.31025, -10.19132, -11.07087, 
    -11.9488, -12.82498, -13.69929, -14.57162, -15.44186, -16.30991, 
    -17.17565, -18.03899, -18.89984, -19.75808, -20.61365, -21.46644, 
    -22.31637, -23.16337, -24.00736, -24.84826, -25.68602, -26.52055, 
    -27.35181, -28.17974, -29.00427, -29.82537, -30.643, -31.45709, 
    -32.26763, -33.07457, -33.87788, -34.67754, -35.47353, -36.26581, 
    -37.05439, -37.83924, -38.62035, -39.39772, -40.17135,
  40.43598, 39.66107, 38.88222, 38.09942, 37.31269, 36.52202, 35.72744, 
    34.92895, 34.12658, 33.32034, 32.51027, 31.6964, 30.87876, 30.05738, 
    29.23232, 28.40361, 27.57131, 26.73548, 25.89616, 25.05343, 24.20735, 
    23.35799, 22.50543, 21.64975, 20.79103, 19.92936, 19.06483, 18.19754, 
    17.32758, 16.45506, 15.58009, 14.70277, 13.82323, 12.94157, 12.05792, 
    11.1724, 10.28514, 9.396269, 8.505915, 7.614214, 6.721301, 5.827315, 
    4.932395, 4.036681, 3.140318, 2.243447, 1.346213, 0.448762, -0.448762, 
    -1.346213, -2.243447, -3.140318, -4.036681, -4.932395, -5.827315, 
    -6.721301, -7.614214, -8.505915, -9.396269, -10.28514, -11.1724, 
    -12.05792, -12.94157, -13.82323, -14.70277, -15.58009, -16.45506, 
    -17.32758, -18.19754, -19.06483, -19.92936, -20.79103, -21.64975, 
    -22.50543, -23.35799, -24.20735, -25.05343, -25.89616, -26.73548, 
    -27.57131, -28.40361, -29.23232, -30.05738, -30.87876, -31.6964, 
    -32.51027, -33.32034, -34.12658, -34.92895, -35.72744, -36.52202, 
    -37.31269, -38.09942, -38.88222, -39.66107, -40.43598,
  40.69355, 39.91746, 39.13723, 38.35286, 37.56434, 36.7717, 35.97494, 
    35.17407, 34.36911, 33.56009, 32.74702, 31.92994, 31.10889, 30.28391, 
    29.45502, 28.6223, 27.78577, 26.94551, 26.10157, 25.25401, 24.40292, 
    23.54835, 22.69039, 21.82912, 20.96463, 20.09701, 19.22636, 18.35277, 
    17.47636, 16.59723, 15.71549, 14.83126, 13.94467, 13.05583, 12.16487, 
    11.27192, 10.37712, 9.480604, 8.582511, 7.682984, 6.782168, 5.880208, 
    4.977254, 4.073455, 3.168964, 2.263932, 1.358514, 0.4528638, -0.4528638, 
    -1.358514, -2.263932, -3.168964, -4.073455, -4.977254, -5.880208, 
    -6.782168, -7.682984, -8.582511, -9.480604, -10.37712, -11.27192, 
    -12.16487, -13.05583, -13.94467, -14.83126, -15.71549, -16.59723, 
    -17.47636, -18.35277, -19.22636, -20.09701, -20.96463, -21.82912, 
    -22.69039, -23.54835, -24.40292, -25.25401, -26.10157, -26.94551, 
    -27.78577, -28.6223, -29.45502, -30.28391, -31.10889, -31.92994, 
    -32.74702, -33.56009, -34.36911, -35.17407, -35.97494, -36.7717, 
    -37.56434, -38.35286, -39.13723, -39.91746, -40.69355,
  40.94394, 40.16676, 39.38524, 38.5994, 37.80922, 37.01471, 36.21589, 
    35.41275, 34.60533, 33.79364, 32.97771, 32.15757, 31.33325, 30.50479, 
    29.67224, 28.83563, 27.99503, 27.1505, 26.30208, 25.44986, 24.5939, 
    23.73428, 22.87107, 22.00438, 21.13428, 20.26088, 19.38427, 18.50457, 
    17.62187, 16.73629, 15.84795, 14.95698, 14.0635, 13.16765, 12.26954, 
    11.36934, 10.46716, 9.563174, 8.657512, 7.750327, 6.841775, 5.93201, 
    5.02119, 4.109474, 3.197022, 2.283998, 1.370563, 0.4568816, -0.4568816, 
    -1.370563, -2.283998, -3.197022, -4.109474, -5.02119, -5.93201, 
    -6.841775, -7.750327, -8.657512, -9.563174, -10.46716, -11.36934, 
    -12.26954, -13.16765, -14.0635, -14.95698, -15.84795, -16.73629, 
    -17.62187, -18.50457, -19.38427, -20.26088, -21.13428, -22.00438, 
    -22.87107, -23.73428, -24.5939, -25.44986, -26.30208, -27.1505, 
    -27.99503, -28.83563, -29.67224, -30.50479, -31.33325, -32.15757, 
    -32.97771, -33.79364, -34.60533, -35.41275, -36.21589, -37.01471, 
    -37.80922, -38.5994, -39.38524, -40.16676, -40.94394,
  41.18702, 40.40884, 39.62614, 38.83891, 38.04717, 37.2509, 36.45013, 
    35.64485, 34.83509, 34.02087, 33.2022, 32.37912, 31.55167, 30.71988, 
    29.88379, 29.04346, 28.19893, 27.35027, 26.49753, 25.6408, 24.78014, 
    23.91562, 23.04734, 22.17539, 21.29985, 20.42083, 19.53844, 18.65277, 
    17.76396, 16.87211, 15.97735, 15.07981, 14.17962, 13.27692, 12.37185, 
    11.46456, 10.55519, 9.643898, 8.730841, 7.816175, 6.900063, 5.982669, 
    5.064158, 4.144701, 3.224465, 2.303623, 1.382348, 0.4608116, -0.4608116, 
    -1.382348, -2.303623, -3.224465, -4.144701, -5.064158, -5.982669, 
    -6.900063, -7.816175, -8.730841, -9.643898, -10.55519, -11.46456, 
    -12.37185, -13.27692, -14.17962, -15.07981, -15.97735, -16.87211, 
    -17.76396, -18.65277, -19.53844, -20.42083, -21.29985, -22.17539, 
    -23.04734, -23.91562, -24.78014, -25.6408, -26.49753, -27.35027, 
    -28.19893, -29.04346, -29.88379, -30.71988, -31.55167, -32.37912, 
    -33.2022, -34.02087, -34.83509, -35.64485, -36.45013, -37.2509, 
    -38.04717, -38.83891, -39.62614, -40.40884, -41.18702,
  41.42268, 40.64358, 39.85978, 39.07127, 38.27806, 37.48015, 36.67753, 
    35.87022, 35.05824, 34.2416, 33.42032, 32.59444, 31.76398, 30.929, 
    30.08952, 29.2456, 28.3973, 27.54466, 26.68777, 25.82668, 24.96147, 
    24.09223, 23.21904, 22.34199, 21.46118, 20.57672, 19.68871, 18.79726, 
    17.9025, 17.00456, 16.10355, 15.19962, 14.2929, 13.38354, 12.47168, 
    11.55748, 10.6411, 9.722692, 8.802423, 7.880459, 6.956971, 6.032131, 
    5.106114, 4.179099, 3.251263, 2.322789, 1.393856, 0.4646493, -0.4646493, 
    -1.393856, -2.322789, -3.251263, -4.179099, -5.106114, -6.032131, 
    -6.956971, -7.880459, -8.802423, -9.722692, -10.6411, -11.55748, 
    -12.47168, -13.38354, -14.2929, -15.19962, -16.10355, -17.00456, 
    -17.9025, -18.79726, -19.68871, -20.57672, -21.46118, -22.34199, 
    -23.21904, -24.09223, -24.96147, -25.82668, -26.68777, -27.54466, 
    -28.3973, -29.2456, -30.08952, -30.929, -31.76398, -32.59444, -33.42032, 
    -34.2416, -35.05824, -35.87022, -36.67753, -37.48015, -38.27806, 
    -39.07127, -39.85978, -40.64358, -41.42268,
  41.65079, 40.87085, 40.08604, 39.29634, 38.50176, 37.70229, 36.89794, 
    36.08871, 35.27462, 34.45568, 33.63192, 32.80336, 31.97004, 31.132, 
    30.28927, 29.44192, 28.58998, 27.73353, 26.87262, 26.00734, 25.13775, 
    24.26394, 23.386, 22.50403, 21.61812, 20.72838, 19.83493, 18.93789, 
    18.03736, 17.1335, 16.22643, 15.31629, 14.40323, 13.48739, 12.56893, 
    11.64802, 10.72481, 9.799476, 8.872184, 7.943112, 7.012438, 6.080344, 
    5.147013, 4.212631, 3.277388, 2.341473, 1.405076, 0.4683909, -0.4683909, 
    -1.405076, -2.341473, -3.277388, -4.212631, -5.147013, -6.080344, 
    -7.012438, -7.943112, -8.872184, -9.799476, -10.72481, -11.64802, 
    -12.56893, -13.48739, -14.40323, -15.31629, -16.22643, -17.1335, 
    -18.03736, -18.93789, -19.83493, -20.72838, -21.61812, -22.50403, 
    -23.386, -24.26394, -25.13775, -26.00734, -26.87262, -27.73353, 
    -28.58998, -29.44192, -30.28927, -31.132, -31.97004, -32.80336, 
    -33.63192, -34.45568, -35.27462, -36.08871, -36.89794, -37.70229, 
    -38.50176, -39.29634, -40.08604, -40.87085, -41.65079,
  41.87124, 41.09053, 40.30479, 39.51399, 38.71813, 37.9172, 37.11122, 
    36.30017, 35.48409, 34.66297, 33.83684, 33.00574, 32.16968, 31.32872, 
    30.48288, 29.63223, 28.77681, 27.91669, 27.05193, 26.18261, 25.3088, 
    24.43059, 23.54808, 22.66135, 21.77052, 20.87569, 19.97698, 19.07451, 
    18.16841, 17.25882, 16.34587, 15.42971, 14.51049, 13.58837, 12.66351, 
    11.73607, 10.80623, 9.874163, 8.940046, 8.004064, 7.066403, 6.127254, 
    5.186808, 4.245261, 3.30281, 2.359655, 1.415995, 0.472032, -0.472032, 
    -1.415995, -2.359655, -3.30281, -4.245261, -5.186808, -6.127254, 
    -7.066403, -8.004064, -8.940046, -9.874163, -10.80623, -11.73607, 
    -12.66351, -13.58837, -14.51049, -15.42971, -16.34587, -17.25882, 
    -18.16841, -19.07451, -19.97698, -20.87569, -21.77052, -22.66135, 
    -23.54808, -24.43059, -25.3088, -26.18261, -27.05193, -27.91669, 
    -28.77681, -29.63223, -30.48288, -31.32872, -32.16968, -33.00574, 
    -33.83684, -34.66297, -35.48409, -36.30017, -37.11122, -37.9172, 
    -38.71813, -39.51399, -40.30479, -41.09053, -41.87124,
  42.08391, 41.30251, 40.51591, 39.72409, 38.92703, 38.12474, 37.31722, 
    36.50447, 35.68649, 34.86331, 34.03494, 33.20141, 32.36275, 31.519, 
    30.6702, 29.81639, 28.95764, 28.094, 27.22555, 26.35234, 25.47448, 
    24.59204, 23.70512, 22.81381, 21.91823, 21.01848, 20.11469, 19.20699, 
    18.2955, 17.38036, 16.46173, 15.53974, 14.61457, 13.68636, 12.75529, 
    11.82154, 10.88527, 9.946671, 9.005934, 8.063247, 7.118805, 6.172808, 
    5.225454, 4.27695, 3.3275, 2.377314, 1.4266, 0.4755684, -0.4755684, 
    -1.4266, -2.377314, -3.3275, -4.27695, -5.225454, -6.172808, -7.118805, 
    -8.063247, -9.005934, -9.946671, -10.88527, -11.82154, -12.75529, 
    -13.68636, -14.61457, -15.53974, -16.46173, -17.38036, -18.2955, 
    -19.20699, -20.11469, -21.01848, -21.91823, -22.81381, -23.70512, 
    -24.59204, -25.47448, -26.35234, -27.22555, -28.094, -28.95764, 
    -29.81639, -30.6702, -31.519, -32.36275, -33.20141, -34.03494, -34.86331, 
    -35.68649, -36.50447, -37.31722, -38.12474, -38.92703, -39.72409, 
    -40.51591, -41.30251, -42.08391,
  42.28868, 41.50666, 40.71927, 39.9265, 39.12834, 38.32478, 37.51582, 
    36.70145, 35.8817, 35.05656, 34.22607, 33.39024, 32.5491, 31.70269, 
    30.85106, 29.99424, 29.1323, 28.2653, 27.3933, 26.51638, 25.63463, 
    24.74813, 23.85697, 22.96125, 22.0611, 21.15662, 20.24794, 19.33519, 
    18.4185, 17.49802, 16.57389, 15.64629, 14.71535, 13.78126, 12.84419, 
    11.90432, 10.96183, 10.01692, 9.069772, 8.120593, 7.169584, 6.216953, 
    5.262908, 4.307662, 3.35143, 2.394429, 1.436878, 0.478996, -0.478996, 
    -1.436878, -2.394429, -3.35143, -4.307662, -5.262908, -6.216953, 
    -7.169584, -8.120593, -9.069772, -10.01692, -10.96183, -11.90432, 
    -12.84419, -13.78126, -14.71535, -15.64629, -16.57389, -17.49802, 
    -18.4185, -19.33519, -20.24794, -21.15662, -22.0611, -22.96125, 
    -23.85697, -24.74813, -25.63463, -26.51638, -27.3933, -28.2653, -29.1323, 
    -29.99424, -30.85106, -31.70269, -32.5491, -33.39024, -34.22607, 
    -35.05656, -35.8817, -36.70145, -37.51582, -38.32478, -39.12834, 
    -39.9265, -40.71927, -41.50666, -42.28868,
  42.48545, 41.70287, 40.91476, 40.12112, 39.32193, 38.51718, 37.70687, 
    36.891, 36.06956, 35.24258, 34.41008, 33.57207, 32.72858, 31.87964, 
    31.02531, 30.16563, 29.30065, 28.43043, 27.55505, 26.67457, 25.78909, 
    24.89869, 24.00347, 23.10353, 22.19899, 21.28997, 20.37659, 19.45897, 
    18.53728, 17.61165, 16.68224, 15.74921, 14.81272, 13.87296, 12.9301, 
    11.98433, 11.03584, 10.08482, 9.131484, 8.176033, 7.218679, 6.259636, 
    5.299122, 4.337358, 3.374569, 2.41098, 1.446817, 0.4823107, -0.4823107, 
    -1.446817, -2.41098, -3.374569, -4.337358, -5.299122, -6.259636, 
    -7.218679, -8.176033, -9.131484, -10.08482, -11.03584, -11.98433, 
    -12.9301, -13.87296, -14.81272, -15.74921, -16.68224, -17.61165, 
    -18.53728, -19.45897, -20.37659, -21.28997, -22.19899, -23.10353, 
    -24.00347, -24.89869, -25.78909, -26.67457, -27.55505, -28.43043, 
    -29.30065, -30.16563, -31.02531, -31.87964, -32.72858, -33.57207, 
    -34.41008, -35.24258, -36.06956, -36.891, -37.70687, -38.51718, 
    -39.32193, -40.12112, -40.91476, -41.70287, -42.48545,
  42.67411, 41.89101, 41.10225, 40.30781, 39.50767, 38.70182, 37.89024, 
    37.07295, 36.24994, 35.42123, 34.58682, 33.74675, 32.90103, 32.0497, 
    31.19281, 30.3304, 29.46252, 28.58924, 27.71063, 26.82676, 25.93772, 
    25.04359, 24.14449, 23.2405, 22.33176, 21.41838, 20.50048, 19.57821, 
    18.65171, 17.72114, 16.78664, 15.8484, 14.90658, 13.96135, 13.01292, 
    12.06147, 11.10719, 10.1503, 9.190996, 8.229501, 7.266029, 6.300805, 
    5.334054, 4.366004, 3.39689, 2.426945, 1.456406, 0.4855082, -0.4855082, 
    -1.456406, -2.426945, -3.39689, -4.366004, -5.334054, -6.300805, 
    -7.266029, -8.229501, -9.190996, -10.1503, -11.10719, -12.06147, 
    -13.01292, -13.96135, -14.90658, -15.8484, -16.78664, -17.72114, 
    -18.65171, -19.57821, -20.50048, -21.41838, -22.33176, -23.2405, 
    -24.14449, -25.04359, -25.93772, -26.82676, -27.71063, -28.58924, 
    -29.46252, -30.3304, -31.19281, -32.0497, -32.90103, -33.74675, 
    -34.58682, -35.42123, -36.24994, -37.07295, -37.89024, -38.70182, 
    -39.50767, -40.30781, -41.10225, -41.89101, -42.67411,
  42.85454, 42.07099, 41.28164, 40.48646, 39.68544, 38.87856, 38.06581, 
    37.2472, 36.42271, 35.59236, 34.75616, 33.91414, 33.06631, 32.21272, 
    31.3534, 30.4884, 29.61777, 28.74158, 27.8599, 26.9728, 26.08036, 
    25.18268, 24.27987, 23.37202, 22.45926, 21.5417, 20.61949, 19.69276, 
    18.76166, 17.82635, 16.88698, 15.94374, 14.99679, 14.04633, 13.09255, 
    12.13564, 11.17581, 10.21327, 9.248235, 8.280929, 7.311576, 6.340407, 
    5.367657, 4.393563, 3.418365, 2.442306, 1.46563, 0.4885846, -0.4885846, 
    -1.46563, -2.442306, -3.418365, -4.393563, -5.367657, -6.340407, 
    -7.311576, -8.280929, -9.248235, -10.21327, -11.17581, -12.13564, 
    -13.09255, -14.04633, -14.99679, -15.94374, -16.88698, -17.82635, 
    -18.76166, -19.69276, -20.61949, -21.5417, -22.45926, -23.37202, 
    -24.27987, -25.18268, -26.08036, -26.9728, -27.8599, -28.74158, 
    -29.61777, -30.4884, -31.3534, -32.21272, -33.06631, -33.91414, 
    -34.75616, -35.59236, -36.42271, -37.2472, -38.06581, -38.87856, 
    -39.68544, -40.48646, -41.28164, -42.07099, -42.85454,
  43.02665, 42.24269, 41.4528, 40.65696, 39.85512, 39.04729, 38.23346, 
    37.4136, 36.58773, 35.75585, 34.91797, 34.07411, 33.2243, 32.36856, 
    31.50695, 30.6395, 29.76627, 28.88731, 28.00271, 27.11254, 26.21687, 
    25.31582, 24.40947, 23.49794, 22.58134, 21.65982, 20.73348, 19.8025, 
    18.867, 17.92716, 16.98314, 16.03511, 15.08327, 14.1278, 13.16889, 
    12.20676, 11.2416, 10.27365, 9.303126, 8.330251, 7.355261, 6.378393, 
    5.399891, 4.419998, 3.438965, 2.457041, 1.47448, 0.4915359, -0.4915359, 
    -1.47448, -2.457041, -3.438965, -4.419998, -5.399891, -6.378393, 
    -7.355261, -8.330251, -9.303126, -10.27365, -11.2416, -12.20676, 
    -13.16889, -14.1278, -15.08327, -16.03511, -16.98314, -17.92716, -18.867, 
    -19.8025, -20.73348, -21.65982, -22.58134, -23.49794, -24.40947, 
    -25.31582, -26.21687, -27.11254, -28.00271, -28.88731, -29.76627, 
    -30.6395, -31.50695, -32.36856, -33.2243, -34.07411, -34.91797, 
    -35.75585, -36.58773, -37.4136, -38.23346, -39.04729, -39.85512, 
    -40.65696, -41.4528, -42.24269, -43.02665,
  43.19033, 42.40602, 41.61564, 40.81918, 40.0166, 39.20789, 38.39304, 
    37.57203, 36.74487, 35.91155, 35.0721, 34.22652, 33.37484, 32.51709, 
    31.65331, 30.78355, 29.90785, 29.02629, 28.13892, 27.24584, 26.34712, 
    25.44285, 24.53315, 23.61813, 22.69789, 21.77258, 20.84233, 19.90729, 
    18.96761, 18.02345, 17.075, 16.12242, 15.1659, 14.20564, 13.24185, 
    12.27472, 11.30449, 10.33138, 9.355601, 8.377405, 7.397027, 6.414712, 
    5.430711, 4.445276, 3.458663, 2.471131, 1.482942, 0.494358, -0.494358, 
    -1.482942, -2.471131, -3.458663, -4.445276, -5.430711, -6.414712, 
    -7.397027, -8.377405, -9.355601, -10.33138, -11.30449, -12.27472, 
    -13.24185, -14.20564, -15.1659, -16.12242, -17.075, -18.02345, -18.96761, 
    -19.90729, -20.84233, -21.77258, -22.69789, -23.61813, -24.53315, 
    -25.44285, -26.34712, -27.24584, -28.13892, -29.02629, -29.90785, 
    -30.78355, -31.65331, -32.51709, -33.37484, -34.22652, -35.0721, 
    -35.91155, -36.74487, -37.57203, -38.39304, -39.20789, -40.0166, 
    -40.81918, -41.61564, -42.40602, -43.19033,
  43.34549, 42.56086, 41.77005, 40.97303, 40.16977, 39.36025, 38.54446, 
    37.72238, 36.89401, 36.05936, 35.21843, 34.37123, 33.5178, 32.65816, 
    31.79235, 30.92041, 30.04239, 29.15837, 28.2684, 27.37256, 26.47095, 
    25.56366, 24.65079, 23.73245, 22.80877, 21.87987, 20.94591, 20.00702, 
    19.06337, 18.11512, 17.16244, 16.20553, 15.24457, 14.27977, 13.31133, 
    12.33946, 11.3644, 10.38636, 9.40559, 8.422327, 7.436818, 6.449316, 
    5.460076, 4.46936, 3.477432, 2.484558, 1.491006, 0.4970472, -0.4970472, 
    -1.491006, -2.484558, -3.477432, -4.46936, -5.460076, -6.449316, 
    -7.436818, -8.422327, -9.40559, -10.38636, -11.3644, -12.33946, 
    -13.31133, -14.27977, -15.24457, -16.20553, -17.16244, -18.11512, 
    -19.06337, -20.00702, -20.94591, -21.87987, -22.80877, -23.73245, 
    -24.65079, -25.56366, -26.47095, -27.37256, -28.2684, -29.15837, 
    -30.04239, -30.92041, -31.79235, -32.65816, -33.5178, -34.37123, 
    -35.21843, -36.05936, -36.89401, -37.72238, -38.54446, -39.36025, 
    -40.16977, -40.97303, -41.77005, -42.56086, -43.34549,
  43.49203, 42.70713, 41.91592, 41.1184, 40.31451, 39.50425, 38.6876, 
    37.86452, 37.03504, 36.19914, 35.35684, 34.50814, 33.65307, 32.79165, 
    31.92393, 31.04995, 30.16976, 29.28342, 28.391, 27.49258, 26.58825, 
    25.6781, 24.76223, 23.84077, 22.91384, 21.98156, 21.04409, 20.10156, 
    19.15416, 18.20203, 17.24537, 16.28436, 15.3192, 14.35008, 13.37724, 
    12.40088, 11.42123, 10.43853, 9.453025, 8.464956, 7.47458, 6.482156, 
    5.487947, 4.49222, 3.495247, 2.497301, 1.49866, 0.4995998, -0.4995998, 
    -1.49866, -2.497301, -3.495247, -4.49222, -5.487947, -6.482156, -7.47458, 
    -8.464956, -9.453025, -10.43853, -11.42123, -12.40088, -13.37724, 
    -14.35008, -15.3192, -16.28436, -17.24537, -18.20203, -19.15416, 
    -20.10156, -21.04409, -21.98156, -22.91384, -23.84077, -24.76223, 
    -25.6781, -26.58825, -27.49258, -28.391, -29.28342, -30.16976, -31.04995, 
    -31.92393, -32.79165, -33.65307, -34.50814, -35.35684, -36.19914, 
    -37.03504, -37.86452, -38.6876, -39.50425, -40.31451, -41.1184, 
    -41.91592, -42.70713, -43.49203,
  43.62987, 42.84472, 42.05317, 41.25519, 40.45074, 39.63979, 38.82234, 
    37.99836, 37.16784, 36.33079, 35.48721, 34.6371, 33.78051, 32.91744, 
    32.04794, 31.17205, 30.28983, 29.40132, 28.50661, 27.60576, 26.69888, 
    25.78605, 24.86737, 23.94298, 23.01299, 22.07753, 21.13675, 20.19081, 
    19.23986, 18.28409, 17.32367, 16.3588, 15.38967, 14.4165, 13.43949, 
    12.45889, 11.47492, 10.48782, 9.49784, 8.505234, 7.510261, 6.513187, 
    5.514283, 4.513822, 3.512082, 2.509345, 1.505893, 0.502012, -0.502012, 
    -1.505893, -2.509345, -3.512082, -4.513822, -5.514283, -6.513187, 
    -7.510261, -8.505234, -9.49784, -10.48782, -11.47492, -12.45889, 
    -13.43949, -14.4165, -15.38967, -16.3588, -17.32367, -18.28409, 
    -19.23986, -20.19081, -21.13675, -22.07753, -23.01299, -23.94298, 
    -24.86737, -25.78605, -26.69888, -27.60576, -28.50661, -29.40132, 
    -30.28983, -31.17205, -32.04794, -32.91744, -33.78051, -34.6371, 
    -35.48721, -36.33079, -37.16784, -37.99836, -38.82234, -39.63979, 
    -40.45074, -41.25519, -42.05317, -42.84472, -43.62987,
  43.75893, 42.97356, 42.18171, 41.38331, 40.57834, 39.76678, 38.94859, 
    38.12377, 37.2923, 36.45418, 35.60942, 34.75802, 33.90001, 33.03541, 
    32.16426, 31.28659, 30.40247, 29.51195, 28.6151, 27.71199, 26.80272, 
    25.88738, 24.96609, 24.03895, 23.10609, 22.16766, 21.22379, 20.27464, 
    19.32038, 18.36119, 17.39725, 16.42875, 15.4559, 14.47891, 13.49801, 
    12.51342, 11.52539, 10.53416, 9.539974, 8.543103, 7.54381, 6.542367, 
    5.539048, 4.534135, 3.527913, 2.52067, 1.512695, 0.5042805, -0.5042805, 
    -1.512695, -2.52067, -3.527913, -4.534135, -5.539048, -6.542367, 
    -7.54381, -8.543103, -9.539974, -10.53416, -11.52539, -12.51342, 
    -13.49801, -14.47891, -15.4559, -16.42875, -17.39725, -18.36119, 
    -19.32038, -20.27464, -21.22379, -22.16766, -23.10609, -24.03895, 
    -24.96609, -25.88738, -26.80272, -27.71199, -28.6151, -29.51195, 
    -30.40247, -31.28659, -32.16426, -33.03541, -33.90001, -34.75802, 
    -35.60942, -36.45418, -37.2923, -38.12377, -38.94859, -39.76678, 
    -40.57834, -41.38331, -42.18171, -42.97356, -43.75893,
  43.87911, 43.09357, 42.30143, 41.50267, 40.69724, 39.88511, 39.06625, 
    38.24066, 37.40832, 36.56922, 35.72337, 34.87078, 34.01146, 33.14545, 
    32.27277, 31.39346, 30.50758, 29.61518, 28.71634, 27.81114, 26.89966, 
    25.98199, 25.05826, 24.12856, 23.19304, 22.25184, 21.30509, 20.35295, 
    19.39561, 18.43323, 17.466, 16.49412, 15.5178, 14.53725, 13.55271, 
    12.5644, 11.57257, 10.57748, 9.579368, 8.578511, 7.57518, 6.56965, 
    5.562205, 4.55313, 3.542717, 2.53126, 1.519056, 0.5064019, -0.5064019, 
    -1.519056, -2.53126, -3.542717, -4.55313, -5.562205, -6.56965, -7.57518, 
    -8.578511, -9.579368, -10.57748, -11.57257, -12.5644, -13.55271, 
    -14.53725, -15.5178, -16.49412, -17.466, -18.43323, -19.39561, -20.35295, 
    -21.30509, -22.25184, -23.19304, -24.12856, -25.05826, -25.98199, 
    -26.89966, -27.81114, -28.71634, -29.61518, -30.50758, -31.39346, 
    -32.27277, -33.14545, -34.01146, -34.87078, -35.72337, -36.56922, 
    -37.40832, -38.24066, -39.06625, -39.88511, -40.69724, -41.50267, 
    -42.30143, -43.09357, -43.87911,
  43.99035, 43.20465, 42.41228, 41.61318, 40.80733, 39.99469, 39.17523, 
    38.34894, 37.5158, 36.67581, 35.82896, 34.97528, 34.11476, 33.24744, 
    32.37335, 31.49253, 30.60504, 29.71092, 28.81025, 27.90311, 26.98958, 
    26.06977, 25.14377, 24.21172, 23.27374, 22.32997, 21.38055, 20.42565, 
    19.46544, 18.50011, 17.52983, 16.55482, 15.57528, 14.59143, 13.60351, 
    12.61175, 11.6164, 10.61772, 9.615962, 8.611405, 7.604323, 6.594999, 
    5.58372, 4.570779, 3.556473, 2.541101, 1.524966, 0.5083731, -0.5083731, 
    -1.524966, -2.541101, -3.556473, -4.570779, -5.58372, -6.594999, 
    -7.604323, -8.611405, -9.615962, -10.61772, -11.6164, -12.61175, 
    -13.60351, -14.59143, -15.57528, -16.55482, -17.52983, -18.50011, 
    -19.46544, -20.42565, -21.38055, -22.32997, -23.27374, -24.21172, 
    -25.14377, -26.06977, -26.98958, -27.90311, -28.81025, -29.71092, 
    -30.60504, -31.49253, -32.37335, -33.24744, -34.11476, -34.97528, 
    -35.82896, -36.67581, -37.5158, -38.34894, -39.17523, -39.99469, 
    -40.80733, -41.61318, -42.41228, -43.20465, -43.99035,
  44.09258, 43.30674, 42.51416, 41.71477, 40.90854, 40.09544, 39.27544, 
    38.44851, 37.61465, 36.77385, 35.9261, 35.07141, 34.20981, 33.3413, 
    32.46593, 31.58372, 30.69475, 29.79905, 28.89671, 27.98779, 27.07239, 
    26.1506, 25.22254, 24.28832, 23.34808, 22.40195, 21.45008, 20.49264, 
    19.5298, 18.56174, 17.58866, 16.61077, 15.62826, 14.64138, 13.65034, 
    12.6554, 11.65681, 10.65482, 9.649706, 8.641738, 7.631198, 6.618376, 
    5.603562, 4.587056, 3.569159, 2.550177, 1.530417, 0.510191, -0.510191, 
    -1.530417, -2.550177, -3.569159, -4.587056, -5.603562, -6.618376, 
    -7.631198, -8.641738, -9.649706, -10.65482, -11.65681, -12.6554, 
    -13.65034, -14.64138, -15.62826, -16.61077, -17.58866, -18.56174, 
    -19.5298, -20.49264, -21.45008, -22.40195, -23.34808, -24.28832, 
    -25.22254, -26.1506, -27.07239, -27.98779, -28.89671, -29.79905, 
    -30.69475, -31.58372, -32.46593, -33.3413, -34.20981, -35.07141, 
    -35.9261, -36.77385, -37.61465, -38.44851, -39.27544, -40.09544, 
    -40.90854, -41.71477, -42.51416, -43.30674, -44.09258,
  44.18572, 43.39978, 42.60701, 41.80736, 41.0008, 40.18729, 39.3668, 
    38.53931, 37.7048, 36.86326, 36.01469, 35.15911, 34.29651, 33.42693, 
    32.55039, 31.66694, 30.77662, 29.87949, 28.97562, 28.06509, 27.14798, 
    26.2244, 25.29446, 24.35827, 23.41596, 22.46768, 21.51358, 20.55383, 
    19.58859, 18.61805, 17.64242, 16.66188, 15.67667, 14.68701, 13.69314, 
    12.6953, 11.69374, 10.68873, 9.680549, 8.669463, 7.655765, 6.639744, 
    5.6217, 4.601935, 3.580756, 2.558473, 1.535401, 0.511853, -0.511853, 
    -1.535401, -2.558473, -3.580756, -4.601935, -5.6217, -6.639744, 
    -7.655765, -8.669463, -9.680549, -10.68873, -11.69374, -12.6953, 
    -13.69314, -14.68701, -15.67667, -16.66188, -17.64242, -18.61805, 
    -19.58859, -20.55383, -21.51358, -22.46768, -23.41596, -24.35827, 
    -25.29446, -26.2244, -27.14798, -28.06509, -28.97562, -29.87949, 
    -30.77662, -31.66694, -32.55039, -33.42693, -34.29651, -35.15911, 
    -36.01469, -36.86326, -37.7048, -38.53931, -39.3668, -40.18729, -41.0008, 
    -41.80736, -42.60701, -43.39978, -44.18572,
  44.26973, 43.48369, 42.69076, 41.89089, 41.08404, 40.27016, 39.44924, 
    38.62124, 37.78615, 36.94396, 36.09467, 35.23827, 34.37479, 33.50424, 
    32.62666, 31.74208, 30.85055, 29.95214, 29.0469, 28.13491, 27.21628, 
    26.29108, 25.35944, 24.42147, 23.47731, 22.52709, 21.57098, 20.60913, 
    19.64173, 18.66896, 17.69101, 16.7081, 15.72045, 14.72828, 13.73184, 
    12.73137, 11.72714, 10.7194, 9.708443, 8.69454, 7.677984, 6.659072, 
    5.638107, 4.615394, 3.591246, 2.565979, 1.539908, 0.5133564, -0.5133564, 
    -1.539908, -2.565979, -3.591246, -4.615394, -5.638107, -6.659072, 
    -7.677984, -8.69454, -9.708443, -10.7194, -11.72714, -12.73137, 
    -13.73184, -14.72828, -15.72045, -16.7081, -17.69101, -18.66896, 
    -19.64173, -20.60913, -21.57098, -22.52709, -23.47731, -24.42147, 
    -25.35944, -26.29108, -27.21628, -28.13491, -29.0469, -29.95214, 
    -30.85055, -31.74208, -32.62666, -33.50424, -34.37479, -35.23827, 
    -36.09467, -36.94396, -37.78615, -38.62124, -39.44924, -40.27016, 
    -41.08404, -41.89089, -42.69076, -43.48369, -44.26973,
  44.34454, 43.55843, 42.76536, 41.96529, 41.15818, 40.34399, 39.52269, 
    38.69425, 37.85865, 37.01588, 36.16594, 35.30883, 34.44456, 33.57316, 
    32.69466, 31.80908, 30.91648, 30.01692, 29.11047, 28.19719, 27.27719, 
    26.35056, 25.41741, 24.47786, 23.53204, 22.5801, 21.6222, 20.65849, 
    19.68916, 18.71439, 17.73438, 16.74936, 15.75952, 14.76512, 13.76639, 
    12.76358, 11.75696, 10.74679, 9.733348, 8.716929, 7.697824, 6.676331, 
    5.652757, 4.627412, 3.600614, 2.57268, 1.543934, 0.5146989, -0.5146989, 
    -1.543934, -2.57268, -3.600614, -4.627412, -5.652757, -6.676331, 
    -7.697824, -8.716929, -9.733348, -10.74679, -11.75696, -12.76358, 
    -13.76639, -14.76512, -15.75952, -16.74936, -17.73438, -18.71439, 
    -19.68916, -20.65849, -21.6222, -22.5801, -23.53204, -24.47786, 
    -25.41741, -26.35056, -27.27719, -28.19719, -29.11047, -30.01692, 
    -30.91648, -31.80908, -32.69466, -33.57316, -34.44456, -35.30883, 
    -36.16594, -37.01588, -37.85865, -38.69425, -39.52269, -40.34399, 
    -41.15818, -41.96529, -42.76536, -43.55843, -44.34454,
  44.41011, 43.62393, 42.83075, 42.03052, 41.22319, 40.40873, 39.58709, 
    38.75827, 37.92222, 37.07895, 36.22845, 35.37072, 34.50577, 33.63363, 
    32.75431, 31.86786, 30.97433, 30.07377, 29.16625, 28.25185, 27.33065, 
    26.40276, 25.46829, 24.52736, 23.58009, 22.62664, 21.66716, 20.70182, 
    19.7308, 18.75428, 17.77247, 16.78558, 15.79384, 14.79747, 13.79673, 
    12.79187, 11.78315, 10.77084, 9.755226, 8.736598, 7.715252, 6.691492, 
    5.665627, 4.63797, 3.608843, 2.578568, 1.54747, 0.5158784, -0.5158784, 
    -1.54747, -2.578568, -3.608843, -4.63797, -5.665627, -6.691492, 
    -7.715252, -8.736598, -9.755226, -10.77084, -11.78315, -12.79187, 
    -13.79673, -14.79747, -15.79384, -16.78558, -17.77247, -18.75428, 
    -19.7308, -20.70182, -21.66716, -22.62664, -23.58009, -24.52736, 
    -25.46829, -26.40276, -27.33065, -28.25185, -29.16625, -30.07377, 
    -30.97433, -31.86786, -32.75431, -33.63363, -34.50577, -35.37072, 
    -36.22845, -37.07895, -37.92222, -38.75827, -39.58709, -40.40873, 
    -41.22319, -42.03052, -42.83075, -43.62393, -44.41011,
  44.46639, 43.68016, 42.88689, 42.08652, 41.279, 40.46431, 39.6424, 
    38.81324, 37.97682, 37.13312, 36.28214, 35.42388, 34.55835, 33.68556, 
    32.80555, 31.91836, 31.02403, 30.12261, 29.21418, 28.29881, 27.3766, 
    26.44763, 25.51202, 24.5699, 23.62139, 22.66665, 21.70582, 20.73908, 
    19.7666, 18.78858, 17.80522, 16.81673, 15.82335, 14.8253, 13.82283, 
    12.8162, 11.80567, 10.79152, 9.774042, 8.753514, 7.730243, 6.704533, 
    5.676696, 4.647052, 3.615922, 2.583632, 1.550512, 0.5168929, -0.5168929, 
    -1.550512, -2.583632, -3.615922, -4.647052, -5.676696, -6.704533, 
    -7.730243, -8.753514, -9.774042, -10.79152, -11.80567, -12.8162, 
    -13.82283, -14.8253, -15.82335, -16.81673, -17.80522, -18.78858, 
    -19.7666, -20.73908, -21.70582, -22.66665, -23.62139, -24.5699, 
    -25.51202, -26.44763, -27.3766, -28.29881, -29.21418, -30.12261, 
    -31.02403, -31.91836, -32.80555, -33.68556, -34.55835, -35.42388, 
    -36.28214, -37.13312, -37.97682, -38.81324, -39.6424, -40.46431, -41.279, 
    -42.08652, -42.88689, -43.68016, -44.46639,
  44.51335, 43.72708, 42.93373, 42.13324, 41.32558, 40.51069, 39.68855, 
    38.85912, 38.02239, 37.17834, 36.32696, 35.46826, 34.60224, 33.72892, 
    32.84834, 31.96053, 31.06553, 30.1634, 29.25421, 28.33804, 27.41497, 
    26.4851, 25.54855, 24.60544, 23.6559, 22.70007, 21.73811, 20.7702, 
    19.79651, 18.81724, 17.83258, 16.84276, 15.84801, 14.84855, 13.84463, 
    12.83653, 11.8245, 10.80881, 9.789767, 8.767653, 7.742771, 6.715432, 
    5.685948, 4.654643, 3.621838, 2.587865, 1.553055, 0.5177408, -0.5177408, 
    -1.553055, -2.587865, -3.621838, -4.654643, -5.685948, -6.715432, 
    -7.742771, -8.767653, -9.789767, -10.80881, -11.8245, -12.83653, 
    -13.84463, -14.84855, -15.84801, -16.84276, -17.83258, -18.81724, 
    -19.79651, -20.7702, -21.73811, -22.70007, -23.6559, -24.60544, 
    -25.54855, -26.4851, -27.41497, -28.33804, -29.25421, -30.1634, 
    -31.06553, -31.96053, -32.84834, -33.72892, -34.60224, -35.46826, 
    -36.32696, -37.17834, -38.02239, -38.85912, -39.68855, -40.51069, 
    -41.32558, -42.13324, -42.93373, -43.72708, -44.51335,
  44.55096, 43.76466, 42.97124, 42.17067, 41.36288, 40.54784, 39.72552, 
    38.89588, 38.0589, 37.21456, 36.36287, 35.50381, 34.63741, 33.76367, 
    32.88263, 31.99432, 31.09879, 30.19609, 29.28629, 28.36947, 27.44572, 
    26.51514, 25.57783, 24.63392, 23.68355, 22.72686, 21.764, 20.79515, 
    19.82049, 18.84021, 17.85452, 16.86363, 15.86777, 14.86719, 13.86212, 
    12.85283, 11.83959, 10.82268, 9.802377, 8.77899, 7.752818, 6.724172, 
    5.693368, 4.660729, 3.626583, 2.59126, 1.555094, 0.5184209, -0.5184209, 
    -1.555094, -2.59126, -3.626583, -4.660729, -5.693368, -6.724172, 
    -7.752818, -8.77899, -9.802377, -10.82268, -11.83959, -12.85283, 
    -13.86212, -14.86719, -15.86777, -16.86363, -17.85452, -18.84021, 
    -19.82049, -20.79515, -21.764, -22.72686, -23.68355, -24.63392, 
    -25.57783, -26.51514, -27.44572, -28.36947, -29.28629, -30.19609, 
    -31.09879, -31.99432, -32.88263, -33.76367, -34.63741, -35.50381, 
    -36.36287, -37.21456, -38.0589, -38.89588, -39.72552, -40.54784, 
    -41.36288, -42.17067, -42.97124, -43.76466, -44.55096,
  44.57919, 43.79286, 42.9994, 42.19876, 41.39089, 40.57574, 39.75327, 
    38.92347, 38.0863, 37.24176, 36.38982, 35.53051, 34.66381, 33.78976, 
    32.90837, 32.01969, 31.12376, 30.22064, 29.31038, 28.39308, 27.46882, 
    26.5377, 25.59982, 24.65532, 23.70432, 22.74698, 21.78345, 20.81389, 
    19.8385, 18.85747, 17.871, 16.87931, 15.88263, 14.88119, 13.87526, 
    12.86508, 11.85093, 10.83309, 9.811852, 8.787509, 7.760367, 6.73074, 
    5.698944, 4.665304, 3.630148, 2.593811, 1.556626, 0.5189319, -0.5189319, 
    -1.556626, -2.593811, -3.630148, -4.665304, -5.698944, -6.73074, 
    -7.760367, -8.787509, -9.811852, -10.83309, -11.85093, -12.86508, 
    -13.87526, -14.88119, -15.88263, -16.87931, -17.871, -18.85747, -19.8385, 
    -20.81389, -21.78345, -22.74698, -23.70432, -24.65532, -25.59982, 
    -26.5377, -27.46882, -28.39308, -29.31038, -30.22064, -31.12376, 
    -32.01969, -32.90837, -33.78976, -34.66381, -35.53051, -36.38982, 
    -37.24176, -38.0863, -38.92347, -39.75327, -40.57574, -41.39089, 
    -42.19876, -42.9994, -43.79286, -44.57919,
  44.59801, 43.81168, 43.01819, 42.2175, 41.40957, 40.59435, 39.77179, 
    38.94188, 38.10459, 37.2599, 36.40781, 35.54832, 34.68143, 33.80717, 
    32.92555, 32.03662, 31.14043, 30.23702, 29.32646, 28.40884, 27.48424, 
    26.55275, 25.6145, 24.6696, 23.71819, 22.76041, 21.79643, 20.8264, 
    19.85053, 18.86899, 17.882, 16.88978, 15.89254, 14.89054, 13.88403, 
    12.87325, 11.8585, 10.84004, 9.818177, 8.793196, 7.765407, 6.735124, 
    5.702665, 4.668357, 3.632529, 2.595514, 1.557649, 0.519273, -0.519273, 
    -1.557649, -2.595514, -3.632529, -4.668357, -5.702665, -6.735124, 
    -7.765407, -8.793196, -9.818177, -10.84004, -11.8585, -12.87325, 
    -13.88403, -14.89054, -15.89254, -16.88978, -17.882, -18.86899, 
    -19.85053, -20.8264, -21.79643, -22.76041, -23.71819, -24.6696, -25.6145, 
    -26.55275, -27.48424, -28.40884, -29.32646, -30.23702, -31.14043, 
    -32.03662, -32.92555, -33.80717, -34.68143, -35.54832, -36.40781, 
    -37.2599, -38.10459, -38.94188, -39.77179, -40.59435, -41.40957, 
    -42.2175, -43.01819, -43.81168, -44.59801,
  44.60743, 43.82109, 43.02758, 42.22688, 41.41891, 40.60365, 39.78105, 
    38.95109, 38.11374, 37.26898, 36.41681, 35.55723, 34.69025, 33.81588, 
    32.93415, 32.04509, 31.14876, 30.24521, 29.33451, 28.41672, 27.49195, 
    26.56029, 25.62184, 24.67674, 23.72513, 22.76713, 21.80292, 20.83266, 
    19.85655, 18.87476, 17.88751, 16.89501, 15.8975, 14.89522, 13.88841, 
    12.87735, 11.86229, 10.84352, 9.821342, 8.796041, 7.767929, 6.737318, 
    5.704528, 4.669885, 3.63372, 2.596366, 1.55816, 0.5194437, -0.5194437, 
    -1.55816, -2.596366, -3.63372, -4.669885, -5.704528, -6.737318, 
    -7.767929, -8.796041, -9.821342, -10.84352, -11.86229, -12.87735, 
    -13.88841, -14.89522, -15.8975, -16.89501, -17.88751, -18.87476, 
    -19.85655, -20.83266, -21.80292, -22.76713, -23.72513, -24.67674, 
    -25.62184, -26.56029, -27.49195, -28.41672, -29.33451, -30.24521, 
    -31.14876, -32.04509, -32.93415, -33.81588, -34.69025, -35.55723, 
    -36.41681, -37.26898, -38.11374, -38.95109, -39.78105, -40.60365, 
    -41.41891, -42.22688, -43.02758, -43.82109, -44.60743,
  44.60743, 43.82109, 43.02758, 42.22688, 41.41891, 40.60365, 39.78105, 
    38.95109, 38.11374, 37.26898, 36.41681, 35.55723, 34.69025, 33.81588, 
    32.93415, 32.04509, 31.14876, 30.24521, 29.33451, 28.41672, 27.49195, 
    26.56029, 25.62184, 24.67674, 23.72513, 22.76713, 21.80292, 20.83266, 
    19.85655, 18.87476, 17.88751, 16.89501, 15.8975, 14.89522, 13.88841, 
    12.87735, 11.86229, 10.84352, 9.821342, 8.796041, 7.767929, 6.737318, 
    5.704528, 4.669885, 3.63372, 2.596366, 1.55816, 0.5194437, -0.5194437, 
    -1.55816, -2.596366, -3.63372, -4.669885, -5.704528, -6.737318, 
    -7.767929, -8.796041, -9.821342, -10.84352, -11.86229, -12.87735, 
    -13.88841, -14.89522, -15.8975, -16.89501, -17.88751, -18.87476, 
    -19.85655, -20.83266, -21.80292, -22.76713, -23.72513, -24.67674, 
    -25.62184, -26.56029, -27.49195, -28.41672, -29.33451, -30.24521, 
    -31.14876, -32.04509, -32.93415, -33.81588, -34.69025, -35.55723, 
    -36.41681, -37.26898, -38.11374, -38.95109, -39.78105, -40.60365, 
    -41.41891, -42.22688, -43.02758, -43.82109, -44.60743,
  44.59801, 43.81168, 43.01819, 42.2175, 41.40957, 40.59435, 39.77179, 
    38.94188, 38.10459, 37.2599, 36.40781, 35.54832, 34.68143, 33.80717, 
    32.92555, 32.03662, 31.14043, 30.23702, 29.32646, 28.40884, 27.48424, 
    26.55275, 25.6145, 24.6696, 23.71819, 22.76041, 21.79643, 20.8264, 
    19.85053, 18.86899, 17.882, 16.88978, 15.89254, 14.89054, 13.88403, 
    12.87325, 11.8585, 10.84004, 9.818177, 8.793196, 7.765407, 6.735124, 
    5.702665, 4.668357, 3.632529, 2.595514, 1.557649, 0.519273, -0.519273, 
    -1.557649, -2.595514, -3.632529, -4.668357, -5.702665, -6.735124, 
    -7.765407, -8.793196, -9.818177, -10.84004, -11.8585, -12.87325, 
    -13.88403, -14.89054, -15.89254, -16.88978, -17.882, -18.86899, 
    -19.85053, -20.8264, -21.79643, -22.76041, -23.71819, -24.6696, -25.6145, 
    -26.55275, -27.48424, -28.40884, -29.32646, -30.23702, -31.14043, 
    -32.03662, -32.92555, -33.80717, -34.68143, -35.54832, -36.40781, 
    -37.2599, -38.10459, -38.94188, -39.77179, -40.59435, -41.40957, 
    -42.2175, -43.01819, -43.81168, -44.59801,
  44.57919, 43.79286, 42.9994, 42.19876, 41.39089, 40.57574, 39.75327, 
    38.92347, 38.0863, 37.24176, 36.38982, 35.53051, 34.66381, 33.78976, 
    32.90837, 32.01969, 31.12376, 30.22064, 29.31038, 28.39308, 27.46882, 
    26.5377, 25.59982, 24.65532, 23.70432, 22.74698, 21.78345, 20.81389, 
    19.8385, 18.85747, 17.871, 16.87931, 15.88263, 14.88119, 13.87526, 
    12.86508, 11.85093, 10.83309, 9.811852, 8.787509, 7.760367, 6.73074, 
    5.698944, 4.665304, 3.630148, 2.593811, 1.556626, 0.5189319, -0.5189319, 
    -1.556626, -2.593811, -3.630148, -4.665304, -5.698944, -6.73074, 
    -7.760367, -8.787509, -9.811852, -10.83309, -11.85093, -12.86508, 
    -13.87526, -14.88119, -15.88263, -16.87931, -17.871, -18.85747, -19.8385, 
    -20.81389, -21.78345, -22.74698, -23.70432, -24.65532, -25.59982, 
    -26.5377, -27.46882, -28.39308, -29.31038, -30.22064, -31.12376, 
    -32.01969, -32.90837, -33.78976, -34.66381, -35.53051, -36.38982, 
    -37.24176, -38.0863, -38.92347, -39.75327, -40.57574, -41.39089, 
    -42.19876, -42.9994, -43.79286, -44.57919,
  44.55096, 43.76466, 42.97124, 42.17067, 41.36288, 40.54784, 39.72552, 
    38.89588, 38.0589, 37.21456, 36.36287, 35.50381, 34.63741, 33.76367, 
    32.88263, 31.99432, 31.09879, 30.19609, 29.28629, 28.36947, 27.44572, 
    26.51514, 25.57783, 24.63392, 23.68355, 22.72686, 21.764, 20.79515, 
    19.82049, 18.84021, 17.85452, 16.86363, 15.86777, 14.86719, 13.86212, 
    12.85283, 11.83959, 10.82268, 9.802377, 8.77899, 7.752818, 6.724172, 
    5.693368, 4.660729, 3.626583, 2.59126, 1.555094, 0.5184209, -0.5184209, 
    -1.555094, -2.59126, -3.626583, -4.660729, -5.693368, -6.724172, 
    -7.752818, -8.77899, -9.802377, -10.82268, -11.83959, -12.85283, 
    -13.86212, -14.86719, -15.86777, -16.86363, -17.85452, -18.84021, 
    -19.82049, -20.79515, -21.764, -22.72686, -23.68355, -24.63392, 
    -25.57783, -26.51514, -27.44572, -28.36947, -29.28629, -30.19609, 
    -31.09879, -31.99432, -32.88263, -33.76367, -34.63741, -35.50381, 
    -36.36287, -37.21456, -38.0589, -38.89588, -39.72552, -40.54784, 
    -41.36288, -42.17067, -42.97124, -43.76466, -44.55096,
  44.51335, 43.72708, 42.93373, 42.13324, 41.32558, 40.51069, 39.68855, 
    38.85912, 38.02239, 37.17834, 36.32696, 35.46826, 34.60224, 33.72892, 
    32.84834, 31.96053, 31.06553, 30.1634, 29.25421, 28.33804, 27.41497, 
    26.4851, 25.54855, 24.60544, 23.6559, 22.70007, 21.73811, 20.7702, 
    19.79651, 18.81724, 17.83258, 16.84276, 15.84801, 14.84855, 13.84463, 
    12.83653, 11.8245, 10.80881, 9.789767, 8.767653, 7.742771, 6.715432, 
    5.685948, 4.654643, 3.621838, 2.587865, 1.553055, 0.5177408, -0.5177408, 
    -1.553055, -2.587865, -3.621838, -4.654643, -5.685948, -6.715432, 
    -7.742771, -8.767653, -9.789767, -10.80881, -11.8245, -12.83653, 
    -13.84463, -14.84855, -15.84801, -16.84276, -17.83258, -18.81724, 
    -19.79651, -20.7702, -21.73811, -22.70007, -23.6559, -24.60544, 
    -25.54855, -26.4851, -27.41497, -28.33804, -29.25421, -30.1634, 
    -31.06553, -31.96053, -32.84834, -33.72892, -34.60224, -35.46826, 
    -36.32696, -37.17834, -38.02239, -38.85912, -39.68855, -40.51069, 
    -41.32558, -42.13324, -42.93373, -43.72708, -44.51335,
  44.46639, 43.68016, 42.88689, 42.08652, 41.279, 40.46431, 39.6424, 
    38.81324, 37.97682, 37.13312, 36.28214, 35.42388, 34.55835, 33.68556, 
    32.80555, 31.91836, 31.02403, 30.12261, 29.21418, 28.29881, 27.3766, 
    26.44763, 25.51202, 24.5699, 23.62139, 22.66665, 21.70582, 20.73908, 
    19.7666, 18.78858, 17.80522, 16.81673, 15.82335, 14.8253, 13.82283, 
    12.8162, 11.80567, 10.79152, 9.774042, 8.753514, 7.730243, 6.704533, 
    5.676696, 4.647052, 3.615922, 2.583632, 1.550512, 0.5168929, -0.5168929, 
    -1.550512, -2.583632, -3.615922, -4.647052, -5.676696, -6.704533, 
    -7.730243, -8.753514, -9.774042, -10.79152, -11.80567, -12.8162, 
    -13.82283, -14.8253, -15.82335, -16.81673, -17.80522, -18.78858, 
    -19.7666, -20.73908, -21.70582, -22.66665, -23.62139, -24.5699, 
    -25.51202, -26.44763, -27.3766, -28.29881, -29.21418, -30.12261, 
    -31.02403, -31.91836, -32.80555, -33.68556, -34.55835, -35.42388, 
    -36.28214, -37.13312, -37.97682, -38.81324, -39.6424, -40.46431, -41.279, 
    -42.08652, -42.88689, -43.68016, -44.46639,
  44.41011, 43.62393, 42.83075, 42.03052, 41.22319, 40.40873, 39.58709, 
    38.75827, 37.92222, 37.07895, 36.22845, 35.37072, 34.50577, 33.63363, 
    32.75431, 31.86786, 30.97433, 30.07377, 29.16625, 28.25185, 27.33065, 
    26.40276, 25.46829, 24.52736, 23.58009, 22.62664, 21.66716, 20.70182, 
    19.7308, 18.75428, 17.77247, 16.78558, 15.79384, 14.79747, 13.79673, 
    12.79187, 11.78315, 10.77084, 9.755226, 8.736598, 7.715252, 6.691492, 
    5.665627, 4.63797, 3.608843, 2.578568, 1.54747, 0.5158784, -0.5158784, 
    -1.54747, -2.578568, -3.608843, -4.63797, -5.665627, -6.691492, 
    -7.715252, -8.736598, -9.755226, -10.77084, -11.78315, -12.79187, 
    -13.79673, -14.79747, -15.79384, -16.78558, -17.77247, -18.75428, 
    -19.7308, -20.70182, -21.66716, -22.62664, -23.58009, -24.52736, 
    -25.46829, -26.40276, -27.33065, -28.25185, -29.16625, -30.07377, 
    -30.97433, -31.86786, -32.75431, -33.63363, -34.50577, -35.37072, 
    -36.22845, -37.07895, -37.92222, -38.75827, -39.58709, -40.40873, 
    -41.22319, -42.03052, -42.83075, -43.62393, -44.41011,
  44.34454, 43.55843, 42.76536, 41.96529, 41.15818, 40.34399, 39.52269, 
    38.69425, 37.85865, 37.01588, 36.16594, 35.30883, 34.44456, 33.57316, 
    32.69466, 31.80908, 30.91648, 30.01692, 29.11047, 28.19719, 27.27719, 
    26.35056, 25.41741, 24.47786, 23.53204, 22.5801, 21.6222, 20.65849, 
    19.68916, 18.71439, 17.73438, 16.74936, 15.75952, 14.76512, 13.76639, 
    12.76358, 11.75696, 10.74679, 9.733348, 8.716929, 7.697824, 6.676331, 
    5.652757, 4.627412, 3.600614, 2.57268, 1.543934, 0.5146989, -0.5146989, 
    -1.543934, -2.57268, -3.600614, -4.627412, -5.652757, -6.676331, 
    -7.697824, -8.716929, -9.733348, -10.74679, -11.75696, -12.76358, 
    -13.76639, -14.76512, -15.75952, -16.74936, -17.73438, -18.71439, 
    -19.68916, -20.65849, -21.6222, -22.5801, -23.53204, -24.47786, 
    -25.41741, -26.35056, -27.27719, -28.19719, -29.11047, -30.01692, 
    -30.91648, -31.80908, -32.69466, -33.57316, -34.44456, -35.30883, 
    -36.16594, -37.01588, -37.85865, -38.69425, -39.52269, -40.34399, 
    -41.15818, -41.96529, -42.76536, -43.55843, -44.34454,
  44.26973, 43.48369, 42.69076, 41.89089, 41.08404, 40.27016, 39.44924, 
    38.62124, 37.78615, 36.94396, 36.09467, 35.23827, 34.37479, 33.50424, 
    32.62666, 31.74208, 30.85055, 29.95214, 29.0469, 28.13491, 27.21628, 
    26.29108, 25.35944, 24.42147, 23.47731, 22.52709, 21.57098, 20.60913, 
    19.64173, 18.66896, 17.69101, 16.7081, 15.72045, 14.72828, 13.73184, 
    12.73137, 11.72714, 10.7194, 9.708443, 8.69454, 7.677984, 6.659072, 
    5.638107, 4.615394, 3.591246, 2.565979, 1.539908, 0.5133564, -0.5133564, 
    -1.539908, -2.565979, -3.591246, -4.615394, -5.638107, -6.659072, 
    -7.677984, -8.69454, -9.708443, -10.7194, -11.72714, -12.73137, 
    -13.73184, -14.72828, -15.72045, -16.7081, -17.69101, -18.66896, 
    -19.64173, -20.60913, -21.57098, -22.52709, -23.47731, -24.42147, 
    -25.35944, -26.29108, -27.21628, -28.13491, -29.0469, -29.95214, 
    -30.85055, -31.74208, -32.62666, -33.50424, -34.37479, -35.23827, 
    -36.09467, -36.94396, -37.78615, -38.62124, -39.44924, -40.27016, 
    -41.08404, -41.89089, -42.69076, -43.48369, -44.26973,
  44.18572, 43.39978, 42.60701, 41.80736, 41.0008, 40.18729, 39.3668, 
    38.53931, 37.7048, 36.86326, 36.01469, 35.15911, 34.29651, 33.42693, 
    32.55039, 31.66694, 30.77662, 29.87949, 28.97562, 28.06509, 27.14798, 
    26.2244, 25.29446, 24.35827, 23.41596, 22.46768, 21.51358, 20.55383, 
    19.58859, 18.61805, 17.64242, 16.66188, 15.67667, 14.68701, 13.69314, 
    12.6953, 11.69374, 10.68873, 9.680549, 8.669463, 7.655765, 6.639744, 
    5.6217, 4.601935, 3.580756, 2.558473, 1.535401, 0.511853, -0.511853, 
    -1.535401, -2.558473, -3.580756, -4.601935, -5.6217, -6.639744, 
    -7.655765, -8.669463, -9.680549, -10.68873, -11.69374, -12.6953, 
    -13.69314, -14.68701, -15.67667, -16.66188, -17.64242, -18.61805, 
    -19.58859, -20.55383, -21.51358, -22.46768, -23.41596, -24.35827, 
    -25.29446, -26.2244, -27.14798, -28.06509, -28.97562, -29.87949, 
    -30.77662, -31.66694, -32.55039, -33.42693, -34.29651, -35.15911, 
    -36.01469, -36.86326, -37.7048, -38.53931, -39.3668, -40.18729, -41.0008, 
    -41.80736, -42.60701, -43.39978, -44.18572,
  44.09258, 43.30674, 42.51416, 41.71477, 40.90854, 40.09544, 39.27544, 
    38.44851, 37.61465, 36.77385, 35.9261, 35.07141, 34.20981, 33.3413, 
    32.46593, 31.58372, 30.69475, 29.79905, 28.89671, 27.98779, 27.07239, 
    26.1506, 25.22254, 24.28832, 23.34808, 22.40195, 21.45008, 20.49264, 
    19.5298, 18.56174, 17.58866, 16.61077, 15.62826, 14.64138, 13.65034, 
    12.6554, 11.65681, 10.65482, 9.649706, 8.641738, 7.631198, 6.618376, 
    5.603562, 4.587056, 3.569159, 2.550177, 1.530417, 0.510191, -0.510191, 
    -1.530417, -2.550177, -3.569159, -4.587056, -5.603562, -6.618376, 
    -7.631198, -8.641738, -9.649706, -10.65482, -11.65681, -12.6554, 
    -13.65034, -14.64138, -15.62826, -16.61077, -17.58866, -18.56174, 
    -19.5298, -20.49264, -21.45008, -22.40195, -23.34808, -24.28832, 
    -25.22254, -26.1506, -27.07239, -27.98779, -28.89671, -29.79905, 
    -30.69475, -31.58372, -32.46593, -33.3413, -34.20981, -35.07141, 
    -35.9261, -36.77385, -37.61465, -38.44851, -39.27544, -40.09544, 
    -40.90854, -41.71477, -42.51416, -43.30674, -44.09258,
  43.99035, 43.20465, 42.41228, 41.61318, 40.80733, 39.99469, 39.17523, 
    38.34894, 37.5158, 36.67581, 35.82896, 34.97528, 34.11476, 33.24744, 
    32.37335, 31.49253, 30.60504, 29.71092, 28.81025, 27.90311, 26.98958, 
    26.06977, 25.14377, 24.21172, 23.27374, 22.32997, 21.38055, 20.42565, 
    19.46544, 18.50011, 17.52983, 16.55482, 15.57528, 14.59143, 13.60351, 
    12.61175, 11.6164, 10.61772, 9.615962, 8.611405, 7.604323, 6.594999, 
    5.58372, 4.570779, 3.556473, 2.541101, 1.524966, 0.5083731, -0.5083731, 
    -1.524966, -2.541101, -3.556473, -4.570779, -5.58372, -6.594999, 
    -7.604323, -8.611405, -9.615962, -10.61772, -11.6164, -12.61175, 
    -13.60351, -14.59143, -15.57528, -16.55482, -17.52983, -18.50011, 
    -19.46544, -20.42565, -21.38055, -22.32997, -23.27374, -24.21172, 
    -25.14377, -26.06977, -26.98958, -27.90311, -28.81025, -29.71092, 
    -30.60504, -31.49253, -32.37335, -33.24744, -34.11476, -34.97528, 
    -35.82896, -36.67581, -37.5158, -38.34894, -39.17523, -39.99469, 
    -40.80733, -41.61318, -42.41228, -43.20465, -43.99035,
  43.87911, 43.09357, 42.30143, 41.50267, 40.69724, 39.88511, 39.06625, 
    38.24066, 37.40832, 36.56922, 35.72337, 34.87078, 34.01146, 33.14545, 
    32.27277, 31.39346, 30.50758, 29.61518, 28.71634, 27.81114, 26.89966, 
    25.98199, 25.05826, 24.12856, 23.19304, 22.25184, 21.30509, 20.35295, 
    19.39561, 18.43323, 17.466, 16.49412, 15.5178, 14.53725, 13.55271, 
    12.5644, 11.57257, 10.57748, 9.579368, 8.578511, 7.57518, 6.56965, 
    5.562205, 4.55313, 3.542717, 2.53126, 1.519056, 0.5064019, -0.5064019, 
    -1.519056, -2.53126, -3.542717, -4.55313, -5.562205, -6.56965, -7.57518, 
    -8.578511, -9.579368, -10.57748, -11.57257, -12.5644, -13.55271, 
    -14.53725, -15.5178, -16.49412, -17.466, -18.43323, -19.39561, -20.35295, 
    -21.30509, -22.25184, -23.19304, -24.12856, -25.05826, -25.98199, 
    -26.89966, -27.81114, -28.71634, -29.61518, -30.50758, -31.39346, 
    -32.27277, -33.14545, -34.01146, -34.87078, -35.72337, -36.56922, 
    -37.40832, -38.24066, -39.06625, -39.88511, -40.69724, -41.50267, 
    -42.30143, -43.09357, -43.87911,
  43.75893, 42.97356, 42.18171, 41.38331, 40.57834, 39.76678, 38.94859, 
    38.12377, 37.2923, 36.45418, 35.60942, 34.75802, 33.90001, 33.03541, 
    32.16426, 31.28659, 30.40247, 29.51195, 28.6151, 27.71199, 26.80272, 
    25.88738, 24.96609, 24.03895, 23.10609, 22.16766, 21.22379, 20.27464, 
    19.32038, 18.36119, 17.39725, 16.42875, 15.4559, 14.47891, 13.49801, 
    12.51342, 11.52539, 10.53416, 9.539974, 8.543103, 7.54381, 6.542367, 
    5.539048, 4.534135, 3.527913, 2.52067, 1.512695, 0.5042805, -0.5042805, 
    -1.512695, -2.52067, -3.527913, -4.534135, -5.539048, -6.542367, 
    -7.54381, -8.543103, -9.539974, -10.53416, -11.52539, -12.51342, 
    -13.49801, -14.47891, -15.4559, -16.42875, -17.39725, -18.36119, 
    -19.32038, -20.27464, -21.22379, -22.16766, -23.10609, -24.03895, 
    -24.96609, -25.88738, -26.80272, -27.71199, -28.6151, -29.51195, 
    -30.40247, -31.28659, -32.16426, -33.03541, -33.90001, -34.75802, 
    -35.60942, -36.45418, -37.2923, -38.12377, -38.94859, -39.76678, 
    -40.57834, -41.38331, -42.18171, -42.97356, -43.75893,
  43.62987, 42.84472, 42.05317, 41.25519, 40.45074, 39.63979, 38.82234, 
    37.99836, 37.16784, 36.33079, 35.48721, 34.6371, 33.78051, 32.91744, 
    32.04794, 31.17205, 30.28983, 29.40132, 28.50661, 27.60576, 26.69888, 
    25.78605, 24.86737, 23.94298, 23.01299, 22.07753, 21.13675, 20.19081, 
    19.23986, 18.28409, 17.32367, 16.3588, 15.38967, 14.4165, 13.43949, 
    12.45889, 11.47492, 10.48782, 9.49784, 8.505234, 7.510261, 6.513187, 
    5.514283, 4.513822, 3.512082, 2.509345, 1.505893, 0.502012, -0.502012, 
    -1.505893, -2.509345, -3.512082, -4.513822, -5.514283, -6.513187, 
    -7.510261, -8.505234, -9.49784, -10.48782, -11.47492, -12.45889, 
    -13.43949, -14.4165, -15.38967, -16.3588, -17.32367, -18.28409, 
    -19.23986, -20.19081, -21.13675, -22.07753, -23.01299, -23.94298, 
    -24.86737, -25.78605, -26.69888, -27.60576, -28.50661, -29.40132, 
    -30.28983, -31.17205, -32.04794, -32.91744, -33.78051, -34.6371, 
    -35.48721, -36.33079, -37.16784, -37.99836, -38.82234, -39.63979, 
    -40.45074, -41.25519, -42.05317, -42.84472, -43.62987,
  43.49203, 42.70713, 41.91592, 41.1184, 40.31451, 39.50425, 38.6876, 
    37.86452, 37.03504, 36.19914, 35.35684, 34.50814, 33.65307, 32.79165, 
    31.92393, 31.04995, 30.16976, 29.28342, 28.391, 27.49258, 26.58825, 
    25.6781, 24.76223, 23.84077, 22.91384, 21.98156, 21.04409, 20.10156, 
    19.15416, 18.20203, 17.24537, 16.28436, 15.3192, 14.35008, 13.37724, 
    12.40088, 11.42123, 10.43853, 9.453025, 8.464956, 7.47458, 6.482156, 
    5.487947, 4.49222, 3.495247, 2.497301, 1.49866, 0.4995998, -0.4995998, 
    -1.49866, -2.497301, -3.495247, -4.49222, -5.487947, -6.482156, -7.47458, 
    -8.464956, -9.453025, -10.43853, -11.42123, -12.40088, -13.37724, 
    -14.35008, -15.3192, -16.28436, -17.24537, -18.20203, -19.15416, 
    -20.10156, -21.04409, -21.98156, -22.91384, -23.84077, -24.76223, 
    -25.6781, -26.58825, -27.49258, -28.391, -29.28342, -30.16976, -31.04995, 
    -31.92393, -32.79165, -33.65307, -34.50814, -35.35684, -36.19914, 
    -37.03504, -37.86452, -38.6876, -39.50425, -40.31451, -41.1184, 
    -41.91592, -42.70713, -43.49203,
  43.34549, 42.56086, 41.77005, 40.97303, 40.16977, 39.36025, 38.54446, 
    37.72238, 36.89401, 36.05936, 35.21843, 34.37123, 33.5178, 32.65816, 
    31.79235, 30.92041, 30.04239, 29.15837, 28.2684, 27.37256, 26.47095, 
    25.56366, 24.65079, 23.73245, 22.80877, 21.87987, 20.94591, 20.00702, 
    19.06337, 18.11512, 17.16244, 16.20553, 15.24457, 14.27977, 13.31133, 
    12.33946, 11.3644, 10.38636, 9.40559, 8.422327, 7.436818, 6.449316, 
    5.460076, 4.46936, 3.477432, 2.484558, 1.491006, 0.4970472, -0.4970472, 
    -1.491006, -2.484558, -3.477432, -4.46936, -5.460076, -6.449316, 
    -7.436818, -8.422327, -9.40559, -10.38636, -11.3644, -12.33946, 
    -13.31133, -14.27977, -15.24457, -16.20553, -17.16244, -18.11512, 
    -19.06337, -20.00702, -20.94591, -21.87987, -22.80877, -23.73245, 
    -24.65079, -25.56366, -26.47095, -27.37256, -28.2684, -29.15837, 
    -30.04239, -30.92041, -31.79235, -32.65816, -33.5178, -34.37123, 
    -35.21843, -36.05936, -36.89401, -37.72238, -38.54446, -39.36025, 
    -40.16977, -40.97303, -41.77005, -42.56086, -43.34549,
  43.19033, 42.40602, 41.61564, 40.81918, 40.0166, 39.20789, 38.39304, 
    37.57203, 36.74487, 35.91155, 35.0721, 34.22652, 33.37484, 32.51709, 
    31.65331, 30.78355, 29.90785, 29.02629, 28.13892, 27.24584, 26.34712, 
    25.44285, 24.53315, 23.61813, 22.69789, 21.77258, 20.84233, 19.90729, 
    18.96761, 18.02345, 17.075, 16.12242, 15.1659, 14.20564, 13.24185, 
    12.27472, 11.30449, 10.33138, 9.355601, 8.377405, 7.397027, 6.414712, 
    5.430711, 4.445276, 3.458663, 2.471131, 1.482942, 0.494358, -0.494358, 
    -1.482942, -2.471131, -3.458663, -4.445276, -5.430711, -6.414712, 
    -7.397027, -8.377405, -9.355601, -10.33138, -11.30449, -12.27472, 
    -13.24185, -14.20564, -15.1659, -16.12242, -17.075, -18.02345, -18.96761, 
    -19.90729, -20.84233, -21.77258, -22.69789, -23.61813, -24.53315, 
    -25.44285, -26.34712, -27.24584, -28.13892, -29.02629, -29.90785, 
    -30.78355, -31.65331, -32.51709, -33.37484, -34.22652, -35.0721, 
    -35.91155, -36.74487, -37.57203, -38.39304, -39.20789, -40.0166, 
    -40.81918, -41.61564, -42.40602, -43.19033,
  43.02665, 42.24269, 41.4528, 40.65696, 39.85512, 39.04729, 38.23346, 
    37.4136, 36.58773, 35.75585, 34.91797, 34.07411, 33.2243, 32.36856, 
    31.50695, 30.6395, 29.76627, 28.88731, 28.00271, 27.11254, 26.21687, 
    25.31582, 24.40947, 23.49794, 22.58134, 21.65982, 20.73348, 19.8025, 
    18.867, 17.92716, 16.98314, 16.03511, 15.08327, 14.1278, 13.16889, 
    12.20676, 11.2416, 10.27365, 9.303126, 8.330251, 7.355261, 6.378393, 
    5.399891, 4.419998, 3.438965, 2.457041, 1.47448, 0.4915359, -0.4915359, 
    -1.47448, -2.457041, -3.438965, -4.419998, -5.399891, -6.378393, 
    -7.355261, -8.330251, -9.303126, -10.27365, -11.2416, -12.20676, 
    -13.16889, -14.1278, -15.08327, -16.03511, -16.98314, -17.92716, -18.867, 
    -19.8025, -20.73348, -21.65982, -22.58134, -23.49794, -24.40947, 
    -25.31582, -26.21687, -27.11254, -28.00271, -28.88731, -29.76627, 
    -30.6395, -31.50695, -32.36856, -33.2243, -34.07411, -34.91797, 
    -35.75585, -36.58773, -37.4136, -38.23346, -39.04729, -39.85512, 
    -40.65696, -41.4528, -42.24269, -43.02665,
  42.85454, 42.07099, 41.28164, 40.48646, 39.68544, 38.87856, 38.06581, 
    37.2472, 36.42271, 35.59236, 34.75616, 33.91414, 33.06631, 32.21272, 
    31.3534, 30.4884, 29.61777, 28.74158, 27.8599, 26.9728, 26.08036, 
    25.18268, 24.27987, 23.37202, 22.45926, 21.5417, 20.61949, 19.69276, 
    18.76166, 17.82635, 16.88698, 15.94374, 14.99679, 14.04633, 13.09255, 
    12.13564, 11.17581, 10.21327, 9.248235, 8.280929, 7.311576, 6.340407, 
    5.367657, 4.393563, 3.418365, 2.442306, 1.46563, 0.4885846, -0.4885846, 
    -1.46563, -2.442306, -3.418365, -4.393563, -5.367657, -6.340407, 
    -7.311576, -8.280929, -9.248235, -10.21327, -11.17581, -12.13564, 
    -13.09255, -14.04633, -14.99679, -15.94374, -16.88698, -17.82635, 
    -18.76166, -19.69276, -20.61949, -21.5417, -22.45926, -23.37202, 
    -24.27987, -25.18268, -26.08036, -26.9728, -27.8599, -28.74158, 
    -29.61777, -30.4884, -31.3534, -32.21272, -33.06631, -33.91414, 
    -34.75616, -35.59236, -36.42271, -37.2472, -38.06581, -38.87856, 
    -39.68544, -40.48646, -41.28164, -42.07099, -42.85454,
  42.67411, 41.89101, 41.10225, 40.30781, 39.50767, 38.70182, 37.89024, 
    37.07295, 36.24994, 35.42123, 34.58682, 33.74675, 32.90103, 32.0497, 
    31.19281, 30.3304, 29.46252, 28.58924, 27.71063, 26.82676, 25.93772, 
    25.04359, 24.14449, 23.2405, 22.33176, 21.41838, 20.50048, 19.57821, 
    18.65171, 17.72114, 16.78664, 15.8484, 14.90658, 13.96135, 13.01292, 
    12.06147, 11.10719, 10.1503, 9.190996, 8.229501, 7.266029, 6.300805, 
    5.334054, 4.366004, 3.39689, 2.426945, 1.456406, 0.4855082, -0.4855082, 
    -1.456406, -2.426945, -3.39689, -4.366004, -5.334054, -6.300805, 
    -7.266029, -8.229501, -9.190996, -10.1503, -11.10719, -12.06147, 
    -13.01292, -13.96135, -14.90658, -15.8484, -16.78664, -17.72114, 
    -18.65171, -19.57821, -20.50048, -21.41838, -22.33176, -23.2405, 
    -24.14449, -25.04359, -25.93772, -26.82676, -27.71063, -28.58924, 
    -29.46252, -30.3304, -31.19281, -32.0497, -32.90103, -33.74675, 
    -34.58682, -35.42123, -36.24994, -37.07295, -37.89024, -38.70182, 
    -39.50767, -40.30781, -41.10225, -41.89101, -42.67411,
  42.48545, 41.70287, 40.91476, 40.12112, 39.32193, 38.51718, 37.70687, 
    36.891, 36.06956, 35.24258, 34.41008, 33.57207, 32.72858, 31.87964, 
    31.02531, 30.16563, 29.30065, 28.43043, 27.55505, 26.67457, 25.78909, 
    24.89869, 24.00347, 23.10353, 22.19899, 21.28997, 20.37659, 19.45897, 
    18.53728, 17.61165, 16.68224, 15.74921, 14.81272, 13.87296, 12.9301, 
    11.98433, 11.03584, 10.08482, 9.131484, 8.176033, 7.218679, 6.259636, 
    5.299122, 4.337358, 3.374569, 2.41098, 1.446817, 0.4823107, -0.4823107, 
    -1.446817, -2.41098, -3.374569, -4.337358, -5.299122, -6.259636, 
    -7.218679, -8.176033, -9.131484, -10.08482, -11.03584, -11.98433, 
    -12.9301, -13.87296, -14.81272, -15.74921, -16.68224, -17.61165, 
    -18.53728, -19.45897, -20.37659, -21.28997, -22.19899, -23.10353, 
    -24.00347, -24.89869, -25.78909, -26.67457, -27.55505, -28.43043, 
    -29.30065, -30.16563, -31.02531, -31.87964, -32.72858, -33.57207, 
    -34.41008, -35.24258, -36.06956, -36.891, -37.70687, -38.51718, 
    -39.32193, -40.12112, -40.91476, -41.70287, -42.48545,
  42.28868, 41.50666, 40.71927, 39.9265, 39.12834, 38.32478, 37.51582, 
    36.70145, 35.8817, 35.05656, 34.22607, 33.39024, 32.5491, 31.70269, 
    30.85106, 29.99424, 29.1323, 28.2653, 27.3933, 26.51638, 25.63463, 
    24.74813, 23.85697, 22.96125, 22.0611, 21.15662, 20.24794, 19.33519, 
    18.4185, 17.49802, 16.57389, 15.64629, 14.71535, 13.78126, 12.84419, 
    11.90432, 10.96183, 10.01692, 9.069772, 8.120593, 7.169584, 6.216953, 
    5.262908, 4.307662, 3.35143, 2.394429, 1.436878, 0.478996, -0.478996, 
    -1.436878, -2.394429, -3.35143, -4.307662, -5.262908, -6.216953, 
    -7.169584, -8.120593, -9.069772, -10.01692, -10.96183, -11.90432, 
    -12.84419, -13.78126, -14.71535, -15.64629, -16.57389, -17.49802, 
    -18.4185, -19.33519, -20.24794, -21.15662, -22.0611, -22.96125, 
    -23.85697, -24.74813, -25.63463, -26.51638, -27.3933, -28.2653, -29.1323, 
    -29.99424, -30.85106, -31.70269, -32.5491, -33.39024, -34.22607, 
    -35.05656, -35.8817, -36.70145, -37.51582, -38.32478, -39.12834, 
    -39.9265, -40.71927, -41.50666, -42.28868,
  42.08391, 41.30251, 40.51591, 39.72409, 38.92703, 38.12474, 37.31722, 
    36.50447, 35.68649, 34.86331, 34.03494, 33.20141, 32.36275, 31.519, 
    30.6702, 29.81639, 28.95764, 28.094, 27.22555, 26.35234, 25.47448, 
    24.59204, 23.70512, 22.81381, 21.91823, 21.01848, 20.11469, 19.20699, 
    18.2955, 17.38036, 16.46173, 15.53974, 14.61457, 13.68636, 12.75529, 
    11.82154, 10.88527, 9.946671, 9.005934, 8.063247, 7.118805, 6.172808, 
    5.225454, 4.27695, 3.3275, 2.377314, 1.4266, 0.4755684, -0.4755684, 
    -1.4266, -2.377314, -3.3275, -4.27695, -5.225454, -6.172808, -7.118805, 
    -8.063247, -9.005934, -9.946671, -10.88527, -11.82154, -12.75529, 
    -13.68636, -14.61457, -15.53974, -16.46173, -17.38036, -18.2955, 
    -19.20699, -20.11469, -21.01848, -21.91823, -22.81381, -23.70512, 
    -24.59204, -25.47448, -26.35234, -27.22555, -28.094, -28.95764, 
    -29.81639, -30.6702, -31.519, -32.36275, -33.20141, -34.03494, -34.86331, 
    -35.68649, -36.50447, -37.31722, -38.12474, -38.92703, -39.72409, 
    -40.51591, -41.30251, -42.08391,
  41.87124, 41.09053, 40.30479, 39.51399, 38.71813, 37.9172, 37.11122, 
    36.30017, 35.48409, 34.66297, 33.83684, 33.00574, 32.16968, 31.32872, 
    30.48288, 29.63223, 28.77681, 27.91669, 27.05193, 26.18261, 25.3088, 
    24.43059, 23.54808, 22.66135, 21.77052, 20.87569, 19.97698, 19.07451, 
    18.16841, 17.25882, 16.34587, 15.42971, 14.51049, 13.58837, 12.66351, 
    11.73607, 10.80623, 9.874163, 8.940046, 8.004064, 7.066403, 6.127254, 
    5.186808, 4.245261, 3.30281, 2.359655, 1.415995, 0.472032, -0.472032, 
    -1.415995, -2.359655, -3.30281, -4.245261, -5.186808, -6.127254, 
    -7.066403, -8.004064, -8.940046, -9.874163, -10.80623, -11.73607, 
    -12.66351, -13.58837, -14.51049, -15.42971, -16.34587, -17.25882, 
    -18.16841, -19.07451, -19.97698, -20.87569, -21.77052, -22.66135, 
    -23.54808, -24.43059, -25.3088, -26.18261, -27.05193, -27.91669, 
    -28.77681, -29.63223, -30.48288, -31.32872, -32.16968, -33.00574, 
    -33.83684, -34.66297, -35.48409, -36.30017, -37.11122, -37.9172, 
    -38.71813, -39.51399, -40.30479, -41.09053, -41.87124,
  41.65079, 40.87085, 40.08604, 39.29634, 38.50176, 37.70229, 36.89794, 
    36.08871, 35.27462, 34.45568, 33.63192, 32.80336, 31.97004, 31.132, 
    30.28927, 29.44192, 28.58998, 27.73353, 26.87262, 26.00734, 25.13775, 
    24.26394, 23.386, 22.50403, 21.61812, 20.72838, 19.83493, 18.93789, 
    18.03736, 17.1335, 16.22643, 15.31629, 14.40323, 13.48739, 12.56893, 
    11.64802, 10.72481, 9.799476, 8.872184, 7.943112, 7.012438, 6.080344, 
    5.147013, 4.212631, 3.277388, 2.341473, 1.405076, 0.4683909, -0.4683909, 
    -1.405076, -2.341473, -3.277388, -4.212631, -5.147013, -6.080344, 
    -7.012438, -7.943112, -8.872184, -9.799476, -10.72481, -11.64802, 
    -12.56893, -13.48739, -14.40323, -15.31629, -16.22643, -17.1335, 
    -18.03736, -18.93789, -19.83493, -20.72838, -21.61812, -22.50403, 
    -23.386, -24.26394, -25.13775, -26.00734, -26.87262, -27.73353, 
    -28.58998, -29.44192, -30.28927, -31.132, -31.97004, -32.80336, 
    -33.63192, -34.45568, -35.27462, -36.08871, -36.89794, -37.70229, 
    -38.50176, -39.29634, -40.08604, -40.87085, -41.65079,
  41.42268, 40.64358, 39.85978, 39.07127, 38.27806, 37.48015, 36.67753, 
    35.87022, 35.05824, 34.2416, 33.42032, 32.59444, 31.76398, 30.929, 
    30.08952, 29.2456, 28.3973, 27.54466, 26.68777, 25.82668, 24.96147, 
    24.09223, 23.21904, 22.34199, 21.46118, 20.57672, 19.68871, 18.79726, 
    17.9025, 17.00456, 16.10355, 15.19962, 14.2929, 13.38354, 12.47168, 
    11.55748, 10.6411, 9.722692, 8.802423, 7.880459, 6.956971, 6.032131, 
    5.106114, 4.179099, 3.251263, 2.322789, 1.393856, 0.4646493, -0.4646493, 
    -1.393856, -2.322789, -3.251263, -4.179099, -5.106114, -6.032131, 
    -6.956971, -7.880459, -8.802423, -9.722692, -10.6411, -11.55748, 
    -12.47168, -13.38354, -14.2929, -15.19962, -16.10355, -17.00456, 
    -17.9025, -18.79726, -19.68871, -20.57672, -21.46118, -22.34199, 
    -23.21904, -24.09223, -24.96147, -25.82668, -26.68777, -27.54466, 
    -28.3973, -29.2456, -30.08952, -30.929, -31.76398, -32.59444, -33.42032, 
    -34.2416, -35.05824, -35.87022, -36.67753, -37.48015, -38.27806, 
    -39.07127, -39.85978, -40.64358, -41.42268,
  41.18702, 40.40884, 39.62614, 38.83891, 38.04717, 37.2509, 36.45013, 
    35.64485, 34.83509, 34.02087, 33.2022, 32.37912, 31.55167, 30.71988, 
    29.88379, 29.04346, 28.19893, 27.35027, 26.49753, 25.6408, 24.78014, 
    23.91562, 23.04734, 22.17539, 21.29985, 20.42083, 19.53844, 18.65277, 
    17.76396, 16.87211, 15.97735, 15.07981, 14.17962, 13.27692, 12.37185, 
    11.46456, 10.55519, 9.643898, 8.730841, 7.816175, 6.900063, 5.982669, 
    5.064158, 4.144701, 3.224465, 2.303623, 1.382348, 0.4608116, -0.4608116, 
    -1.382348, -2.303623, -3.224465, -4.144701, -5.064158, -5.982669, 
    -6.900063, -7.816175, -8.730841, -9.643898, -10.55519, -11.46456, 
    -12.37185, -13.27692, -14.17962, -15.07981, -15.97735, -16.87211, 
    -17.76396, -18.65277, -19.53844, -20.42083, -21.29985, -22.17539, 
    -23.04734, -23.91562, -24.78014, -25.6408, -26.49753, -27.35027, 
    -28.19893, -29.04346, -29.88379, -30.71988, -31.55167, -32.37912, 
    -33.2022, -34.02087, -34.83509, -35.64485, -36.45013, -37.2509, 
    -38.04717, -38.83891, -39.62614, -40.40884, -41.18702,
  40.94394, 40.16676, 39.38524, 38.5994, 37.80922, 37.01471, 36.21589, 
    35.41275, 34.60533, 33.79364, 32.97771, 32.15757, 31.33325, 30.50479, 
    29.67224, 28.83563, 27.99503, 27.1505, 26.30208, 25.44986, 24.5939, 
    23.73428, 22.87107, 22.00438, 21.13428, 20.26088, 19.38427, 18.50457, 
    17.62187, 16.73629, 15.84795, 14.95698, 14.0635, 13.16765, 12.26954, 
    11.36934, 10.46716, 9.563174, 8.657512, 7.750327, 6.841775, 5.93201, 
    5.02119, 4.109474, 3.197022, 2.283998, 1.370563, 0.4568816, -0.4568816, 
    -1.370563, -2.283998, -3.197022, -4.109474, -5.02119, -5.93201, 
    -6.841775, -7.750327, -8.657512, -9.563174, -10.46716, -11.36934, 
    -12.26954, -13.16765, -14.0635, -14.95698, -15.84795, -16.73629, 
    -17.62187, -18.50457, -19.38427, -20.26088, -21.13428, -22.00438, 
    -22.87107, -23.73428, -24.5939, -25.44986, -26.30208, -27.1505, 
    -27.99503, -28.83563, -29.67224, -30.50479, -31.33325, -32.15757, 
    -32.97771, -33.79364, -34.60533, -35.41275, -36.21589, -37.01471, 
    -37.80922, -38.5994, -39.38524, -40.16676, -40.94394,
  40.69355, 39.91746, 39.13723, 38.35286, 37.56434, 36.7717, 35.97494, 
    35.17407, 34.36911, 33.56009, 32.74702, 31.92994, 31.10889, 30.28391, 
    29.45502, 28.6223, 27.78577, 26.94551, 26.10157, 25.25401, 24.40292, 
    23.54835, 22.69039, 21.82912, 20.96463, 20.09701, 19.22636, 18.35277, 
    17.47636, 16.59723, 15.71549, 14.83126, 13.94467, 13.05583, 12.16487, 
    11.27192, 10.37712, 9.480604, 8.582511, 7.682984, 6.782168, 5.880208, 
    4.977254, 4.073455, 3.168964, 2.263932, 1.358514, 0.4528638, -0.4528638, 
    -1.358514, -2.263932, -3.168964, -4.073455, -4.977254, -5.880208, 
    -6.782168, -7.682984, -8.582511, -9.480604, -10.37712, -11.27192, 
    -12.16487, -13.05583, -13.94467, -14.83126, -15.71549, -16.59723, 
    -17.47636, -18.35277, -19.22636, -20.09701, -20.96463, -21.82912, 
    -22.69039, -23.54835, -24.40292, -25.25401, -26.10157, -26.94551, 
    -27.78577, -28.6223, -29.45502, -30.28391, -31.10889, -31.92994, 
    -32.74702, -33.56009, -34.36911, -35.17407, -35.97494, -36.7717, 
    -37.56434, -38.35286, -39.13723, -39.91746, -40.69355,
  40.43598, 39.66107, 38.88222, 38.09942, 37.31269, 36.52202, 35.72744, 
    34.92895, 34.12658, 33.32034, 32.51027, 31.6964, 30.87876, 30.05738, 
    29.23232, 28.40361, 27.57131, 26.73548, 25.89616, 25.05343, 24.20735, 
    23.35799, 22.50543, 21.64975, 20.79103, 19.92936, 19.06483, 18.19754, 
    17.32758, 16.45506, 15.58009, 14.70277, 13.82323, 12.94157, 12.05792, 
    11.1724, 10.28514, 9.396269, 8.505915, 7.614214, 6.721301, 5.827315, 
    4.932395, 4.036681, 3.140318, 2.243447, 1.346213, 0.448762, -0.448762, 
    -1.346213, -2.243447, -3.140318, -4.036681, -4.932395, -5.827315, 
    -6.721301, -7.614214, -8.505915, -9.396269, -10.28514, -11.1724, 
    -12.05792, -12.94157, -13.82323, -14.70277, -15.58009, -16.45506, 
    -17.32758, -18.19754, -19.06483, -19.92936, -20.79103, -21.64975, 
    -22.50543, -23.35799, -24.20735, -25.05343, -25.89616, -26.73548, 
    -27.57131, -28.40361, -29.23232, -30.05738, -30.87876, -31.6964, 
    -32.51027, -33.32034, -34.12658, -34.92895, -35.72744, -36.52202, 
    -37.31269, -38.09942, -38.88222, -39.66107, -40.43598,
  40.17135, 39.39772, 38.62035, 37.83924, 37.05439, 36.26581, 35.47353, 
    34.67754, 33.87788, 33.07457, 32.26763, 31.45709, 30.643, 29.82537, 
    29.00427, 28.17974, 27.35181, 26.52055, 25.68602, 24.84826, 24.00736, 
    23.16337, 22.31637, 21.46644, 20.61365, 19.75808, 18.89984, 18.03899, 
    17.17565, 16.30991, 15.44186, 14.57162, 13.69929, 12.82498, 11.9488, 
    11.07087, 10.19132, 9.31025, 8.427797, 7.544083, 6.659235, 5.773382, 
    4.886656, 3.999188, 3.111113, 2.222563, 1.333673, 0.4445804, -0.4445804, 
    -1.333673, -2.222563, -3.111113, -3.999188, -4.886656, -5.773382, 
    -6.659235, -7.544083, -8.427797, -9.31025, -10.19132, -11.07087, 
    -11.9488, -12.82498, -13.69929, -14.57162, -15.44186, -16.30991, 
    -17.17565, -18.03899, -18.89984, -19.75808, -20.61365, -21.46644, 
    -22.31637, -23.16337, -24.00736, -24.84826, -25.68602, -26.52055, 
    -27.35181, -28.17974, -29.00427, -29.82537, -30.643, -31.45709, 
    -32.26763, -33.07457, -33.87788, -34.67754, -35.47353, -36.26581, 
    -37.05439, -37.83924, -38.62035, -39.39772, -40.17135,
  39.89979, 39.12755, 38.35176, 37.57244, 36.78959, 36.00322, 35.21335, 
    34.42, 33.62318, 32.82292, 32.01924, 31.21218, 30.40177, 29.58805, 
    28.77106, 27.95084, 27.12744, 26.30091, 25.4713, 24.63868, 23.8031, 
    22.96464, 22.12335, 21.27932, 20.43262, 19.58332, 18.73152, 17.87728, 
    17.02072, 16.1619, 15.30094, 14.43793, 13.57297, 12.70616, 11.83762, 
    10.96744, 10.09574, 9.222629, 8.34823, 7.472656, 6.596026, 5.718461, 
    4.840082, 3.961012, 3.081377, 2.201299, 1.320906, 0.4403231, -0.4403231, 
    -1.320906, -2.201299, -3.081377, -3.961012, -4.840082, -5.718461, 
    -6.596026, -7.472656, -8.34823, -9.222629, -10.09574, -10.96744, 
    -11.83762, -12.70616, -13.57297, -14.43793, -15.30094, -16.1619, 
    -17.02072, -17.87728, -18.73152, -19.58332, -20.43262, -21.27932, 
    -22.12335, -22.96464, -23.8031, -24.63868, -25.4713, -26.30091, 
    -27.12744, -27.95084, -28.77106, -29.58805, -30.40177, -31.21218, 
    -32.01924, -32.82292, -33.62318, -34.42, -35.21335, -36.00322, -36.78959, 
    -37.57244, -38.35176, -39.12755, -39.89979,
  39.62142, 38.85067, 38.07658, 37.29916, 36.51843, 35.73439, 34.94707, 
    34.15647, 33.36263, 32.56555, 31.76528, 30.96183, 30.15525, 29.34557, 
    28.53283, 27.71707, 26.89834, 26.07669, 25.25217, 24.42483, 23.59474, 
    22.76195, 21.92654, 21.08856, 20.2481, 19.40522, 18.56001, 17.71254, 
    16.8629, 16.01117, 15.15745, 14.30182, 13.44438, 12.58523, 11.72446, 
    10.86218, 9.998483, 9.133484, 8.267286, 7.4, 6.531734, 5.662601, 
    4.792715, 3.922188, 3.051136, 2.179676, 1.307923, 0.4359938, -0.4359938, 
    -1.307923, -2.179676, -3.051136, -3.922188, -4.792715, -5.662601, 
    -6.531734, -7.4, -8.267286, -9.133484, -9.998483, -10.86218, -11.72446, 
    -12.58523, -13.44438, -14.30182, -15.15745, -16.01117, -16.8629, 
    -17.71254, -18.56001, -19.40522, -20.2481, -21.08856, -21.92654, 
    -22.76195, -23.59474, -24.42483, -25.25217, -26.07669, -26.89834, 
    -27.71707, -28.53283, -29.34557, -30.15525, -30.96183, -31.76528, 
    -32.56555, -33.36263, -34.15647, -34.94707, -35.73439, -36.51843, 
    -37.29916, -38.07658, -38.85067, -39.62142,
  39.33637, 38.56721, 37.79493, 37.01954, 36.24105, 35.45947, 34.67482, 
    33.88711, 33.09637, 32.30262, 31.50589, 30.7062, 29.90359, 29.0981, 
    28.28975, 27.47861, 26.6647, 25.84807, 25.02878, 24.20688, 23.38242, 
    22.55546, 21.72607, 20.8943, 20.06023, 19.22392, 18.38545, 17.5449, 
    16.70233, 15.85784, 15.0115, 14.1634, 13.31363, 12.46228, 11.60943, 
    10.75519, 9.899641, 9.042892, 8.185037, 7.326178, 6.466415, 5.605854, 
    4.744597, 3.88275, 3.02042, 2.157712, 1.294735, 0.4315965, -0.4315965, 
    -1.294735, -2.157712, -3.02042, -3.88275, -4.744597, -5.605854, 
    -6.466415, -7.326178, -8.185037, -9.042892, -9.899641, -10.75519, 
    -11.60943, -12.46228, -13.31363, -14.1634, -15.0115, -15.85784, 
    -16.70233, -17.5449, -18.38545, -19.22392, -20.06023, -20.8943, 
    -21.72607, -22.55546, -23.38242, -24.20688, -25.02878, -25.84807, 
    -26.6647, -27.47861, -28.28975, -29.0981, -29.90359, -30.7062, -31.50589, 
    -32.30262, -33.09637, -33.88711, -34.67482, -35.45947, -36.24105, 
    -37.01954, -37.79493, -38.56721, -39.33637,
  39.04476, 38.27731, 37.50697, 36.73372, 35.9576, 35.1786, 34.39675, 
    33.61207, 32.82457, 32.03428, 31.24123, 30.44544, 29.64695, 28.84579, 
    28.04199, 27.2356, 26.42666, 25.61521, 24.8013, 23.98498, 23.1663, 
    22.34532, 21.52209, 20.69669, 19.86915, 19.03956, 18.20799, 17.37449, 
    16.53915, 15.70203, 14.86322, 14.02279, 13.18083, 12.33741, 11.49262, 
    10.64656, 9.799295, 8.95093, 8.101551, 7.251252, 6.400125, 5.548265, 
    4.695769, 3.842732, 2.989253, 2.135427, 1.281355, 0.4271349, -0.4271349, 
    -1.281355, -2.135427, -2.989253, -3.842732, -4.695769, -5.548265, 
    -6.400125, -7.251252, -8.101551, -8.95093, -9.799295, -10.64656, 
    -11.49262, -12.33741, -13.18083, -14.02279, -14.86322, -15.70203, 
    -16.53915, -17.37449, -18.20799, -19.03956, -19.86915, -20.69669, 
    -21.52209, -22.34532, -23.1663, -23.98498, -24.8013, -25.61521, 
    -26.42666, -27.2356, -28.04199, -28.84579, -29.64695, -30.44544, 
    -31.24123, -32.03428, -32.82457, -33.61207, -34.39675, -35.1786, 
    -35.9576, -36.73372, -37.50697, -38.27731, -39.04476,
  38.74672, 37.9811, 37.21281, 36.44184, 35.66821, 34.89193, 34.11302, 
    33.33149, 32.54737, 31.76069, 30.97146, 30.17971, 29.38548, 28.5888, 
    27.78969, 26.98821, 26.18438, 25.37826, 24.56988, 23.75929, 22.94654, 
    22.13168, 21.31477, 20.49586, 19.67501, 18.85229, 18.02774, 17.20144, 
    16.37346, 15.54386, 14.71272, 13.88009, 13.04607, 12.21073, 11.37413, 
    10.53637, 9.697527, 8.857674, 8.016898, 7.175284, 6.332918, 5.489884, 
    4.646272, 3.802168, 2.957661, 2.112839, 1.267794, 0.4226128, -0.4226128, 
    -1.267794, -2.112839, -2.957661, -3.802168, -4.646272, -5.489884, 
    -6.332918, -7.175284, -8.016898, -8.857674, -9.697527, -10.53637, 
    -11.37413, -12.21073, -13.04607, -13.88009, -14.71272, -15.54386, 
    -16.37346, -17.20144, -18.02774, -18.85229, -19.67501, -20.49586, 
    -21.31477, -22.13168, -22.94654, -23.75929, -24.56988, -25.37826, 
    -26.18438, -26.98821, -27.78969, -28.5888, -29.38548, -30.17971, 
    -30.97146, -31.76069, -32.54737, -33.33149, -34.11302, -34.89193, 
    -35.66821, -36.44184, -37.21281, -37.9811, -38.74672,
  38.44237, 37.67871, 36.91259, 36.14403, 35.37302, 34.59959, 33.82376, 
    33.04553, 32.26494, 31.482, 30.69673, 29.90917, 29.11935, 28.32729, 
    27.53302, 26.73659, 25.93803, 25.13737, 24.33467, 23.52995, 22.72328, 
    21.91469, 21.10424, 20.29198, 19.47795, 18.66223, 17.84485, 17.02589, 
    16.20541, 15.38346, 14.56011, 13.73542, 12.90947, 12.08233, 11.25405, 
    10.42472, 9.594414, 8.763195, 7.931143, 7.098334, 6.264847, 5.430757, 
    4.596145, 3.761089, 2.925669, 2.089966, 1.254061, 0.4180338, -0.4180338, 
    -1.254061, -2.089966, -2.925669, -3.761089, -4.596145, -5.430757, 
    -6.264847, -7.098334, -7.931143, -8.763195, -9.594414, -10.42472, 
    -11.25405, -12.08233, -12.90947, -13.73542, -14.56011, -15.38346, 
    -16.20541, -17.02589, -17.84485, -18.66223, -19.47795, -20.29198, 
    -21.10424, -21.91469, -22.72328, -23.52995, -24.33467, -25.13737, 
    -25.93803, -26.73659, -27.53302, -28.32729, -29.11935, -29.90917, 
    -30.69673, -31.482, -32.26494, -33.04553, -33.82376, -34.59959, 
    -35.37302, -36.14403, -36.91259, -37.67871, -38.44237,
  38.13184, 37.37026, 36.60646, 35.84042, 35.07218, 34.30174, 33.52912, 
    32.75434, 31.97741, 31.19835, 30.4172, 29.63398, 28.84871, 28.06141, 
    27.27213, 26.4809, 25.68774, 24.89271, 24.09582, 23.29713, 22.49667, 
    21.6945, 20.89065, 20.08517, 19.2781, 18.46952, 17.65945, 16.84796, 
    16.0351, 15.22093, 14.4055, 13.58888, 12.77113, 11.9523, 11.13247, 
    10.31169, 9.490034, 8.667565, 7.844352, 7.020462, 6.195964, 5.370928, 
    4.545426, 3.719527, 2.893303, 2.066826, 1.240168, 0.4134014, -0.4134014, 
    -1.240168, -2.066826, -2.893303, -3.719527, -4.545426, -5.370928, 
    -6.195964, -7.020462, -7.844352, -8.667565, -9.490034, -10.31169, 
    -11.13247, -11.9523, -12.77113, -13.58888, -14.4055, -15.22093, -16.0351, 
    -16.84796, -17.65945, -18.46952, -19.2781, -20.08517, -20.89065, 
    -21.6945, -22.49667, -23.29713, -24.09582, -24.89271, -25.68774, 
    -26.4809, -27.27213, -28.06141, -28.84871, -29.63398, -30.4172, 
    -31.19835, -31.97741, -32.75434, -33.52912, -34.30174, -35.07218, 
    -35.84042, -36.60646, -37.37026, -38.13184,
  37.81525, 37.05589, 36.29453, 35.53117, 34.76583, 33.99852, 33.22925, 
    32.45805, 31.68493, 30.90992, 30.13302, 29.35428, 28.5737, 27.79133, 
    27.00718, 26.22129, 25.43369, 24.64441, 23.85349, 23.06096, 22.26687, 
    21.47124, 20.67413, 19.87557, 19.07561, 18.27429, 17.47165, 16.66776, 
    15.86266, 15.05639, 14.24901, 13.44058, 12.63114, 11.82075, 11.00947, 
    10.19736, 9.384465, 8.570855, 7.756588, 6.941722, 6.12632, 5.310442, 
    4.494153, 3.677513, 2.860586, 2.043435, 1.226125, 0.4087191, -0.4087191, 
    -1.226125, -2.043435, -2.860586, -3.677513, -4.494153, -5.310442, 
    -6.12632, -6.941722, -7.756588, -8.570855, -9.384465, -10.19736, 
    -11.00947, -11.82075, -12.63114, -13.44058, -14.24901, -15.05639, 
    -15.86266, -16.66776, -17.47165, -18.27429, -19.07561, -19.87557, 
    -20.67413, -21.47124, -22.26687, -23.06096, -23.85349, -24.64441, 
    -25.43369, -26.22129, -27.00718, -27.79133, -28.5737, -29.35428, 
    -30.13302, -30.90992, -31.68493, -32.45805, -33.22925, -33.99852, 
    -34.76583, -35.53117, -36.29453, -37.05589, -37.81525,
  37.49273, 36.73572, 35.97694, 35.2164, 34.4541, 33.69006, 32.9243, 
    32.15683, 31.38766, 30.61683, 29.84434, 29.07022, 28.29449, 27.51719, 
    26.73832, 25.95792, 25.17602, 24.39264, 23.60783, 22.8216, 22.034, 
    21.24507, 20.45482, 19.66332, 18.87058, 18.07666, 17.2816, 16.48543, 
    15.6882, 14.88996, 14.09074, 13.29061, 12.4896, 11.68776, 10.88514, 
    10.0818, 9.277779, 8.473132, 7.667912, 6.862171, 6.055964, 5.249342, 
    4.442361, 3.635076, 2.827541, 2.019811, 1.211942, 0.40399, -0.40399, 
    -1.211942, -2.019811, -2.827541, -3.635076, -4.442361, -5.249342, 
    -6.055964, -6.862171, -7.667912, -8.473132, -9.277779, -10.0818, 
    -10.88514, -11.68776, -12.4896, -13.29061, -14.09074, -14.88996, 
    -15.6882, -16.48543, -17.2816, -18.07666, -18.87058, -19.66332, 
    -20.45482, -21.24507, -22.034, -22.8216, -23.60783, -24.39264, -25.17602, 
    -25.95792, -26.73832, -27.51719, -28.29449, -29.07022, -29.84434, 
    -30.61683, -31.38766, -32.15683, -32.9243, -33.69006, -34.4541, -35.2164, 
    -35.97694, -36.73572, -37.49273,
  37.1644, 36.40988, 35.65382, 34.89624, 34.13713, 33.37651, 32.6144, 
    31.8508, 31.08575, 30.31924, 29.55131, 28.78197, 28.01123, 27.23913, 
    26.46569, 25.69092, 24.91487, 24.13754, 23.35897, 22.57919, 21.79822, 
    21.01611, 20.23287, 19.44855, 18.66317, 17.87678, 17.0894, 16.30107, 
    15.51184, 14.72173, 13.9308, 13.13908, 12.3466, 11.55342, 10.75957, 
    9.965097, 9.170046, 8.37446, 7.578384, 6.781863, 5.984942, 5.187668, 
    4.390087, 3.592245, 2.79419, 1.995969, 1.197629, 0.3992176, -0.3992176, 
    -1.197629, -1.995969, -2.79419, -3.592245, -4.390087, -5.187668, 
    -5.984942, -6.781863, -7.578384, -8.37446, -9.170046, -9.965097, 
    -10.75957, -11.55342, -12.3466, -13.13908, -13.9308, -14.72173, 
    -15.51184, -16.30107, -17.0894, -17.87678, -18.66317, -19.44855, 
    -20.23287, -21.01611, -21.79822, -22.57919, -23.35897, -24.13754, 
    -24.91487, -25.69092, -26.46569, -27.23913, -28.01123, -28.78197, 
    -29.55131, -30.31924, -31.08575, -31.8508, -32.6144, -33.37651, 
    -34.13713, -34.89624, -35.65382, -36.40988, -37.1644,
  36.83038, 36.0785, 35.32531, 34.57083, 33.81506, 33.05801, 32.29969, 
    31.54013, 30.77932, 30.0173, 29.25407, 28.48965, 27.72406, 26.95732, 
    26.18944, 25.42046, 24.65038, 23.87924, 23.10706, 22.33386, 21.55966, 
    20.7845, 20.0084, 19.23139, 18.45349, 17.67474, 16.89517, 16.11481, 
    15.33368, 14.55183, 13.76928, 12.98607, 12.20224, 11.41781, 10.63283, 
    9.847324, 9.061338, 8.274905, 7.488063, 6.70085, 5.913303, 5.125462, 
    4.337364, 3.549049, 2.760556, 1.971925, 1.183195, 0.3944048, -0.3944048, 
    -1.183195, -1.971925, -2.760556, -3.549049, -4.337364, -5.125462, 
    -5.913303, -6.70085, -7.488063, -8.274905, -9.061338, -9.847324, 
    -10.63283, -11.41781, -12.20224, -12.98607, -13.76928, -14.55183, 
    -15.33368, -16.11481, -16.89517, -17.67474, -18.45349, -19.23139, 
    -20.0084, -20.7845, -21.55966, -22.33386, -23.10706, -23.87924, 
    -24.65038, -25.42046, -26.18944, -26.95732, -27.72406, -28.48965, 
    -29.25407, -30.0173, -30.77932, -31.54013, -32.29969, -33.05801, 
    -33.81506, -34.57083, -35.32531, -36.0785, -36.83038,
  36.4908, 35.7417, 34.99154, 34.2403, 33.48802, 32.73469, 31.98032, 
    31.22494, 30.46854, 29.71115, 28.95277, 28.19342, 27.43312, 26.67189, 
    25.90973, 25.14667, 24.38272, 23.6179, 22.85224, 22.08575, 21.31846, 
    20.55038, 19.78154, 19.01196, 18.24167, 17.47068, 16.69903, 15.92674, 
    15.15383, 14.38034, 13.60628, 12.83169, 12.05659, 11.28102, 10.505, 
    9.728554, 8.951721, 8.174527, 7.397004, 6.619181, 5.84109, 5.06276, 
    4.284225, 3.505514, 2.72666, 1.947694, 1.168648, 0.3895547, -0.3895547, 
    -1.168648, -1.947694, -2.72666, -3.505514, -4.284225, -5.06276, -5.84109, 
    -6.619181, -7.397004, -8.174527, -8.951721, -9.728554, -10.505, 
    -11.28102, -12.05659, -12.83169, -13.60628, -14.38034, -15.15383, 
    -15.92674, -16.69903, -17.47068, -18.24167, -19.01196, -19.78154, 
    -20.55038, -21.31846, -22.08575, -22.85224, -23.6179, -24.38272, 
    -25.14667, -25.90973, -26.67189, -27.43312, -28.19342, -28.95277, 
    -29.71115, -30.46854, -31.22494, -31.98032, -32.73469, -33.48802, 
    -34.2403, -34.99154, -35.7417, -36.4908,
  36.14578, 35.39962, 34.65261, 33.90479, 33.15614, 32.40669, 31.65643, 
    30.90537, 30.15354, 29.40093, 28.64755, 27.89343, 27.13857, 26.38298, 
    25.62668, 24.86968, 24.112, 23.35365, 22.59464, 21.835, 21.07474, 
    20.31387, 19.55242, 18.79039, 18.02782, 17.26471, 16.50109, 15.73699, 
    14.9724, 14.20737, 13.4419, 12.67602, 11.90976, 11.14313, 10.37615, 
    9.608856, 8.84126, 8.073387, 7.305261, 6.536906, 5.768345, 4.999602, 
    4.230701, 3.461666, 2.692521, 1.92329, 1.153999, 0.3846703, -0.3846703, 
    -1.153999, -1.92329, -2.692521, -3.461666, -4.230701, -4.999602, 
    -5.768345, -6.536906, -7.305261, -8.073387, -8.84126, -9.608856, 
    -10.37615, -11.14313, -11.90976, -12.67602, -13.4419, -14.20737, 
    -14.9724, -15.73699, -16.50109, -17.26471, -18.02782, -18.79039, 
    -19.55242, -20.31387, -21.07474, -21.835, -22.59464, -23.35365, -24.112, 
    -24.86968, -25.62668, -26.38298, -27.13857, -27.89343, -28.64755, 
    -29.40093, -30.15354, -30.90537, -31.65643, -32.40669, -33.15614, 
    -33.90479, -34.65261, -35.39962, -36.14578,
  35.79544, 35.05236, 34.30869, 33.56442, 32.81957, 32.07414, 31.32814, 
    30.58158, 29.83445, 29.08677, 28.33856, 27.58981, 26.84053, 26.09074, 
    25.34044, 24.58965, 23.83837, 23.08662, 22.33441, 21.58174, 20.82863, 
    20.0751, 19.32115, 18.5668, 17.81206, 17.05695, 16.30147, 15.54564, 
    14.78949, 14.03301, 13.27623, 12.51916, 11.76182, 11.00421, 10.24637, 
    9.488298, 8.730017, 7.971541, 7.212887, 6.454072, 5.695111, 4.936023, 
    4.176824, 3.41753, 2.658159, 1.898728, 1.139254, 0.3797542, -0.3797542, 
    -1.139254, -1.898728, -2.658159, -3.41753, -4.176824, -4.936023, 
    -5.695111, -6.454072, -7.212887, -7.971541, -8.730017, -9.488298, 
    -10.24637, -11.00421, -11.76182, -12.51916, -13.27623, -14.03301, 
    -14.78949, -15.54564, -16.30147, -17.05695, -17.81206, -18.5668, 
    -19.32115, -20.0751, -20.82863, -21.58174, -22.33441, -23.08662, 
    -23.83837, -24.58965, -25.34044, -26.09074, -26.84053, -27.58981, 
    -28.33856, -29.08677, -29.83445, -30.58158, -31.32814, -32.07414, 
    -32.81957, -33.56442, -34.30869, -35.05236, -35.79544,
  35.43988, 34.70005, 33.95987, 33.21932, 32.47842, 31.73718, 30.9956, 
    30.25368, 29.51142, 28.76883, 28.02592, 27.28269, 26.53915, 25.7953, 
    25.05115, 24.3067, 23.56197, 22.81695, 22.07165, 21.32609, 20.58027, 
    19.83419, 19.08786, 18.3413, 17.59451, 16.84749, 16.10026, 15.35282, 
    14.60518, 13.85736, 13.10935, 12.36118, 11.61284, 10.86435, 10.11571, 
    9.366945, 8.618052, 7.869044, 7.119931, 6.370722, 5.621428, 4.872057, 
    4.122622, 3.37313, 2.623593, 1.87402, 1.124422, 0.3748092, -0.3748092, 
    -1.124422, -1.87402, -2.623593, -3.37313, -4.122622, -4.872057, 
    -5.621428, -6.370722, -7.119931, -7.869044, -8.618052, -9.366945, 
    -10.11571, -10.86435, -11.61284, -12.36118, -13.10935, -13.85736, 
    -14.60518, -15.35282, -16.10026, -16.84749, -17.59451, -18.3413, 
    -19.08786, -19.83419, -20.58027, -21.32609, -22.07165, -22.81695, 
    -23.56197, -24.3067, -25.05115, -25.7953, -26.53915, -27.28269, 
    -28.02592, -28.76883, -29.51142, -30.25368, -30.9956, -31.73718, 
    -32.47842, -33.21932, -33.95987, -34.70005, -35.43988,
  35.07925, 34.34282, 33.60628, 32.86962, 32.13284, 31.39594, 30.65893, 
    29.92181, 29.18457, 28.44723, 27.70978, 26.97222, 26.23456, 25.4968, 
    24.75893, 24.02097, 23.28291, 22.54476, 21.80651, 21.06818, 20.32976, 
    19.59126, 18.85267, 18.114, 17.37526, 16.63645, 15.89756, 15.15861, 
    14.41959, 13.6805, 12.94136, 12.20216, 11.46291, 10.72361, 9.984256, 
    9.244861, 8.505425, 7.765951, 7.026442, 6.286901, 5.547333, 4.807739, 
    4.068124, 3.32849, 2.588841, 1.849181, 1.109512, 0.3698378, -0.3698378, 
    -1.109512, -1.849181, -2.588841, -3.32849, -4.068124, -4.807739, 
    -5.547333, -6.286901, -7.026442, -7.765951, -8.505425, -9.244861, 
    -9.984256, -10.72361, -11.46291, -12.20216, -12.94136, -13.6805, 
    -14.41959, -15.15861, -15.89756, -16.63645, -17.37526, -18.114, 
    -18.85267, -19.59126, -20.32976, -21.06818, -21.80651, -22.54476, 
    -23.28291, -24.02097, -24.75893, -25.4968, -26.23456, -26.97222, 
    -27.70978, -28.44723, -29.18457, -29.92181, -30.65893, -31.39594, 
    -32.13284, -32.86962, -33.60628, -34.34282, -35.07925 ;

 area =
  5.832426e+09, 5.885548e+09, 5.937712e+09, 5.988909e+09, 6.039129e+09, 
    6.088361e+09, 6.136596e+09, 6.183825e+09, 6.230037e+09, 6.275223e+09, 
    6.319373e+09, 6.362479e+09, 6.404531e+09, 6.445522e+09, 6.485442e+09, 
    6.524282e+09, 6.562035e+09, 6.598693e+09, 6.634248e+09, 6.668692e+09, 
    6.702019e+09, 6.734221e+09, 6.76529e+09, 6.795221e+09, 6.824007e+09, 
    6.851641e+09, 6.878117e+09, 6.903431e+09, 6.927576e+09, 6.950547e+09, 
    6.972339e+09, 6.992947e+09, 7.012366e+09, 7.030593e+09, 7.047623e+09, 
    7.063453e+09, 7.078078e+09, 7.091497e+09, 7.103705e+09, 7.1147e+09, 
    7.124479e+09, 7.133041e+09, 7.140384e+09, 7.146505e+09, 7.151404e+09, 
    7.155078e+09, 7.157529e+09, 7.158754e+09, 7.158754e+09, 7.157529e+09, 
    7.155078e+09, 7.151404e+09, 7.146505e+09, 7.140384e+09, 7.133041e+09, 
    7.124479e+09, 7.1147e+09, 7.103705e+09, 7.091497e+09, 7.078078e+09, 
    7.063453e+09, 7.047623e+09, 7.030593e+09, 7.012366e+09, 6.992947e+09, 
    6.972339e+09, 6.950547e+09, 6.927576e+09, 6.903431e+09, 6.878117e+09, 
    6.851641e+09, 6.824007e+09, 6.795221e+09, 6.76529e+09, 6.734221e+09, 
    6.702019e+09, 6.668692e+09, 6.634248e+09, 6.598693e+09, 6.562035e+09, 
    6.524282e+09, 6.485442e+09, 6.445522e+09, 6.404531e+09, 6.362479e+09, 
    6.319373e+09, 6.275223e+09, 6.230037e+09, 6.183825e+09, 6.136596e+09, 
    6.088361e+09, 6.039129e+09, 5.988909e+09, 5.937712e+09, 5.885548e+09, 
    5.832426e+09,
  5.885548e+09, 5.942029e+09, 5.99757e+09, 6.052155e+09, 6.105772e+09, 
    6.158404e+09, 6.210038e+09, 6.260659e+09, 6.310255e+09, 6.35881e+09, 
    6.406312e+09, 6.452746e+09, 6.4981e+09, 6.54236e+09, 6.585513e+09, 
    6.627547e+09, 6.668449e+09, 6.708208e+09, 6.74681e+09, 6.784244e+09, 
    6.8205e+09, 6.855565e+09, 6.889429e+09, 6.922081e+09, 6.953512e+09, 
    6.98371e+09, 7.012667e+09, 7.040374e+09, 7.066821e+09, 7.092e+09, 
    7.115902e+09, 7.138521e+09, 7.159848e+09, 7.179877e+09, 7.198601e+09, 
    7.216014e+09, 7.23211e+09, 7.246883e+09, 7.260329e+09, 7.272444e+09, 
    7.283223e+09, 7.292662e+09, 7.30076e+09, 7.307511e+09, 7.312915e+09, 
    7.316969e+09, 7.319673e+09, 7.321026e+09, 7.321026e+09, 7.319673e+09, 
    7.316969e+09, 7.312915e+09, 7.307511e+09, 7.30076e+09, 7.292662e+09, 
    7.283223e+09, 7.272444e+09, 7.260329e+09, 7.246883e+09, 7.23211e+09, 
    7.216014e+09, 7.198601e+09, 7.179877e+09, 7.159848e+09, 7.138521e+09, 
    7.115902e+09, 7.092e+09, 7.066821e+09, 7.040374e+09, 7.012667e+09, 
    6.98371e+09, 6.953512e+09, 6.922081e+09, 6.889429e+09, 6.855565e+09, 
    6.8205e+09, 6.784244e+09, 6.74681e+09, 6.708208e+09, 6.668449e+09, 
    6.627547e+09, 6.585513e+09, 6.54236e+09, 6.4981e+09, 6.452746e+09, 
    6.406312e+09, 6.35881e+09, 6.310255e+09, 6.260659e+09, 6.210038e+09, 
    6.158404e+09, 6.105772e+09, 6.052155e+09, 5.99757e+09, 5.942029e+09, 
    5.885548e+09,
  5.937712e+09, 5.99757e+09, 6.056508e+09, 6.114508e+09, 6.171552e+09, 
    6.227619e+09, 6.282692e+09, 6.336752e+09, 6.38978e+09, 6.441759e+09, 
    6.492669e+09, 6.542493e+09, 6.591213e+09, 6.638811e+09, 6.685269e+09, 
    6.730571e+09, 6.774699e+09, 6.817636e+09, 6.859367e+09, 6.899874e+09, 
    6.939143e+09, 6.977157e+09, 7.013901e+09, 7.049361e+09, 7.083523e+09, 
    7.116371e+09, 7.147894e+09, 7.178077e+09, 7.206909e+09, 7.234377e+09, 
    7.260469e+09, 7.285175e+09, 7.308484e+09, 7.330385e+09, 7.350871e+09, 
    7.36993e+09, 7.387556e+09, 7.403741e+09, 7.418477e+09, 7.431758e+09, 
    7.443579e+09, 7.453934e+09, 7.462817e+09, 7.470226e+09, 7.476158e+09, 
    7.480609e+09, 7.483577e+09, 7.485062e+09, 7.485062e+09, 7.483577e+09, 
    7.480609e+09, 7.476158e+09, 7.470226e+09, 7.462817e+09, 7.453934e+09, 
    7.443579e+09, 7.431758e+09, 7.418477e+09, 7.403741e+09, 7.387556e+09, 
    7.36993e+09, 7.350871e+09, 7.330385e+09, 7.308484e+09, 7.285175e+09, 
    7.260469e+09, 7.234377e+09, 7.206909e+09, 7.178077e+09, 7.147894e+09, 
    7.116371e+09, 7.083523e+09, 7.049361e+09, 7.013901e+09, 6.977157e+09, 
    6.939143e+09, 6.899874e+09, 6.859367e+09, 6.817636e+09, 6.774699e+09, 
    6.730571e+09, 6.685269e+09, 6.638811e+09, 6.591213e+09, 6.542493e+09, 
    6.492669e+09, 6.441759e+09, 6.38978e+09, 6.336752e+09, 6.282692e+09, 
    6.227619e+09, 6.171552e+09, 6.114508e+09, 6.056508e+09, 5.99757e+09, 
    5.937712e+09,
  5.988909e+09, 6.052155e+09, 6.114508e+09, 6.175945e+09, 6.236442e+09, 
    6.295976e+09, 6.354524e+09, 6.412062e+09, 6.468569e+09, 6.52402e+09, 
    6.578392e+09, 6.631664e+09, 6.683811e+09, 6.734811e+09, 6.784643e+09, 
    6.833284e+09, 6.880711e+09, 6.926904e+09, 6.971842e+09, 7.015503e+09, 
    7.057866e+09, 7.098912e+09, 7.13862e+09, 7.176973e+09, 7.21395e+09, 
    7.249533e+09, 7.283705e+09, 7.316448e+09, 7.347746e+09, 7.377583e+09, 
    7.405943e+09, 7.432813e+09, 7.458176e+09, 7.482021e+09, 7.504335e+09, 
    7.525106e+09, 7.544322e+09, 7.561974e+09, 7.578052e+09, 7.592547e+09, 
    7.605452e+09, 7.616759e+09, 7.626462e+09, 7.634556e+09, 7.641037e+09, 
    7.645901e+09, 7.649145e+09, 7.650767e+09, 7.650767e+09, 7.649145e+09, 
    7.645901e+09, 7.641037e+09, 7.634556e+09, 7.626462e+09, 7.616759e+09, 
    7.605452e+09, 7.592547e+09, 7.578052e+09, 7.561974e+09, 7.544322e+09, 
    7.525106e+09, 7.504335e+09, 7.482021e+09, 7.458176e+09, 7.432813e+09, 
    7.405943e+09, 7.377583e+09, 7.347746e+09, 7.316448e+09, 7.283705e+09, 
    7.249533e+09, 7.21395e+09, 7.176973e+09, 7.13862e+09, 7.098912e+09, 
    7.057866e+09, 7.015503e+09, 6.971842e+09, 6.926904e+09, 6.880711e+09, 
    6.833284e+09, 6.784643e+09, 6.734811e+09, 6.683811e+09, 6.631664e+09, 
    6.578392e+09, 6.52402e+09, 6.468569e+09, 6.412062e+09, 6.354524e+09, 
    6.295976e+09, 6.236442e+09, 6.175945e+09, 6.114508e+09, 6.052155e+09, 
    5.988909e+09,
  6.039129e+09, 6.105772e+09, 6.171552e+09, 6.236442e+09, 6.300414e+09, 
    6.363442e+09, 6.425497e+09, 6.486551e+09, 6.546576e+09, 6.605544e+09, 
    6.663429e+09, 6.720201e+09, 6.775833e+09, 6.830297e+09, 6.883567e+09, 
    6.935614e+09, 6.986412e+09, 7.035934e+09, 7.084154e+09, 7.131045e+09, 
    7.176583e+09, 7.220742e+09, 7.263496e+09, 7.304823e+09, 7.344698e+09, 
    7.383099e+09, 7.420003e+09, 7.455388e+09, 7.489233e+09, 7.521518e+09, 
    7.552224e+09, 7.581331e+09, 7.608822e+09, 7.634681e+09, 7.65889e+09, 
    7.681435e+09, 7.702302e+09, 7.721477e+09, 7.738948e+09, 7.754704e+09, 
    7.768736e+09, 7.781033e+09, 7.791588e+09, 7.800395e+09, 7.807448e+09, 
    7.812741e+09, 7.816271e+09, 7.818037e+09, 7.818037e+09, 7.816271e+09, 
    7.812741e+09, 7.807448e+09, 7.800395e+09, 7.791588e+09, 7.781033e+09, 
    7.768736e+09, 7.754704e+09, 7.738948e+09, 7.721477e+09, 7.702302e+09, 
    7.681435e+09, 7.65889e+09, 7.634681e+09, 7.608822e+09, 7.581331e+09, 
    7.552224e+09, 7.521518e+09, 7.489233e+09, 7.455388e+09, 7.420003e+09, 
    7.383099e+09, 7.344698e+09, 7.304823e+09, 7.263496e+09, 7.220742e+09, 
    7.176583e+09, 7.131045e+09, 7.084154e+09, 7.035934e+09, 6.986412e+09, 
    6.935614e+09, 6.883567e+09, 6.830297e+09, 6.775833e+09, 6.720201e+09, 
    6.663429e+09, 6.605544e+09, 6.546576e+09, 6.486551e+09, 6.425497e+09, 
    6.363442e+09, 6.300414e+09, 6.236442e+09, 6.171552e+09, 6.105772e+09, 
    6.039129e+09,
  6.088361e+09, 6.158404e+09, 6.227619e+09, 6.295976e+09, 6.363442e+09, 
    6.429985e+09, 6.495574e+09, 6.560175e+09, 6.623755e+09, 6.686283e+09, 
    6.747724e+09, 6.808046e+09, 6.867216e+09, 6.925201e+09, 6.981969e+09, 
    7.037487e+09, 7.091722e+09, 7.144643e+09, 7.196217e+09, 7.246414e+09, 
    7.295202e+09, 7.342552e+09, 7.388432e+09, 7.432814e+09, 7.475667e+09, 
    7.516966e+09, 7.556683e+09, 7.594789e+09, 7.631261e+09, 7.666072e+09, 
    7.699199e+09, 7.73062e+09, 7.760311e+09, 7.788252e+09, 7.814423e+09, 
    7.838806e+09, 7.861382e+09, 7.882135e+09, 7.901051e+09, 7.918115e+09, 
    7.933316e+09, 7.946641e+09, 7.958081e+09, 7.967627e+09, 7.975273e+09, 
    7.981012e+09, 7.984841e+09, 7.986756e+09, 7.986756e+09, 7.984841e+09, 
    7.981012e+09, 7.975273e+09, 7.967627e+09, 7.958081e+09, 7.946641e+09, 
    7.933316e+09, 7.918115e+09, 7.901051e+09, 7.882135e+09, 7.861382e+09, 
    7.838806e+09, 7.814423e+09, 7.788252e+09, 7.760311e+09, 7.73062e+09, 
    7.699199e+09, 7.666072e+09, 7.631261e+09, 7.594789e+09, 7.556683e+09, 
    7.516966e+09, 7.475667e+09, 7.432814e+09, 7.388432e+09, 7.342552e+09, 
    7.295202e+09, 7.246414e+09, 7.196217e+09, 7.144643e+09, 7.091722e+09, 
    7.037487e+09, 6.981969e+09, 6.925201e+09, 6.867216e+09, 6.808046e+09, 
    6.747724e+09, 6.686283e+09, 6.623755e+09, 6.560175e+09, 6.495574e+09, 
    6.429985e+09, 6.363442e+09, 6.295976e+09, 6.227619e+09, 6.158404e+09, 
    6.088361e+09,
  6.136596e+09, 6.210038e+09, 6.282692e+09, 6.354524e+09, 6.425497e+09, 
    6.495574e+09, 6.564719e+09, 6.632894e+09, 6.700061e+09, 6.766183e+09, 
    6.831222e+09, 6.895139e+09, 6.957896e+09, 7.019455e+09, 7.079777e+09, 
    7.138825e+09, 7.196561e+09, 7.252946e+09, 7.307944e+09, 7.361518e+09, 
    7.41363e+09, 7.464245e+09, 7.513327e+09, 7.56084e+09, 7.606751e+09, 
    7.651027e+09, 7.693634e+09, 7.734541e+09, 7.773715e+09, 7.811129e+09, 
    7.846753e+09, 7.880559e+09, 7.912521e+09, 7.942612e+09, 7.970811e+09, 
    7.997093e+09, 8.021437e+09, 8.043825e+09, 8.064236e+09, 8.082655e+09, 
    8.099066e+09, 8.113456e+09, 8.125813e+09, 8.136126e+09, 8.144387e+09, 
    8.150589e+09, 8.154726e+09, 8.156796e+09, 8.156796e+09, 8.154726e+09, 
    8.150589e+09, 8.144387e+09, 8.136126e+09, 8.125813e+09, 8.113456e+09, 
    8.099066e+09, 8.082655e+09, 8.064236e+09, 8.043825e+09, 8.021437e+09, 
    7.997093e+09, 7.970811e+09, 7.942612e+09, 7.912521e+09, 7.880559e+09, 
    7.846753e+09, 7.811129e+09, 7.773715e+09, 7.734541e+09, 7.693634e+09, 
    7.651027e+09, 7.606751e+09, 7.56084e+09, 7.513327e+09, 7.464245e+09, 
    7.41363e+09, 7.361518e+09, 7.307944e+09, 7.252946e+09, 7.196561e+09, 
    7.138825e+09, 7.079777e+09, 7.019455e+09, 6.957896e+09, 6.895139e+09, 
    6.831222e+09, 6.766183e+09, 6.700061e+09, 6.632894e+09, 6.564719e+09, 
    6.495574e+09, 6.425497e+09, 6.354524e+09, 6.282692e+09, 6.210038e+09, 
    6.136596e+09,
  6.183825e+09, 6.260659e+09, 6.336752e+09, 6.412062e+09, 6.486551e+09, 
    6.560175e+09, 6.632894e+09, 6.704666e+09, 6.775447e+09, 6.845195e+09, 
    6.913867e+09, 6.981418e+09, 7.047806e+09, 7.112987e+09, 7.176916e+09, 
    7.23955e+09, 7.300845e+09, 7.360757e+09, 7.419243e+09, 7.47626e+09, 
    7.531766e+09, 7.585717e+09, 7.638074e+09, 7.688794e+09, 7.737838e+09, 
    7.785166e+09, 7.830739e+09, 7.874522e+09, 7.916475e+09, 7.956566e+09, 
    7.994759e+09, 8.031022e+09, 8.065324e+09, 8.097633e+09, 8.127923e+09, 
    8.156166e+09, 8.182336e+09, 8.20641e+09, 8.228367e+09, 8.248187e+09, 
    8.26585e+09, 8.281342e+09, 8.294647e+09, 8.305754e+09, 8.314652e+09, 
    8.321333e+09, 8.32579e+09, 8.32802e+09, 8.32802e+09, 8.32579e+09, 
    8.321333e+09, 8.314652e+09, 8.305754e+09, 8.294647e+09, 8.281342e+09, 
    8.26585e+09, 8.248187e+09, 8.228367e+09, 8.20641e+09, 8.182336e+09, 
    8.156166e+09, 8.127923e+09, 8.097633e+09, 8.065324e+09, 8.031022e+09, 
    7.994759e+09, 7.956566e+09, 7.916475e+09, 7.874522e+09, 7.830739e+09, 
    7.785166e+09, 7.737838e+09, 7.688794e+09, 7.638074e+09, 7.585717e+09, 
    7.531766e+09, 7.47626e+09, 7.419243e+09, 7.360757e+09, 7.300845e+09, 
    7.23955e+09, 7.176916e+09, 7.112987e+09, 7.047806e+09, 6.981418e+09, 
    6.913867e+09, 6.845195e+09, 6.775447e+09, 6.704666e+09, 6.632894e+09, 
    6.560175e+09, 6.486551e+09, 6.412062e+09, 6.336752e+09, 6.260659e+09, 
    6.183825e+09,
  6.230037e+09, 6.310255e+09, 6.38978e+09, 6.468569e+09, 6.546576e+09, 
    6.623755e+09, 6.700061e+09, 6.775447e+09, 6.849864e+09, 6.923265e+09, 
    6.9956e+09, 7.066822e+09, 7.136881e+09, 7.205726e+09, 7.273309e+09, 
    7.339579e+09, 7.404488e+09, 7.467984e+09, 7.530018e+09, 7.590542e+09, 
    7.649507e+09, 7.706863e+09, 7.762563e+09, 7.816561e+09, 7.868808e+09, 
    7.919261e+09, 7.967875e+09, 8.014606e+09, 8.059411e+09, 8.10225e+09, 
    8.143084e+09, 8.181873e+09, 8.218582e+09, 8.253174e+09, 8.285618e+09, 
    8.31588e+09, 8.343933e+09, 8.369748e+09, 8.3933e+09, 8.414565e+09, 
    8.433522e+09, 8.450151e+09, 8.464436e+09, 8.476363e+09, 8.485919e+09, 
    8.493095e+09, 8.497883e+09, 8.500278e+09, 8.500278e+09, 8.497883e+09, 
    8.493095e+09, 8.485919e+09, 8.476363e+09, 8.464436e+09, 8.450151e+09, 
    8.433522e+09, 8.414565e+09, 8.3933e+09, 8.369748e+09, 8.343933e+09, 
    8.31588e+09, 8.285618e+09, 8.253174e+09, 8.218582e+09, 8.181873e+09, 
    8.143084e+09, 8.10225e+09, 8.059411e+09, 8.014606e+09, 7.967875e+09, 
    7.919261e+09, 7.868808e+09, 7.816561e+09, 7.762563e+09, 7.706863e+09, 
    7.649507e+09, 7.590542e+09, 7.530018e+09, 7.467984e+09, 7.404488e+09, 
    7.339579e+09, 7.273309e+09, 7.205726e+09, 7.136881e+09, 7.066822e+09, 
    6.9956e+09, 6.923265e+09, 6.849864e+09, 6.775447e+09, 6.700061e+09, 
    6.623755e+09, 6.546576e+09, 6.468569e+09, 6.38978e+09, 6.310255e+09, 
    6.230037e+09,
  6.275223e+09, 6.35881e+09, 6.441759e+09, 6.52402e+09, 6.605544e+09, 
    6.686283e+09, 6.766183e+09, 6.845195e+09, 6.923265e+09, 7.000339e+09, 
    7.076365e+09, 7.151286e+09, 7.225049e+09, 7.297597e+09, 7.368877e+09, 
    7.438829e+09, 7.5074e+09, 7.574533e+09, 7.640172e+09, 7.704261e+09, 
    7.766745e+09, 7.827569e+09, 7.886679e+09, 7.94402e+09, 7.99954e+09, 
    8.053188e+09, 8.10491e+09, 8.15466e+09, 8.202386e+09, 8.248043e+09, 
    8.291585e+09, 8.332967e+09, 8.372148e+09, 8.409087e+09, 8.443745e+09, 
    8.476086e+09, 8.506077e+09, 8.533684e+09, 8.558878e+09, 8.581632e+09, 
    8.601922e+09, 8.619724e+09, 8.63502e+09, 8.647793e+09, 8.658028e+09, 
    8.665715e+09, 8.670843e+09, 8.673409e+09, 8.673409e+09, 8.670843e+09, 
    8.665715e+09, 8.658028e+09, 8.647793e+09, 8.63502e+09, 8.619724e+09, 
    8.601922e+09, 8.581632e+09, 8.558878e+09, 8.533684e+09, 8.506077e+09, 
    8.476086e+09, 8.443745e+09, 8.409087e+09, 8.372148e+09, 8.332967e+09, 
    8.291585e+09, 8.248043e+09, 8.202386e+09, 8.15466e+09, 8.10491e+09, 
    8.053188e+09, 7.99954e+09, 7.94402e+09, 7.886679e+09, 7.827569e+09, 
    7.766745e+09, 7.704261e+09, 7.640172e+09, 7.574533e+09, 7.5074e+09, 
    7.438829e+09, 7.368877e+09, 7.297597e+09, 7.225049e+09, 7.151286e+09, 
    7.076365e+09, 7.000339e+09, 6.923265e+09, 6.845195e+09, 6.766183e+09, 
    6.686283e+09, 6.605544e+09, 6.52402e+09, 6.441759e+09, 6.35881e+09, 
    6.275223e+09,
  6.319373e+09, 6.406312e+09, 6.492669e+09, 6.578392e+09, 6.663429e+09, 
    6.747724e+09, 6.831222e+09, 6.913867e+09, 6.9956e+09, 7.076365e+09, 
    7.1561e+09, 7.234745e+09, 7.312241e+09, 7.388526e+09, 7.463537e+09, 
    7.537212e+09, 7.60949e+09, 7.680307e+09, 7.749601e+09, 7.817309e+09, 
    7.883369e+09, 7.94772e+09, 8.010299e+09, 8.071048e+09, 8.129904e+09, 
    8.186811e+09, 8.241709e+09, 8.294543e+09, 8.345257e+09, 8.393798e+09, 
    8.440113e+09, 8.484152e+09, 8.525868e+09, 8.565214e+09, 8.602145e+09, 
    8.636621e+09, 8.668601e+09, 8.698051e+09, 8.724934e+09, 8.749221e+09, 
    8.770882e+09, 8.789891e+09, 8.806228e+09, 8.819871e+09, 8.830806e+09, 
    8.839017e+09, 8.844498e+09, 8.84724e+09, 8.84724e+09, 8.844498e+09, 
    8.839017e+09, 8.830806e+09, 8.819871e+09, 8.806228e+09, 8.789891e+09, 
    8.770882e+09, 8.749221e+09, 8.724934e+09, 8.698051e+09, 8.668601e+09, 
    8.636621e+09, 8.602145e+09, 8.565214e+09, 8.525868e+09, 8.484152e+09, 
    8.440113e+09, 8.393798e+09, 8.345257e+09, 8.294543e+09, 8.241709e+09, 
    8.186811e+09, 8.129904e+09, 8.071048e+09, 8.010299e+09, 7.94772e+09, 
    7.883369e+09, 7.817309e+09, 7.749601e+09, 7.680307e+09, 7.60949e+09, 
    7.537212e+09, 7.463537e+09, 7.388526e+09, 7.312241e+09, 7.234745e+09, 
    7.1561e+09, 7.076365e+09, 6.9956e+09, 6.913867e+09, 6.831222e+09, 
    6.747724e+09, 6.663429e+09, 6.578392e+09, 6.492669e+09, 6.406312e+09, 
    6.319373e+09,
  6.362479e+09, 6.452746e+09, 6.542493e+09, 6.631664e+09, 6.720201e+09, 
    6.808046e+09, 6.895139e+09, 6.981418e+09, 7.066822e+09, 7.151286e+09, 
    7.234745e+09, 7.317134e+09, 7.398386e+09, 7.478433e+09, 7.557208e+09, 
    7.634641e+09, 7.710664e+09, 7.785207e+09, 7.858201e+09, 7.929576e+09, 
    7.999264e+09, 8.067195e+09, 8.133301e+09, 8.197513e+09, 8.259766e+09, 
    8.319992e+09, 8.378128e+09, 8.434108e+09, 8.487873e+09, 8.539359e+09, 
    8.58851e+09, 8.635267e+09, 8.679578e+09, 8.721389e+09, 8.760649e+09, 
    8.797313e+09, 8.831335e+09, 8.862674e+09, 8.891291e+09, 8.917151e+09, 
    8.940219e+09, 8.96047e+09, 8.977876e+09, 8.992415e+09, 9.004068e+09, 
    9.012821e+09, 9.018663e+09, 9.021585e+09, 9.021585e+09, 9.018663e+09, 
    9.012821e+09, 9.004068e+09, 8.992415e+09, 8.977876e+09, 8.96047e+09, 
    8.940219e+09, 8.917151e+09, 8.891291e+09, 8.862674e+09, 8.831335e+09, 
    8.797313e+09, 8.760649e+09, 8.721389e+09, 8.679578e+09, 8.635267e+09, 
    8.58851e+09, 8.539359e+09, 8.487873e+09, 8.434108e+09, 8.378128e+09, 
    8.319992e+09, 8.259766e+09, 8.197513e+09, 8.133301e+09, 8.067195e+09, 
    7.999264e+09, 7.929576e+09, 7.858201e+09, 7.785207e+09, 7.710664e+09, 
    7.634641e+09, 7.557208e+09, 7.478433e+09, 7.398386e+09, 7.317134e+09, 
    7.234745e+09, 7.151286e+09, 7.066822e+09, 6.981418e+09, 6.895139e+09, 
    6.808046e+09, 6.720201e+09, 6.631664e+09, 6.542493e+09, 6.452746e+09, 
    6.362479e+09,
  6.404531e+09, 6.4981e+09, 6.591213e+09, 6.683811e+09, 6.775833e+09, 
    6.867216e+09, 6.957896e+09, 7.047806e+09, 7.136881e+09, 7.225049e+09, 
    7.312241e+09, 7.398386e+09, 7.483411e+09, 7.567242e+09, 7.649805e+09, 
    7.731025e+09, 7.810825e+09, 7.889131e+09, 7.965864e+09, 8.04095e+09, 
    8.11431e+09, 8.18587e+09, 8.255552e+09, 8.323282e+09, 8.388985e+09, 
    8.452588e+09, 8.514017e+09, 8.573202e+09, 8.630074e+09, 8.684566e+09, 
    8.736609e+09, 8.786142e+09, 8.833104e+09, 8.877434e+09, 8.919077e+09, 
    8.95798e+09, 8.994092e+09, 9.027367e+09, 9.05776e+09, 9.085231e+09, 
    9.109745e+09, 9.131267e+09, 9.14977e+09, 9.165227e+09, 9.177618e+09, 
    9.186927e+09, 9.193139e+09, 9.196247e+09, 9.196247e+09, 9.193139e+09, 
    9.186927e+09, 9.177618e+09, 9.165227e+09, 9.14977e+09, 9.131267e+09, 
    9.109745e+09, 9.085231e+09, 9.05776e+09, 9.027367e+09, 8.994092e+09, 
    8.95798e+09, 8.919077e+09, 8.877434e+09, 8.833104e+09, 8.786142e+09, 
    8.736609e+09, 8.684566e+09, 8.630074e+09, 8.573202e+09, 8.514017e+09, 
    8.452588e+09, 8.388985e+09, 8.323282e+09, 8.255552e+09, 8.18587e+09, 
    8.11431e+09, 8.04095e+09, 7.965864e+09, 7.889131e+09, 7.810825e+09, 
    7.731025e+09, 7.649805e+09, 7.567242e+09, 7.483411e+09, 7.398386e+09, 
    7.312241e+09, 7.225049e+09, 7.136881e+09, 7.047806e+09, 6.957896e+09, 
    6.867216e+09, 6.775833e+09, 6.683811e+09, 6.591213e+09, 6.4981e+09, 
    6.404531e+09,
  6.445522e+09, 6.54236e+09, 6.638811e+09, 6.734811e+09, 6.830297e+09, 
    6.925201e+09, 7.019455e+09, 7.112987e+09, 7.205726e+09, 7.297597e+09, 
    7.388526e+09, 7.478433e+09, 7.567242e+09, 7.654872e+09, 7.741242e+09, 
    7.826271e+09, 7.909876e+09, 7.991974e+09, 8.072481e+09, 8.151313e+09, 
    8.228386e+09, 8.303616e+09, 8.37692e+09, 8.448214e+09, 8.517416e+09, 
    8.584445e+09, 8.649221e+09, 8.711665e+09, 8.771699e+09, 8.829247e+09, 
    8.884238e+09, 8.936601e+09, 8.986266e+09, 9.033167e+09, 9.077242e+09, 
    9.118431e+09, 9.156679e+09, 9.191932e+09, 9.224142e+09, 9.253263e+09, 
    9.279254e+09, 9.302078e+09, 9.321703e+09, 9.338102e+09, 9.351248e+09, 
    9.361125e+09, 9.367718e+09, 9.371016e+09, 9.371016e+09, 9.367718e+09, 
    9.361125e+09, 9.351248e+09, 9.338102e+09, 9.321703e+09, 9.302078e+09, 
    9.279254e+09, 9.253263e+09, 9.224142e+09, 9.191932e+09, 9.156679e+09, 
    9.118431e+09, 9.077242e+09, 9.033167e+09, 8.986266e+09, 8.936601e+09, 
    8.884238e+09, 8.829247e+09, 8.771699e+09, 8.711665e+09, 8.649221e+09, 
    8.584445e+09, 8.517416e+09, 8.448214e+09, 8.37692e+09, 8.303616e+09, 
    8.228386e+09, 8.151313e+09, 8.072481e+09, 7.991974e+09, 7.909876e+09, 
    7.826271e+09, 7.741242e+09, 7.654872e+09, 7.567242e+09, 7.478433e+09, 
    7.388526e+09, 7.297597e+09, 7.205726e+09, 7.112987e+09, 7.019455e+09, 
    6.925201e+09, 6.830297e+09, 6.734811e+09, 6.638811e+09, 6.54236e+09, 
    6.445522e+09,
  6.485442e+09, 6.585513e+09, 6.685269e+09, 6.784643e+09, 6.883567e+09, 
    6.981969e+09, 7.079777e+09, 7.176916e+09, 7.273309e+09, 7.368877e+09, 
    7.463537e+09, 7.557208e+09, 7.649805e+09, 7.741242e+09, 7.831433e+09, 
    7.920287e+09, 8.007716e+09, 8.093629e+09, 8.177936e+09, 8.260545e+09, 
    8.341364e+09, 8.420301e+09, 8.497266e+09, 8.572165e+09, 8.64491e+09, 
    8.715411e+09, 8.78358e+09, 8.849328e+09, 8.912572e+09, 8.973229e+09, 
    9.031216e+09, 9.086456e+09, 9.138871e+09, 9.188391e+09, 9.234944e+09, 
    9.278465e+09, 9.318892e+09, 9.356163e+09, 9.390226e+09, 9.421031e+09, 
    9.448532e+09, 9.472687e+09, 9.49346e+09, 9.510819e+09, 9.524738e+09, 
    9.535196e+09, 9.542177e+09, 9.54567e+09, 9.54567e+09, 9.542177e+09, 
    9.535196e+09, 9.524738e+09, 9.510819e+09, 9.49346e+09, 9.472687e+09, 
    9.448532e+09, 9.421031e+09, 9.390226e+09, 9.356163e+09, 9.318892e+09, 
    9.278465e+09, 9.234944e+09, 9.188391e+09, 9.138871e+09, 9.086456e+09, 
    9.031216e+09, 8.973229e+09, 8.912572e+09, 8.849328e+09, 8.78358e+09, 
    8.715411e+09, 8.64491e+09, 8.572165e+09, 8.497266e+09, 8.420301e+09, 
    8.341364e+09, 8.260545e+09, 8.177936e+09, 8.093629e+09, 8.007716e+09, 
    7.920287e+09, 7.831433e+09, 7.741242e+09, 7.649805e+09, 7.557208e+09, 
    7.463537e+09, 7.368877e+09, 7.273309e+09, 7.176916e+09, 7.079777e+09, 
    6.981969e+09, 6.883567e+09, 6.784643e+09, 6.685269e+09, 6.585513e+09, 
    6.485442e+09,
  6.524282e+09, 6.627547e+09, 6.730571e+09, 6.833284e+09, 6.935614e+09, 
    7.037487e+09, 7.138825e+09, 7.23955e+09, 7.339579e+09, 7.438829e+09, 
    7.537212e+09, 7.634641e+09, 7.731025e+09, 7.826271e+09, 7.920287e+09, 
    8.012976e+09, 8.104243e+09, 8.193989e+09, 8.282116e+09, 8.368525e+09, 
    8.453116e+09, 8.53579e+09, 8.616447e+09, 8.694987e+09, 8.771312e+09, 
    8.845323e+09, 8.916924e+09, 8.986021e+09, 9.052518e+09, 9.116325e+09, 
    9.177352e+09, 9.235513e+09, 9.290724e+09, 9.342905e+09, 9.391978e+09, 
    9.437871e+09, 9.480515e+09, 9.519842e+09, 9.555794e+09, 9.588315e+09, 
    9.617354e+09, 9.642865e+09, 9.664807e+09, 9.683147e+09, 9.697854e+09, 
    9.708905e+09, 9.716282e+09, 9.719975e+09, 9.719975e+09, 9.716282e+09, 
    9.708905e+09, 9.697854e+09, 9.683147e+09, 9.664807e+09, 9.642865e+09, 
    9.617354e+09, 9.588315e+09, 9.555794e+09, 9.519842e+09, 9.480515e+09, 
    9.437871e+09, 9.391978e+09, 9.342905e+09, 9.290724e+09, 9.235513e+09, 
    9.177352e+09, 9.116325e+09, 9.052518e+09, 8.986021e+09, 8.916924e+09, 
    8.845323e+09, 8.771312e+09, 8.694987e+09, 8.616447e+09, 8.53579e+09, 
    8.453116e+09, 8.368525e+09, 8.282116e+09, 8.193989e+09, 8.104243e+09, 
    8.012976e+09, 7.920287e+09, 7.826271e+09, 7.731025e+09, 7.634641e+09, 
    7.537212e+09, 7.438829e+09, 7.339579e+09, 7.23955e+09, 7.138825e+09, 
    7.037487e+09, 6.935614e+09, 6.833284e+09, 6.730571e+09, 6.627547e+09, 
    6.524282e+09,
  6.562035e+09, 6.668449e+09, 6.774699e+09, 6.880711e+09, 6.986412e+09, 
    7.091722e+09, 7.196561e+09, 7.300845e+09, 7.404488e+09, 7.5074e+09, 
    7.60949e+09, 7.710664e+09, 7.810825e+09, 7.909876e+09, 8.007716e+09, 
    8.104243e+09, 8.199353e+09, 8.292941e+09, 8.384902e+09, 8.475127e+09, 
    8.563511e+09, 8.649944e+09, 8.734319e+09, 8.816526e+09, 8.896461e+09, 
    8.974015e+09, 9.049084e+09, 9.121564e+09, 9.191351e+09, 9.258346e+09, 
    9.322452e+09, 9.383574e+09, 9.441618e+09, 9.496498e+09, 9.548129e+09, 
    9.596429e+09, 9.641325e+09, 9.68274e+09, 9.720613e+09, 9.754878e+09, 
    9.785482e+09, 9.812372e+09, 9.835507e+09, 9.854844e+09, 9.870353e+09, 
    9.882009e+09, 9.88979e+09, 9.893683e+09, 9.893683e+09, 9.88979e+09, 
    9.882009e+09, 9.870353e+09, 9.854844e+09, 9.835507e+09, 9.812372e+09, 
    9.785482e+09, 9.754878e+09, 9.720613e+09, 9.68274e+09, 9.641325e+09, 
    9.596429e+09, 9.548129e+09, 9.496498e+09, 9.441618e+09, 9.383574e+09, 
    9.322452e+09, 9.258346e+09, 9.191351e+09, 9.121564e+09, 9.049084e+09, 
    8.974015e+09, 8.896461e+09, 8.816526e+09, 8.734319e+09, 8.649944e+09, 
    8.563511e+09, 8.475127e+09, 8.384902e+09, 8.292941e+09, 8.199353e+09, 
    8.104243e+09, 8.007716e+09, 7.909876e+09, 7.810825e+09, 7.710664e+09, 
    7.60949e+09, 7.5074e+09, 7.404488e+09, 7.300845e+09, 7.196561e+09, 
    7.091722e+09, 6.986412e+09, 6.880711e+09, 6.774699e+09, 6.668449e+09, 
    6.562035e+09,
  6.598693e+09, 6.708208e+09, 6.817636e+09, 6.926904e+09, 7.035934e+09, 
    7.144643e+09, 7.252946e+09, 7.360757e+09, 7.467984e+09, 7.574533e+09, 
    7.680307e+09, 7.785207e+09, 7.889131e+09, 7.991974e+09, 8.093629e+09, 
    8.193989e+09, 8.292941e+09, 8.390374e+09, 8.486173e+09, 8.580225e+09, 
    8.672412e+09, 8.762619e+09, 8.85073e+09, 8.936627e+09, 9.020195e+09, 
    9.101317e+09, 9.17988e+09, 9.255772e+09, 9.32888e+09, 9.399095e+09, 
    9.466312e+09, 9.530426e+09, 9.591338e+09, 9.64895e+09, 9.703171e+09, 
    9.753911e+09, 9.801088e+09, 9.844622e+09, 9.884442e+09, 9.920478e+09, 
    9.95267e+09, 9.980962e+09, 1.00053e+10, 1.002566e+10, 1.004198e+10, 
    1.005425e+10, 1.006244e+10, 1.006654e+10, 1.006654e+10, 1.006244e+10, 
    1.005425e+10, 1.004198e+10, 1.002566e+10, 1.00053e+10, 9.980962e+09, 
    9.95267e+09, 9.920478e+09, 9.884442e+09, 9.844622e+09, 9.801088e+09, 
    9.753911e+09, 9.703171e+09, 9.64895e+09, 9.591338e+09, 9.530426e+09, 
    9.466312e+09, 9.399095e+09, 9.32888e+09, 9.255772e+09, 9.17988e+09, 
    9.101317e+09, 9.020195e+09, 8.936627e+09, 8.85073e+09, 8.762619e+09, 
    8.672412e+09, 8.580225e+09, 8.486173e+09, 8.390374e+09, 8.292941e+09, 
    8.193989e+09, 8.093629e+09, 7.991974e+09, 7.889131e+09, 7.785207e+09, 
    7.680307e+09, 7.574533e+09, 7.467984e+09, 7.360757e+09, 7.252946e+09, 
    7.144643e+09, 7.035934e+09, 6.926904e+09, 6.817636e+09, 6.708208e+09, 
    6.598693e+09,
  6.634248e+09, 6.74681e+09, 6.859367e+09, 6.971842e+09, 7.084154e+09, 
    7.196217e+09, 7.307944e+09, 7.419243e+09, 7.530018e+09, 7.640172e+09, 
    7.749601e+09, 7.858201e+09, 7.965864e+09, 8.072481e+09, 8.177936e+09, 
    8.282116e+09, 8.384902e+09, 8.486173e+09, 8.585809e+09, 8.683688e+09, 
    8.779684e+09, 8.873673e+09, 8.96553e+09, 9.055129e+09, 9.142345e+09, 
    9.227054e+09, 9.309132e+09, 9.388457e+09, 9.464909e+09, 9.53837e+09, 
    9.608722e+09, 9.675857e+09, 9.739662e+09, 9.800034e+09, 9.856871e+09, 
    9.910078e+09, 9.959563e+09, 1.000524e+10, 1.004703e+10, 1.008486e+10, 
    1.011866e+10, 1.014837e+10, 1.017394e+10, 1.019532e+10, 1.021247e+10, 
    1.022536e+10, 1.023397e+10, 1.023827e+10, 1.023827e+10, 1.023397e+10, 
    1.022536e+10, 1.021247e+10, 1.019532e+10, 1.017394e+10, 1.014837e+10, 
    1.011866e+10, 1.008486e+10, 1.004703e+10, 1.000524e+10, 9.959563e+09, 
    9.910078e+09, 9.856871e+09, 9.800034e+09, 9.739662e+09, 9.675857e+09, 
    9.608722e+09, 9.53837e+09, 9.464909e+09, 9.388457e+09, 9.309132e+09, 
    9.227054e+09, 9.142345e+09, 9.055129e+09, 8.96553e+09, 8.873673e+09, 
    8.779684e+09, 8.683688e+09, 8.585809e+09, 8.486173e+09, 8.384902e+09, 
    8.282116e+09, 8.177936e+09, 8.072481e+09, 7.965864e+09, 7.858201e+09, 
    7.749601e+09, 7.640172e+09, 7.530018e+09, 7.419243e+09, 7.307944e+09, 
    7.196217e+09, 7.084154e+09, 6.971842e+09, 6.859367e+09, 6.74681e+09, 
    6.634248e+09,
  6.668692e+09, 6.784244e+09, 6.899874e+09, 7.015503e+09, 7.131045e+09, 
    7.246414e+09, 7.361518e+09, 7.47626e+09, 7.590542e+09, 7.704261e+09, 
    7.817309e+09, 7.929576e+09, 8.04095e+09, 8.151313e+09, 8.260545e+09, 
    8.368525e+09, 8.475127e+09, 8.580225e+09, 8.683688e+09, 8.785385e+09, 
    8.885187e+09, 8.982957e+09, 9.078562e+09, 9.171869e+09, 9.262742e+09, 
    9.351046e+09, 9.436652e+09, 9.519426e+09, 9.599237e+09, 9.67596e+09, 
    9.749469e+09, 9.819643e+09, 9.886363e+09, 9.949515e+09, 1.000899e+10, 
    1.006469e+10, 1.01165e+10, 1.016434e+10, 1.020812e+10, 1.024776e+10, 
    1.028319e+10, 1.031433e+10, 1.034114e+10, 1.036355e+10, 1.038154e+10, 
    1.039506e+10, 1.040409e+10, 1.040861e+10, 1.040861e+10, 1.040409e+10, 
    1.039506e+10, 1.038154e+10, 1.036355e+10, 1.034114e+10, 1.031433e+10, 
    1.028319e+10, 1.024776e+10, 1.020812e+10, 1.016434e+10, 1.01165e+10, 
    1.006469e+10, 1.000899e+10, 9.949515e+09, 9.886363e+09, 9.819643e+09, 
    9.749469e+09, 9.67596e+09, 9.599237e+09, 9.519426e+09, 9.436652e+09, 
    9.351046e+09, 9.262742e+09, 9.171869e+09, 9.078562e+09, 8.982957e+09, 
    8.885187e+09, 8.785385e+09, 8.683688e+09, 8.580225e+09, 8.475127e+09, 
    8.368525e+09, 8.260545e+09, 8.151313e+09, 8.04095e+09, 7.929576e+09, 
    7.817309e+09, 7.704261e+09, 7.590542e+09, 7.47626e+09, 7.361518e+09, 
    7.246414e+09, 7.131045e+09, 7.015503e+09, 6.899874e+09, 6.784244e+09, 
    6.668692e+09,
  6.702019e+09, 6.8205e+09, 6.939143e+09, 7.057866e+09, 7.176583e+09, 
    7.295202e+09, 7.41363e+09, 7.531766e+09, 7.649507e+09, 7.766745e+09, 
    7.883369e+09, 7.999264e+09, 8.11431e+09, 8.228386e+09, 8.341364e+09, 
    8.453116e+09, 8.563511e+09, 8.672412e+09, 8.779684e+09, 8.885187e+09, 
    8.988781e+09, 9.090322e+09, 9.18967e+09, 9.286681e+09, 9.381209e+09, 
    9.473112e+09, 9.562249e+09, 9.648477e+09, 9.731658e+09, 9.811654e+09, 
    9.88833e+09, 9.961556e+09, 1.00312e+10, 1.009715e+10, 1.015928e+10, 
    1.021748e+10, 1.027164e+10, 1.032166e+10, 1.036744e+10, 1.040891e+10, 
    1.044597e+10, 1.047856e+10, 1.050662e+10, 1.053008e+10, 1.054891e+10, 
    1.056306e+10, 1.057252e+10, 1.057725e+10, 1.057725e+10, 1.057252e+10, 
    1.056306e+10, 1.054891e+10, 1.053008e+10, 1.050662e+10, 1.047856e+10, 
    1.044597e+10, 1.040891e+10, 1.036744e+10, 1.032166e+10, 1.027164e+10, 
    1.021748e+10, 1.015928e+10, 1.009715e+10, 1.00312e+10, 9.961556e+09, 
    9.88833e+09, 9.811654e+09, 9.731658e+09, 9.648477e+09, 9.562249e+09, 
    9.473112e+09, 9.381209e+09, 9.286681e+09, 9.18967e+09, 9.090322e+09, 
    8.988781e+09, 8.885187e+09, 8.779684e+09, 8.672412e+09, 8.563511e+09, 
    8.453116e+09, 8.341364e+09, 8.228386e+09, 8.11431e+09, 7.999264e+09, 
    7.883369e+09, 7.766745e+09, 7.649507e+09, 7.531766e+09, 7.41363e+09, 
    7.295202e+09, 7.176583e+09, 7.057866e+09, 6.939143e+09, 6.8205e+09, 
    6.702019e+09,
  6.734221e+09, 6.855565e+09, 6.977157e+09, 7.098912e+09, 7.220742e+09, 
    7.342552e+09, 7.464245e+09, 7.585717e+09, 7.706863e+09, 7.827569e+09, 
    7.94772e+09, 8.067195e+09, 8.18587e+09, 8.303616e+09, 8.420301e+09, 
    8.53579e+09, 8.649944e+09, 8.762619e+09, 8.873673e+09, 8.982957e+09, 
    9.090322e+09, 9.195619e+09, 9.298694e+09, 9.399396e+09, 9.497571e+09, 
    9.593066e+09, 9.68573e+09, 9.775411e+09, 9.861961e+09, 9.945231e+09, 
    1.002508e+10, 1.010136e+10, 1.017395e+10, 1.02427e+10, 1.030749e+10, 
    1.03682e+10, 1.042471e+10, 1.047692e+10, 1.052472e+10, 1.056802e+10, 
    1.060673e+10, 1.064077e+10, 1.067009e+10, 1.06946e+10, 1.071428e+10, 
    1.072907e+10, 1.073895e+10, 1.07439e+10, 1.07439e+10, 1.073895e+10, 
    1.072907e+10, 1.071428e+10, 1.06946e+10, 1.067009e+10, 1.064077e+10, 
    1.060673e+10, 1.056802e+10, 1.052472e+10, 1.047692e+10, 1.042471e+10, 
    1.03682e+10, 1.030749e+10, 1.02427e+10, 1.017395e+10, 1.010136e+10, 
    1.002508e+10, 9.945231e+09, 9.861961e+09, 9.775411e+09, 9.68573e+09, 
    9.593066e+09, 9.497571e+09, 9.399396e+09, 9.298694e+09, 9.195619e+09, 
    9.090322e+09, 8.982957e+09, 8.873673e+09, 8.762619e+09, 8.649944e+09, 
    8.53579e+09, 8.420301e+09, 8.303616e+09, 8.18587e+09, 8.067195e+09, 
    7.94772e+09, 7.827569e+09, 7.706863e+09, 7.585717e+09, 7.464245e+09, 
    7.342552e+09, 7.220742e+09, 7.098912e+09, 6.977157e+09, 6.855565e+09, 
    6.734221e+09,
  6.76529e+09, 6.889429e+09, 7.013901e+09, 7.13862e+09, 7.263496e+09, 
    7.388432e+09, 7.513327e+09, 7.638074e+09, 7.762563e+09, 7.886679e+09, 
    8.010299e+09, 8.133301e+09, 8.255552e+09, 8.37692e+09, 8.497266e+09, 
    8.616447e+09, 8.734319e+09, 8.85073e+09, 8.96553e+09, 9.078562e+09, 
    9.18967e+09, 9.298694e+09, 9.405474e+09, 9.509846e+09, 9.61165e+09, 
    9.710721e+09, 9.806899e+09, 9.900023e+09, 9.989933e+09, 1.007647e+10, 
    1.015949e+10, 1.023883e+10, 1.031435e+10, 1.03859e+10, 1.045336e+10, 
    1.051658e+10, 1.057545e+10, 1.062985e+10, 1.067967e+10, 1.07248e+10, 
    1.076517e+10, 1.080067e+10, 1.083124e+10, 1.085682e+10, 1.087735e+10, 
    1.089278e+10, 1.090309e+10, 1.090825e+10, 1.090825e+10, 1.090309e+10, 
    1.089278e+10, 1.087735e+10, 1.085682e+10, 1.083124e+10, 1.080067e+10, 
    1.076517e+10, 1.07248e+10, 1.067967e+10, 1.062985e+10, 1.057545e+10, 
    1.051658e+10, 1.045336e+10, 1.03859e+10, 1.031435e+10, 1.023883e+10, 
    1.015949e+10, 1.007647e+10, 9.989933e+09, 9.900023e+09, 9.806899e+09, 
    9.710721e+09, 9.61165e+09, 9.509846e+09, 9.405474e+09, 9.298694e+09, 
    9.18967e+09, 9.078562e+09, 8.96553e+09, 8.85073e+09, 8.734319e+09, 
    8.616447e+09, 8.497266e+09, 8.37692e+09, 8.255552e+09, 8.133301e+09, 
    8.010299e+09, 7.886679e+09, 7.762563e+09, 7.638074e+09, 7.513327e+09, 
    7.388432e+09, 7.263496e+09, 7.13862e+09, 7.013901e+09, 6.889429e+09, 
    6.76529e+09,
  6.795221e+09, 6.922081e+09, 7.049361e+09, 7.176973e+09, 7.304823e+09, 
    7.432814e+09, 7.56084e+09, 7.688794e+09, 7.816561e+09, 7.94402e+09, 
    8.071048e+09, 8.197513e+09, 8.323282e+09, 8.448214e+09, 8.572165e+09, 
    8.694987e+09, 8.816526e+09, 8.936627e+09, 9.055129e+09, 9.171869e+09, 
    9.286681e+09, 9.399396e+09, 9.509846e+09, 9.61786e+09, 9.723264e+09, 
    9.825887e+09, 9.925557e+09, 1.00221e+10, 1.011536e+10, 1.020515e+10, 
    1.029132e+10, 1.037371e+10, 1.045215e+10, 1.05265e+10, 1.059662e+10, 
    1.066235e+10, 1.072358e+10, 1.078017e+10, 1.0832e+10, 1.087898e+10, 
    1.092099e+10, 1.095795e+10, 1.098979e+10, 1.101642e+10, 1.10378e+10, 
    1.105388e+10, 1.106461e+10, 1.106999e+10, 1.106999e+10, 1.106461e+10, 
    1.105388e+10, 1.10378e+10, 1.101642e+10, 1.098979e+10, 1.095795e+10, 
    1.092099e+10, 1.087898e+10, 1.0832e+10, 1.078017e+10, 1.072358e+10, 
    1.066235e+10, 1.059662e+10, 1.05265e+10, 1.045215e+10, 1.037371e+10, 
    1.029132e+10, 1.020515e+10, 1.011536e+10, 1.00221e+10, 9.925557e+09, 
    9.825887e+09, 9.723264e+09, 9.61786e+09, 9.509846e+09, 9.399396e+09, 
    9.286681e+09, 9.171869e+09, 9.055129e+09, 8.936627e+09, 8.816526e+09, 
    8.694987e+09, 8.572165e+09, 8.448214e+09, 8.323282e+09, 8.197513e+09, 
    8.071048e+09, 7.94402e+09, 7.816561e+09, 7.688794e+09, 7.56084e+09, 
    7.432814e+09, 7.304823e+09, 7.176973e+09, 7.049361e+09, 6.922081e+09, 
    6.795221e+09,
  6.824007e+09, 6.953512e+09, 7.083523e+09, 7.21395e+09, 7.344698e+09, 
    7.475667e+09, 7.606751e+09, 7.737838e+09, 7.868808e+09, 7.99954e+09, 
    8.129904e+09, 8.259766e+09, 8.388985e+09, 8.517416e+09, 8.64491e+09, 
    8.771312e+09, 8.896461e+09, 9.020195e+09, 9.142345e+09, 9.262742e+09, 
    9.381209e+09, 9.497571e+09, 9.61165e+09, 9.723264e+09, 9.832232e+09, 
    9.938373e+09, 1.00415e+10, 1.014144e+10, 1.023802e+10, 1.033104e+10, 
    1.042034e+10, 1.050575e+10, 1.058711e+10, 1.066424e+10, 1.0737e+10, 
    1.080523e+10, 1.08688e+10, 1.092757e+10, 1.098142e+10, 1.103023e+10, 
    1.107389e+10, 1.111231e+10, 1.11454e+10, 1.117309e+10, 1.119532e+10, 
    1.121203e+10, 1.12232e+10, 1.122879e+10, 1.122879e+10, 1.12232e+10, 
    1.121203e+10, 1.119532e+10, 1.117309e+10, 1.11454e+10, 1.111231e+10, 
    1.107389e+10, 1.103023e+10, 1.098142e+10, 1.092757e+10, 1.08688e+10, 
    1.080523e+10, 1.0737e+10, 1.066424e+10, 1.058711e+10, 1.050575e+10, 
    1.042034e+10, 1.033104e+10, 1.023802e+10, 1.014144e+10, 1.00415e+10, 
    9.938373e+09, 9.832232e+09, 9.723264e+09, 9.61165e+09, 9.497571e+09, 
    9.381209e+09, 9.262742e+09, 9.142345e+09, 9.020195e+09, 8.896461e+09, 
    8.771312e+09, 8.64491e+09, 8.517416e+09, 8.388985e+09, 8.259766e+09, 
    8.129904e+09, 7.99954e+09, 7.868808e+09, 7.737838e+09, 7.606751e+09, 
    7.475667e+09, 7.344698e+09, 7.21395e+09, 7.083523e+09, 6.953512e+09, 
    6.824007e+09,
  6.851641e+09, 6.98371e+09, 7.116371e+09, 7.249533e+09, 7.383099e+09, 
    7.516966e+09, 7.651027e+09, 7.785166e+09, 7.919261e+09, 8.053188e+09, 
    8.186811e+09, 8.319992e+09, 8.452588e+09, 8.584445e+09, 8.715411e+09, 
    8.845323e+09, 8.974015e+09, 9.101317e+09, 9.227054e+09, 9.351046e+09, 
    9.473112e+09, 9.593066e+09, 9.710721e+09, 9.825887e+09, 9.938373e+09, 
    1.004799e+10, 1.015454e+10, 1.025783e+10, 1.035769e+10, 1.045391e+10, 
    1.054631e+10, 1.063472e+10, 1.071896e+10, 1.079885e+10, 1.087423e+10, 
    1.094495e+10, 1.101085e+10, 1.107179e+10, 1.112763e+10, 1.117826e+10, 
    1.122356e+10, 1.126342e+10, 1.129776e+10, 1.13265e+10, 1.134958e+10, 
    1.136693e+10, 1.137852e+10, 1.138432e+10, 1.138432e+10, 1.137852e+10, 
    1.136693e+10, 1.134958e+10, 1.13265e+10, 1.129776e+10, 1.126342e+10, 
    1.122356e+10, 1.117826e+10, 1.112763e+10, 1.107179e+10, 1.101085e+10, 
    1.094495e+10, 1.087423e+10, 1.079885e+10, 1.071896e+10, 1.063472e+10, 
    1.054631e+10, 1.045391e+10, 1.035769e+10, 1.025783e+10, 1.015454e+10, 
    1.004799e+10, 9.938373e+09, 9.825887e+09, 9.710721e+09, 9.593066e+09, 
    9.473112e+09, 9.351046e+09, 9.227054e+09, 9.101317e+09, 8.974015e+09, 
    8.845323e+09, 8.715411e+09, 8.584445e+09, 8.452588e+09, 8.319992e+09, 
    8.186811e+09, 8.053188e+09, 7.919261e+09, 7.785166e+09, 7.651027e+09, 
    7.516966e+09, 7.383099e+09, 7.249533e+09, 7.116371e+09, 6.98371e+09, 
    6.851641e+09,
  6.878117e+09, 7.012667e+09, 7.147894e+09, 7.283705e+09, 7.420003e+09, 
    7.556683e+09, 7.693634e+09, 7.830739e+09, 7.967875e+09, 8.10491e+09, 
    8.241709e+09, 8.378128e+09, 8.514017e+09, 8.649221e+09, 8.78358e+09, 
    8.916924e+09, 9.049084e+09, 9.17988e+09, 9.309132e+09, 9.436652e+09, 
    9.562249e+09, 9.68573e+09, 9.806899e+09, 9.925557e+09, 1.00415e+10, 
    1.015454e+10, 1.026446e+10, 1.037106e+10, 1.047415e+10, 1.057352e+10, 
    1.066899e+10, 1.076036e+10, 1.084745e+10, 1.093007e+10, 1.100805e+10, 
    1.108122e+10, 1.114942e+10, 1.12125e+10, 1.127033e+10, 1.132276e+10, 
    1.136968e+10, 1.141097e+10, 1.144656e+10, 1.147634e+10, 1.150025e+10, 
    1.151823e+10, 1.153025e+10, 1.153626e+10, 1.153626e+10, 1.153025e+10, 
    1.151823e+10, 1.150025e+10, 1.147634e+10, 1.144656e+10, 1.141097e+10, 
    1.136968e+10, 1.132276e+10, 1.127033e+10, 1.12125e+10, 1.114942e+10, 
    1.108122e+10, 1.100805e+10, 1.093007e+10, 1.084745e+10, 1.076036e+10, 
    1.066899e+10, 1.057352e+10, 1.047415e+10, 1.037106e+10, 1.026446e+10, 
    1.015454e+10, 1.00415e+10, 9.925557e+09, 9.806899e+09, 9.68573e+09, 
    9.562249e+09, 9.436652e+09, 9.309132e+09, 9.17988e+09, 9.049084e+09, 
    8.916924e+09, 8.78358e+09, 8.649221e+09, 8.514017e+09, 8.378128e+09, 
    8.241709e+09, 8.10491e+09, 7.967875e+09, 7.830739e+09, 7.693634e+09, 
    7.556683e+09, 7.420003e+09, 7.283705e+09, 7.147894e+09, 7.012667e+09, 
    6.878117e+09,
  6.903431e+09, 7.040374e+09, 7.178077e+09, 7.316448e+09, 7.455388e+09, 
    7.594789e+09, 7.734541e+09, 7.874522e+09, 8.014606e+09, 8.15466e+09, 
    8.294543e+09, 8.434108e+09, 8.573202e+09, 8.711665e+09, 8.849328e+09, 
    8.986021e+09, 9.121564e+09, 9.255772e+09, 9.388457e+09, 9.519426e+09, 
    9.648477e+09, 9.775411e+09, 9.900023e+09, 1.00221e+10, 1.014144e+10, 
    1.025783e+10, 1.037106e+10, 1.048091e+10, 1.058718e+10, 1.068966e+10, 
    1.078814e+10, 1.088243e+10, 1.097232e+10, 1.105763e+10, 1.113816e+10, 
    1.121375e+10, 1.128423e+10, 1.134943e+10, 1.14092e+10, 1.146341e+10, 
    1.151193e+10, 1.155465e+10, 1.159146e+10, 1.162227e+10, 1.164701e+10, 
    1.166561e+10, 1.167804e+10, 1.168427e+10, 1.168427e+10, 1.167804e+10, 
    1.166561e+10, 1.164701e+10, 1.162227e+10, 1.159146e+10, 1.155465e+10, 
    1.151193e+10, 1.146341e+10, 1.14092e+10, 1.134943e+10, 1.128423e+10, 
    1.121375e+10, 1.113816e+10, 1.105763e+10, 1.097232e+10, 1.088243e+10, 
    1.078814e+10, 1.068966e+10, 1.058718e+10, 1.048091e+10, 1.037106e+10, 
    1.025783e+10, 1.014144e+10, 1.00221e+10, 9.900023e+09, 9.775411e+09, 
    9.648477e+09, 9.519426e+09, 9.388457e+09, 9.255772e+09, 9.121564e+09, 
    8.986021e+09, 8.849328e+09, 8.711665e+09, 8.573202e+09, 8.434108e+09, 
    8.294543e+09, 8.15466e+09, 8.014606e+09, 7.874522e+09, 7.734541e+09, 
    7.594789e+09, 7.455388e+09, 7.316448e+09, 7.178077e+09, 7.040374e+09, 
    6.903431e+09,
  6.927576e+09, 7.066821e+09, 7.206909e+09, 7.347746e+09, 7.489233e+09, 
    7.631261e+09, 7.773715e+09, 7.916475e+09, 8.059411e+09, 8.202386e+09, 
    8.345257e+09, 8.487873e+09, 8.630074e+09, 8.771699e+09, 8.912572e+09, 
    9.052518e+09, 9.191351e+09, 9.32888e+09, 9.464909e+09, 9.599237e+09, 
    9.731658e+09, 9.861961e+09, 9.989933e+09, 1.011536e+10, 1.023802e+10, 
    1.035769e+10, 1.047415e+10, 1.058718e+10, 1.069657e+10, 1.080209e+10, 
    1.090352e+10, 1.100067e+10, 1.109331e+10, 1.118125e+10, 1.12643e+10, 
    1.134227e+10, 1.141498e+10, 1.148226e+10, 1.154395e+10, 1.159992e+10, 
    1.165001e+10, 1.169412e+10, 1.173213e+10, 1.176396e+10, 1.178951e+10, 
    1.180873e+10, 1.182158e+10, 1.1828e+10, 1.1828e+10, 1.182158e+10, 
    1.180873e+10, 1.178951e+10, 1.176396e+10, 1.173213e+10, 1.169412e+10, 
    1.165001e+10, 1.159992e+10, 1.154395e+10, 1.148226e+10, 1.141498e+10, 
    1.134227e+10, 1.12643e+10, 1.118125e+10, 1.109331e+10, 1.100067e+10, 
    1.090352e+10, 1.080209e+10, 1.069657e+10, 1.058718e+10, 1.047415e+10, 
    1.035769e+10, 1.023802e+10, 1.011536e+10, 9.989933e+09, 9.861961e+09, 
    9.731658e+09, 9.599237e+09, 9.464909e+09, 9.32888e+09, 9.191351e+09, 
    9.052518e+09, 8.912572e+09, 8.771699e+09, 8.630074e+09, 8.487873e+09, 
    8.345257e+09, 8.202386e+09, 8.059411e+09, 7.916475e+09, 7.773715e+09, 
    7.631261e+09, 7.489233e+09, 7.347746e+09, 7.206909e+09, 7.066821e+09, 
    6.927576e+09,
  6.950547e+09, 7.092e+09, 7.234377e+09, 7.377583e+09, 7.521518e+09, 
    7.666072e+09, 7.811129e+09, 7.956566e+09, 8.10225e+09, 8.248043e+09, 
    8.393798e+09, 8.539359e+09, 8.684566e+09, 8.829247e+09, 8.973229e+09, 
    9.116325e+09, 9.258346e+09, 9.399095e+09, 9.53837e+09, 9.67596e+09, 
    9.811654e+09, 9.945231e+09, 1.007647e+10, 1.020515e+10, 1.033104e+10, 
    1.045391e+10, 1.057352e+10, 1.068966e+10, 1.080209e+10, 1.091057e+10, 
    1.10149e+10, 1.111483e+10, 1.121017e+10, 1.130069e+10, 1.13862e+10, 
    1.146649e+10, 1.154138e+10, 1.16107e+10, 1.167428e+10, 1.173195e+10, 
    1.17836e+10, 1.182907e+10, 1.186826e+10, 1.190108e+10, 1.192743e+10, 
    1.194726e+10, 1.19605e+10, 1.196713e+10, 1.196713e+10, 1.19605e+10, 
    1.194726e+10, 1.192743e+10, 1.190108e+10, 1.186826e+10, 1.182907e+10, 
    1.17836e+10, 1.173195e+10, 1.167428e+10, 1.16107e+10, 1.154138e+10, 
    1.146649e+10, 1.13862e+10, 1.130069e+10, 1.121017e+10, 1.111483e+10, 
    1.10149e+10, 1.091057e+10, 1.080209e+10, 1.068966e+10, 1.057352e+10, 
    1.045391e+10, 1.033104e+10, 1.020515e+10, 1.007647e+10, 9.945231e+09, 
    9.811654e+09, 9.67596e+09, 9.53837e+09, 9.399095e+09, 9.258346e+09, 
    9.116325e+09, 8.973229e+09, 8.829247e+09, 8.684566e+09, 8.539359e+09, 
    8.393798e+09, 8.248043e+09, 8.10225e+09, 7.956566e+09, 7.811129e+09, 
    7.666072e+09, 7.521518e+09, 7.377583e+09, 7.234377e+09, 7.092e+09, 
    6.950547e+09,
  6.972339e+09, 7.115902e+09, 7.260469e+09, 7.405943e+09, 7.552224e+09, 
    7.699199e+09, 7.846753e+09, 7.994759e+09, 8.143084e+09, 8.291585e+09, 
    8.440113e+09, 8.58851e+09, 8.736609e+09, 8.884238e+09, 9.031216e+09, 
    9.177352e+09, 9.322452e+09, 9.466312e+09, 9.608722e+09, 9.749469e+09, 
    9.88833e+09, 1.002508e+10, 1.015949e+10, 1.029132e+10, 1.042034e+10, 
    1.054631e+10, 1.066899e+10, 1.078814e+10, 1.090352e+10, 1.10149e+10, 
    1.112203e+10, 1.122468e+10, 1.132264e+10, 1.141567e+10, 1.150357e+10, 
    1.158613e+10, 1.166315e+10, 1.173446e+10, 1.179987e+10, 1.185922e+10, 
    1.191237e+10, 1.195917e+10, 1.199952e+10, 1.203331e+10, 1.206044e+10, 
    1.208085e+10, 1.209449e+10, 1.210132e+10, 1.210132e+10, 1.209449e+10, 
    1.208085e+10, 1.206044e+10, 1.203331e+10, 1.199952e+10, 1.195917e+10, 
    1.191237e+10, 1.185922e+10, 1.179987e+10, 1.173446e+10, 1.166315e+10, 
    1.158613e+10, 1.150357e+10, 1.141567e+10, 1.132264e+10, 1.122468e+10, 
    1.112203e+10, 1.10149e+10, 1.090352e+10, 1.078814e+10, 1.066899e+10, 
    1.054631e+10, 1.042034e+10, 1.029132e+10, 1.015949e+10, 1.002508e+10, 
    9.88833e+09, 9.749469e+09, 9.608722e+09, 9.466312e+09, 9.322452e+09, 
    9.177352e+09, 9.031216e+09, 8.884238e+09, 8.736609e+09, 8.58851e+09, 
    8.440113e+09, 8.291585e+09, 8.143084e+09, 7.994759e+09, 7.846753e+09, 
    7.699199e+09, 7.552224e+09, 7.405943e+09, 7.260469e+09, 7.115902e+09, 
    6.972339e+09,
  6.992947e+09, 7.138521e+09, 7.285175e+09, 7.432813e+09, 7.581331e+09, 
    7.73062e+09, 7.880559e+09, 8.031022e+09, 8.181873e+09, 8.332967e+09, 
    8.484152e+09, 8.635267e+09, 8.786142e+09, 8.936601e+09, 9.086456e+09, 
    9.235513e+09, 9.383574e+09, 9.530426e+09, 9.675857e+09, 9.819643e+09, 
    9.961556e+09, 1.010136e+10, 1.023883e+10, 1.037371e+10, 1.050575e+10, 
    1.063472e+10, 1.076036e+10, 1.088243e+10, 1.100067e+10, 1.111483e+10, 
    1.122468e+10, 1.132997e+10, 1.143046e+10, 1.152593e+10, 1.161615e+10, 
    1.170091e+10, 1.178001e+10, 1.185324e+10, 1.192043e+10, 1.198141e+10, 
    1.203602e+10, 1.208412e+10, 1.212559e+10, 1.216031e+10, 1.218821e+10, 
    1.220919e+10, 1.222321e+10, 1.223023e+10, 1.223023e+10, 1.222321e+10, 
    1.220919e+10, 1.218821e+10, 1.216031e+10, 1.212559e+10, 1.208412e+10, 
    1.203602e+10, 1.198141e+10, 1.192043e+10, 1.185324e+10, 1.178001e+10, 
    1.170091e+10, 1.161615e+10, 1.152593e+10, 1.143046e+10, 1.132997e+10, 
    1.122468e+10, 1.111483e+10, 1.100067e+10, 1.088243e+10, 1.076036e+10, 
    1.063472e+10, 1.050575e+10, 1.037371e+10, 1.023883e+10, 1.010136e+10, 
    9.961556e+09, 9.819643e+09, 9.675857e+09, 9.530426e+09, 9.383574e+09, 
    9.235513e+09, 9.086456e+09, 8.936601e+09, 8.786142e+09, 8.635267e+09, 
    8.484152e+09, 8.332967e+09, 8.181873e+09, 8.031022e+09, 7.880559e+09, 
    7.73062e+09, 7.581331e+09, 7.432813e+09, 7.285175e+09, 7.138521e+09, 
    6.992947e+09,
  7.012366e+09, 7.159848e+09, 7.308484e+09, 7.458176e+09, 7.608822e+09, 
    7.760311e+09, 7.912521e+09, 8.065324e+09, 8.218582e+09, 8.372148e+09, 
    8.525868e+09, 8.679578e+09, 8.833104e+09, 8.986266e+09, 9.138871e+09, 
    9.290724e+09, 9.441618e+09, 9.591338e+09, 9.739662e+09, 9.886363e+09, 
    1.00312e+10, 1.017395e+10, 1.031435e+10, 1.045215e+10, 1.058711e+10, 
    1.071896e+10, 1.084745e+10, 1.097232e+10, 1.109331e+10, 1.121017e+10, 
    1.132264e+10, 1.143046e+10, 1.153341e+10, 1.163122e+10, 1.172369e+10, 
    1.181057e+10, 1.189166e+10, 1.196675e+10, 1.203567e+10, 1.209821e+10, 
    1.215424e+10, 1.220359e+10, 1.224615e+10, 1.228178e+10, 1.231041e+10, 
    1.233195e+10, 1.234634e+10, 1.235355e+10, 1.235355e+10, 1.234634e+10, 
    1.233195e+10, 1.231041e+10, 1.228178e+10, 1.224615e+10, 1.220359e+10, 
    1.215424e+10, 1.209821e+10, 1.203567e+10, 1.196675e+10, 1.189166e+10, 
    1.181057e+10, 1.172369e+10, 1.163122e+10, 1.153341e+10, 1.143046e+10, 
    1.132264e+10, 1.121017e+10, 1.109331e+10, 1.097232e+10, 1.084745e+10, 
    1.071896e+10, 1.058711e+10, 1.045215e+10, 1.031435e+10, 1.017395e+10, 
    1.00312e+10, 9.886363e+09, 9.739662e+09, 9.591338e+09, 9.441618e+09, 
    9.290724e+09, 9.138871e+09, 8.986266e+09, 8.833104e+09, 8.679578e+09, 
    8.525868e+09, 8.372148e+09, 8.218582e+09, 8.065324e+09, 7.912521e+09, 
    7.760311e+09, 7.608822e+09, 7.458176e+09, 7.308484e+09, 7.159848e+09, 
    7.012366e+09,
  7.030593e+09, 7.179877e+09, 7.330385e+09, 7.482021e+09, 7.634681e+09, 
    7.788252e+09, 7.942612e+09, 8.097633e+09, 8.253174e+09, 8.409087e+09, 
    8.565214e+09, 8.721389e+09, 8.877434e+09, 9.033167e+09, 9.188391e+09, 
    9.342905e+09, 9.496498e+09, 9.64895e+09, 9.800034e+09, 9.949515e+09, 
    1.009715e+10, 1.02427e+10, 1.03859e+10, 1.05265e+10, 1.066424e+10, 
    1.079885e+10, 1.093007e+10, 1.105763e+10, 1.118125e+10, 1.130069e+10, 
    1.141567e+10, 1.152593e+10, 1.163122e+10, 1.17313e+10, 1.182591e+10, 
    1.191483e+10, 1.199784e+10, 1.207473e+10, 1.214529e+10, 1.220935e+10, 
    1.226673e+10, 1.231729e+10, 1.236089e+10, 1.23974e+10, 1.242673e+10, 
    1.24488e+10, 1.246355e+10, 1.247093e+10, 1.247093e+10, 1.246355e+10, 
    1.24488e+10, 1.242673e+10, 1.23974e+10, 1.236089e+10, 1.231729e+10, 
    1.226673e+10, 1.220935e+10, 1.214529e+10, 1.207473e+10, 1.199784e+10, 
    1.191483e+10, 1.182591e+10, 1.17313e+10, 1.163122e+10, 1.152593e+10, 
    1.141567e+10, 1.130069e+10, 1.118125e+10, 1.105763e+10, 1.093007e+10, 
    1.079885e+10, 1.066424e+10, 1.05265e+10, 1.03859e+10, 1.02427e+10, 
    1.009715e+10, 9.949515e+09, 9.800034e+09, 9.64895e+09, 9.496498e+09, 
    9.342905e+09, 9.188391e+09, 9.033167e+09, 8.877434e+09, 8.721389e+09, 
    8.565214e+09, 8.409087e+09, 8.253174e+09, 8.097633e+09, 7.942612e+09, 
    7.788252e+09, 7.634681e+09, 7.482021e+09, 7.330385e+09, 7.179877e+09, 
    7.030593e+09,
  7.047623e+09, 7.198601e+09, 7.350871e+09, 7.504335e+09, 7.65889e+09, 
    7.814423e+09, 7.970811e+09, 8.127923e+09, 8.285618e+09, 8.443745e+09, 
    8.602145e+09, 8.760649e+09, 8.919077e+09, 9.077242e+09, 9.234944e+09, 
    9.391978e+09, 9.548129e+09, 9.703171e+09, 9.856871e+09, 1.000899e+10, 
    1.015928e+10, 1.030749e+10, 1.045336e+10, 1.059662e+10, 1.0737e+10, 
    1.087423e+10, 1.100805e+10, 1.113816e+10, 1.12643e+10, 1.13862e+10, 
    1.150357e+10, 1.161615e+10, 1.172369e+10, 1.182591e+10, 1.192258e+10, 
    1.201345e+10, 1.209829e+10, 1.217688e+10, 1.224902e+10, 1.231452e+10, 
    1.237321e+10, 1.242492e+10, 1.246951e+10, 1.250686e+10, 1.253687e+10, 
    1.255944e+10, 1.257453e+10, 1.258209e+10, 1.258209e+10, 1.257453e+10, 
    1.255944e+10, 1.253687e+10, 1.250686e+10, 1.246951e+10, 1.242492e+10, 
    1.237321e+10, 1.231452e+10, 1.224902e+10, 1.217688e+10, 1.209829e+10, 
    1.201345e+10, 1.192258e+10, 1.182591e+10, 1.172369e+10, 1.161615e+10, 
    1.150357e+10, 1.13862e+10, 1.12643e+10, 1.113816e+10, 1.100805e+10, 
    1.087423e+10, 1.0737e+10, 1.059662e+10, 1.045336e+10, 1.030749e+10, 
    1.015928e+10, 1.000899e+10, 9.856871e+09, 9.703171e+09, 9.548129e+09, 
    9.391978e+09, 9.234944e+09, 9.077242e+09, 8.919077e+09, 8.760649e+09, 
    8.602145e+09, 8.443745e+09, 8.285618e+09, 8.127923e+09, 7.970811e+09, 
    7.814423e+09, 7.65889e+09, 7.504335e+09, 7.350871e+09, 7.198601e+09, 
    7.047623e+09,
  7.063453e+09, 7.216014e+09, 7.36993e+09, 7.525106e+09, 7.681435e+09, 
    7.838806e+09, 7.997093e+09, 8.156166e+09, 8.31588e+09, 8.476086e+09, 
    8.636621e+09, 8.797313e+09, 8.95798e+09, 9.118431e+09, 9.278465e+09, 
    9.437871e+09, 9.596429e+09, 9.753911e+09, 9.910078e+09, 1.006469e+10, 
    1.021748e+10, 1.03682e+10, 1.051658e+10, 1.066235e+10, 1.080523e+10, 
    1.094495e+10, 1.108122e+10, 1.121375e+10, 1.134227e+10, 1.146649e+10, 
    1.158613e+10, 1.170091e+10, 1.181057e+10, 1.191483e+10, 1.201345e+10, 
    1.210616e+10, 1.219274e+10, 1.227295e+10, 1.234659e+10, 1.241347e+10, 
    1.247338e+10, 1.252618e+10, 1.257172e+10, 1.260987e+10, 1.264052e+10, 
    1.266358e+10, 1.267899e+10, 1.268671e+10, 1.268671e+10, 1.267899e+10, 
    1.266358e+10, 1.264052e+10, 1.260987e+10, 1.257172e+10, 1.252618e+10, 
    1.247338e+10, 1.241347e+10, 1.234659e+10, 1.227295e+10, 1.219274e+10, 
    1.210616e+10, 1.201345e+10, 1.191483e+10, 1.181057e+10, 1.170091e+10, 
    1.158613e+10, 1.146649e+10, 1.134227e+10, 1.121375e+10, 1.108122e+10, 
    1.094495e+10, 1.080523e+10, 1.066235e+10, 1.051658e+10, 1.03682e+10, 
    1.021748e+10, 1.006469e+10, 9.910078e+09, 9.753911e+09, 9.596429e+09, 
    9.437871e+09, 9.278465e+09, 9.118431e+09, 8.95798e+09, 8.797313e+09, 
    8.636621e+09, 8.476086e+09, 8.31588e+09, 8.156166e+09, 7.997093e+09, 
    7.838806e+09, 7.681435e+09, 7.525106e+09, 7.36993e+09, 7.216014e+09, 
    7.063453e+09,
  7.078078e+09, 7.23211e+09, 7.387556e+09, 7.544322e+09, 7.702302e+09, 
    7.861382e+09, 8.021437e+09, 8.182336e+09, 8.343933e+09, 8.506077e+09, 
    8.668601e+09, 8.831335e+09, 8.994092e+09, 9.156679e+09, 9.318892e+09, 
    9.480515e+09, 9.641325e+09, 9.801088e+09, 9.959563e+09, 1.01165e+10, 
    1.027164e+10, 1.042471e+10, 1.057545e+10, 1.072358e+10, 1.08688e+10, 
    1.101085e+10, 1.114942e+10, 1.128423e+10, 1.141498e+10, 1.154138e+10, 
    1.166315e+10, 1.178001e+10, 1.189166e+10, 1.199784e+10, 1.209829e+10, 
    1.219274e+10, 1.228095e+10, 1.236269e+10, 1.243775e+10, 1.250591e+10, 
    1.256699e+10, 1.262082e+10, 1.266725e+10, 1.270614e+10, 1.273739e+10, 
    1.276091e+10, 1.277663e+10, 1.27845e+10, 1.27845e+10, 1.277663e+10, 
    1.276091e+10, 1.273739e+10, 1.270614e+10, 1.266725e+10, 1.262082e+10, 
    1.256699e+10, 1.250591e+10, 1.243775e+10, 1.236269e+10, 1.228095e+10, 
    1.219274e+10, 1.209829e+10, 1.199784e+10, 1.189166e+10, 1.178001e+10, 
    1.166315e+10, 1.154138e+10, 1.141498e+10, 1.128423e+10, 1.114942e+10, 
    1.101085e+10, 1.08688e+10, 1.072358e+10, 1.057545e+10, 1.042471e+10, 
    1.027164e+10, 1.01165e+10, 9.959563e+09, 9.801088e+09, 9.641325e+09, 
    9.480515e+09, 9.318892e+09, 9.156679e+09, 8.994092e+09, 8.831335e+09, 
    8.668601e+09, 8.506077e+09, 8.343933e+09, 8.182336e+09, 8.021437e+09, 
    7.861382e+09, 7.702302e+09, 7.544322e+09, 7.387556e+09, 7.23211e+09, 
    7.078078e+09,
  7.091497e+09, 7.246883e+09, 7.403741e+09, 7.561974e+09, 7.721477e+09, 
    7.882135e+09, 8.043825e+09, 8.20641e+09, 8.369748e+09, 8.533684e+09, 
    8.698051e+09, 8.862674e+09, 9.027367e+09, 9.191932e+09, 9.356163e+09, 
    9.519842e+09, 9.68274e+09, 9.844622e+09, 1.000524e+10, 1.016434e+10, 
    1.032166e+10, 1.047692e+10, 1.062985e+10, 1.078017e+10, 1.092757e+10, 
    1.107179e+10, 1.12125e+10, 1.134943e+10, 1.148226e+10, 1.16107e+10, 
    1.173446e+10, 1.185324e+10, 1.196675e+10, 1.207473e+10, 1.217688e+10, 
    1.227295e+10, 1.236269e+10, 1.244586e+10, 1.252223e+10, 1.25916e+10, 
    1.265377e+10, 1.270856e+10, 1.275582e+10, 1.279542e+10, 1.282723e+10, 
    1.285118e+10, 1.286718e+10, 1.287519e+10, 1.287519e+10, 1.286718e+10, 
    1.285118e+10, 1.282723e+10, 1.279542e+10, 1.275582e+10, 1.270856e+10, 
    1.265377e+10, 1.25916e+10, 1.252223e+10, 1.244586e+10, 1.236269e+10, 
    1.227295e+10, 1.217688e+10, 1.207473e+10, 1.196675e+10, 1.185324e+10, 
    1.173446e+10, 1.16107e+10, 1.148226e+10, 1.134943e+10, 1.12125e+10, 
    1.107179e+10, 1.092757e+10, 1.078017e+10, 1.062985e+10, 1.047692e+10, 
    1.032166e+10, 1.016434e+10, 1.000524e+10, 9.844622e+09, 9.68274e+09, 
    9.519842e+09, 9.356163e+09, 9.191932e+09, 9.027367e+09, 8.862674e+09, 
    8.698051e+09, 8.533684e+09, 8.369748e+09, 8.20641e+09, 8.043825e+09, 
    7.882135e+09, 7.721477e+09, 7.561974e+09, 7.403741e+09, 7.246883e+09, 
    7.091497e+09,
  7.103705e+09, 7.260329e+09, 7.418477e+09, 7.578052e+09, 7.738948e+09, 
    7.901051e+09, 8.064236e+09, 8.228367e+09, 8.3933e+09, 8.558878e+09, 
    8.724934e+09, 8.891291e+09, 9.05776e+09, 9.224142e+09, 9.390226e+09, 
    9.555794e+09, 9.720613e+09, 9.884442e+09, 1.004703e+10, 1.020812e+10, 
    1.036744e+10, 1.052472e+10, 1.067967e+10, 1.0832e+10, 1.098142e+10, 
    1.112763e+10, 1.127033e+10, 1.14092e+10, 1.154395e+10, 1.167428e+10, 
    1.179987e+10, 1.192043e+10, 1.203567e+10, 1.214529e+10, 1.224902e+10, 
    1.234659e+10, 1.243775e+10, 1.252223e+10, 1.259983e+10, 1.267031e+10, 
    1.273348e+10, 1.278916e+10, 1.283719e+10, 1.287743e+10, 1.290977e+10, 
    1.293411e+10, 1.295038e+10, 1.295852e+10, 1.295852e+10, 1.295038e+10, 
    1.293411e+10, 1.290977e+10, 1.287743e+10, 1.283719e+10, 1.278916e+10, 
    1.273348e+10, 1.267031e+10, 1.259983e+10, 1.252223e+10, 1.243775e+10, 
    1.234659e+10, 1.224902e+10, 1.214529e+10, 1.203567e+10, 1.192043e+10, 
    1.179987e+10, 1.167428e+10, 1.154395e+10, 1.14092e+10, 1.127033e+10, 
    1.112763e+10, 1.098142e+10, 1.0832e+10, 1.067967e+10, 1.052472e+10, 
    1.036744e+10, 1.020812e+10, 1.004703e+10, 9.884442e+09, 9.720613e+09, 
    9.555794e+09, 9.390226e+09, 9.224142e+09, 9.05776e+09, 8.891291e+09, 
    8.724934e+09, 8.558878e+09, 8.3933e+09, 8.228367e+09, 8.064236e+09, 
    7.901051e+09, 7.738948e+09, 7.578052e+09, 7.418477e+09, 7.260329e+09, 
    7.103705e+09,
  7.1147e+09, 7.272444e+09, 7.431758e+09, 7.592547e+09, 7.754704e+09, 
    7.918115e+09, 8.082655e+09, 8.248187e+09, 8.414565e+09, 8.581632e+09, 
    8.749221e+09, 8.917151e+09, 9.085231e+09, 9.253263e+09, 9.421031e+09, 
    9.588315e+09, 9.754878e+09, 9.920478e+09, 1.008486e+10, 1.024776e+10, 
    1.040891e+10, 1.056802e+10, 1.07248e+10, 1.087898e+10, 1.103023e+10, 
    1.117826e+10, 1.132276e+10, 1.146341e+10, 1.159992e+10, 1.173195e+10, 
    1.185922e+10, 1.198141e+10, 1.209821e+10, 1.220935e+10, 1.231452e+10, 
    1.241347e+10, 1.250591e+10, 1.25916e+10, 1.267031e+10, 1.27418e+10, 
    1.280589e+10, 1.286239e+10, 1.291113e+10, 1.295196e+10, 1.298478e+10, 
    1.300948e+10, 1.302599e+10, 1.303425e+10, 1.303425e+10, 1.302599e+10, 
    1.300948e+10, 1.298478e+10, 1.295196e+10, 1.291113e+10, 1.286239e+10, 
    1.280589e+10, 1.27418e+10, 1.267031e+10, 1.25916e+10, 1.250591e+10, 
    1.241347e+10, 1.231452e+10, 1.220935e+10, 1.209821e+10, 1.198141e+10, 
    1.185922e+10, 1.173195e+10, 1.159992e+10, 1.146341e+10, 1.132276e+10, 
    1.117826e+10, 1.103023e+10, 1.087898e+10, 1.07248e+10, 1.056802e+10, 
    1.040891e+10, 1.024776e+10, 1.008486e+10, 9.920478e+09, 9.754878e+09, 
    9.588315e+09, 9.421031e+09, 9.253263e+09, 9.085231e+09, 8.917151e+09, 
    8.749221e+09, 8.581632e+09, 8.414565e+09, 8.248187e+09, 8.082655e+09, 
    7.918115e+09, 7.754704e+09, 7.592547e+09, 7.431758e+09, 7.272444e+09, 
    7.1147e+09,
  7.124479e+09, 7.283223e+09, 7.443579e+09, 7.605452e+09, 7.768736e+09, 
    7.933316e+09, 8.099066e+09, 8.26585e+09, 8.433522e+09, 8.601922e+09, 
    8.770882e+09, 8.940219e+09, 9.109745e+09, 9.279254e+09, 9.448532e+09, 
    9.617354e+09, 9.785482e+09, 9.95267e+09, 1.011866e+10, 1.028319e+10, 
    1.044597e+10, 1.060673e+10, 1.076517e+10, 1.092099e+10, 1.107389e+10, 
    1.122356e+10, 1.136968e+10, 1.151193e+10, 1.165001e+10, 1.17836e+10, 
    1.191237e+10, 1.203602e+10, 1.215424e+10, 1.226673e+10, 1.237321e+10, 
    1.247338e+10, 1.256699e+10, 1.265377e+10, 1.273348e+10, 1.280589e+10, 
    1.287081e+10, 1.292804e+10, 1.297741e+10, 1.301878e+10, 1.305203e+10, 
    1.307706e+10, 1.309378e+10, 1.310215e+10, 1.310215e+10, 1.309378e+10, 
    1.307706e+10, 1.305203e+10, 1.301878e+10, 1.297741e+10, 1.292804e+10, 
    1.287081e+10, 1.280589e+10, 1.273348e+10, 1.265377e+10, 1.256699e+10, 
    1.247338e+10, 1.237321e+10, 1.226673e+10, 1.215424e+10, 1.203602e+10, 
    1.191237e+10, 1.17836e+10, 1.165001e+10, 1.151193e+10, 1.136968e+10, 
    1.122356e+10, 1.107389e+10, 1.092099e+10, 1.076517e+10, 1.060673e+10, 
    1.044597e+10, 1.028319e+10, 1.011866e+10, 9.95267e+09, 9.785482e+09, 
    9.617354e+09, 9.448532e+09, 9.279254e+09, 9.109745e+09, 8.940219e+09, 
    8.770882e+09, 8.601922e+09, 8.433522e+09, 8.26585e+09, 8.099066e+09, 
    7.933316e+09, 7.768736e+09, 7.605452e+09, 7.443579e+09, 7.283223e+09, 
    7.124479e+09,
  7.133041e+09, 7.292662e+09, 7.453934e+09, 7.616759e+09, 7.781033e+09, 
    7.946641e+09, 8.113456e+09, 8.281342e+09, 8.450151e+09, 8.619724e+09, 
    8.789891e+09, 8.96047e+09, 9.131267e+09, 9.302078e+09, 9.472687e+09, 
    9.642865e+09, 9.812372e+09, 9.980962e+09, 1.014837e+10, 1.031433e+10, 
    1.047856e+10, 1.064077e+10, 1.080067e+10, 1.095795e+10, 1.111231e+10, 
    1.126342e+10, 1.141097e+10, 1.155465e+10, 1.169412e+10, 1.182907e+10, 
    1.195917e+10, 1.208412e+10, 1.220359e+10, 1.231729e+10, 1.242492e+10, 
    1.252618e+10, 1.262082e+10, 1.270856e+10, 1.278916e+10, 1.286239e+10, 
    1.292804e+10, 1.298592e+10, 1.303585e+10, 1.30777e+10, 1.311133e+10, 
    1.313664e+10, 1.315356e+10, 1.316203e+10, 1.316203e+10, 1.315356e+10, 
    1.313664e+10, 1.311133e+10, 1.30777e+10, 1.303585e+10, 1.298592e+10, 
    1.292804e+10, 1.286239e+10, 1.278916e+10, 1.270856e+10, 1.262082e+10, 
    1.252618e+10, 1.242492e+10, 1.231729e+10, 1.220359e+10, 1.208412e+10, 
    1.195917e+10, 1.182907e+10, 1.169412e+10, 1.155465e+10, 1.141097e+10, 
    1.126342e+10, 1.111231e+10, 1.095795e+10, 1.080067e+10, 1.064077e+10, 
    1.047856e+10, 1.031433e+10, 1.014837e+10, 9.980962e+09, 9.812372e+09, 
    9.642865e+09, 9.472687e+09, 9.302078e+09, 9.131267e+09, 8.96047e+09, 
    8.789891e+09, 8.619724e+09, 8.450151e+09, 8.281342e+09, 8.113456e+09, 
    7.946641e+09, 7.781033e+09, 7.616759e+09, 7.453934e+09, 7.292662e+09, 
    7.133041e+09,
  7.140384e+09, 7.30076e+09, 7.462817e+09, 7.626462e+09, 7.791588e+09, 
    7.958081e+09, 8.125813e+09, 8.294647e+09, 8.464436e+09, 8.63502e+09, 
    8.806228e+09, 8.977876e+09, 9.14977e+09, 9.321703e+09, 9.49346e+09, 
    9.664807e+09, 9.835507e+09, 1.00053e+10, 1.017394e+10, 1.034114e+10, 
    1.050662e+10, 1.067009e+10, 1.083124e+10, 1.098979e+10, 1.11454e+10, 
    1.129776e+10, 1.144656e+10, 1.159146e+10, 1.173213e+10, 1.186826e+10, 
    1.199952e+10, 1.212559e+10, 1.224615e+10, 1.236089e+10, 1.246951e+10, 
    1.257172e+10, 1.266725e+10, 1.275582e+10, 1.283719e+10, 1.291113e+10, 
    1.297741e+10, 1.303585e+10, 1.308628e+10, 1.312854e+10, 1.316249e+10, 
    1.318806e+10, 1.320514e+10, 1.32137e+10, 1.32137e+10, 1.320514e+10, 
    1.318806e+10, 1.316249e+10, 1.312854e+10, 1.308628e+10, 1.303585e+10, 
    1.297741e+10, 1.291113e+10, 1.283719e+10, 1.275582e+10, 1.266725e+10, 
    1.257172e+10, 1.246951e+10, 1.236089e+10, 1.224615e+10, 1.212559e+10, 
    1.199952e+10, 1.186826e+10, 1.173213e+10, 1.159146e+10, 1.144656e+10, 
    1.129776e+10, 1.11454e+10, 1.098979e+10, 1.083124e+10, 1.067009e+10, 
    1.050662e+10, 1.034114e+10, 1.017394e+10, 1.00053e+10, 9.835507e+09, 
    9.664807e+09, 9.49346e+09, 9.321703e+09, 9.14977e+09, 8.977876e+09, 
    8.806228e+09, 8.63502e+09, 8.464436e+09, 8.294647e+09, 8.125813e+09, 
    7.958081e+09, 7.791588e+09, 7.626462e+09, 7.462817e+09, 7.30076e+09, 
    7.140384e+09,
  7.146505e+09, 7.307511e+09, 7.470226e+09, 7.634556e+09, 7.800395e+09, 
    7.967627e+09, 8.136126e+09, 8.305754e+09, 8.476363e+09, 8.647793e+09, 
    8.819871e+09, 8.992415e+09, 9.165227e+09, 9.338102e+09, 9.510819e+09, 
    9.683147e+09, 9.854844e+09, 1.002566e+10, 1.019532e+10, 1.036355e+10, 
    1.053008e+10, 1.06946e+10, 1.085682e+10, 1.101642e+10, 1.117309e+10, 
    1.13265e+10, 1.147634e+10, 1.162227e+10, 1.176396e+10, 1.190108e+10, 
    1.203331e+10, 1.216031e+10, 1.228178e+10, 1.23974e+10, 1.250686e+10, 
    1.260987e+10, 1.270614e+10, 1.279542e+10, 1.287743e+10, 1.295196e+10, 
    1.301878e+10, 1.30777e+10, 1.312854e+10, 1.317114e+10, 1.320537e+10, 
    1.323115e+10, 1.324837e+10, 1.3257e+10, 1.3257e+10, 1.324837e+10, 
    1.323115e+10, 1.320537e+10, 1.317114e+10, 1.312854e+10, 1.30777e+10, 
    1.301878e+10, 1.295196e+10, 1.287743e+10, 1.279542e+10, 1.270614e+10, 
    1.260987e+10, 1.250686e+10, 1.23974e+10, 1.228178e+10, 1.216031e+10, 
    1.203331e+10, 1.190108e+10, 1.176396e+10, 1.162227e+10, 1.147634e+10, 
    1.13265e+10, 1.117309e+10, 1.101642e+10, 1.085682e+10, 1.06946e+10, 
    1.053008e+10, 1.036355e+10, 1.019532e+10, 1.002566e+10, 9.854844e+09, 
    9.683147e+09, 9.510819e+09, 9.338102e+09, 9.165227e+09, 8.992415e+09, 
    8.819871e+09, 8.647793e+09, 8.476363e+09, 8.305754e+09, 8.136126e+09, 
    7.967627e+09, 7.800395e+09, 7.634556e+09, 7.470226e+09, 7.307511e+09, 
    7.146505e+09,
  7.151404e+09, 7.312915e+09, 7.476158e+09, 7.641037e+09, 7.807448e+09, 
    7.975273e+09, 8.144387e+09, 8.314652e+09, 8.485919e+09, 8.658028e+09, 
    8.830806e+09, 9.004068e+09, 9.177618e+09, 9.351248e+09, 9.524738e+09, 
    9.697854e+09, 9.870353e+09, 1.004198e+10, 1.021247e+10, 1.038154e+10, 
    1.054891e+10, 1.071428e+10, 1.087735e+10, 1.10378e+10, 1.119532e+10, 
    1.134958e+10, 1.150025e+10, 1.164701e+10, 1.178951e+10, 1.192743e+10, 
    1.206044e+10, 1.218821e+10, 1.231041e+10, 1.242673e+10, 1.253687e+10, 
    1.264052e+10, 1.273739e+10, 1.282723e+10, 1.290977e+10, 1.298478e+10, 
    1.305203e+10, 1.311133e+10, 1.316249e+10, 1.320537e+10, 1.323984e+10, 
    1.326578e+10, 1.328312e+10, 1.32918e+10, 1.32918e+10, 1.328312e+10, 
    1.326578e+10, 1.323984e+10, 1.320537e+10, 1.316249e+10, 1.311133e+10, 
    1.305203e+10, 1.298478e+10, 1.290977e+10, 1.282723e+10, 1.273739e+10, 
    1.264052e+10, 1.253687e+10, 1.242673e+10, 1.231041e+10, 1.218821e+10, 
    1.206044e+10, 1.192743e+10, 1.178951e+10, 1.164701e+10, 1.150025e+10, 
    1.134958e+10, 1.119532e+10, 1.10378e+10, 1.087735e+10, 1.071428e+10, 
    1.054891e+10, 1.038154e+10, 1.021247e+10, 1.004198e+10, 9.870353e+09, 
    9.697854e+09, 9.524738e+09, 9.351248e+09, 9.177618e+09, 9.004068e+09, 
    8.830806e+09, 8.658028e+09, 8.485919e+09, 8.314652e+09, 8.144387e+09, 
    7.975273e+09, 7.807448e+09, 7.641037e+09, 7.476158e+09, 7.312915e+09, 
    7.151404e+09,
  7.155078e+09, 7.316969e+09, 7.480609e+09, 7.645901e+09, 7.812741e+09, 
    7.981012e+09, 8.150589e+09, 8.321333e+09, 8.493095e+09, 8.665715e+09, 
    8.839017e+09, 9.012821e+09, 9.186927e+09, 9.361125e+09, 9.535196e+09, 
    9.708905e+09, 9.882009e+09, 1.005425e+10, 1.022536e+10, 1.039506e+10, 
    1.056306e+10, 1.072907e+10, 1.089278e+10, 1.105388e+10, 1.121203e+10, 
    1.136693e+10, 1.151823e+10, 1.166561e+10, 1.180873e+10, 1.194726e+10, 
    1.208085e+10, 1.220919e+10, 1.233195e+10, 1.24488e+10, 1.255944e+10, 
    1.266358e+10, 1.276091e+10, 1.285118e+10, 1.293411e+10, 1.300948e+10, 
    1.307706e+10, 1.313664e+10, 1.318806e+10, 1.323115e+10, 1.326578e+10, 
    1.329185e+10, 1.330927e+10, 1.3318e+10, 1.3318e+10, 1.330927e+10, 
    1.329185e+10, 1.326578e+10, 1.323115e+10, 1.318806e+10, 1.313664e+10, 
    1.307706e+10, 1.300948e+10, 1.293411e+10, 1.285118e+10, 1.276091e+10, 
    1.266358e+10, 1.255944e+10, 1.24488e+10, 1.233195e+10, 1.220919e+10, 
    1.208085e+10, 1.194726e+10, 1.180873e+10, 1.166561e+10, 1.151823e+10, 
    1.136693e+10, 1.121203e+10, 1.105388e+10, 1.089278e+10, 1.072907e+10, 
    1.056306e+10, 1.039506e+10, 1.022536e+10, 1.005425e+10, 9.882009e+09, 
    9.708905e+09, 9.535196e+09, 9.361125e+09, 9.186927e+09, 9.012821e+09, 
    8.839017e+09, 8.665715e+09, 8.493095e+09, 8.321333e+09, 8.150589e+09, 
    7.981012e+09, 7.812741e+09, 7.645901e+09, 7.480609e+09, 7.316969e+09, 
    7.155078e+09,
  7.157529e+09, 7.319673e+09, 7.483577e+09, 7.649145e+09, 7.816271e+09, 
    7.984841e+09, 8.154726e+09, 8.32579e+09, 8.497883e+09, 8.670843e+09, 
    8.844498e+09, 9.018663e+09, 9.193139e+09, 9.367718e+09, 9.542177e+09, 
    9.716282e+09, 9.88979e+09, 1.006244e+10, 1.023397e+10, 1.040409e+10, 
    1.057252e+10, 1.073895e+10, 1.090309e+10, 1.106461e+10, 1.12232e+10, 
    1.137852e+10, 1.153025e+10, 1.167804e+10, 1.182158e+10, 1.19605e+10, 
    1.209449e+10, 1.222321e+10, 1.234634e+10, 1.246355e+10, 1.257453e+10, 
    1.267899e+10, 1.277663e+10, 1.286718e+10, 1.295038e+10, 1.302599e+10, 
    1.309378e+10, 1.315356e+10, 1.320514e+10, 1.324837e+10, 1.328312e+10, 
    1.330927e+10, 1.332675e+10, 1.333551e+10, 1.333551e+10, 1.332675e+10, 
    1.330927e+10, 1.328312e+10, 1.324837e+10, 1.320514e+10, 1.315356e+10, 
    1.309378e+10, 1.302599e+10, 1.295038e+10, 1.286718e+10, 1.277663e+10, 
    1.267899e+10, 1.257453e+10, 1.246355e+10, 1.234634e+10, 1.222321e+10, 
    1.209449e+10, 1.19605e+10, 1.182158e+10, 1.167804e+10, 1.153025e+10, 
    1.137852e+10, 1.12232e+10, 1.106461e+10, 1.090309e+10, 1.073895e+10, 
    1.057252e+10, 1.040409e+10, 1.023397e+10, 1.006244e+10, 9.88979e+09, 
    9.716282e+09, 9.542177e+09, 9.367718e+09, 9.193139e+09, 9.018663e+09, 
    8.844498e+09, 8.670843e+09, 8.497883e+09, 8.32579e+09, 8.154726e+09, 
    7.984841e+09, 7.816271e+09, 7.649145e+09, 7.483577e+09, 7.319673e+09, 
    7.157529e+09,
  7.158754e+09, 7.321026e+09, 7.485062e+09, 7.650767e+09, 7.818037e+09, 
    7.986756e+09, 8.156796e+09, 8.32802e+09, 8.500278e+09, 8.673409e+09, 
    8.84724e+09, 9.021585e+09, 9.196247e+09, 9.371016e+09, 9.54567e+09, 
    9.719975e+09, 9.893683e+09, 1.006654e+10, 1.023827e+10, 1.040861e+10, 
    1.057725e+10, 1.07439e+10, 1.090825e+10, 1.106999e+10, 1.122879e+10, 
    1.138432e+10, 1.153626e+10, 1.168427e+10, 1.1828e+10, 1.196713e+10, 
    1.210132e+10, 1.223023e+10, 1.235355e+10, 1.247093e+10, 1.258209e+10, 
    1.268671e+10, 1.27845e+10, 1.287519e+10, 1.295852e+10, 1.303425e+10, 
    1.310215e+10, 1.316203e+10, 1.32137e+10, 1.3257e+10, 1.32918e+10, 
    1.3318e+10, 1.333551e+10, 1.334428e+10, 1.334428e+10, 1.333551e+10, 
    1.3318e+10, 1.32918e+10, 1.3257e+10, 1.32137e+10, 1.316203e+10, 
    1.310215e+10, 1.303425e+10, 1.295852e+10, 1.287519e+10, 1.27845e+10, 
    1.268671e+10, 1.258209e+10, 1.247093e+10, 1.235355e+10, 1.223023e+10, 
    1.210132e+10, 1.196713e+10, 1.1828e+10, 1.168427e+10, 1.153626e+10, 
    1.138432e+10, 1.122879e+10, 1.106999e+10, 1.090825e+10, 1.07439e+10, 
    1.057725e+10, 1.040861e+10, 1.023827e+10, 1.006654e+10, 9.893683e+09, 
    9.719975e+09, 9.54567e+09, 9.371016e+09, 9.196247e+09, 9.021585e+09, 
    8.84724e+09, 8.673409e+09, 8.500278e+09, 8.32802e+09, 8.156796e+09, 
    7.986756e+09, 7.818037e+09, 7.650767e+09, 7.485062e+09, 7.321026e+09, 
    7.158754e+09,
  7.158754e+09, 7.321026e+09, 7.485062e+09, 7.650767e+09, 7.818037e+09, 
    7.986756e+09, 8.156796e+09, 8.32802e+09, 8.500278e+09, 8.673409e+09, 
    8.84724e+09, 9.021585e+09, 9.196247e+09, 9.371016e+09, 9.54567e+09, 
    9.719975e+09, 9.893683e+09, 1.006654e+10, 1.023827e+10, 1.040861e+10, 
    1.057725e+10, 1.07439e+10, 1.090825e+10, 1.106999e+10, 1.122879e+10, 
    1.138432e+10, 1.153626e+10, 1.168427e+10, 1.1828e+10, 1.196713e+10, 
    1.210132e+10, 1.223023e+10, 1.235355e+10, 1.247093e+10, 1.258209e+10, 
    1.268671e+10, 1.27845e+10, 1.287519e+10, 1.295852e+10, 1.303425e+10, 
    1.310215e+10, 1.316203e+10, 1.32137e+10, 1.3257e+10, 1.32918e+10, 
    1.3318e+10, 1.333551e+10, 1.334428e+10, 1.334428e+10, 1.333551e+10, 
    1.3318e+10, 1.32918e+10, 1.3257e+10, 1.32137e+10, 1.316203e+10, 
    1.310215e+10, 1.303425e+10, 1.295852e+10, 1.287519e+10, 1.27845e+10, 
    1.268671e+10, 1.258209e+10, 1.247093e+10, 1.235355e+10, 1.223023e+10, 
    1.210132e+10, 1.196713e+10, 1.1828e+10, 1.168427e+10, 1.153626e+10, 
    1.138432e+10, 1.122879e+10, 1.106999e+10, 1.090825e+10, 1.07439e+10, 
    1.057725e+10, 1.040861e+10, 1.023827e+10, 1.006654e+10, 9.893683e+09, 
    9.719975e+09, 9.54567e+09, 9.371016e+09, 9.196247e+09, 9.021585e+09, 
    8.84724e+09, 8.673409e+09, 8.500278e+09, 8.32802e+09, 8.156796e+09, 
    7.986756e+09, 7.818037e+09, 7.650767e+09, 7.485062e+09, 7.321026e+09, 
    7.158754e+09,
  7.157529e+09, 7.319673e+09, 7.483577e+09, 7.649145e+09, 7.816271e+09, 
    7.984841e+09, 8.154726e+09, 8.32579e+09, 8.497883e+09, 8.670843e+09, 
    8.844498e+09, 9.018663e+09, 9.193139e+09, 9.367718e+09, 9.542177e+09, 
    9.716282e+09, 9.88979e+09, 1.006244e+10, 1.023397e+10, 1.040409e+10, 
    1.057252e+10, 1.073895e+10, 1.090309e+10, 1.106461e+10, 1.12232e+10, 
    1.137852e+10, 1.153025e+10, 1.167804e+10, 1.182158e+10, 1.19605e+10, 
    1.209449e+10, 1.222321e+10, 1.234634e+10, 1.246355e+10, 1.257453e+10, 
    1.267899e+10, 1.277663e+10, 1.286718e+10, 1.295038e+10, 1.302599e+10, 
    1.309378e+10, 1.315356e+10, 1.320514e+10, 1.324837e+10, 1.328312e+10, 
    1.330927e+10, 1.332675e+10, 1.333551e+10, 1.333551e+10, 1.332675e+10, 
    1.330927e+10, 1.328312e+10, 1.324837e+10, 1.320514e+10, 1.315356e+10, 
    1.309378e+10, 1.302599e+10, 1.295038e+10, 1.286718e+10, 1.277663e+10, 
    1.267899e+10, 1.257453e+10, 1.246355e+10, 1.234634e+10, 1.222321e+10, 
    1.209449e+10, 1.19605e+10, 1.182158e+10, 1.167804e+10, 1.153025e+10, 
    1.137852e+10, 1.12232e+10, 1.106461e+10, 1.090309e+10, 1.073895e+10, 
    1.057252e+10, 1.040409e+10, 1.023397e+10, 1.006244e+10, 9.88979e+09, 
    9.716282e+09, 9.542177e+09, 9.367718e+09, 9.193139e+09, 9.018663e+09, 
    8.844498e+09, 8.670843e+09, 8.497883e+09, 8.32579e+09, 8.154726e+09, 
    7.984841e+09, 7.816271e+09, 7.649145e+09, 7.483577e+09, 7.319673e+09, 
    7.157529e+09,
  7.155078e+09, 7.316969e+09, 7.480609e+09, 7.645901e+09, 7.812741e+09, 
    7.981012e+09, 8.150589e+09, 8.321333e+09, 8.493095e+09, 8.665715e+09, 
    8.839017e+09, 9.012821e+09, 9.186927e+09, 9.361125e+09, 9.535196e+09, 
    9.708905e+09, 9.882009e+09, 1.005425e+10, 1.022536e+10, 1.039506e+10, 
    1.056306e+10, 1.072907e+10, 1.089278e+10, 1.105388e+10, 1.121203e+10, 
    1.136693e+10, 1.151823e+10, 1.166561e+10, 1.180873e+10, 1.194726e+10, 
    1.208085e+10, 1.220919e+10, 1.233195e+10, 1.24488e+10, 1.255944e+10, 
    1.266358e+10, 1.276091e+10, 1.285118e+10, 1.293411e+10, 1.300948e+10, 
    1.307706e+10, 1.313664e+10, 1.318806e+10, 1.323115e+10, 1.326578e+10, 
    1.329185e+10, 1.330927e+10, 1.3318e+10, 1.3318e+10, 1.330927e+10, 
    1.329185e+10, 1.326578e+10, 1.323115e+10, 1.318806e+10, 1.313664e+10, 
    1.307706e+10, 1.300948e+10, 1.293411e+10, 1.285118e+10, 1.276091e+10, 
    1.266358e+10, 1.255944e+10, 1.24488e+10, 1.233195e+10, 1.220919e+10, 
    1.208085e+10, 1.194726e+10, 1.180873e+10, 1.166561e+10, 1.151823e+10, 
    1.136693e+10, 1.121203e+10, 1.105388e+10, 1.089278e+10, 1.072907e+10, 
    1.056306e+10, 1.039506e+10, 1.022536e+10, 1.005425e+10, 9.882009e+09, 
    9.708905e+09, 9.535196e+09, 9.361125e+09, 9.186927e+09, 9.012821e+09, 
    8.839017e+09, 8.665715e+09, 8.493095e+09, 8.321333e+09, 8.150589e+09, 
    7.981012e+09, 7.812741e+09, 7.645901e+09, 7.480609e+09, 7.316969e+09, 
    7.155078e+09,
  7.151404e+09, 7.312915e+09, 7.476158e+09, 7.641037e+09, 7.807448e+09, 
    7.975273e+09, 8.144387e+09, 8.314652e+09, 8.485919e+09, 8.658028e+09, 
    8.830806e+09, 9.004068e+09, 9.177618e+09, 9.351248e+09, 9.524738e+09, 
    9.697854e+09, 9.870353e+09, 1.004198e+10, 1.021247e+10, 1.038154e+10, 
    1.054891e+10, 1.071428e+10, 1.087735e+10, 1.10378e+10, 1.119532e+10, 
    1.134958e+10, 1.150025e+10, 1.164701e+10, 1.178951e+10, 1.192743e+10, 
    1.206044e+10, 1.218821e+10, 1.231041e+10, 1.242673e+10, 1.253687e+10, 
    1.264052e+10, 1.273739e+10, 1.282723e+10, 1.290977e+10, 1.298478e+10, 
    1.305203e+10, 1.311133e+10, 1.316249e+10, 1.320537e+10, 1.323984e+10, 
    1.326578e+10, 1.328312e+10, 1.32918e+10, 1.32918e+10, 1.328312e+10, 
    1.326578e+10, 1.323984e+10, 1.320537e+10, 1.316249e+10, 1.311133e+10, 
    1.305203e+10, 1.298478e+10, 1.290977e+10, 1.282723e+10, 1.273739e+10, 
    1.264052e+10, 1.253687e+10, 1.242673e+10, 1.231041e+10, 1.218821e+10, 
    1.206044e+10, 1.192743e+10, 1.178951e+10, 1.164701e+10, 1.150025e+10, 
    1.134958e+10, 1.119532e+10, 1.10378e+10, 1.087735e+10, 1.071428e+10, 
    1.054891e+10, 1.038154e+10, 1.021247e+10, 1.004198e+10, 9.870353e+09, 
    9.697854e+09, 9.524738e+09, 9.351248e+09, 9.177618e+09, 9.004068e+09, 
    8.830806e+09, 8.658028e+09, 8.485919e+09, 8.314652e+09, 8.144387e+09, 
    7.975273e+09, 7.807448e+09, 7.641037e+09, 7.476158e+09, 7.312915e+09, 
    7.151404e+09,
  7.146505e+09, 7.307511e+09, 7.470226e+09, 7.634556e+09, 7.800395e+09, 
    7.967627e+09, 8.136126e+09, 8.305754e+09, 8.476363e+09, 8.647793e+09, 
    8.819871e+09, 8.992415e+09, 9.165227e+09, 9.338102e+09, 9.510819e+09, 
    9.683147e+09, 9.854844e+09, 1.002566e+10, 1.019532e+10, 1.036355e+10, 
    1.053008e+10, 1.06946e+10, 1.085682e+10, 1.101642e+10, 1.117309e+10, 
    1.13265e+10, 1.147634e+10, 1.162227e+10, 1.176396e+10, 1.190108e+10, 
    1.203331e+10, 1.216031e+10, 1.228178e+10, 1.23974e+10, 1.250686e+10, 
    1.260987e+10, 1.270614e+10, 1.279542e+10, 1.287743e+10, 1.295196e+10, 
    1.301878e+10, 1.30777e+10, 1.312854e+10, 1.317114e+10, 1.320537e+10, 
    1.323115e+10, 1.324837e+10, 1.3257e+10, 1.3257e+10, 1.324837e+10, 
    1.323115e+10, 1.320537e+10, 1.317114e+10, 1.312854e+10, 1.30777e+10, 
    1.301878e+10, 1.295196e+10, 1.287743e+10, 1.279542e+10, 1.270614e+10, 
    1.260987e+10, 1.250686e+10, 1.23974e+10, 1.228178e+10, 1.216031e+10, 
    1.203331e+10, 1.190108e+10, 1.176396e+10, 1.162227e+10, 1.147634e+10, 
    1.13265e+10, 1.117309e+10, 1.101642e+10, 1.085682e+10, 1.06946e+10, 
    1.053008e+10, 1.036355e+10, 1.019532e+10, 1.002566e+10, 9.854844e+09, 
    9.683147e+09, 9.510819e+09, 9.338102e+09, 9.165227e+09, 8.992415e+09, 
    8.819871e+09, 8.647793e+09, 8.476363e+09, 8.305754e+09, 8.136126e+09, 
    7.967627e+09, 7.800395e+09, 7.634556e+09, 7.470226e+09, 7.307511e+09, 
    7.146505e+09,
  7.140384e+09, 7.30076e+09, 7.462817e+09, 7.626462e+09, 7.791588e+09, 
    7.958081e+09, 8.125813e+09, 8.294647e+09, 8.464436e+09, 8.63502e+09, 
    8.806228e+09, 8.977876e+09, 9.14977e+09, 9.321703e+09, 9.49346e+09, 
    9.664807e+09, 9.835507e+09, 1.00053e+10, 1.017394e+10, 1.034114e+10, 
    1.050662e+10, 1.067009e+10, 1.083124e+10, 1.098979e+10, 1.11454e+10, 
    1.129776e+10, 1.144656e+10, 1.159146e+10, 1.173213e+10, 1.186826e+10, 
    1.199952e+10, 1.212559e+10, 1.224615e+10, 1.236089e+10, 1.246951e+10, 
    1.257172e+10, 1.266725e+10, 1.275582e+10, 1.283719e+10, 1.291113e+10, 
    1.297741e+10, 1.303585e+10, 1.308628e+10, 1.312854e+10, 1.316249e+10, 
    1.318806e+10, 1.320514e+10, 1.32137e+10, 1.32137e+10, 1.320514e+10, 
    1.318806e+10, 1.316249e+10, 1.312854e+10, 1.308628e+10, 1.303585e+10, 
    1.297741e+10, 1.291113e+10, 1.283719e+10, 1.275582e+10, 1.266725e+10, 
    1.257172e+10, 1.246951e+10, 1.236089e+10, 1.224615e+10, 1.212559e+10, 
    1.199952e+10, 1.186826e+10, 1.173213e+10, 1.159146e+10, 1.144656e+10, 
    1.129776e+10, 1.11454e+10, 1.098979e+10, 1.083124e+10, 1.067009e+10, 
    1.050662e+10, 1.034114e+10, 1.017394e+10, 1.00053e+10, 9.835507e+09, 
    9.664807e+09, 9.49346e+09, 9.321703e+09, 9.14977e+09, 8.977876e+09, 
    8.806228e+09, 8.63502e+09, 8.464436e+09, 8.294647e+09, 8.125813e+09, 
    7.958081e+09, 7.791588e+09, 7.626462e+09, 7.462817e+09, 7.30076e+09, 
    7.140384e+09,
  7.133041e+09, 7.292662e+09, 7.453934e+09, 7.616759e+09, 7.781033e+09, 
    7.946641e+09, 8.113456e+09, 8.281342e+09, 8.450151e+09, 8.619724e+09, 
    8.789891e+09, 8.96047e+09, 9.131267e+09, 9.302078e+09, 9.472687e+09, 
    9.642865e+09, 9.812372e+09, 9.980962e+09, 1.014837e+10, 1.031433e+10, 
    1.047856e+10, 1.064077e+10, 1.080067e+10, 1.095795e+10, 1.111231e+10, 
    1.126342e+10, 1.141097e+10, 1.155465e+10, 1.169412e+10, 1.182907e+10, 
    1.195917e+10, 1.208412e+10, 1.220359e+10, 1.231729e+10, 1.242492e+10, 
    1.252618e+10, 1.262082e+10, 1.270856e+10, 1.278916e+10, 1.286239e+10, 
    1.292804e+10, 1.298592e+10, 1.303585e+10, 1.30777e+10, 1.311133e+10, 
    1.313664e+10, 1.315356e+10, 1.316203e+10, 1.316203e+10, 1.315356e+10, 
    1.313664e+10, 1.311133e+10, 1.30777e+10, 1.303585e+10, 1.298592e+10, 
    1.292804e+10, 1.286239e+10, 1.278916e+10, 1.270856e+10, 1.262082e+10, 
    1.252618e+10, 1.242492e+10, 1.231729e+10, 1.220359e+10, 1.208412e+10, 
    1.195917e+10, 1.182907e+10, 1.169412e+10, 1.155465e+10, 1.141097e+10, 
    1.126342e+10, 1.111231e+10, 1.095795e+10, 1.080067e+10, 1.064077e+10, 
    1.047856e+10, 1.031433e+10, 1.014837e+10, 9.980962e+09, 9.812372e+09, 
    9.642865e+09, 9.472687e+09, 9.302078e+09, 9.131267e+09, 8.96047e+09, 
    8.789891e+09, 8.619724e+09, 8.450151e+09, 8.281342e+09, 8.113456e+09, 
    7.946641e+09, 7.781033e+09, 7.616759e+09, 7.453934e+09, 7.292662e+09, 
    7.133041e+09,
  7.124479e+09, 7.283223e+09, 7.443579e+09, 7.605452e+09, 7.768736e+09, 
    7.933316e+09, 8.099066e+09, 8.26585e+09, 8.433522e+09, 8.601922e+09, 
    8.770882e+09, 8.940219e+09, 9.109745e+09, 9.279254e+09, 9.448532e+09, 
    9.617354e+09, 9.785482e+09, 9.95267e+09, 1.011866e+10, 1.028319e+10, 
    1.044597e+10, 1.060673e+10, 1.076517e+10, 1.092099e+10, 1.107389e+10, 
    1.122356e+10, 1.136968e+10, 1.151193e+10, 1.165001e+10, 1.17836e+10, 
    1.191237e+10, 1.203602e+10, 1.215424e+10, 1.226673e+10, 1.237321e+10, 
    1.247338e+10, 1.256699e+10, 1.265377e+10, 1.273348e+10, 1.280589e+10, 
    1.287081e+10, 1.292804e+10, 1.297741e+10, 1.301878e+10, 1.305203e+10, 
    1.307706e+10, 1.309378e+10, 1.310215e+10, 1.310215e+10, 1.309378e+10, 
    1.307706e+10, 1.305203e+10, 1.301878e+10, 1.297741e+10, 1.292804e+10, 
    1.287081e+10, 1.280589e+10, 1.273348e+10, 1.265377e+10, 1.256699e+10, 
    1.247338e+10, 1.237321e+10, 1.226673e+10, 1.215424e+10, 1.203602e+10, 
    1.191237e+10, 1.17836e+10, 1.165001e+10, 1.151193e+10, 1.136968e+10, 
    1.122356e+10, 1.107389e+10, 1.092099e+10, 1.076517e+10, 1.060673e+10, 
    1.044597e+10, 1.028319e+10, 1.011866e+10, 9.95267e+09, 9.785482e+09, 
    9.617354e+09, 9.448532e+09, 9.279254e+09, 9.109745e+09, 8.940219e+09, 
    8.770882e+09, 8.601922e+09, 8.433522e+09, 8.26585e+09, 8.099066e+09, 
    7.933316e+09, 7.768736e+09, 7.605452e+09, 7.443579e+09, 7.283223e+09, 
    7.124479e+09,
  7.1147e+09, 7.272444e+09, 7.431758e+09, 7.592547e+09, 7.754704e+09, 
    7.918115e+09, 8.082655e+09, 8.248187e+09, 8.414565e+09, 8.581632e+09, 
    8.749221e+09, 8.917151e+09, 9.085231e+09, 9.253263e+09, 9.421031e+09, 
    9.588315e+09, 9.754878e+09, 9.920478e+09, 1.008486e+10, 1.024776e+10, 
    1.040891e+10, 1.056802e+10, 1.07248e+10, 1.087898e+10, 1.103023e+10, 
    1.117826e+10, 1.132276e+10, 1.146341e+10, 1.159992e+10, 1.173195e+10, 
    1.185922e+10, 1.198141e+10, 1.209821e+10, 1.220935e+10, 1.231452e+10, 
    1.241347e+10, 1.250591e+10, 1.25916e+10, 1.267031e+10, 1.27418e+10, 
    1.280589e+10, 1.286239e+10, 1.291113e+10, 1.295196e+10, 1.298478e+10, 
    1.300948e+10, 1.302599e+10, 1.303425e+10, 1.303425e+10, 1.302599e+10, 
    1.300948e+10, 1.298478e+10, 1.295196e+10, 1.291113e+10, 1.286239e+10, 
    1.280589e+10, 1.27418e+10, 1.267031e+10, 1.25916e+10, 1.250591e+10, 
    1.241347e+10, 1.231452e+10, 1.220935e+10, 1.209821e+10, 1.198141e+10, 
    1.185922e+10, 1.173195e+10, 1.159992e+10, 1.146341e+10, 1.132276e+10, 
    1.117826e+10, 1.103023e+10, 1.087898e+10, 1.07248e+10, 1.056802e+10, 
    1.040891e+10, 1.024776e+10, 1.008486e+10, 9.920478e+09, 9.754878e+09, 
    9.588315e+09, 9.421031e+09, 9.253263e+09, 9.085231e+09, 8.917151e+09, 
    8.749221e+09, 8.581632e+09, 8.414565e+09, 8.248187e+09, 8.082655e+09, 
    7.918115e+09, 7.754704e+09, 7.592547e+09, 7.431758e+09, 7.272444e+09, 
    7.1147e+09,
  7.103705e+09, 7.260329e+09, 7.418477e+09, 7.578052e+09, 7.738948e+09, 
    7.901051e+09, 8.064236e+09, 8.228367e+09, 8.3933e+09, 8.558878e+09, 
    8.724934e+09, 8.891291e+09, 9.05776e+09, 9.224142e+09, 9.390226e+09, 
    9.555794e+09, 9.720613e+09, 9.884442e+09, 1.004703e+10, 1.020812e+10, 
    1.036744e+10, 1.052472e+10, 1.067967e+10, 1.0832e+10, 1.098142e+10, 
    1.112763e+10, 1.127033e+10, 1.14092e+10, 1.154395e+10, 1.167428e+10, 
    1.179987e+10, 1.192043e+10, 1.203567e+10, 1.214529e+10, 1.224902e+10, 
    1.234659e+10, 1.243775e+10, 1.252223e+10, 1.259983e+10, 1.267031e+10, 
    1.273348e+10, 1.278916e+10, 1.283719e+10, 1.287743e+10, 1.290977e+10, 
    1.293411e+10, 1.295038e+10, 1.295852e+10, 1.295852e+10, 1.295038e+10, 
    1.293411e+10, 1.290977e+10, 1.287743e+10, 1.283719e+10, 1.278916e+10, 
    1.273348e+10, 1.267031e+10, 1.259983e+10, 1.252223e+10, 1.243775e+10, 
    1.234659e+10, 1.224902e+10, 1.214529e+10, 1.203567e+10, 1.192043e+10, 
    1.179987e+10, 1.167428e+10, 1.154395e+10, 1.14092e+10, 1.127033e+10, 
    1.112763e+10, 1.098142e+10, 1.0832e+10, 1.067967e+10, 1.052472e+10, 
    1.036744e+10, 1.020812e+10, 1.004703e+10, 9.884442e+09, 9.720613e+09, 
    9.555794e+09, 9.390226e+09, 9.224142e+09, 9.05776e+09, 8.891291e+09, 
    8.724934e+09, 8.558878e+09, 8.3933e+09, 8.228367e+09, 8.064236e+09, 
    7.901051e+09, 7.738948e+09, 7.578052e+09, 7.418477e+09, 7.260329e+09, 
    7.103705e+09,
  7.091497e+09, 7.246883e+09, 7.403741e+09, 7.561974e+09, 7.721477e+09, 
    7.882135e+09, 8.043825e+09, 8.20641e+09, 8.369748e+09, 8.533684e+09, 
    8.698051e+09, 8.862674e+09, 9.027367e+09, 9.191932e+09, 9.356163e+09, 
    9.519842e+09, 9.68274e+09, 9.844622e+09, 1.000524e+10, 1.016434e+10, 
    1.032166e+10, 1.047692e+10, 1.062985e+10, 1.078017e+10, 1.092757e+10, 
    1.107179e+10, 1.12125e+10, 1.134943e+10, 1.148226e+10, 1.16107e+10, 
    1.173446e+10, 1.185324e+10, 1.196675e+10, 1.207473e+10, 1.217688e+10, 
    1.227295e+10, 1.236269e+10, 1.244586e+10, 1.252223e+10, 1.25916e+10, 
    1.265377e+10, 1.270856e+10, 1.275582e+10, 1.279542e+10, 1.282723e+10, 
    1.285118e+10, 1.286718e+10, 1.287519e+10, 1.287519e+10, 1.286718e+10, 
    1.285118e+10, 1.282723e+10, 1.279542e+10, 1.275582e+10, 1.270856e+10, 
    1.265377e+10, 1.25916e+10, 1.252223e+10, 1.244586e+10, 1.236269e+10, 
    1.227295e+10, 1.217688e+10, 1.207473e+10, 1.196675e+10, 1.185324e+10, 
    1.173446e+10, 1.16107e+10, 1.148226e+10, 1.134943e+10, 1.12125e+10, 
    1.107179e+10, 1.092757e+10, 1.078017e+10, 1.062985e+10, 1.047692e+10, 
    1.032166e+10, 1.016434e+10, 1.000524e+10, 9.844622e+09, 9.68274e+09, 
    9.519842e+09, 9.356163e+09, 9.191932e+09, 9.027367e+09, 8.862674e+09, 
    8.698051e+09, 8.533684e+09, 8.369748e+09, 8.20641e+09, 8.043825e+09, 
    7.882135e+09, 7.721477e+09, 7.561974e+09, 7.403741e+09, 7.246883e+09, 
    7.091497e+09,
  7.078078e+09, 7.23211e+09, 7.387556e+09, 7.544322e+09, 7.702302e+09, 
    7.861382e+09, 8.021437e+09, 8.182336e+09, 8.343933e+09, 8.506077e+09, 
    8.668601e+09, 8.831335e+09, 8.994092e+09, 9.156679e+09, 9.318892e+09, 
    9.480515e+09, 9.641325e+09, 9.801088e+09, 9.959563e+09, 1.01165e+10, 
    1.027164e+10, 1.042471e+10, 1.057545e+10, 1.072358e+10, 1.08688e+10, 
    1.101085e+10, 1.114942e+10, 1.128423e+10, 1.141498e+10, 1.154138e+10, 
    1.166315e+10, 1.178001e+10, 1.189166e+10, 1.199784e+10, 1.209829e+10, 
    1.219274e+10, 1.228095e+10, 1.236269e+10, 1.243775e+10, 1.250591e+10, 
    1.256699e+10, 1.262082e+10, 1.266725e+10, 1.270614e+10, 1.273739e+10, 
    1.276091e+10, 1.277663e+10, 1.27845e+10, 1.27845e+10, 1.277663e+10, 
    1.276091e+10, 1.273739e+10, 1.270614e+10, 1.266725e+10, 1.262082e+10, 
    1.256699e+10, 1.250591e+10, 1.243775e+10, 1.236269e+10, 1.228095e+10, 
    1.219274e+10, 1.209829e+10, 1.199784e+10, 1.189166e+10, 1.178001e+10, 
    1.166315e+10, 1.154138e+10, 1.141498e+10, 1.128423e+10, 1.114942e+10, 
    1.101085e+10, 1.08688e+10, 1.072358e+10, 1.057545e+10, 1.042471e+10, 
    1.027164e+10, 1.01165e+10, 9.959563e+09, 9.801088e+09, 9.641325e+09, 
    9.480515e+09, 9.318892e+09, 9.156679e+09, 8.994092e+09, 8.831335e+09, 
    8.668601e+09, 8.506077e+09, 8.343933e+09, 8.182336e+09, 8.021437e+09, 
    7.861382e+09, 7.702302e+09, 7.544322e+09, 7.387556e+09, 7.23211e+09, 
    7.078078e+09,
  7.063453e+09, 7.216014e+09, 7.36993e+09, 7.525106e+09, 7.681435e+09, 
    7.838806e+09, 7.997093e+09, 8.156166e+09, 8.31588e+09, 8.476086e+09, 
    8.636621e+09, 8.797313e+09, 8.95798e+09, 9.118431e+09, 9.278465e+09, 
    9.437871e+09, 9.596429e+09, 9.753911e+09, 9.910078e+09, 1.006469e+10, 
    1.021748e+10, 1.03682e+10, 1.051658e+10, 1.066235e+10, 1.080523e+10, 
    1.094495e+10, 1.108122e+10, 1.121375e+10, 1.134227e+10, 1.146649e+10, 
    1.158613e+10, 1.170091e+10, 1.181057e+10, 1.191483e+10, 1.201345e+10, 
    1.210616e+10, 1.219274e+10, 1.227295e+10, 1.234659e+10, 1.241347e+10, 
    1.247338e+10, 1.252618e+10, 1.257172e+10, 1.260987e+10, 1.264052e+10, 
    1.266358e+10, 1.267899e+10, 1.268671e+10, 1.268671e+10, 1.267899e+10, 
    1.266358e+10, 1.264052e+10, 1.260987e+10, 1.257172e+10, 1.252618e+10, 
    1.247338e+10, 1.241347e+10, 1.234659e+10, 1.227295e+10, 1.219274e+10, 
    1.210616e+10, 1.201345e+10, 1.191483e+10, 1.181057e+10, 1.170091e+10, 
    1.158613e+10, 1.146649e+10, 1.134227e+10, 1.121375e+10, 1.108122e+10, 
    1.094495e+10, 1.080523e+10, 1.066235e+10, 1.051658e+10, 1.03682e+10, 
    1.021748e+10, 1.006469e+10, 9.910078e+09, 9.753911e+09, 9.596429e+09, 
    9.437871e+09, 9.278465e+09, 9.118431e+09, 8.95798e+09, 8.797313e+09, 
    8.636621e+09, 8.476086e+09, 8.31588e+09, 8.156166e+09, 7.997093e+09, 
    7.838806e+09, 7.681435e+09, 7.525106e+09, 7.36993e+09, 7.216014e+09, 
    7.063453e+09,
  7.047623e+09, 7.198601e+09, 7.350871e+09, 7.504335e+09, 7.65889e+09, 
    7.814423e+09, 7.970811e+09, 8.127923e+09, 8.285618e+09, 8.443745e+09, 
    8.602145e+09, 8.760649e+09, 8.919077e+09, 9.077242e+09, 9.234944e+09, 
    9.391978e+09, 9.548129e+09, 9.703171e+09, 9.856871e+09, 1.000899e+10, 
    1.015928e+10, 1.030749e+10, 1.045336e+10, 1.059662e+10, 1.0737e+10, 
    1.087423e+10, 1.100805e+10, 1.113816e+10, 1.12643e+10, 1.13862e+10, 
    1.150357e+10, 1.161615e+10, 1.172369e+10, 1.182591e+10, 1.192258e+10, 
    1.201345e+10, 1.209829e+10, 1.217688e+10, 1.224902e+10, 1.231452e+10, 
    1.237321e+10, 1.242492e+10, 1.246951e+10, 1.250686e+10, 1.253687e+10, 
    1.255944e+10, 1.257453e+10, 1.258209e+10, 1.258209e+10, 1.257453e+10, 
    1.255944e+10, 1.253687e+10, 1.250686e+10, 1.246951e+10, 1.242492e+10, 
    1.237321e+10, 1.231452e+10, 1.224902e+10, 1.217688e+10, 1.209829e+10, 
    1.201345e+10, 1.192258e+10, 1.182591e+10, 1.172369e+10, 1.161615e+10, 
    1.150357e+10, 1.13862e+10, 1.12643e+10, 1.113816e+10, 1.100805e+10, 
    1.087423e+10, 1.0737e+10, 1.059662e+10, 1.045336e+10, 1.030749e+10, 
    1.015928e+10, 1.000899e+10, 9.856871e+09, 9.703171e+09, 9.548129e+09, 
    9.391978e+09, 9.234944e+09, 9.077242e+09, 8.919077e+09, 8.760649e+09, 
    8.602145e+09, 8.443745e+09, 8.285618e+09, 8.127923e+09, 7.970811e+09, 
    7.814423e+09, 7.65889e+09, 7.504335e+09, 7.350871e+09, 7.198601e+09, 
    7.047623e+09,
  7.030593e+09, 7.179877e+09, 7.330385e+09, 7.482021e+09, 7.634681e+09, 
    7.788252e+09, 7.942612e+09, 8.097633e+09, 8.253174e+09, 8.409087e+09, 
    8.565214e+09, 8.721389e+09, 8.877434e+09, 9.033167e+09, 9.188391e+09, 
    9.342905e+09, 9.496498e+09, 9.64895e+09, 9.800034e+09, 9.949515e+09, 
    1.009715e+10, 1.02427e+10, 1.03859e+10, 1.05265e+10, 1.066424e+10, 
    1.079885e+10, 1.093007e+10, 1.105763e+10, 1.118125e+10, 1.130069e+10, 
    1.141567e+10, 1.152593e+10, 1.163122e+10, 1.17313e+10, 1.182591e+10, 
    1.191483e+10, 1.199784e+10, 1.207473e+10, 1.214529e+10, 1.220935e+10, 
    1.226673e+10, 1.231729e+10, 1.236089e+10, 1.23974e+10, 1.242673e+10, 
    1.24488e+10, 1.246355e+10, 1.247093e+10, 1.247093e+10, 1.246355e+10, 
    1.24488e+10, 1.242673e+10, 1.23974e+10, 1.236089e+10, 1.231729e+10, 
    1.226673e+10, 1.220935e+10, 1.214529e+10, 1.207473e+10, 1.199784e+10, 
    1.191483e+10, 1.182591e+10, 1.17313e+10, 1.163122e+10, 1.152593e+10, 
    1.141567e+10, 1.130069e+10, 1.118125e+10, 1.105763e+10, 1.093007e+10, 
    1.079885e+10, 1.066424e+10, 1.05265e+10, 1.03859e+10, 1.02427e+10, 
    1.009715e+10, 9.949515e+09, 9.800034e+09, 9.64895e+09, 9.496498e+09, 
    9.342905e+09, 9.188391e+09, 9.033167e+09, 8.877434e+09, 8.721389e+09, 
    8.565214e+09, 8.409087e+09, 8.253174e+09, 8.097633e+09, 7.942612e+09, 
    7.788252e+09, 7.634681e+09, 7.482021e+09, 7.330385e+09, 7.179877e+09, 
    7.030593e+09,
  7.012366e+09, 7.159848e+09, 7.308484e+09, 7.458176e+09, 7.608822e+09, 
    7.760311e+09, 7.912521e+09, 8.065324e+09, 8.218582e+09, 8.372148e+09, 
    8.525868e+09, 8.679578e+09, 8.833104e+09, 8.986266e+09, 9.138871e+09, 
    9.290724e+09, 9.441618e+09, 9.591338e+09, 9.739662e+09, 9.886363e+09, 
    1.00312e+10, 1.017395e+10, 1.031435e+10, 1.045215e+10, 1.058711e+10, 
    1.071896e+10, 1.084745e+10, 1.097232e+10, 1.109331e+10, 1.121017e+10, 
    1.132264e+10, 1.143046e+10, 1.153341e+10, 1.163122e+10, 1.172369e+10, 
    1.181057e+10, 1.189166e+10, 1.196675e+10, 1.203567e+10, 1.209821e+10, 
    1.215424e+10, 1.220359e+10, 1.224615e+10, 1.228178e+10, 1.231041e+10, 
    1.233195e+10, 1.234634e+10, 1.235355e+10, 1.235355e+10, 1.234634e+10, 
    1.233195e+10, 1.231041e+10, 1.228178e+10, 1.224615e+10, 1.220359e+10, 
    1.215424e+10, 1.209821e+10, 1.203567e+10, 1.196675e+10, 1.189166e+10, 
    1.181057e+10, 1.172369e+10, 1.163122e+10, 1.153341e+10, 1.143046e+10, 
    1.132264e+10, 1.121017e+10, 1.109331e+10, 1.097232e+10, 1.084745e+10, 
    1.071896e+10, 1.058711e+10, 1.045215e+10, 1.031435e+10, 1.017395e+10, 
    1.00312e+10, 9.886363e+09, 9.739662e+09, 9.591338e+09, 9.441618e+09, 
    9.290724e+09, 9.138871e+09, 8.986266e+09, 8.833104e+09, 8.679578e+09, 
    8.525868e+09, 8.372148e+09, 8.218582e+09, 8.065324e+09, 7.912521e+09, 
    7.760311e+09, 7.608822e+09, 7.458176e+09, 7.308484e+09, 7.159848e+09, 
    7.012366e+09,
  6.992947e+09, 7.138521e+09, 7.285175e+09, 7.432813e+09, 7.581331e+09, 
    7.73062e+09, 7.880559e+09, 8.031022e+09, 8.181873e+09, 8.332967e+09, 
    8.484152e+09, 8.635267e+09, 8.786142e+09, 8.936601e+09, 9.086456e+09, 
    9.235513e+09, 9.383574e+09, 9.530426e+09, 9.675857e+09, 9.819643e+09, 
    9.961556e+09, 1.010136e+10, 1.023883e+10, 1.037371e+10, 1.050575e+10, 
    1.063472e+10, 1.076036e+10, 1.088243e+10, 1.100067e+10, 1.111483e+10, 
    1.122468e+10, 1.132997e+10, 1.143046e+10, 1.152593e+10, 1.161615e+10, 
    1.170091e+10, 1.178001e+10, 1.185324e+10, 1.192043e+10, 1.198141e+10, 
    1.203602e+10, 1.208412e+10, 1.212559e+10, 1.216031e+10, 1.218821e+10, 
    1.220919e+10, 1.222321e+10, 1.223023e+10, 1.223023e+10, 1.222321e+10, 
    1.220919e+10, 1.218821e+10, 1.216031e+10, 1.212559e+10, 1.208412e+10, 
    1.203602e+10, 1.198141e+10, 1.192043e+10, 1.185324e+10, 1.178001e+10, 
    1.170091e+10, 1.161615e+10, 1.152593e+10, 1.143046e+10, 1.132997e+10, 
    1.122468e+10, 1.111483e+10, 1.100067e+10, 1.088243e+10, 1.076036e+10, 
    1.063472e+10, 1.050575e+10, 1.037371e+10, 1.023883e+10, 1.010136e+10, 
    9.961556e+09, 9.819643e+09, 9.675857e+09, 9.530426e+09, 9.383574e+09, 
    9.235513e+09, 9.086456e+09, 8.936601e+09, 8.786142e+09, 8.635267e+09, 
    8.484152e+09, 8.332967e+09, 8.181873e+09, 8.031022e+09, 7.880559e+09, 
    7.73062e+09, 7.581331e+09, 7.432813e+09, 7.285175e+09, 7.138521e+09, 
    6.992947e+09,
  6.972339e+09, 7.115902e+09, 7.260469e+09, 7.405943e+09, 7.552224e+09, 
    7.699199e+09, 7.846753e+09, 7.994759e+09, 8.143084e+09, 8.291585e+09, 
    8.440113e+09, 8.58851e+09, 8.736609e+09, 8.884238e+09, 9.031216e+09, 
    9.177352e+09, 9.322452e+09, 9.466312e+09, 9.608722e+09, 9.749469e+09, 
    9.88833e+09, 1.002508e+10, 1.015949e+10, 1.029132e+10, 1.042034e+10, 
    1.054631e+10, 1.066899e+10, 1.078814e+10, 1.090352e+10, 1.10149e+10, 
    1.112203e+10, 1.122468e+10, 1.132264e+10, 1.141567e+10, 1.150357e+10, 
    1.158613e+10, 1.166315e+10, 1.173446e+10, 1.179987e+10, 1.185922e+10, 
    1.191237e+10, 1.195917e+10, 1.199952e+10, 1.203331e+10, 1.206044e+10, 
    1.208085e+10, 1.209449e+10, 1.210132e+10, 1.210132e+10, 1.209449e+10, 
    1.208085e+10, 1.206044e+10, 1.203331e+10, 1.199952e+10, 1.195917e+10, 
    1.191237e+10, 1.185922e+10, 1.179987e+10, 1.173446e+10, 1.166315e+10, 
    1.158613e+10, 1.150357e+10, 1.141567e+10, 1.132264e+10, 1.122468e+10, 
    1.112203e+10, 1.10149e+10, 1.090352e+10, 1.078814e+10, 1.066899e+10, 
    1.054631e+10, 1.042034e+10, 1.029132e+10, 1.015949e+10, 1.002508e+10, 
    9.88833e+09, 9.749469e+09, 9.608722e+09, 9.466312e+09, 9.322452e+09, 
    9.177352e+09, 9.031216e+09, 8.884238e+09, 8.736609e+09, 8.58851e+09, 
    8.440113e+09, 8.291585e+09, 8.143084e+09, 7.994759e+09, 7.846753e+09, 
    7.699199e+09, 7.552224e+09, 7.405943e+09, 7.260469e+09, 7.115902e+09, 
    6.972339e+09,
  6.950547e+09, 7.092e+09, 7.234377e+09, 7.377583e+09, 7.521518e+09, 
    7.666072e+09, 7.811129e+09, 7.956566e+09, 8.10225e+09, 8.248043e+09, 
    8.393798e+09, 8.539359e+09, 8.684566e+09, 8.829247e+09, 8.973229e+09, 
    9.116325e+09, 9.258346e+09, 9.399095e+09, 9.53837e+09, 9.67596e+09, 
    9.811654e+09, 9.945231e+09, 1.007647e+10, 1.020515e+10, 1.033104e+10, 
    1.045391e+10, 1.057352e+10, 1.068966e+10, 1.080209e+10, 1.091057e+10, 
    1.10149e+10, 1.111483e+10, 1.121017e+10, 1.130069e+10, 1.13862e+10, 
    1.146649e+10, 1.154138e+10, 1.16107e+10, 1.167428e+10, 1.173195e+10, 
    1.17836e+10, 1.182907e+10, 1.186826e+10, 1.190108e+10, 1.192743e+10, 
    1.194726e+10, 1.19605e+10, 1.196713e+10, 1.196713e+10, 1.19605e+10, 
    1.194726e+10, 1.192743e+10, 1.190108e+10, 1.186826e+10, 1.182907e+10, 
    1.17836e+10, 1.173195e+10, 1.167428e+10, 1.16107e+10, 1.154138e+10, 
    1.146649e+10, 1.13862e+10, 1.130069e+10, 1.121017e+10, 1.111483e+10, 
    1.10149e+10, 1.091057e+10, 1.080209e+10, 1.068966e+10, 1.057352e+10, 
    1.045391e+10, 1.033104e+10, 1.020515e+10, 1.007647e+10, 9.945231e+09, 
    9.811654e+09, 9.67596e+09, 9.53837e+09, 9.399095e+09, 9.258346e+09, 
    9.116325e+09, 8.973229e+09, 8.829247e+09, 8.684566e+09, 8.539359e+09, 
    8.393798e+09, 8.248043e+09, 8.10225e+09, 7.956566e+09, 7.811129e+09, 
    7.666072e+09, 7.521518e+09, 7.377583e+09, 7.234377e+09, 7.092e+09, 
    6.950547e+09,
  6.927576e+09, 7.066821e+09, 7.206909e+09, 7.347746e+09, 7.489233e+09, 
    7.631261e+09, 7.773715e+09, 7.916475e+09, 8.059411e+09, 8.202386e+09, 
    8.345257e+09, 8.487873e+09, 8.630074e+09, 8.771699e+09, 8.912572e+09, 
    9.052518e+09, 9.191351e+09, 9.32888e+09, 9.464909e+09, 9.599237e+09, 
    9.731658e+09, 9.861961e+09, 9.989933e+09, 1.011536e+10, 1.023802e+10, 
    1.035769e+10, 1.047415e+10, 1.058718e+10, 1.069657e+10, 1.080209e+10, 
    1.090352e+10, 1.100067e+10, 1.109331e+10, 1.118125e+10, 1.12643e+10, 
    1.134227e+10, 1.141498e+10, 1.148226e+10, 1.154395e+10, 1.159992e+10, 
    1.165001e+10, 1.169412e+10, 1.173213e+10, 1.176396e+10, 1.178951e+10, 
    1.180873e+10, 1.182158e+10, 1.1828e+10, 1.1828e+10, 1.182158e+10, 
    1.180873e+10, 1.178951e+10, 1.176396e+10, 1.173213e+10, 1.169412e+10, 
    1.165001e+10, 1.159992e+10, 1.154395e+10, 1.148226e+10, 1.141498e+10, 
    1.134227e+10, 1.12643e+10, 1.118125e+10, 1.109331e+10, 1.100067e+10, 
    1.090352e+10, 1.080209e+10, 1.069657e+10, 1.058718e+10, 1.047415e+10, 
    1.035769e+10, 1.023802e+10, 1.011536e+10, 9.989933e+09, 9.861961e+09, 
    9.731658e+09, 9.599237e+09, 9.464909e+09, 9.32888e+09, 9.191351e+09, 
    9.052518e+09, 8.912572e+09, 8.771699e+09, 8.630074e+09, 8.487873e+09, 
    8.345257e+09, 8.202386e+09, 8.059411e+09, 7.916475e+09, 7.773715e+09, 
    7.631261e+09, 7.489233e+09, 7.347746e+09, 7.206909e+09, 7.066821e+09, 
    6.927576e+09,
  6.903431e+09, 7.040374e+09, 7.178077e+09, 7.316448e+09, 7.455388e+09, 
    7.594789e+09, 7.734541e+09, 7.874522e+09, 8.014606e+09, 8.15466e+09, 
    8.294543e+09, 8.434108e+09, 8.573202e+09, 8.711665e+09, 8.849328e+09, 
    8.986021e+09, 9.121564e+09, 9.255772e+09, 9.388457e+09, 9.519426e+09, 
    9.648477e+09, 9.775411e+09, 9.900023e+09, 1.00221e+10, 1.014144e+10, 
    1.025783e+10, 1.037106e+10, 1.048091e+10, 1.058718e+10, 1.068966e+10, 
    1.078814e+10, 1.088243e+10, 1.097232e+10, 1.105763e+10, 1.113816e+10, 
    1.121375e+10, 1.128423e+10, 1.134943e+10, 1.14092e+10, 1.146341e+10, 
    1.151193e+10, 1.155465e+10, 1.159146e+10, 1.162227e+10, 1.164701e+10, 
    1.166561e+10, 1.167804e+10, 1.168427e+10, 1.168427e+10, 1.167804e+10, 
    1.166561e+10, 1.164701e+10, 1.162227e+10, 1.159146e+10, 1.155465e+10, 
    1.151193e+10, 1.146341e+10, 1.14092e+10, 1.134943e+10, 1.128423e+10, 
    1.121375e+10, 1.113816e+10, 1.105763e+10, 1.097232e+10, 1.088243e+10, 
    1.078814e+10, 1.068966e+10, 1.058718e+10, 1.048091e+10, 1.037106e+10, 
    1.025783e+10, 1.014144e+10, 1.00221e+10, 9.900023e+09, 9.775411e+09, 
    9.648477e+09, 9.519426e+09, 9.388457e+09, 9.255772e+09, 9.121564e+09, 
    8.986021e+09, 8.849328e+09, 8.711665e+09, 8.573202e+09, 8.434108e+09, 
    8.294543e+09, 8.15466e+09, 8.014606e+09, 7.874522e+09, 7.734541e+09, 
    7.594789e+09, 7.455388e+09, 7.316448e+09, 7.178077e+09, 7.040374e+09, 
    6.903431e+09,
  6.878117e+09, 7.012667e+09, 7.147894e+09, 7.283705e+09, 7.420003e+09, 
    7.556683e+09, 7.693634e+09, 7.830739e+09, 7.967875e+09, 8.10491e+09, 
    8.241709e+09, 8.378128e+09, 8.514017e+09, 8.649221e+09, 8.78358e+09, 
    8.916924e+09, 9.049084e+09, 9.17988e+09, 9.309132e+09, 9.436652e+09, 
    9.562249e+09, 9.68573e+09, 9.806899e+09, 9.925557e+09, 1.00415e+10, 
    1.015454e+10, 1.026446e+10, 1.037106e+10, 1.047415e+10, 1.057352e+10, 
    1.066899e+10, 1.076036e+10, 1.084745e+10, 1.093007e+10, 1.100805e+10, 
    1.108122e+10, 1.114942e+10, 1.12125e+10, 1.127033e+10, 1.132276e+10, 
    1.136968e+10, 1.141097e+10, 1.144656e+10, 1.147634e+10, 1.150025e+10, 
    1.151823e+10, 1.153025e+10, 1.153626e+10, 1.153626e+10, 1.153025e+10, 
    1.151823e+10, 1.150025e+10, 1.147634e+10, 1.144656e+10, 1.141097e+10, 
    1.136968e+10, 1.132276e+10, 1.127033e+10, 1.12125e+10, 1.114942e+10, 
    1.108122e+10, 1.100805e+10, 1.093007e+10, 1.084745e+10, 1.076036e+10, 
    1.066899e+10, 1.057352e+10, 1.047415e+10, 1.037106e+10, 1.026446e+10, 
    1.015454e+10, 1.00415e+10, 9.925557e+09, 9.806899e+09, 9.68573e+09, 
    9.562249e+09, 9.436652e+09, 9.309132e+09, 9.17988e+09, 9.049084e+09, 
    8.916924e+09, 8.78358e+09, 8.649221e+09, 8.514017e+09, 8.378128e+09, 
    8.241709e+09, 8.10491e+09, 7.967875e+09, 7.830739e+09, 7.693634e+09, 
    7.556683e+09, 7.420003e+09, 7.283705e+09, 7.147894e+09, 7.012667e+09, 
    6.878117e+09,
  6.851641e+09, 6.98371e+09, 7.116371e+09, 7.249533e+09, 7.383099e+09, 
    7.516966e+09, 7.651027e+09, 7.785166e+09, 7.919261e+09, 8.053188e+09, 
    8.186811e+09, 8.319992e+09, 8.452588e+09, 8.584445e+09, 8.715411e+09, 
    8.845323e+09, 8.974015e+09, 9.101317e+09, 9.227054e+09, 9.351046e+09, 
    9.473112e+09, 9.593066e+09, 9.710721e+09, 9.825887e+09, 9.938373e+09, 
    1.004799e+10, 1.015454e+10, 1.025783e+10, 1.035769e+10, 1.045391e+10, 
    1.054631e+10, 1.063472e+10, 1.071896e+10, 1.079885e+10, 1.087423e+10, 
    1.094495e+10, 1.101085e+10, 1.107179e+10, 1.112763e+10, 1.117826e+10, 
    1.122356e+10, 1.126342e+10, 1.129776e+10, 1.13265e+10, 1.134958e+10, 
    1.136693e+10, 1.137852e+10, 1.138432e+10, 1.138432e+10, 1.137852e+10, 
    1.136693e+10, 1.134958e+10, 1.13265e+10, 1.129776e+10, 1.126342e+10, 
    1.122356e+10, 1.117826e+10, 1.112763e+10, 1.107179e+10, 1.101085e+10, 
    1.094495e+10, 1.087423e+10, 1.079885e+10, 1.071896e+10, 1.063472e+10, 
    1.054631e+10, 1.045391e+10, 1.035769e+10, 1.025783e+10, 1.015454e+10, 
    1.004799e+10, 9.938373e+09, 9.825887e+09, 9.710721e+09, 9.593066e+09, 
    9.473112e+09, 9.351046e+09, 9.227054e+09, 9.101317e+09, 8.974015e+09, 
    8.845323e+09, 8.715411e+09, 8.584445e+09, 8.452588e+09, 8.319992e+09, 
    8.186811e+09, 8.053188e+09, 7.919261e+09, 7.785166e+09, 7.651027e+09, 
    7.516966e+09, 7.383099e+09, 7.249533e+09, 7.116371e+09, 6.98371e+09, 
    6.851641e+09,
  6.824007e+09, 6.953512e+09, 7.083523e+09, 7.21395e+09, 7.344698e+09, 
    7.475667e+09, 7.606751e+09, 7.737838e+09, 7.868808e+09, 7.99954e+09, 
    8.129904e+09, 8.259766e+09, 8.388985e+09, 8.517416e+09, 8.64491e+09, 
    8.771312e+09, 8.896461e+09, 9.020195e+09, 9.142345e+09, 9.262742e+09, 
    9.381209e+09, 9.497571e+09, 9.61165e+09, 9.723264e+09, 9.832232e+09, 
    9.938373e+09, 1.00415e+10, 1.014144e+10, 1.023802e+10, 1.033104e+10, 
    1.042034e+10, 1.050575e+10, 1.058711e+10, 1.066424e+10, 1.0737e+10, 
    1.080523e+10, 1.08688e+10, 1.092757e+10, 1.098142e+10, 1.103023e+10, 
    1.107389e+10, 1.111231e+10, 1.11454e+10, 1.117309e+10, 1.119532e+10, 
    1.121203e+10, 1.12232e+10, 1.122879e+10, 1.122879e+10, 1.12232e+10, 
    1.121203e+10, 1.119532e+10, 1.117309e+10, 1.11454e+10, 1.111231e+10, 
    1.107389e+10, 1.103023e+10, 1.098142e+10, 1.092757e+10, 1.08688e+10, 
    1.080523e+10, 1.0737e+10, 1.066424e+10, 1.058711e+10, 1.050575e+10, 
    1.042034e+10, 1.033104e+10, 1.023802e+10, 1.014144e+10, 1.00415e+10, 
    9.938373e+09, 9.832232e+09, 9.723264e+09, 9.61165e+09, 9.497571e+09, 
    9.381209e+09, 9.262742e+09, 9.142345e+09, 9.020195e+09, 8.896461e+09, 
    8.771312e+09, 8.64491e+09, 8.517416e+09, 8.388985e+09, 8.259766e+09, 
    8.129904e+09, 7.99954e+09, 7.868808e+09, 7.737838e+09, 7.606751e+09, 
    7.475667e+09, 7.344698e+09, 7.21395e+09, 7.083523e+09, 6.953512e+09, 
    6.824007e+09,
  6.795221e+09, 6.922081e+09, 7.049361e+09, 7.176973e+09, 7.304823e+09, 
    7.432814e+09, 7.56084e+09, 7.688794e+09, 7.816561e+09, 7.94402e+09, 
    8.071048e+09, 8.197513e+09, 8.323282e+09, 8.448214e+09, 8.572165e+09, 
    8.694987e+09, 8.816526e+09, 8.936627e+09, 9.055129e+09, 9.171869e+09, 
    9.286681e+09, 9.399396e+09, 9.509846e+09, 9.61786e+09, 9.723264e+09, 
    9.825887e+09, 9.925557e+09, 1.00221e+10, 1.011536e+10, 1.020515e+10, 
    1.029132e+10, 1.037371e+10, 1.045215e+10, 1.05265e+10, 1.059662e+10, 
    1.066235e+10, 1.072358e+10, 1.078017e+10, 1.0832e+10, 1.087898e+10, 
    1.092099e+10, 1.095795e+10, 1.098979e+10, 1.101642e+10, 1.10378e+10, 
    1.105388e+10, 1.106461e+10, 1.106999e+10, 1.106999e+10, 1.106461e+10, 
    1.105388e+10, 1.10378e+10, 1.101642e+10, 1.098979e+10, 1.095795e+10, 
    1.092099e+10, 1.087898e+10, 1.0832e+10, 1.078017e+10, 1.072358e+10, 
    1.066235e+10, 1.059662e+10, 1.05265e+10, 1.045215e+10, 1.037371e+10, 
    1.029132e+10, 1.020515e+10, 1.011536e+10, 1.00221e+10, 9.925557e+09, 
    9.825887e+09, 9.723264e+09, 9.61786e+09, 9.509846e+09, 9.399396e+09, 
    9.286681e+09, 9.171869e+09, 9.055129e+09, 8.936627e+09, 8.816526e+09, 
    8.694987e+09, 8.572165e+09, 8.448214e+09, 8.323282e+09, 8.197513e+09, 
    8.071048e+09, 7.94402e+09, 7.816561e+09, 7.688794e+09, 7.56084e+09, 
    7.432814e+09, 7.304823e+09, 7.176973e+09, 7.049361e+09, 6.922081e+09, 
    6.795221e+09,
  6.76529e+09, 6.889429e+09, 7.013901e+09, 7.13862e+09, 7.263496e+09, 
    7.388432e+09, 7.513327e+09, 7.638074e+09, 7.762563e+09, 7.886679e+09, 
    8.010299e+09, 8.133301e+09, 8.255552e+09, 8.37692e+09, 8.497266e+09, 
    8.616447e+09, 8.734319e+09, 8.85073e+09, 8.96553e+09, 9.078562e+09, 
    9.18967e+09, 9.298694e+09, 9.405474e+09, 9.509846e+09, 9.61165e+09, 
    9.710721e+09, 9.806899e+09, 9.900023e+09, 9.989933e+09, 1.007647e+10, 
    1.015949e+10, 1.023883e+10, 1.031435e+10, 1.03859e+10, 1.045336e+10, 
    1.051658e+10, 1.057545e+10, 1.062985e+10, 1.067967e+10, 1.07248e+10, 
    1.076517e+10, 1.080067e+10, 1.083124e+10, 1.085682e+10, 1.087735e+10, 
    1.089278e+10, 1.090309e+10, 1.090825e+10, 1.090825e+10, 1.090309e+10, 
    1.089278e+10, 1.087735e+10, 1.085682e+10, 1.083124e+10, 1.080067e+10, 
    1.076517e+10, 1.07248e+10, 1.067967e+10, 1.062985e+10, 1.057545e+10, 
    1.051658e+10, 1.045336e+10, 1.03859e+10, 1.031435e+10, 1.023883e+10, 
    1.015949e+10, 1.007647e+10, 9.989933e+09, 9.900023e+09, 9.806899e+09, 
    9.710721e+09, 9.61165e+09, 9.509846e+09, 9.405474e+09, 9.298694e+09, 
    9.18967e+09, 9.078562e+09, 8.96553e+09, 8.85073e+09, 8.734319e+09, 
    8.616447e+09, 8.497266e+09, 8.37692e+09, 8.255552e+09, 8.133301e+09, 
    8.010299e+09, 7.886679e+09, 7.762563e+09, 7.638074e+09, 7.513327e+09, 
    7.388432e+09, 7.263496e+09, 7.13862e+09, 7.013901e+09, 6.889429e+09, 
    6.76529e+09,
  6.734221e+09, 6.855565e+09, 6.977157e+09, 7.098912e+09, 7.220742e+09, 
    7.342552e+09, 7.464245e+09, 7.585717e+09, 7.706863e+09, 7.827569e+09, 
    7.94772e+09, 8.067195e+09, 8.18587e+09, 8.303616e+09, 8.420301e+09, 
    8.53579e+09, 8.649944e+09, 8.762619e+09, 8.873673e+09, 8.982957e+09, 
    9.090322e+09, 9.195619e+09, 9.298694e+09, 9.399396e+09, 9.497571e+09, 
    9.593066e+09, 9.68573e+09, 9.775411e+09, 9.861961e+09, 9.945231e+09, 
    1.002508e+10, 1.010136e+10, 1.017395e+10, 1.02427e+10, 1.030749e+10, 
    1.03682e+10, 1.042471e+10, 1.047692e+10, 1.052472e+10, 1.056802e+10, 
    1.060673e+10, 1.064077e+10, 1.067009e+10, 1.06946e+10, 1.071428e+10, 
    1.072907e+10, 1.073895e+10, 1.07439e+10, 1.07439e+10, 1.073895e+10, 
    1.072907e+10, 1.071428e+10, 1.06946e+10, 1.067009e+10, 1.064077e+10, 
    1.060673e+10, 1.056802e+10, 1.052472e+10, 1.047692e+10, 1.042471e+10, 
    1.03682e+10, 1.030749e+10, 1.02427e+10, 1.017395e+10, 1.010136e+10, 
    1.002508e+10, 9.945231e+09, 9.861961e+09, 9.775411e+09, 9.68573e+09, 
    9.593066e+09, 9.497571e+09, 9.399396e+09, 9.298694e+09, 9.195619e+09, 
    9.090322e+09, 8.982957e+09, 8.873673e+09, 8.762619e+09, 8.649944e+09, 
    8.53579e+09, 8.420301e+09, 8.303616e+09, 8.18587e+09, 8.067195e+09, 
    7.94772e+09, 7.827569e+09, 7.706863e+09, 7.585717e+09, 7.464245e+09, 
    7.342552e+09, 7.220742e+09, 7.098912e+09, 6.977157e+09, 6.855565e+09, 
    6.734221e+09,
  6.702019e+09, 6.8205e+09, 6.939143e+09, 7.057866e+09, 7.176583e+09, 
    7.295202e+09, 7.41363e+09, 7.531766e+09, 7.649507e+09, 7.766745e+09, 
    7.883369e+09, 7.999264e+09, 8.11431e+09, 8.228386e+09, 8.341364e+09, 
    8.453116e+09, 8.563511e+09, 8.672412e+09, 8.779684e+09, 8.885187e+09, 
    8.988781e+09, 9.090322e+09, 9.18967e+09, 9.286681e+09, 9.381209e+09, 
    9.473112e+09, 9.562249e+09, 9.648477e+09, 9.731658e+09, 9.811654e+09, 
    9.88833e+09, 9.961556e+09, 1.00312e+10, 1.009715e+10, 1.015928e+10, 
    1.021748e+10, 1.027164e+10, 1.032166e+10, 1.036744e+10, 1.040891e+10, 
    1.044597e+10, 1.047856e+10, 1.050662e+10, 1.053008e+10, 1.054891e+10, 
    1.056306e+10, 1.057252e+10, 1.057725e+10, 1.057725e+10, 1.057252e+10, 
    1.056306e+10, 1.054891e+10, 1.053008e+10, 1.050662e+10, 1.047856e+10, 
    1.044597e+10, 1.040891e+10, 1.036744e+10, 1.032166e+10, 1.027164e+10, 
    1.021748e+10, 1.015928e+10, 1.009715e+10, 1.00312e+10, 9.961556e+09, 
    9.88833e+09, 9.811654e+09, 9.731658e+09, 9.648477e+09, 9.562249e+09, 
    9.473112e+09, 9.381209e+09, 9.286681e+09, 9.18967e+09, 9.090322e+09, 
    8.988781e+09, 8.885187e+09, 8.779684e+09, 8.672412e+09, 8.563511e+09, 
    8.453116e+09, 8.341364e+09, 8.228386e+09, 8.11431e+09, 7.999264e+09, 
    7.883369e+09, 7.766745e+09, 7.649507e+09, 7.531766e+09, 7.41363e+09, 
    7.295202e+09, 7.176583e+09, 7.057866e+09, 6.939143e+09, 6.8205e+09, 
    6.702019e+09,
  6.668692e+09, 6.784244e+09, 6.899874e+09, 7.015503e+09, 7.131045e+09, 
    7.246414e+09, 7.361518e+09, 7.47626e+09, 7.590542e+09, 7.704261e+09, 
    7.817309e+09, 7.929576e+09, 8.04095e+09, 8.151313e+09, 8.260545e+09, 
    8.368525e+09, 8.475127e+09, 8.580225e+09, 8.683688e+09, 8.785385e+09, 
    8.885187e+09, 8.982957e+09, 9.078562e+09, 9.171869e+09, 9.262742e+09, 
    9.351046e+09, 9.436652e+09, 9.519426e+09, 9.599237e+09, 9.67596e+09, 
    9.749469e+09, 9.819643e+09, 9.886363e+09, 9.949515e+09, 1.000899e+10, 
    1.006469e+10, 1.01165e+10, 1.016434e+10, 1.020812e+10, 1.024776e+10, 
    1.028319e+10, 1.031433e+10, 1.034114e+10, 1.036355e+10, 1.038154e+10, 
    1.039506e+10, 1.040409e+10, 1.040861e+10, 1.040861e+10, 1.040409e+10, 
    1.039506e+10, 1.038154e+10, 1.036355e+10, 1.034114e+10, 1.031433e+10, 
    1.028319e+10, 1.024776e+10, 1.020812e+10, 1.016434e+10, 1.01165e+10, 
    1.006469e+10, 1.000899e+10, 9.949515e+09, 9.886363e+09, 9.819643e+09, 
    9.749469e+09, 9.67596e+09, 9.599237e+09, 9.519426e+09, 9.436652e+09, 
    9.351046e+09, 9.262742e+09, 9.171869e+09, 9.078562e+09, 8.982957e+09, 
    8.885187e+09, 8.785385e+09, 8.683688e+09, 8.580225e+09, 8.475127e+09, 
    8.368525e+09, 8.260545e+09, 8.151313e+09, 8.04095e+09, 7.929576e+09, 
    7.817309e+09, 7.704261e+09, 7.590542e+09, 7.47626e+09, 7.361518e+09, 
    7.246414e+09, 7.131045e+09, 7.015503e+09, 6.899874e+09, 6.784244e+09, 
    6.668692e+09,
  6.634248e+09, 6.74681e+09, 6.859367e+09, 6.971842e+09, 7.084154e+09, 
    7.196217e+09, 7.307944e+09, 7.419243e+09, 7.530018e+09, 7.640172e+09, 
    7.749601e+09, 7.858201e+09, 7.965864e+09, 8.072481e+09, 8.177936e+09, 
    8.282116e+09, 8.384902e+09, 8.486173e+09, 8.585809e+09, 8.683688e+09, 
    8.779684e+09, 8.873673e+09, 8.96553e+09, 9.055129e+09, 9.142345e+09, 
    9.227054e+09, 9.309132e+09, 9.388457e+09, 9.464909e+09, 9.53837e+09, 
    9.608722e+09, 9.675857e+09, 9.739662e+09, 9.800034e+09, 9.856871e+09, 
    9.910078e+09, 9.959563e+09, 1.000524e+10, 1.004703e+10, 1.008486e+10, 
    1.011866e+10, 1.014837e+10, 1.017394e+10, 1.019532e+10, 1.021247e+10, 
    1.022536e+10, 1.023397e+10, 1.023827e+10, 1.023827e+10, 1.023397e+10, 
    1.022536e+10, 1.021247e+10, 1.019532e+10, 1.017394e+10, 1.014837e+10, 
    1.011866e+10, 1.008486e+10, 1.004703e+10, 1.000524e+10, 9.959563e+09, 
    9.910078e+09, 9.856871e+09, 9.800034e+09, 9.739662e+09, 9.675857e+09, 
    9.608722e+09, 9.53837e+09, 9.464909e+09, 9.388457e+09, 9.309132e+09, 
    9.227054e+09, 9.142345e+09, 9.055129e+09, 8.96553e+09, 8.873673e+09, 
    8.779684e+09, 8.683688e+09, 8.585809e+09, 8.486173e+09, 8.384902e+09, 
    8.282116e+09, 8.177936e+09, 8.072481e+09, 7.965864e+09, 7.858201e+09, 
    7.749601e+09, 7.640172e+09, 7.530018e+09, 7.419243e+09, 7.307944e+09, 
    7.196217e+09, 7.084154e+09, 6.971842e+09, 6.859367e+09, 6.74681e+09, 
    6.634248e+09,
  6.598693e+09, 6.708208e+09, 6.817636e+09, 6.926904e+09, 7.035934e+09, 
    7.144643e+09, 7.252946e+09, 7.360757e+09, 7.467984e+09, 7.574533e+09, 
    7.680307e+09, 7.785207e+09, 7.889131e+09, 7.991974e+09, 8.093629e+09, 
    8.193989e+09, 8.292941e+09, 8.390374e+09, 8.486173e+09, 8.580225e+09, 
    8.672412e+09, 8.762619e+09, 8.85073e+09, 8.936627e+09, 9.020195e+09, 
    9.101317e+09, 9.17988e+09, 9.255772e+09, 9.32888e+09, 9.399095e+09, 
    9.466312e+09, 9.530426e+09, 9.591338e+09, 9.64895e+09, 9.703171e+09, 
    9.753911e+09, 9.801088e+09, 9.844622e+09, 9.884442e+09, 9.920478e+09, 
    9.95267e+09, 9.980962e+09, 1.00053e+10, 1.002566e+10, 1.004198e+10, 
    1.005425e+10, 1.006244e+10, 1.006654e+10, 1.006654e+10, 1.006244e+10, 
    1.005425e+10, 1.004198e+10, 1.002566e+10, 1.00053e+10, 9.980962e+09, 
    9.95267e+09, 9.920478e+09, 9.884442e+09, 9.844622e+09, 9.801088e+09, 
    9.753911e+09, 9.703171e+09, 9.64895e+09, 9.591338e+09, 9.530426e+09, 
    9.466312e+09, 9.399095e+09, 9.32888e+09, 9.255772e+09, 9.17988e+09, 
    9.101317e+09, 9.020195e+09, 8.936627e+09, 8.85073e+09, 8.762619e+09, 
    8.672412e+09, 8.580225e+09, 8.486173e+09, 8.390374e+09, 8.292941e+09, 
    8.193989e+09, 8.093629e+09, 7.991974e+09, 7.889131e+09, 7.785207e+09, 
    7.680307e+09, 7.574533e+09, 7.467984e+09, 7.360757e+09, 7.252946e+09, 
    7.144643e+09, 7.035934e+09, 6.926904e+09, 6.817636e+09, 6.708208e+09, 
    6.598693e+09,
  6.562035e+09, 6.668449e+09, 6.774699e+09, 6.880711e+09, 6.986412e+09, 
    7.091722e+09, 7.196561e+09, 7.300845e+09, 7.404488e+09, 7.5074e+09, 
    7.60949e+09, 7.710664e+09, 7.810825e+09, 7.909876e+09, 8.007716e+09, 
    8.104243e+09, 8.199353e+09, 8.292941e+09, 8.384902e+09, 8.475127e+09, 
    8.563511e+09, 8.649944e+09, 8.734319e+09, 8.816526e+09, 8.896461e+09, 
    8.974015e+09, 9.049084e+09, 9.121564e+09, 9.191351e+09, 9.258346e+09, 
    9.322452e+09, 9.383574e+09, 9.441618e+09, 9.496498e+09, 9.548129e+09, 
    9.596429e+09, 9.641325e+09, 9.68274e+09, 9.720613e+09, 9.754878e+09, 
    9.785482e+09, 9.812372e+09, 9.835507e+09, 9.854844e+09, 9.870353e+09, 
    9.882009e+09, 9.88979e+09, 9.893683e+09, 9.893683e+09, 9.88979e+09, 
    9.882009e+09, 9.870353e+09, 9.854844e+09, 9.835507e+09, 9.812372e+09, 
    9.785482e+09, 9.754878e+09, 9.720613e+09, 9.68274e+09, 9.641325e+09, 
    9.596429e+09, 9.548129e+09, 9.496498e+09, 9.441618e+09, 9.383574e+09, 
    9.322452e+09, 9.258346e+09, 9.191351e+09, 9.121564e+09, 9.049084e+09, 
    8.974015e+09, 8.896461e+09, 8.816526e+09, 8.734319e+09, 8.649944e+09, 
    8.563511e+09, 8.475127e+09, 8.384902e+09, 8.292941e+09, 8.199353e+09, 
    8.104243e+09, 8.007716e+09, 7.909876e+09, 7.810825e+09, 7.710664e+09, 
    7.60949e+09, 7.5074e+09, 7.404488e+09, 7.300845e+09, 7.196561e+09, 
    7.091722e+09, 6.986412e+09, 6.880711e+09, 6.774699e+09, 6.668449e+09, 
    6.562035e+09,
  6.524282e+09, 6.627547e+09, 6.730571e+09, 6.833284e+09, 6.935614e+09, 
    7.037487e+09, 7.138825e+09, 7.23955e+09, 7.339579e+09, 7.438829e+09, 
    7.537212e+09, 7.634641e+09, 7.731025e+09, 7.826271e+09, 7.920287e+09, 
    8.012976e+09, 8.104243e+09, 8.193989e+09, 8.282116e+09, 8.368525e+09, 
    8.453116e+09, 8.53579e+09, 8.616447e+09, 8.694987e+09, 8.771312e+09, 
    8.845323e+09, 8.916924e+09, 8.986021e+09, 9.052518e+09, 9.116325e+09, 
    9.177352e+09, 9.235513e+09, 9.290724e+09, 9.342905e+09, 9.391978e+09, 
    9.437871e+09, 9.480515e+09, 9.519842e+09, 9.555794e+09, 9.588315e+09, 
    9.617354e+09, 9.642865e+09, 9.664807e+09, 9.683147e+09, 9.697854e+09, 
    9.708905e+09, 9.716282e+09, 9.719975e+09, 9.719975e+09, 9.716282e+09, 
    9.708905e+09, 9.697854e+09, 9.683147e+09, 9.664807e+09, 9.642865e+09, 
    9.617354e+09, 9.588315e+09, 9.555794e+09, 9.519842e+09, 9.480515e+09, 
    9.437871e+09, 9.391978e+09, 9.342905e+09, 9.290724e+09, 9.235513e+09, 
    9.177352e+09, 9.116325e+09, 9.052518e+09, 8.986021e+09, 8.916924e+09, 
    8.845323e+09, 8.771312e+09, 8.694987e+09, 8.616447e+09, 8.53579e+09, 
    8.453116e+09, 8.368525e+09, 8.282116e+09, 8.193989e+09, 8.104243e+09, 
    8.012976e+09, 7.920287e+09, 7.826271e+09, 7.731025e+09, 7.634641e+09, 
    7.537212e+09, 7.438829e+09, 7.339579e+09, 7.23955e+09, 7.138825e+09, 
    7.037487e+09, 6.935614e+09, 6.833284e+09, 6.730571e+09, 6.627547e+09, 
    6.524282e+09,
  6.485442e+09, 6.585513e+09, 6.685269e+09, 6.784643e+09, 6.883567e+09, 
    6.981969e+09, 7.079777e+09, 7.176916e+09, 7.273309e+09, 7.368877e+09, 
    7.463537e+09, 7.557208e+09, 7.649805e+09, 7.741242e+09, 7.831433e+09, 
    7.920287e+09, 8.007716e+09, 8.093629e+09, 8.177936e+09, 8.260545e+09, 
    8.341364e+09, 8.420301e+09, 8.497266e+09, 8.572165e+09, 8.64491e+09, 
    8.715411e+09, 8.78358e+09, 8.849328e+09, 8.912572e+09, 8.973229e+09, 
    9.031216e+09, 9.086456e+09, 9.138871e+09, 9.188391e+09, 9.234944e+09, 
    9.278465e+09, 9.318892e+09, 9.356163e+09, 9.390226e+09, 9.421031e+09, 
    9.448532e+09, 9.472687e+09, 9.49346e+09, 9.510819e+09, 9.524738e+09, 
    9.535196e+09, 9.542177e+09, 9.54567e+09, 9.54567e+09, 9.542177e+09, 
    9.535196e+09, 9.524738e+09, 9.510819e+09, 9.49346e+09, 9.472687e+09, 
    9.448532e+09, 9.421031e+09, 9.390226e+09, 9.356163e+09, 9.318892e+09, 
    9.278465e+09, 9.234944e+09, 9.188391e+09, 9.138871e+09, 9.086456e+09, 
    9.031216e+09, 8.973229e+09, 8.912572e+09, 8.849328e+09, 8.78358e+09, 
    8.715411e+09, 8.64491e+09, 8.572165e+09, 8.497266e+09, 8.420301e+09, 
    8.341364e+09, 8.260545e+09, 8.177936e+09, 8.093629e+09, 8.007716e+09, 
    7.920287e+09, 7.831433e+09, 7.741242e+09, 7.649805e+09, 7.557208e+09, 
    7.463537e+09, 7.368877e+09, 7.273309e+09, 7.176916e+09, 7.079777e+09, 
    6.981969e+09, 6.883567e+09, 6.784643e+09, 6.685269e+09, 6.585513e+09, 
    6.485442e+09,
  6.445522e+09, 6.54236e+09, 6.638811e+09, 6.734811e+09, 6.830297e+09, 
    6.925201e+09, 7.019455e+09, 7.112987e+09, 7.205726e+09, 7.297597e+09, 
    7.388526e+09, 7.478433e+09, 7.567242e+09, 7.654872e+09, 7.741242e+09, 
    7.826271e+09, 7.909876e+09, 7.991974e+09, 8.072481e+09, 8.151313e+09, 
    8.228386e+09, 8.303616e+09, 8.37692e+09, 8.448214e+09, 8.517416e+09, 
    8.584445e+09, 8.649221e+09, 8.711665e+09, 8.771699e+09, 8.829247e+09, 
    8.884238e+09, 8.936601e+09, 8.986266e+09, 9.033167e+09, 9.077242e+09, 
    9.118431e+09, 9.156679e+09, 9.191932e+09, 9.224142e+09, 9.253263e+09, 
    9.279254e+09, 9.302078e+09, 9.321703e+09, 9.338102e+09, 9.351248e+09, 
    9.361125e+09, 9.367718e+09, 9.371016e+09, 9.371016e+09, 9.367718e+09, 
    9.361125e+09, 9.351248e+09, 9.338102e+09, 9.321703e+09, 9.302078e+09, 
    9.279254e+09, 9.253263e+09, 9.224142e+09, 9.191932e+09, 9.156679e+09, 
    9.118431e+09, 9.077242e+09, 9.033167e+09, 8.986266e+09, 8.936601e+09, 
    8.884238e+09, 8.829247e+09, 8.771699e+09, 8.711665e+09, 8.649221e+09, 
    8.584445e+09, 8.517416e+09, 8.448214e+09, 8.37692e+09, 8.303616e+09, 
    8.228386e+09, 8.151313e+09, 8.072481e+09, 7.991974e+09, 7.909876e+09, 
    7.826271e+09, 7.741242e+09, 7.654872e+09, 7.567242e+09, 7.478433e+09, 
    7.388526e+09, 7.297597e+09, 7.205726e+09, 7.112987e+09, 7.019455e+09, 
    6.925201e+09, 6.830297e+09, 6.734811e+09, 6.638811e+09, 6.54236e+09, 
    6.445522e+09,
  6.404531e+09, 6.4981e+09, 6.591213e+09, 6.683811e+09, 6.775833e+09, 
    6.867216e+09, 6.957896e+09, 7.047806e+09, 7.136881e+09, 7.225049e+09, 
    7.312241e+09, 7.398386e+09, 7.483411e+09, 7.567242e+09, 7.649805e+09, 
    7.731025e+09, 7.810825e+09, 7.889131e+09, 7.965864e+09, 8.04095e+09, 
    8.11431e+09, 8.18587e+09, 8.255552e+09, 8.323282e+09, 8.388985e+09, 
    8.452588e+09, 8.514017e+09, 8.573202e+09, 8.630074e+09, 8.684566e+09, 
    8.736609e+09, 8.786142e+09, 8.833104e+09, 8.877434e+09, 8.919077e+09, 
    8.95798e+09, 8.994092e+09, 9.027367e+09, 9.05776e+09, 9.085231e+09, 
    9.109745e+09, 9.131267e+09, 9.14977e+09, 9.165227e+09, 9.177618e+09, 
    9.186927e+09, 9.193139e+09, 9.196247e+09, 9.196247e+09, 9.193139e+09, 
    9.186927e+09, 9.177618e+09, 9.165227e+09, 9.14977e+09, 9.131267e+09, 
    9.109745e+09, 9.085231e+09, 9.05776e+09, 9.027367e+09, 8.994092e+09, 
    8.95798e+09, 8.919077e+09, 8.877434e+09, 8.833104e+09, 8.786142e+09, 
    8.736609e+09, 8.684566e+09, 8.630074e+09, 8.573202e+09, 8.514017e+09, 
    8.452588e+09, 8.388985e+09, 8.323282e+09, 8.255552e+09, 8.18587e+09, 
    8.11431e+09, 8.04095e+09, 7.965864e+09, 7.889131e+09, 7.810825e+09, 
    7.731025e+09, 7.649805e+09, 7.567242e+09, 7.483411e+09, 7.398386e+09, 
    7.312241e+09, 7.225049e+09, 7.136881e+09, 7.047806e+09, 6.957896e+09, 
    6.867216e+09, 6.775833e+09, 6.683811e+09, 6.591213e+09, 6.4981e+09, 
    6.404531e+09,
  6.362479e+09, 6.452746e+09, 6.542493e+09, 6.631664e+09, 6.720201e+09, 
    6.808046e+09, 6.895139e+09, 6.981418e+09, 7.066822e+09, 7.151286e+09, 
    7.234745e+09, 7.317134e+09, 7.398386e+09, 7.478433e+09, 7.557208e+09, 
    7.634641e+09, 7.710664e+09, 7.785207e+09, 7.858201e+09, 7.929576e+09, 
    7.999264e+09, 8.067195e+09, 8.133301e+09, 8.197513e+09, 8.259766e+09, 
    8.319992e+09, 8.378128e+09, 8.434108e+09, 8.487873e+09, 8.539359e+09, 
    8.58851e+09, 8.635267e+09, 8.679578e+09, 8.721389e+09, 8.760649e+09, 
    8.797313e+09, 8.831335e+09, 8.862674e+09, 8.891291e+09, 8.917151e+09, 
    8.940219e+09, 8.96047e+09, 8.977876e+09, 8.992415e+09, 9.004068e+09, 
    9.012821e+09, 9.018663e+09, 9.021585e+09, 9.021585e+09, 9.018663e+09, 
    9.012821e+09, 9.004068e+09, 8.992415e+09, 8.977876e+09, 8.96047e+09, 
    8.940219e+09, 8.917151e+09, 8.891291e+09, 8.862674e+09, 8.831335e+09, 
    8.797313e+09, 8.760649e+09, 8.721389e+09, 8.679578e+09, 8.635267e+09, 
    8.58851e+09, 8.539359e+09, 8.487873e+09, 8.434108e+09, 8.378128e+09, 
    8.319992e+09, 8.259766e+09, 8.197513e+09, 8.133301e+09, 8.067195e+09, 
    7.999264e+09, 7.929576e+09, 7.858201e+09, 7.785207e+09, 7.710664e+09, 
    7.634641e+09, 7.557208e+09, 7.478433e+09, 7.398386e+09, 7.317134e+09, 
    7.234745e+09, 7.151286e+09, 7.066822e+09, 6.981418e+09, 6.895139e+09, 
    6.808046e+09, 6.720201e+09, 6.631664e+09, 6.542493e+09, 6.452746e+09, 
    6.362479e+09,
  6.319373e+09, 6.406312e+09, 6.492669e+09, 6.578392e+09, 6.663429e+09, 
    6.747724e+09, 6.831222e+09, 6.913867e+09, 6.9956e+09, 7.076365e+09, 
    7.1561e+09, 7.234745e+09, 7.312241e+09, 7.388526e+09, 7.463537e+09, 
    7.537212e+09, 7.60949e+09, 7.680307e+09, 7.749601e+09, 7.817309e+09, 
    7.883369e+09, 7.94772e+09, 8.010299e+09, 8.071048e+09, 8.129904e+09, 
    8.186811e+09, 8.241709e+09, 8.294543e+09, 8.345257e+09, 8.393798e+09, 
    8.440113e+09, 8.484152e+09, 8.525868e+09, 8.565214e+09, 8.602145e+09, 
    8.636621e+09, 8.668601e+09, 8.698051e+09, 8.724934e+09, 8.749221e+09, 
    8.770882e+09, 8.789891e+09, 8.806228e+09, 8.819871e+09, 8.830806e+09, 
    8.839017e+09, 8.844498e+09, 8.84724e+09, 8.84724e+09, 8.844498e+09, 
    8.839017e+09, 8.830806e+09, 8.819871e+09, 8.806228e+09, 8.789891e+09, 
    8.770882e+09, 8.749221e+09, 8.724934e+09, 8.698051e+09, 8.668601e+09, 
    8.636621e+09, 8.602145e+09, 8.565214e+09, 8.525868e+09, 8.484152e+09, 
    8.440113e+09, 8.393798e+09, 8.345257e+09, 8.294543e+09, 8.241709e+09, 
    8.186811e+09, 8.129904e+09, 8.071048e+09, 8.010299e+09, 7.94772e+09, 
    7.883369e+09, 7.817309e+09, 7.749601e+09, 7.680307e+09, 7.60949e+09, 
    7.537212e+09, 7.463537e+09, 7.388526e+09, 7.312241e+09, 7.234745e+09, 
    7.1561e+09, 7.076365e+09, 6.9956e+09, 6.913867e+09, 6.831222e+09, 
    6.747724e+09, 6.663429e+09, 6.578392e+09, 6.492669e+09, 6.406312e+09, 
    6.319373e+09,
  6.275223e+09, 6.35881e+09, 6.441759e+09, 6.52402e+09, 6.605544e+09, 
    6.686283e+09, 6.766183e+09, 6.845195e+09, 6.923265e+09, 7.000339e+09, 
    7.076365e+09, 7.151286e+09, 7.225049e+09, 7.297597e+09, 7.368877e+09, 
    7.438829e+09, 7.5074e+09, 7.574533e+09, 7.640172e+09, 7.704261e+09, 
    7.766745e+09, 7.827569e+09, 7.886679e+09, 7.94402e+09, 7.99954e+09, 
    8.053188e+09, 8.10491e+09, 8.15466e+09, 8.202386e+09, 8.248043e+09, 
    8.291585e+09, 8.332967e+09, 8.372148e+09, 8.409087e+09, 8.443745e+09, 
    8.476086e+09, 8.506077e+09, 8.533684e+09, 8.558878e+09, 8.581632e+09, 
    8.601922e+09, 8.619724e+09, 8.63502e+09, 8.647793e+09, 8.658028e+09, 
    8.665715e+09, 8.670843e+09, 8.673409e+09, 8.673409e+09, 8.670843e+09, 
    8.665715e+09, 8.658028e+09, 8.647793e+09, 8.63502e+09, 8.619724e+09, 
    8.601922e+09, 8.581632e+09, 8.558878e+09, 8.533684e+09, 8.506077e+09, 
    8.476086e+09, 8.443745e+09, 8.409087e+09, 8.372148e+09, 8.332967e+09, 
    8.291585e+09, 8.248043e+09, 8.202386e+09, 8.15466e+09, 8.10491e+09, 
    8.053188e+09, 7.99954e+09, 7.94402e+09, 7.886679e+09, 7.827569e+09, 
    7.766745e+09, 7.704261e+09, 7.640172e+09, 7.574533e+09, 7.5074e+09, 
    7.438829e+09, 7.368877e+09, 7.297597e+09, 7.225049e+09, 7.151286e+09, 
    7.076365e+09, 7.000339e+09, 6.923265e+09, 6.845195e+09, 6.766183e+09, 
    6.686283e+09, 6.605544e+09, 6.52402e+09, 6.441759e+09, 6.35881e+09, 
    6.275223e+09,
  6.230037e+09, 6.310255e+09, 6.38978e+09, 6.468569e+09, 6.546576e+09, 
    6.623755e+09, 6.700061e+09, 6.775447e+09, 6.849864e+09, 6.923265e+09, 
    6.9956e+09, 7.066822e+09, 7.136881e+09, 7.205726e+09, 7.273309e+09, 
    7.339579e+09, 7.404488e+09, 7.467984e+09, 7.530018e+09, 7.590542e+09, 
    7.649507e+09, 7.706863e+09, 7.762563e+09, 7.816561e+09, 7.868808e+09, 
    7.919261e+09, 7.967875e+09, 8.014606e+09, 8.059411e+09, 8.10225e+09, 
    8.143084e+09, 8.181873e+09, 8.218582e+09, 8.253174e+09, 8.285618e+09, 
    8.31588e+09, 8.343933e+09, 8.369748e+09, 8.3933e+09, 8.414565e+09, 
    8.433522e+09, 8.450151e+09, 8.464436e+09, 8.476363e+09, 8.485919e+09, 
    8.493095e+09, 8.497883e+09, 8.500278e+09, 8.500278e+09, 8.497883e+09, 
    8.493095e+09, 8.485919e+09, 8.476363e+09, 8.464436e+09, 8.450151e+09, 
    8.433522e+09, 8.414565e+09, 8.3933e+09, 8.369748e+09, 8.343933e+09, 
    8.31588e+09, 8.285618e+09, 8.253174e+09, 8.218582e+09, 8.181873e+09, 
    8.143084e+09, 8.10225e+09, 8.059411e+09, 8.014606e+09, 7.967875e+09, 
    7.919261e+09, 7.868808e+09, 7.816561e+09, 7.762563e+09, 7.706863e+09, 
    7.649507e+09, 7.590542e+09, 7.530018e+09, 7.467984e+09, 7.404488e+09, 
    7.339579e+09, 7.273309e+09, 7.205726e+09, 7.136881e+09, 7.066822e+09, 
    6.9956e+09, 6.923265e+09, 6.849864e+09, 6.775447e+09, 6.700061e+09, 
    6.623755e+09, 6.546576e+09, 6.468569e+09, 6.38978e+09, 6.310255e+09, 
    6.230037e+09,
  6.183825e+09, 6.260659e+09, 6.336752e+09, 6.412062e+09, 6.486551e+09, 
    6.560175e+09, 6.632894e+09, 6.704666e+09, 6.775447e+09, 6.845195e+09, 
    6.913867e+09, 6.981418e+09, 7.047806e+09, 7.112987e+09, 7.176916e+09, 
    7.23955e+09, 7.300845e+09, 7.360757e+09, 7.419243e+09, 7.47626e+09, 
    7.531766e+09, 7.585717e+09, 7.638074e+09, 7.688794e+09, 7.737838e+09, 
    7.785166e+09, 7.830739e+09, 7.874522e+09, 7.916475e+09, 7.956566e+09, 
    7.994759e+09, 8.031022e+09, 8.065324e+09, 8.097633e+09, 8.127923e+09, 
    8.156166e+09, 8.182336e+09, 8.20641e+09, 8.228367e+09, 8.248187e+09, 
    8.26585e+09, 8.281342e+09, 8.294647e+09, 8.305754e+09, 8.314652e+09, 
    8.321333e+09, 8.32579e+09, 8.32802e+09, 8.32802e+09, 8.32579e+09, 
    8.321333e+09, 8.314652e+09, 8.305754e+09, 8.294647e+09, 8.281342e+09, 
    8.26585e+09, 8.248187e+09, 8.228367e+09, 8.20641e+09, 8.182336e+09, 
    8.156166e+09, 8.127923e+09, 8.097633e+09, 8.065324e+09, 8.031022e+09, 
    7.994759e+09, 7.956566e+09, 7.916475e+09, 7.874522e+09, 7.830739e+09, 
    7.785166e+09, 7.737838e+09, 7.688794e+09, 7.638074e+09, 7.585717e+09, 
    7.531766e+09, 7.47626e+09, 7.419243e+09, 7.360757e+09, 7.300845e+09, 
    7.23955e+09, 7.176916e+09, 7.112987e+09, 7.047806e+09, 6.981418e+09, 
    6.913867e+09, 6.845195e+09, 6.775447e+09, 6.704666e+09, 6.632894e+09, 
    6.560175e+09, 6.486551e+09, 6.412062e+09, 6.336752e+09, 6.260659e+09, 
    6.183825e+09,
  6.136596e+09, 6.210038e+09, 6.282692e+09, 6.354524e+09, 6.425497e+09, 
    6.495574e+09, 6.564719e+09, 6.632894e+09, 6.700061e+09, 6.766183e+09, 
    6.831222e+09, 6.895139e+09, 6.957896e+09, 7.019455e+09, 7.079777e+09, 
    7.138825e+09, 7.196561e+09, 7.252946e+09, 7.307944e+09, 7.361518e+09, 
    7.41363e+09, 7.464245e+09, 7.513327e+09, 7.56084e+09, 7.606751e+09, 
    7.651027e+09, 7.693634e+09, 7.734541e+09, 7.773715e+09, 7.811129e+09, 
    7.846753e+09, 7.880559e+09, 7.912521e+09, 7.942612e+09, 7.970811e+09, 
    7.997093e+09, 8.021437e+09, 8.043825e+09, 8.064236e+09, 8.082655e+09, 
    8.099066e+09, 8.113456e+09, 8.125813e+09, 8.136126e+09, 8.144387e+09, 
    8.150589e+09, 8.154726e+09, 8.156796e+09, 8.156796e+09, 8.154726e+09, 
    8.150589e+09, 8.144387e+09, 8.136126e+09, 8.125813e+09, 8.113456e+09, 
    8.099066e+09, 8.082655e+09, 8.064236e+09, 8.043825e+09, 8.021437e+09, 
    7.997093e+09, 7.970811e+09, 7.942612e+09, 7.912521e+09, 7.880559e+09, 
    7.846753e+09, 7.811129e+09, 7.773715e+09, 7.734541e+09, 7.693634e+09, 
    7.651027e+09, 7.606751e+09, 7.56084e+09, 7.513327e+09, 7.464245e+09, 
    7.41363e+09, 7.361518e+09, 7.307944e+09, 7.252946e+09, 7.196561e+09, 
    7.138825e+09, 7.079777e+09, 7.019455e+09, 6.957896e+09, 6.895139e+09, 
    6.831222e+09, 6.766183e+09, 6.700061e+09, 6.632894e+09, 6.564719e+09, 
    6.495574e+09, 6.425497e+09, 6.354524e+09, 6.282692e+09, 6.210038e+09, 
    6.136596e+09,
  6.088361e+09, 6.158404e+09, 6.227619e+09, 6.295976e+09, 6.363442e+09, 
    6.429985e+09, 6.495574e+09, 6.560175e+09, 6.623755e+09, 6.686283e+09, 
    6.747724e+09, 6.808046e+09, 6.867216e+09, 6.925201e+09, 6.981969e+09, 
    7.037487e+09, 7.091722e+09, 7.144643e+09, 7.196217e+09, 7.246414e+09, 
    7.295202e+09, 7.342552e+09, 7.388432e+09, 7.432814e+09, 7.475667e+09, 
    7.516966e+09, 7.556683e+09, 7.594789e+09, 7.631261e+09, 7.666072e+09, 
    7.699199e+09, 7.73062e+09, 7.760311e+09, 7.788252e+09, 7.814423e+09, 
    7.838806e+09, 7.861382e+09, 7.882135e+09, 7.901051e+09, 7.918115e+09, 
    7.933316e+09, 7.946641e+09, 7.958081e+09, 7.967627e+09, 7.975273e+09, 
    7.981012e+09, 7.984841e+09, 7.986756e+09, 7.986756e+09, 7.984841e+09, 
    7.981012e+09, 7.975273e+09, 7.967627e+09, 7.958081e+09, 7.946641e+09, 
    7.933316e+09, 7.918115e+09, 7.901051e+09, 7.882135e+09, 7.861382e+09, 
    7.838806e+09, 7.814423e+09, 7.788252e+09, 7.760311e+09, 7.73062e+09, 
    7.699199e+09, 7.666072e+09, 7.631261e+09, 7.594789e+09, 7.556683e+09, 
    7.516966e+09, 7.475667e+09, 7.432814e+09, 7.388432e+09, 7.342552e+09, 
    7.295202e+09, 7.246414e+09, 7.196217e+09, 7.144643e+09, 7.091722e+09, 
    7.037487e+09, 6.981969e+09, 6.925201e+09, 6.867216e+09, 6.808046e+09, 
    6.747724e+09, 6.686283e+09, 6.623755e+09, 6.560175e+09, 6.495574e+09, 
    6.429985e+09, 6.363442e+09, 6.295976e+09, 6.227619e+09, 6.158404e+09, 
    6.088361e+09,
  6.039129e+09, 6.105772e+09, 6.171552e+09, 6.236442e+09, 6.300414e+09, 
    6.363442e+09, 6.425497e+09, 6.486551e+09, 6.546576e+09, 6.605544e+09, 
    6.663429e+09, 6.720201e+09, 6.775833e+09, 6.830297e+09, 6.883567e+09, 
    6.935614e+09, 6.986412e+09, 7.035934e+09, 7.084154e+09, 7.131045e+09, 
    7.176583e+09, 7.220742e+09, 7.263496e+09, 7.304823e+09, 7.344698e+09, 
    7.383099e+09, 7.420003e+09, 7.455388e+09, 7.489233e+09, 7.521518e+09, 
    7.552224e+09, 7.581331e+09, 7.608822e+09, 7.634681e+09, 7.65889e+09, 
    7.681435e+09, 7.702302e+09, 7.721477e+09, 7.738948e+09, 7.754704e+09, 
    7.768736e+09, 7.781033e+09, 7.791588e+09, 7.800395e+09, 7.807448e+09, 
    7.812741e+09, 7.816271e+09, 7.818037e+09, 7.818037e+09, 7.816271e+09, 
    7.812741e+09, 7.807448e+09, 7.800395e+09, 7.791588e+09, 7.781033e+09, 
    7.768736e+09, 7.754704e+09, 7.738948e+09, 7.721477e+09, 7.702302e+09, 
    7.681435e+09, 7.65889e+09, 7.634681e+09, 7.608822e+09, 7.581331e+09, 
    7.552224e+09, 7.521518e+09, 7.489233e+09, 7.455388e+09, 7.420003e+09, 
    7.383099e+09, 7.344698e+09, 7.304823e+09, 7.263496e+09, 7.220742e+09, 
    7.176583e+09, 7.131045e+09, 7.084154e+09, 7.035934e+09, 6.986412e+09, 
    6.935614e+09, 6.883567e+09, 6.830297e+09, 6.775833e+09, 6.720201e+09, 
    6.663429e+09, 6.605544e+09, 6.546576e+09, 6.486551e+09, 6.425497e+09, 
    6.363442e+09, 6.300414e+09, 6.236442e+09, 6.171552e+09, 6.105772e+09, 
    6.039129e+09,
  5.988909e+09, 6.052155e+09, 6.114508e+09, 6.175945e+09, 6.236442e+09, 
    6.295976e+09, 6.354524e+09, 6.412062e+09, 6.468569e+09, 6.52402e+09, 
    6.578392e+09, 6.631664e+09, 6.683811e+09, 6.734811e+09, 6.784643e+09, 
    6.833284e+09, 6.880711e+09, 6.926904e+09, 6.971842e+09, 7.015503e+09, 
    7.057866e+09, 7.098912e+09, 7.13862e+09, 7.176973e+09, 7.21395e+09, 
    7.249533e+09, 7.283705e+09, 7.316448e+09, 7.347746e+09, 7.377583e+09, 
    7.405943e+09, 7.432813e+09, 7.458176e+09, 7.482021e+09, 7.504335e+09, 
    7.525106e+09, 7.544322e+09, 7.561974e+09, 7.578052e+09, 7.592547e+09, 
    7.605452e+09, 7.616759e+09, 7.626462e+09, 7.634556e+09, 7.641037e+09, 
    7.645901e+09, 7.649145e+09, 7.650767e+09, 7.650767e+09, 7.649145e+09, 
    7.645901e+09, 7.641037e+09, 7.634556e+09, 7.626462e+09, 7.616759e+09, 
    7.605452e+09, 7.592547e+09, 7.578052e+09, 7.561974e+09, 7.544322e+09, 
    7.525106e+09, 7.504335e+09, 7.482021e+09, 7.458176e+09, 7.432813e+09, 
    7.405943e+09, 7.377583e+09, 7.347746e+09, 7.316448e+09, 7.283705e+09, 
    7.249533e+09, 7.21395e+09, 7.176973e+09, 7.13862e+09, 7.098912e+09, 
    7.057866e+09, 7.015503e+09, 6.971842e+09, 6.926904e+09, 6.880711e+09, 
    6.833284e+09, 6.784643e+09, 6.734811e+09, 6.683811e+09, 6.631664e+09, 
    6.578392e+09, 6.52402e+09, 6.468569e+09, 6.412062e+09, 6.354524e+09, 
    6.295976e+09, 6.236442e+09, 6.175945e+09, 6.114508e+09, 6.052155e+09, 
    5.988909e+09,
  5.937712e+09, 5.99757e+09, 6.056508e+09, 6.114508e+09, 6.171552e+09, 
    6.227619e+09, 6.282692e+09, 6.336752e+09, 6.38978e+09, 6.441759e+09, 
    6.492669e+09, 6.542493e+09, 6.591213e+09, 6.638811e+09, 6.685269e+09, 
    6.730571e+09, 6.774699e+09, 6.817636e+09, 6.859367e+09, 6.899874e+09, 
    6.939143e+09, 6.977157e+09, 7.013901e+09, 7.049361e+09, 7.083523e+09, 
    7.116371e+09, 7.147894e+09, 7.178077e+09, 7.206909e+09, 7.234377e+09, 
    7.260469e+09, 7.285175e+09, 7.308484e+09, 7.330385e+09, 7.350871e+09, 
    7.36993e+09, 7.387556e+09, 7.403741e+09, 7.418477e+09, 7.431758e+09, 
    7.443579e+09, 7.453934e+09, 7.462817e+09, 7.470226e+09, 7.476158e+09, 
    7.480609e+09, 7.483577e+09, 7.485062e+09, 7.485062e+09, 7.483577e+09, 
    7.480609e+09, 7.476158e+09, 7.470226e+09, 7.462817e+09, 7.453934e+09, 
    7.443579e+09, 7.431758e+09, 7.418477e+09, 7.403741e+09, 7.387556e+09, 
    7.36993e+09, 7.350871e+09, 7.330385e+09, 7.308484e+09, 7.285175e+09, 
    7.260469e+09, 7.234377e+09, 7.206909e+09, 7.178077e+09, 7.147894e+09, 
    7.116371e+09, 7.083523e+09, 7.049361e+09, 7.013901e+09, 6.977157e+09, 
    6.939143e+09, 6.899874e+09, 6.859367e+09, 6.817636e+09, 6.774699e+09, 
    6.730571e+09, 6.685269e+09, 6.638811e+09, 6.591213e+09, 6.542493e+09, 
    6.492669e+09, 6.441759e+09, 6.38978e+09, 6.336752e+09, 6.282692e+09, 
    6.227619e+09, 6.171552e+09, 6.114508e+09, 6.056508e+09, 5.99757e+09, 
    5.937712e+09,
  5.885548e+09, 5.942029e+09, 5.99757e+09, 6.052155e+09, 6.105772e+09, 
    6.158404e+09, 6.210038e+09, 6.260659e+09, 6.310255e+09, 6.35881e+09, 
    6.406312e+09, 6.452746e+09, 6.4981e+09, 6.54236e+09, 6.585513e+09, 
    6.627547e+09, 6.668449e+09, 6.708208e+09, 6.74681e+09, 6.784244e+09, 
    6.8205e+09, 6.855565e+09, 6.889429e+09, 6.922081e+09, 6.953512e+09, 
    6.98371e+09, 7.012667e+09, 7.040374e+09, 7.066821e+09, 7.092e+09, 
    7.115902e+09, 7.138521e+09, 7.159848e+09, 7.179877e+09, 7.198601e+09, 
    7.216014e+09, 7.23211e+09, 7.246883e+09, 7.260329e+09, 7.272444e+09, 
    7.283223e+09, 7.292662e+09, 7.30076e+09, 7.307511e+09, 7.312915e+09, 
    7.316969e+09, 7.319673e+09, 7.321026e+09, 7.321026e+09, 7.319673e+09, 
    7.316969e+09, 7.312915e+09, 7.307511e+09, 7.30076e+09, 7.292662e+09, 
    7.283223e+09, 7.272444e+09, 7.260329e+09, 7.246883e+09, 7.23211e+09, 
    7.216014e+09, 7.198601e+09, 7.179877e+09, 7.159848e+09, 7.138521e+09, 
    7.115902e+09, 7.092e+09, 7.066821e+09, 7.040374e+09, 7.012667e+09, 
    6.98371e+09, 6.953512e+09, 6.922081e+09, 6.889429e+09, 6.855565e+09, 
    6.8205e+09, 6.784244e+09, 6.74681e+09, 6.708208e+09, 6.668449e+09, 
    6.627547e+09, 6.585513e+09, 6.54236e+09, 6.4981e+09, 6.452746e+09, 
    6.406312e+09, 6.35881e+09, 6.310255e+09, 6.260659e+09, 6.210038e+09, 
    6.158404e+09, 6.105772e+09, 6.052155e+09, 5.99757e+09, 5.942029e+09, 
    5.885548e+09,
  5.832426e+09, 5.885548e+09, 5.937712e+09, 5.988909e+09, 6.039129e+09, 
    6.088361e+09, 6.136596e+09, 6.183825e+09, 6.230037e+09, 6.275223e+09, 
    6.319373e+09, 6.362479e+09, 6.404531e+09, 6.445522e+09, 6.485442e+09, 
    6.524282e+09, 6.562035e+09, 6.598693e+09, 6.634248e+09, 6.668692e+09, 
    6.702019e+09, 6.734221e+09, 6.76529e+09, 6.795221e+09, 6.824007e+09, 
    6.851641e+09, 6.878117e+09, 6.903431e+09, 6.927576e+09, 6.950547e+09, 
    6.972339e+09, 6.992947e+09, 7.012366e+09, 7.030593e+09, 7.047623e+09, 
    7.063453e+09, 7.078078e+09, 7.091497e+09, 7.103705e+09, 7.1147e+09, 
    7.124479e+09, 7.133041e+09, 7.140384e+09, 7.146505e+09, 7.151404e+09, 
    7.155078e+09, 7.157529e+09, 7.158754e+09, 7.158754e+09, 7.157529e+09, 
    7.155078e+09, 7.151404e+09, 7.146505e+09, 7.140384e+09, 7.133041e+09, 
    7.124479e+09, 7.1147e+09, 7.103705e+09, 7.091497e+09, 7.078078e+09, 
    7.063453e+09, 7.047623e+09, 7.030593e+09, 7.012366e+09, 6.992947e+09, 
    6.972339e+09, 6.950547e+09, 6.927576e+09, 6.903431e+09, 6.878117e+09, 
    6.851641e+09, 6.824007e+09, 6.795221e+09, 6.76529e+09, 6.734221e+09, 
    6.702019e+09, 6.668692e+09, 6.634248e+09, 6.598693e+09, 6.562035e+09, 
    6.524282e+09, 6.485442e+09, 6.445522e+09, 6.404531e+09, 6.362479e+09, 
    6.319373e+09, 6.275223e+09, 6.230037e+09, 6.183825e+09, 6.136596e+09, 
    6.088361e+09, 6.039129e+09, 5.988909e+09, 5.937712e+09, 5.885548e+09, 
    5.832426e+09 ;

 bk = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.01253, 0.04887, 0.10724, 0.18455, 0.27461, 0.36914, 
    0.46103, 0.54623, 0.62305, 0.69099, 0.75016, 0.8011, 0.84453, 0.88125, 
    0.9121, 0.93766, 0.95849, 0.97495, 0.98743, 0.9958, 1 ;

 pk = 1, 2.69722, 5.17136, 8.89455, 14.2479, 22.07157, 33.61283, 50.48096, 
    74.79993, 109.4006, 158.0046, 225.4411, 317.8956, 443.1935, 611.1156, 
    833.7439, 1125.834, 1505.208, 1993.158, 2614.863, 3399.784, 4382.062, 
    5600.87, 7100.731, 8931.782, 11149.97, 13817.17, 17001.21, 20775.82, 
    23967.34, 25527.65, 25671.22, 24609.3, 22640.51, 20147.13, 17477.63, 
    14859.86, 12414.93, 10201.44, 8241.503, 6534.432, 5066.179, 3815.607, 
    2758.603, 1880.646, 1169.339, 618.4799, 225, 10, 0 ;

 sftlf =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0.2418439, 0, 0.1507849, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0.9672335, 0.7867691, 0.8897236, 0.7868192, 0.4295904, 0.103123, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 0.8583792, 0.24312, 0.02330228, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 0.7519304, 0.3075978, 0.05466554, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 0.7495267, 0.07681742, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.8367906, 0.08314215, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.341669, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9609066, 0.3417271, 0.0006489863, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.6232235, 0.1494775, 0.0620707, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.8576373, 0.4441393, 
    0.02198116, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9266944, 0.7165388, 0.8939224, 
    0.5627504, 0.03366798, 0.3162485, 0.02661187, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9785867, 0.3546079, 
    0.001069293, 0.5276027, 0.6956339, 0.8771922, 0.3122943, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.6351135, 0.1552348, 
    0.2120383, 0.6413907, 0.72313, 0.05286491, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.4744368, 
    0.01789349, 0.362444, 0.7183179, 0.6351389, 0.2321099, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.537541, 
    0.02737221, 0.1637618, 0.5896915, 0.6713976, 0.06366118, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.5861796, 
    0.0982726, 0.02536981, 0.1802837, 0.5701141, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.8579165, 
    0.275193, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.91327, 
    0.2402546, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.918274, 0.5621569, 0.0209811, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.588654, 0.3020536, 0.30206, 0.2020797, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 0.9413478, 0.1002747, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 0.6651581, 0.001533675, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 0.3886248, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 0.6325621, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 0.995119, 0.2749188, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 0.6972129, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.9737231, 0.9926948, 1, 1, 1, 1, 0.8642177, 0.08541915, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9564105, 
    0.4497338, 0.407091, 0.4070948, 0.4070986, 0.4071023, 0.2621634, 
    0.3688191, 0.6872182, 0.9677767, 1, 1, 1, 0.4953253, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.2941011, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.2652708, 0.8491837, 1, 1, 0.4804461, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.648157, 0.03258629, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0.4520298, 1, 1, 0.3871183, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9116583, 0.07233045, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1828122, 1, 1, 0.1171441, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.553419, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.08816408, 1, 1, 0.7507677, 0.04885805, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.6228713, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.3365233, 1, 1, 1, 0.5879625, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9385124, 0.1065637, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0.2791502, 0.6271809, 1, 1, 1, 0.9890413, 
    0.2517519, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1216078, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.6900454, 0.06213602, 
    0, 0, 0, 0, 0, 0, 0, 0.1037045, 0.7385923, 0.9886956, 1, 1, 1, 1, 1, 
    0.4103255, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.908018, 0.1728964, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.3633319, 1, 1, 1, 1, 1, 1, 1, 0.7623217, 
    0.0008263012, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.6658352, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.4360288, 0.957324, 0.635229, 0.4226641, 0.2175488, 
    0.3202175, 0.8472205, 1, 0.9694546, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.5564398, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.2841633, 0.1100108, 0, 0, 0, 0, 0.8772225, 1, 0.9926439, 
    0.7188581, 0.01636519, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.6282753, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.9419357, 1, 1, 1, 0.5849457, 0.315834, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9848972, 0.2503584, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01595704, 0.995867, 1, 1, 1, 1, 
    0.9787351, 0.2506236, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.6914676, 0.02198116, 0, 
    0, 0, 0, 0, 0, 0.08334821, 0.1012918, 0, 0, 0, 0, 0, 0.005334743, 
    0.7088248, 1, 1, 1, 0.8540698, 0.9996781, 0.6620048, 0.03839629, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9575872, 0.6579381, 
    0.3669165, 0, 0, 0, 0, 0, 0.5810857, 0.3034903, 0, 0, 0, 0, 0, 0, 
    0.07322878, 0.3065482, 0.1025856, 0.1025909, 0.06481452, 0.2606909, 
    0.8556811, 0.4936866, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9884753, 0.8030674, 
    0.2831464, 0, 0, 0, 0.4692461, 0.05008297, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.2312002, 0.6806778, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.8807496, 0.4964221, 0.118718, 
    0.2605629, 0.7617009, 1, 1, 0.9638987, 0.2762473, 0, 0.01970084, 
    0.866532, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.03466008, 0.9590737, 
    0.3642623, 0, 0, 0, 0, 0, 0, 0, 0.03183588, 0.3728453, 0.1801692, 
    0.07776905, 0.3728562, 0.2684634, 0.07811955, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.825218, 0.1281082, 0, 0, 0, 
    0.05450449, 0.1359098, 0.6320257, 0.6364659, 0.07199212, 0, 0.07605698, 
    0.7873569, 0.08185559, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.5112837, 
    0.5608108, 0.3629351, 0, 0, 0, 0, 0, 0, 0.3923621, 0.8759633, 1, 
    0.9305333, 0.6235623, 1, 0.9620325, 0.6514717, 0.1631414, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.7229308, 0.07197631, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.8089566, 0.1385804, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.718082, 0.0345762, 0, 0, 0, 0, 0, 0, 0.3329219, 0.987651, 1, 1, 1, 1, 
    1, 1, 1, 0.9168873, 0.5666844, 0.05440859, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.8832299, 0.1472945, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.4424467, 0.1988707, 0.007988392, 0.4272325, 0.7964597, 0.1058136, 0, 
    0.1016413, 0.03233812, 0, 0, 0, 0, 0, 0, 0, 0, 0.4837731, 0.6387944, 
    0.2020133, 0, 0, 0, 0.0193575, 0.5679138, 0.9483995, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 0.8473101, 0.6221716, 0.1199134, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9533704, 0.1238984, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.1078062, 4.039702e-05, 0.02094627, 0.7635151, 0.6279824, 0, 
    0.4214649, 0.03240846, 0, 0, 0, 0, 0, 0, 0, 0, 0.1298708, 0.9593522, 
    0.8726715, 0.6254805, 0.6615382, 0.6156211, 0.7938948, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 0.8723933, 0.576844, 0.1146775, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  1, 1, 1, 0.9439595, 0.8502378, 0.4763551, 0.4259781, 0.7869197, 0.754113, 
    0.2165837, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.483312, 
    0.5854645, 0, 0.1202012, 0, 0, 0, 0, 0, 0, 0, 0, 0.01637845, 0.6564068, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.859898, 0.7360823, 0.2172089, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 0.6529251, 0.507857, 0.3280367, 0.03502538, 0, 0.1547292, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1886325, 0.4330523, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.4363211, 0.7168808, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.8921524, 0.3981088, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0,
  1, 0.9714789, 0.9004541, 0.4634776, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0.05552825, 0.120399, 0.03792001, 0.00843242, 0, 
    0, 0, 0, 0, 0, 0.07417351, 0.8822758, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.8686383, 0.1390514, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.01985216, 0.09956025, 0.09957455,
  0.9850286, 0.5513424, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.01466178, 0.4497637, 0.01945193, 0, 0, 0, 0, 0, 0, 
    0.2087137, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 0.7150637, 0.00703513, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01038911, 0.03078478, 0.5223621, 
    0.5656272, 0.5656678, 0.6186966, 1, 0.975225,
  0.5147771, 0.2509983, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.01205661, 0.5400833, 0.6323332, 0, 0, 0, 0, 0, 0, 
    0.0640404, 0.8329736, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.5314379, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.06310866, 0.6251156, 1, 1, 1, 1, 1, 
    1, 1,
  0.04331701, 0.004251128, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.7602282, 0.9885215, 0.1360401, 0, 0, 0, 0, 0, 
    0.5068112, 0.1770562, 0.9897748, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9330676, 0.3697935, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.2310756, 0.410401, 0.4104408, 
    0.4104811, 0.4105217, 0.4105628, 0.6770073, 0.9558303, 1, 1, 1, 1, 1, 1, 
    1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.003479148, 0.9392874, 0.5581517, 0.007009166, 0, 0, 0, 0, 0, 0.1731326, 
    0.4696587, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9879944, 0.3274225, 0.317915, 
    0.008586753, 0.1531166, 0.007366235, 0.3192428, 0.3195822, 0.3196146, 
    0.3196478, 0.3314601, 0.8600246, 0.8667862, 0.9326418, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.01336217, 0.6549731, 0.145487, 0, 0, 0, 0, 0, 0, 0.1268012, 0.9062009, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.7842681, 0.8845835, 0.7709545, 0.9917373, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.4637389, 0.1322377, 0, 0, 0, 0, 0, 0, 0.03724731, 0.7512087, 
    0.9969589, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.03823176, 0.9980064, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.1325942, 0.07740931, 0, 0, 0, 0, 0, 0, 0, 0.1540521, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.3038891, 0.04776999, 0, 0, 0, 0, 0, 0, 0, 0.1829891, 0.9730953, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.03913443, 0.0341659, 0, 0, 0, 0, 0, 0, 0, 0, 0.009582857, 0.9771051, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.1451908, 0.07445376, 0, 0, 0, 0, 0, 0, 0, 0, 0.3511962, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0.3498454, 0.9953002, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0.2403926, 0.9019648, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.005788924, 0.01535262, 0, 0, 0, 0, 0, 0.1437764, 0.2917262, 
    0.9888229, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.1149602, 0.1676279, 0, 0, 0, 0, 0, 0.2839805, 0.2067913, 
    0.6178907, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1299978, 0.9375334, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.5485037, 0.9940798, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.4170257, 0.986974, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.8614578, 0.9180768, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0009119348, 0.393558, 0.9921986, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 0.9273752, 0.1889167, 0.7825502, 0.8380716,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0002601096, 0.8132703, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 0.6767043, 0.05085213, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.04240416, 0.8030222, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 0.8947946, 0.0665093,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.2244188, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.5003253 ;

 orog =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01534718, 
    0.004565009, 0.008999515, 0.009599131, 0.0008479413, 0, 0, 0.0007195598, 
    0.004574103, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.7068716, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.003399682, 
    0.0147934, 0.002706561, 0, 0, 0, 0.004826599, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.004755895, 
    0.00314351, 0.002793752, 0, 0, 0, 0.006179405, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.006290677, 
    0.007201957, 0, 0.01463142, 0.003162183, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.008779748, 0, 0, 0, 
    0.00300725, 0.002690252, 0.005241457, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 1.506357, 3.305288, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.007343553, 0, 0.009825814, 0.01535672, 0.006712195, 0, 0, 0.005644962, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19.68891, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.008339305, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.00178691, 18.51452, 0.01244308, 0, 0, 0, 
    0, 0.009080717, 0, 0, 0, 0, 0.006611669, 0.003060021, 0.008406991, 0, 
    0.005074322, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01017599, 
    0, 0, 0, 0.004030156, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.003469607, 0, 0, 0, 0, 0, 0.002995649, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.004560474, 0, 0, 0.01124365, 0.003597797, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.01154227, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.2431989, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.001374771, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.06463672, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.1425494, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  33.14798, 0, 34.79201, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.0004971988, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  668.3605, 750.8135, 625.5392, 386.1679, 158.3386, 2.453814, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1070.732, 1178.2, 1004.681, 772.6516, 403.6846, 150.0447, 26.30301, 
    1.64736, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1507.715, 1421.274, 1144.302, 833.4024, 441.414, 72.99273, 109.9673, 
    184.5779, 220.3756, 0.00647221, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1551.811, 1623.509, 1564.146, 1482.56, 1154.821, 803.4989, 487.0388, 
    202.9149, 268.4435, 226.8269, 46.07853, 0.3954178, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0,
  1557.897, 1671.874, 1696.626, 1635.232, 1700.021, 1734.235, 1559.076, 
    995.3284, 449.7531, 276.2559, 565.8065, 21.12218, 0.8193069, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1468.874, 1600.571, 1614.583, 1414.91, 1396.924, 1757.31, 2173.984, 
    2018.616, 1396.95, 1025.211, 762.0422, 232.5291, 8.014444, 1.140886, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0,
  1326.019, 1541.283, 1555.617, 1480.098, 1514.677, 1689.735, 1982.568, 
    2007.651, 1670.599, 1186.88, 1048.513, 684.1181, 117.3529, 0.1669138, 0, 
    0, 0, 14.15248, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1146.4, 1447.466, 1700.664, 1654.412, 1747.869, 2042.93, 1975.362, 
    1731.381, 1260.238, 1003.032, 874.1664, 965.1847, 711.4643, 390.3766, 
    173.5833, 3.412067, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1373.781, 1329.12, 1740.19, 1867.481, 1919.821, 2046.155, 2020.59, 
    1730.883, 1388.832, 990.3948, 863.0721, 733.3089, 488.1863, 444.3896, 
    642.3708, 630.8365, 208.2363, 11.2473, 0.03753853, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1914.861, 1386.722, 1730.161, 1876.041, 1894.845, 2047.599, 1965.026, 
    1787.49, 1283.865, 1007.386, 831.1433, 589.1078, 291.1984, 130.3001, 
    245.2175, 308.7728, 423.5323, 287.8249, 17.96172, 32.98395, 0.1041703, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.1970985, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  2061.196, 1476.068, 1648.332, 1574.314, 1569.191, 1744.371, 1828.933, 
    1790.968, 1558.644, 1149.688, 1213.996, 906.5831, 504.1509, 233.0578, 
    183.2224, 38.9668, 0.0118664, 233.6236, 272.1967, 144.2618, 56.46022, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  1840.156, 1504.441, 1582.167, 1490.926, 1402.836, 1518.827, 1694.572, 
    2058.519, 1824.339, 1671.718, 1643.01, 1482.167, 815.0604, 396.3656, 
    379.8361, 318.8223, 100.745, 65.86816, 107.3457, 244.7698, 250.1199, 
    15.35586, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0,
  1837.63, 1728.632, 1902.097, 1719.298, 1875.763, 1918.201, 2012.239, 
    2196.799, 2065.854, 1799.648, 1839.158, 1689.026, 1220.946, 556.4898, 
    653.7017, 762.9083, 615.2339, 393.6399, 83.12075, 4.564439, 169.0518, 
    231.0936, 86.59752, 8.810427, 0, 0, 0, 0, 0.004199471, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  2287.553, 2375.422, 2227.182, 2205.671, 2448.729, 2173.713, 2069.91, 
    1804.564, 1718.86, 1645.912, 1760.087, 1774.775, 1588.443, 1158.239, 
    1042.855, 1238.964, 1055.679, 720.4163, 300.8953, 74.61289, 2.083953, 
    10.21264, 134.772, 93.68505, 9.525565, 0, 0, 0, 0.06281511, 3.428892, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  2614.957, 2546.323, 2390.928, 2148.965, 2257.577, 2052.22, 1766.787, 
    1770.134, 1673.074, 1765.732, 1825.648, 1895.919, 1992.829, 1695.072, 
    1362.996, 1422.211, 1302.389, 1040.16, 627.5578, 400.1667, 51.56722, 
    2.257818, 0.1849899, 56.72547, 250.1037, 1.460486, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.967957, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1897.78, 2076.201, 2129.073, 2115.72, 2166.538, 1872.045, 2072.919, 
    1904.649, 2256.727, 1803.393, 1983.677, 2108.663, 2195.764, 2050.119, 
    1605.954, 1432.204, 1511.048, 1487.268, 1426.227, 1196.583, 721.2061, 
    185.3391, 24.12744, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0004704067, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.2958491, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1716.921, 1748.802, 1939.11, 2058.646, 2214.479, 2215.264, 2299.508, 
    2683.908, 2679.552, 2308.606, 2102.935, 2086.155, 2177.915, 2051.186, 
    1598.307, 1383.17, 1438.509, 1773.132, 2076.03, 2118.625, 1700.985, 
    1170.254, 459.9845, 48.66238, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1594.9, 1717.709, 1846.341, 2183, 2416.479, 2646.638, 2920.714, 2901.701, 
    3107.744, 2624.682, 2306.014, 2028.034, 1806.9, 1723.413, 1505.019, 
    1253.708, 1291.276, 1617.983, 1898.304, 2037.906, 2075.454, 2108.36, 
    1570.701, 841.1761, 129.8114, 0.2389687, 3.660637, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1414.581, 1499.586, 1735.549, 1988.982, 2430.141, 2544.231, 2714.589, 
    2826.258, 2566.761, 2620.082, 2419.738, 2052.477, 1891.764, 1767.929, 
    1617.863, 1432.407, 1338.126, 1367.179, 1424.379, 1473.549, 1661.907, 
    2049.929, 2230.574, 1919.274, 1373.336, 316.5095, 39.45748, 94.61289, 
    39.49365, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    7.207365e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1235.553, 1437.662, 1381.895, 1611.005, 1679.951, 1728.312, 1922.424, 
    1964.016, 1953.016, 2112.162, 2098.977, 1710.801, 1526.079, 1414.803, 
    1368.911, 1237.472, 1292.035, 1341.555, 1204.039, 1329.621, 1429.259, 
    1572.953, 1800.086, 2189.089, 2119.821, 1455.417, 1083.626, 1022.557, 
    862.4561, 51.87525, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1174.93, 1228.427, 1291.553, 1290.888, 1424, 1351.69, 1468.16, 1589.555, 
    1427.788, 1689.11, 1630.9, 1414.054, 1334.024, 1248.547, 1122.594, 
    1033.518, 1091.201, 1192.766, 1168.232, 1309.946, 1314.83, 1245.706, 
    1400.043, 1858.552, 2194.833, 2118.342, 1668, 1707.535, 1364.425, 
    595.4224, 15.76594, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  823.5144, 966.8268, 1033.309, 1192.71, 1210.489, 1193.993, 1280.92, 
    1308.805, 1209.215, 1289.174, 1294.622, 1176.932, 1193.732, 1146.91, 
    1025.355, 875.7115, 882.8735, 978.463, 1033.714, 1232.486, 1255.239, 
    1216.565, 1342.363, 1716.272, 2074.805, 2120.552, 2071.005, 1786.363, 
    1785.419, 844.6271, 169.2518, 0.001837272, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  661.3832, 741.7489, 952.168, 1073.759, 1053.268, 1013.894, 1031.548, 
    1062.557, 1014.31, 1013.214, 1007.304, 1006.718, 987.2679, 929.3942, 
    846.1819, 807.7843, 729.1191, 717.0919, 644.5469, 733.0809, 815.4983, 
    1055.672, 1469.535, 1941.911, 2045.901, 2101.024, 2062.683, 2086.129, 
    1883.878, 989.241, 529.9884, 1.092551, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0,
  574.1776, 618.1168, 795.5441, 907.0357, 894.5935, 851.0385, 820.7712, 
    843.4498, 837.6264, 813.8089, 821.1804, 790.303, 694.8225, 637.4512, 
    626.2227, 661.035, 688.275, 597.9715, 427.0944, 299.6628, 342.4961, 
    676.9834, 1214.729, 1706.491, 1881.969, 1649.495, 1733.168, 2044.59, 
    2105.82, 1415.646, 915.3256, 166.6185, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0,
  503.9159, 538.9011, 631.793, 737.8944, 750.1324, 703.1216, 655.9878, 
    654.8143, 672.593, 642.7423, 621.7355, 602.098, 473.79, 425.5311, 
    461.755, 530.6566, 568.3069, 558.3639, 330.7892, 179.9599, 143.326, 
    168.8803, 392.449, 875.6781, 1042.997, 940.2807, 1005.778, 1682.482, 
    2467.645, 1832.106, 1341.977, 441.4869, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0,
  453.9662, 441.7195, 504.0019, 592.8539, 608.1069, 578.1291, 526.2635, 
    513.4938, 532.1535, 479.4901, 447.4254, 444.3315, 379.7191, 325.8571, 
    347.1577, 396.39, 397.7914, 382.2119, 225.9507, 114.7197, 95.74188, 
    70.67721, 57.3841, 157.933, 314.682, 123.271, 156.6136, 1009.174, 
    2106.859, 2219.086, 1513.035, 924.8544, 29.27477, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  503.6515, 465.5753, 433.9768, 478.4191, 482.0991, 473.893, 436.3061, 
    425.1155, 431.4804, 382.6123, 325.8517, 340.3661, 314.822, 260.5178, 
    239.2539, 233.0164, 209.3085, 185.2675, 99.46118, 35.69082, 15.04999, 
    5.81494, 7.321244, 7.285094, 10.49513, 6.034019, 12.30279, 178.9217, 
    1494.86, 1747.576, 1843.446, 1614.362, 380.1558, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  438.2668, 471.7402, 408.1164, 400.8929, 380.3304, 374.7529, 382.5601, 
    372.2382, 382.916, 320.6809, 264.4974, 252.2818, 258.8326, 194.5873, 
    162.8055, 141.8769, 114.3217, 85.31949, 39.80796, 4.830305, 0, 0, 0, 0, 
    0, 0, 0, 0.02132653, 176.2921, 430.069, 932.7458, 1392.24, 747.5593, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  375.052, 414.3507, 415.5859, 381.3595, 361.0887, 329.3397, 313.1617, 
    313.8601, 298.01, 280.3281, 250.9803, 220.6591, 244.4896, 157.4741, 
    126.7682, 118.9209, 91.80339, 46.5208, 11.15798, 0.09899135, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 50.89595, 153.9082, 606.8809, 122.0387, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0,
  304.4448, 364.8189, 357.5074, 352.7218, 337.0601, 318.3467, 277.0119, 
    265.5412, 282.2703, 328.1339, 341.168, 288.7758, 254.3146, 138.1611, 
    97.54157, 97.74657, 73.76514, 23.01658, 0.5496842, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 3.476873, 75.94135, 449.1298, 34.83492, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  306.857, 361.5244, 342.5269, 300.4066, 292.6741, 274.3279, 251.7741, 
    245.3346, 294.167, 380.9618, 372.6419, 271.2439, 204.3829, 99.51021, 
    69.604, 73.45421, 50.67704, 12.05578, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3.512501, 149.8454, 851.515, 526.5105, 5.040119, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  319.7339, 346.4661, 325.2934, 268.1579, 235.2851, 243.1511, 224.0061, 
    242.3429, 319.4263, 334.612, 274.955, 164.2817, 109.9028, 55.26638, 
    47.65622, 41.80495, 35.97699, 2.775469, 0.03288275, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 6.357764, 280.3884, 1031.42, 1222.137, 606.0325, 0.7514994, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.07952388, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  294.8905, 319.0948, 294.4915, 238.6062, 212.2333, 193.6535, 202.8654, 
    221.7048, 288.9077, 248.9493, 137.382, 84.58096, 51.21586, 40.6296, 
    44.39739, 63.04242, 40.62316, 8.783824, 0.268134, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.7404718, 15.12963, 65.80754, 738.6376, 1257.209, 1292.93, 64.7064, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13.92286, 118.2891, 0.07517834, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  313.3622, 298.425, 277.4745, 233.6075, 198.1856, 187.4898, 173.2009, 
    175.6373, 200.6465, 144.9214, 80.57291, 77.81576, 66.51388, 73.39558, 
    92.76784, 95.03912, 61.3536, 3.831983, 0.1158118, 0, 0, 0, 0, 0, 0, 0, 
    0.6463583, 18.92656, 71.69862, 132.442, 95.90388, 289.954, 763.129, 
    1148.201, 229.1096, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.065996, 
    17.50426, 2.459143, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  289.323, 276.3043, 265.5132, 220.7219, 216.1242, 195.0884, 181.3391, 
    143.4675, 147.2648, 111.0426, 110.6656, 125.9561, 122.3719, 105.6208, 
    113.7486, 98.84241, 43.68995, 0.9661562, 0.02680171, 0, 0, 0, 0, 0, 0, 0, 
    3.878528, 38.69389, 97.16181, 132.8956, 207.0652, 216.3446, 424.0393, 
    918.3037, 351.0448, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6.011113, 
    0.1137814, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  230.5823, 241.4872, 225.9881, 214.9098, 207.3458, 206.6044, 173.4783, 
    138.0395, 130.4559, 142.9235, 167.6159, 175.7432, 143.494, 103.3232, 
    73.60364, 63.91725, 27.10206, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10.20466, 
    20.16096, 25.27402, 21.63544, 14.64767, 43.60937, 331.3476, 893.1275, 
    454.1429, 1.288543, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  191.6571, 178.5321, 189.9285, 201.3738, 214.7888, 215.5745, 179.5497, 
    147.2228, 153.1658, 179.6961, 230.3224, 239.8835, 194.1318, 137.8888, 
    87.66043, 69.8594, 27.32165, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6.084438, 
    6.930506, 0.584422, 0.003764597, 0.003457344, 0.4655042, 543.0778, 
    932.6347, 615.3885, 85.28525, 0.2777186, 0, 0, 0, 0, 0, 0.422377, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0,
  231.2289, 207.4846, 224.9596, 237.2916, 248.9516, 252.8323, 212.7034, 
    195.5234, 197.4957, 263.0653, 303.2209, 280.5213, 264.7434, 194.2222, 
    116.7919, 78.11273, 25.05218, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    4.827813, 526.7432, 777.7427, 639.5916, 362.6419, 79.72997, 29.67748, 
    0.912546, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  278.9553, 267.2621, 269.6895, 261.4806, 287.7636, 281.252, 243.8186, 
    240.3938, 298.7545, 342.4502, 399.08, 363.9893, 266.6101, 221.5975, 
    126.7727, 76.75681, 26.75876, 0.9402217, 0, 0, 0, 0, 0, 0, 0, 0.3805751, 
    0, 0, 0, 0, 0, 3.231741, 309.7996, 351.9758, 387.7886, 218.6437, 153.275, 
    263.9878, 54.07672, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  241.8856, 246.4237, 245.6055, 259.1919, 286.3187, 285.9484, 254.3894, 
    280.3928, 369.3888, 439.415, 618.7897, 387.4653, 291.7344, 174.3447, 
    113.5729, 67.22175, 24.12755, 0, 0, 0, 0, 0, 0, 0, 20.0383, 16.96434, 0, 
    0, 0, 0, 0.003687347, 0.00572379, 52.21835, 70.8857, 55.61906, 70.92522, 
    123.4313, 420.684, 636.3296, 6.528507, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  202.4083, 219.8558, 207.086, 261.2129, 295.0167, 264.0109, 249.5903, 
    352.6951, 497.0891, 679.3617, 595.9517, 404.6982, 150.7021, 114.5868, 
    78.8996, 54.99938, 26.96955, 5.426031, 1.965392, 0.1738949, 0, 0, 0, 0, 
    39.73782, 6.958992, 0, 0, 0, 0, 0, 0.0001729098, 1.584328, 6.905681, 
    0.7596173, 0.490705, 0, 84.19572, 863.5649, 289.1957, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  210.9862, 176.5489, 218.8383, 299.7639, 293.6812, 247.376, 300.3907, 
    490.8528, 720.3207, 577.838, 503.2361, 148.1991, 107.7899, 63.81637, 
    42.55847, 31.07135, 27.5754, 28.17957, 28.8343, 16.63614, 2.660592, 0, 
    0.01031376, 0.9608897, 33.86351, 0.509288, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.05132846, 0, 0, 160.5816, 333.4066, 8.909275, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  247.1366, 214.9977, 272.471, 323.8452, 298.5703, 362.521, 537.7053, 
    668.5198, 624.8367, 453.5524, 165.6625, 102.4959, 57.48196, 21.7608, 
    4.573749, 1.787246, 5.738702, 13.79587, 21.61514, 15.3555, 7.805641, 
    1.753023, 0.05135195, 1.186182, 39.27137, 0.8040789, 0, 0.01927231, 
    0.09756799, 0, 0, 0, 0, 0, 0.1619276, 0, 0, 0, 9.406398, 314.6326, 
    92.01137, 0, 0, 0.001729056, 0, 0, 0, 0, 0.6381596, 31.72947, 4.45034, 
    6.862898, 161.6274, 35.41436, 10.87154, 0.005455857, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2.744836, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  229.433, 306.0153, 351.427, 376.3137, 463.0498, 627.9566, 686.7066, 
    565.6674, 405.129, 181.5926, 102.0433, 47.04384, 16.67009, 1.10613, 0, 0, 
    0, 0.09115441, 1.67472, 5.002741, 3.653378, 0.914476, 0.0004763628, 
    1.392298, 81.95518, 36.95679, 0, 0.102858, 0, 0, 0, 0, 0, 7.409501e-05, 
    0, 0, 0, 0, 55.38284, 97.32481, 47.17434, 0, 0, 0, 0, 0, 0.03468706, 
    60.15501, 130.7003, 244.7536, 135.677, 424.9022, 731.8262, 553.5016, 
    151.7469, 15.67891, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.1039039, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  298.4516, 455.0074, 496.0555, 490.0974, 549.4736, 625.2988, 487.0647, 
    277.1122, 157.1025, 104.1153, 47.97492, 9.955524, 1.711641, 0, 0, 0, 0, 
    0, 0, 0.08672119, 0.02051163, 0.0005947647, 0, 0.02029713, 58.99087, 
    18.83587, 0.0248516, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 110.5765, 3.497101, 
    0, 0, 0, 0, 0, 0.05597858, 47.99405, 655.0215, 1362.752, 1510.303, 
    1890.99, 1900.117, 1904.355, 1649.458, 1608.771, 1245.189, 378.5316, 
    4.13827, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 1.282194, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  430.407, 573.2601, 458.0574, 384.715, 322.2038, 270.0156, 169.9159, 
    89.97162, 81.54353, 47.91539, 13.97083, 0.9449826, 0, 0, 0, 0, 0, 0, 
    0.0004252571, 0.3309443, 0.03876647, 1.728635, 0.4185002, 0, 15.5728, 
    39.27885, 1.380751, 0.007368555, 55.84319, 1.191139, 0, 0, 0, 0, 0, 0, 0, 
    0, 115.976, 114.2675, 74.08803, 0, 0, 0, 0.3069585, 74.61648, 1023.105, 
    1976.442, 2391.624, 2180.577, 1604.411, 1326.77, 901.5997, 1351.656, 
    2254.224, 2631.384, 2637.751, 1822.456, 620.1605, 20.8799, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  430.7066, 471.0601, 333.3573, 224.1613, 108.1152, 65.5984, 26.94351, 
    37.64307, 24.10448, 10.83371, 1.795868, 0, 0, 0, 0, 0, 0, 0, 0, 0.421066, 
    0.211959, 0.211567, 0.4754283, 0, 1.457668, 49.35142, 77.70663, 0.225208, 
    177.6199, 27.2492, 0, 0, 0, 0, 0, 0, 0, 0, 16.10499, 144.5139, 247.1739, 
    155.9424, 68.87181, 112.7537, 548.5216, 1326.625, 1537.927, 1522.117, 
    1053.582, 538.7177, 494.4248, 237.3714, 225.9437, 723.8336, 1495.832, 
    2103.182, 2873.699, 3292.384, 3380.365, 2269.825, 515.0248, 4.337821, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0,
  431.9473, 396.6402, 222.4012, 114.462, 25.37888, 7.691118, 6.677791, 
    7.348661, 3.157577, 0.984972, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.3024256, 
    0.2389092, 0.1394803, 0.00746349, 0, 70.57438, 149.7564, 0, 80.11617, 
    0.0417327, 0, 0, 0, 0, 0, 0, 0, 0.01057512, 27.73273, 266.8832, 915.6628, 
    1100.12, 1117.166, 1315.549, 1758.784, 2041.483, 1431.61, 474.8531, 
    232.1502, 208.0247, 196.3371, 166.9769, 139.262, 189.603, 539.9, 
    636.6401, 1134.973, 2116.188, 3255.661, 3725.555, 3525.62, 2041.445, 
    414.1652, 93.96832, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  441.435, 319.8361, 136.8747, 29.58521, 4.141918, 2.825089, 0.08903898, 
    0.08046266, 0.2208437, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.3990609, 
    0.3265876, 0.0633444, 0.05431467, 84.71734, 149.596, 0, 0.04963135, 0, 0, 
    0, 0, 0, 0, 0, 27.05583, 59.55542, 2.632703, 383.2401, 1071.188, 
    1466.155, 1676.46, 1735.292, 1635.764, 1205.279, 587.2426, 204.6946, 
    192.8305, 201.6285, 192.1485, 173.3057, 135.0386, 115.5985, 154.6932, 
    207.6518, 252.7319, 408.4037, 1234.129, 2512.059, 3625.666, 3840.744, 
    2953.312, 1398.119, 200.1961, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  298.2758, 155.1034, 25.55248, 4.920603, 0.003125044, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1279996, 0.02609903, 0.3170911, 0, 23.67887, 
    68.64729, 35.86671, 72.66331, 0, 0, 0, 0, 0, 0, 27.26858, 361.5938, 
    62.6906, 207.8889, 270.3431, 466.9674, 991.8314, 1723.766, 1665.32, 
    1134.25, 697.3764, 239.1669, 204.7155, 192.0341, 177.9332, 167.6514, 
    147.1711, 124.0248, 116.1455, 138.7632, 205.803, 202.1669, 218.9659, 
    445.2673, 918.5952, 2052.283, 3110.208, 3814.63, 3245.299, 1978.916, 
    128.154, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.621783, 0, 0, 1.331606, 2.106077,
  156.3812, 18.64756, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.02620244, 0.1723592, 0.6139864, 0.7052164, 39.91206, 73.66648, 
    34.73109, 0, 0, 0, 0, 0, 0, 103.6746, 970.1916, 637.6611, 308.0594, 
    768.11, 1294.207, 1777.075, 1670.896, 1144.713, 449.2721, 228.4367, 
    250.4818, 226.3325, 198.0396, 169.848, 146.4091, 131.5473, 124.774, 
    133.6427, 162.3437, 232.3307, 229.8633, 231.2848, 277.8121, 478.211, 
    827.6024, 1960.805, 3358.45, 4059.359, 3432.779, 1310.91, 0.5703501, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11.00629, 
    172.8352, 183.9977, 46.27448, 129.1229, 178.4515, 97.62695,
  36.70903, 1.210476, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.226078, 0.04288947, 3.178066, 257.9394, 343.0803, 13.00084, 0, 
    0, 0, 0, 0, 2.137605, 96.99342, 646.0239, 147.4564, 527.7556, 1280.455, 
    1827.782, 1949.41, 1110.227, 192.4001, 183.5117, 228.3509, 244.9112, 
    227.8943, 192.5254, 159.7048, 137.4386, 124.2721, 122.957, 142.0076, 
    164.3923, 198.738, 229.3472, 259.537, 313.7084, 313.5366, 602.6287, 
    1546.649, 3188.223, 4339.325, 4235.496, 2657.681, 348.9787, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15.4312, 110.2107, 
    133.0185, 292.7062, 324.6068, 298.3218, 359.0092, 476.8519, 554.6548,
  1.995229, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.4212663, 0.04588909, 11.18899, 517.642, 542.4244, 51.31382, 0, 0, 0, 0, 
    0, 43.47145, 14.86237, 90.16446, 49.90094, 852.6797, 695.9244, 698.5693, 
    469.248, 149.1092, 136.4317, 196.3584, 211.3587, 231.4343, 214.1757, 
    171.0396, 141.9184, 127.4874, 119.4414, 115.9838, 130.7626, 159.6196, 
    192.4039, 226.2965, 268.5108, 312.2362, 358.5796, 389.9218, 1083.607, 
    2472.518, 4258.277, 4571.348, 3741.117, 2121.892, 269.5249, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 4.388186, 133.4869, 148.3846, 211.8387, 382.2953, 
    257.1787, 180.7228, 149.7092, 212.2956, 459.678, 761.8045, 1055.912, 
    1120.853, 1110.582, 1166.25, 1085.751, 1108.78,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.001913318, 33.17125, 520.3718, 399.8852, 0, 0, 0, 0, 0, 0, 0.8113799, 
    95.28371, 460.3841, 937.3494, 915.1066, 445.8253, 106.3576, 103.3282, 
    112.4795, 164.6748, 183.3819, 200.0266, 220.7052, 195.8168, 166.651, 
    121.4309, 123.9416, 113.4673, 102.3118, 125.9921, 156.5412, 179.7962, 
    206.3467, 238.4389, 260.7508, 315.1216, 328.1903, 360.6142, 1509.248, 
    3565.005, 4402.538, 4396.66, 3602.803, 2091.149, 261.0787, 82.22005, 
    0.2868135, 0, 0.5076911, 60.36261, 183.4623, 519.5708, 450.9728, 
    353.2507, 488.7053, 617.8168, 1421.896, 2045.6, 2299.798, 2328.442, 
    2164.863, 1835.325, 1553.868, 1649.168, 1826.316, 1985.27, 1961.338, 
    1556.79, 1371.403, 1288.084, 1040.601, 1072.717,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5.771062, 165.8212, 28.28846, 0, 0, 0, 0, 0, 0.1610673, 17.69787, 
    260.4066, 714.0234, 586.6948, 462.326, 79.98116, 88.8905, 101.472, 
    127.5234, 151.2906, 172.9191, 187.4914, 183.702, 173.0886, 139.7318, 
    124.8896, 118.3931, 105.5773, 109.4129, 131.1672, 156.9932, 163.0083, 
    184.8383, 204.416, 225.2426, 266.9706, 316.145, 224.5979, 381.9278, 
    2492.509, 3806.261, 4259.841, 4400.584, 3759.828, 2950.103, 2123.126, 
    1457.011, 1071.604, 1158.814, 1261.4, 1360.847, 1651.959, 2091.039, 
    2134.101, 2298.518, 2832.512, 3516.553, 3862.269, 3539.123, 3228.904, 
    3070.49, 3133.28, 3088.744, 2907.435, 2507.032, 2134.26, 1858.328, 
    1274.926, 962.0797, 842.9384, 710.9687, 939.0226,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 51.69876, 6.425387, 0, 0, 0, 0, 0, 0, 2.873953, 169.8395, 449.1624, 
    300.1902, 62.32654, 69.31486, 78.20786, 85.0916, 97.69564, 127.4337, 
    145.2199, 162.7987, 148.36, 126.3364, 126.9805, 112.7666, 113.0274, 
    97.65716, 107.4775, 138.243, 148.1546, 151.6598, 170.6716, 190.0256, 
    201.0505, 226.6755, 261.319, 232.2254, 219.3973, 932.7808, 2511.412, 
    3070.967, 3937.193, 4288.645, 4117.858, 3970.56, 3654.04, 3348.081, 
    3098.408, 2970.42, 2560.729, 2923.75, 3655.134, 3966.941, 4254.809, 
    4391.425, 4123.873, 3285.485, 2428.365, 1895.18, 1763.043, 1610.22, 
    1446.99, 1407.953, 1387.499, 1476.249, 1487.882, 1047.58, 652.7329, 
    528.4442, 542.4118, 917.0056,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.3669669, 0.3634669, 0, 0, 0, 0, 0, 0, 0.6933007, 13.2217, 484.2191, 
    144.2932, 49.07107, 47.2271, 55.1874, 111.1454, 210.9041, 104.5796, 
    116.9778, 131.3689, 115.879, 101.3334, 98.76527, 97.77927, 91.92683, 
    82.82296, 102.0775, 115.0132, 128.6879, 136.6141, 155.6852, 166.7384, 
    172.6179, 192.5376, 207.4939, 206.3573, 175.2231, 245.1321, 792.022, 
    1577.401, 2693.881, 3723.349, 4046.354, 3911.702, 3846.095, 3873.51, 
    4067.074, 4060.027, 3885.769, 3648.284, 4000.79, 4255.121, 4298.765, 
    3941.536, 2986.297, 2167.081, 1555.988, 1086.933, 981.1671, 671.5908, 
    517.9108, 560.5896, 604.6505, 737.5284, 838.4316, 663.5747, 487.8661, 
    405.7701, 432.4994, 598.6184,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 87.07624, 9.664433, 0, 0, 0, 0, 0, 0, 0.1396964, 165.1147, 498.7843, 
    209.5764, 50.07817, 49.66368, 196.0763, 442.8151, 358.6526, 227.8948, 
    104.9866, 105.646, 125.2638, 109.2299, 82.44156, 78.38992, 73.12806, 
    72.46248, 85.68304, 100.9489, 111.212, 121.0391, 131.6541, 139.9958, 
    153.3166, 166.8747, 176.9339, 177.9256, 166.0943, 164.8257, 217.7268, 
    390.218, 1575.724, 3050.704, 3828.212, 3839.21, 3919.247, 3790.678, 
    3970.27, 4419.288, 4398.239, 4177.742, 4184.263, 4184.499, 4041.16, 
    3409.468, 2121.299, 1508.151, 989.2469, 766.4855, 749.4873, 491.5999, 
    500.2154, 587.9318, 432.9168, 407.4583, 403.593, 373.3047, 314.6314, 
    310.2964, 287.6699, 288.7629,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 137.5109, 1.268968, 0, 0, 0, 0, 0, 0, 0.1147682, 82.57735, 311.5683, 
    151.4449, 78.04676, 128.0494, 376.5229, 522.9591, 427.1115, 256.4601, 
    112.6585, 142.7851, 266.511, 196.9078, 88.25249, 66.20465, 58.85111, 
    66.82548, 83.11908, 91.31876, 101.4318, 105.2445, 110.9949, 121.9766, 
    145.8439, 152.8409, 158.7673, 160.5151, 158.0549, 151.2477, 147.5351, 
    168.9152, 567.9518, 1848.487, 3247.352, 3623.287, 3933.537, 4026.396, 
    3815.863, 3989.005, 4117.667, 4075.111, 3740.598, 3347.181, 3151.984, 
    2783.441, 1733.658, 1189.891, 689.3563, 352.485, 479.9682, 518.3051, 
    654.5156, 843.5643, 637.5115, 436.4144, 356.3743, 315.6976, 287.2369, 
    264.154, 245.379, 203.1721,
  0, 0, 0, 0, 0, 0, 0, 0, 0.0005155665, 0.00535053, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 5.954806, 0.008552877, 0, 0, 0, 0, 0, 0, 0, 
    1.392343, 147.5822, 117.1248, 79.08617, 161.021, 478.1805, 672.9123, 
    747.8989, 659.3046, 435.462, 300.6021, 411.5335, 261.7856, 93.77441, 
    56.53286, 59.12653, 61.15051, 76.3445, 85.60712, 87.65303, 86.02962, 
    90.52665, 104.9385, 125.5316, 141.8028, 161.3927, 151.9469, 148.933, 
    141.536, 144.3197, 149.6154, 172.0073, 623.9898, 1684.723, 2641.521, 
    3090.655, 3319.659, 3217.01, 3316.014, 3452.869, 3067.782, 2450.786, 
    1764.937, 1428.371, 1315.265, 759.3845, 608.1971, 375.0185, 229.107, 
    391.8174, 639.2117, 819.7453, 915.3849, 607.8117, 379.9553, 305.7845, 
    306.8441, 298.1168, 286.4967, 240.3828, 184.6151,
  0, 0, 0, 0, 0, 0, 0, 0, 0.121945, 0.03938331, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.3118506, 3.291815, 0.01598853, 0, 0, 0, 0, 0, 0.1340173, 
    4.044582, 143.5697, 233.638, 191.9344, 118.6989, 147.4646, 285.2692, 
    535.5562, 720.2246, 908.1365, 672.2578, 505.0814, 365.3874, 130.3261, 
    44.65852, 61.89712, 58.099, 59.19082, 61.83461, 73.12101, 69.1452, 
    71.91867, 79.77286, 88.05507, 108.2875, 147.0296, 195.7139, 207.4643, 
    157.7728, 145.7407, 144.7948, 163.3843, 160.5329, 192.4493, 810.9302, 
    1566.056, 2149.559, 2256.098, 2102.709, 1810.442, 1541.477, 1113.111, 
    754.5137, 622.1283, 649.4427, 513.0068, 210.115, 259.1717, 228.6151, 
    216.1971, 473.4304, 783.3362, 789.3256, 686.4561, 419.5589, 249.4682, 
    205.099, 202.2573, 216.5917, 217.1671, 199.7617, 132.155,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.005494107, 0.4346767, 0, 0, 0, 0, 0, 0, 0, 9.391527, 298.571, 237.2993, 
    140.6926, 155.2257, 256.6727, 406.4414, 433.8806, 600.3461, 683.2579, 
    620.795, 483.5708, 265.2493, 69.42221, 44.01501, 51.81279, 60.87005, 
    53.39784, 52.44471, 56.40654, 59.58292, 67.88076, 74.34882, 81.33792, 
    95.65347, 148.0806, 236.6955, 255.9585, 205.559, 151.0034, 159.6844, 
    176.646, 199.4624, 204.3659, 270.1312, 848.1915, 1003.153, 1148.617, 
    1003.102, 887.6286, 594.8246, 321.8112, 230.0089, 347.2778, 260.032, 
    255.0762, 190.1423, 159.5509, 136.5862, 182.9312, 271.9562, 310.1284, 
    283.9276, 277.2419, 213.3407, 155.9381, 136.6259, 129.9663, 124.8657, 
    144.5141, 150.6962, 106.1049,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.2010026, 5.480222, 1.905644, 0, 0, 0, 0, 0, 0, 10.41574, 79.70645, 
    33.17719, 101.7773, 211.8761, 328.2486, 519.1068, 687.5656, 568.6201, 
    426.9638, 407.4171, 258.6449, 133.8155, 46.44923, 40.82528, 43.58858, 
    52.29549, 51.97647, 43.10914, 47.15418, 57.30152, 61.27217, 67.14295, 
    78.3484, 97.84009, 141.1024, 209.3585, 245.7221, 223.8985, 178.6274, 
    164.8928, 205.0671, 272.722, 329.3512, 281.3043, 329.6042, 396.7708, 
    453.139, 536.9029, 418.7523, 345.6891, 235.4872, 214.9491, 197.1605, 
    217.0889, 210.202, 187.8262, 155.8819, 114.6811, 108.0696, 103.5813, 
    75.537, 103.2833, 131.8954, 130.8562, 121.067, 118.0025, 105.5169, 
    96.54052, 119.8245, 176.6302, 195.5793,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 1.086443, 9.708963, 25.8066, 0, 0, 0, 0.6762983, 7.368328, 15.26273, 
    7.240432, 15.79535, 109.3353, 221.0537, 269.0515, 704.3265, 939.6818, 
    701.0948, 330.6563, 190.7539, 178.3714, 105.7215, 59.61247, 39.14966, 
    45.20544, 46.21466, 48.67001, 35.86091, 46.08049, 52.98456, 62.92745, 
    69.35141, 85.43824, 110.8834, 142.6441, 180.2906, 238.7265, 252.6595, 
    239.7324, 184.5832, 228.8213, 276.7168, 392.7193, 388.6469, 296.1601, 
    280.3641, 341.4388, 353.615, 317.2159, 244.4351, 223.8407, 201.6992, 
    183.6967, 176.9333, 172.614, 165.7017, 145.3332, 110.9088, 80.85966, 
    70.93066, 76.48385, 91.80798, 97.15785, 91.67457, 100.7875, 107.6938, 
    96.9532, 86.08794, 101.3551, 185.22, 281.0552,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 2.485921, 26.4163, 34.1476, 13.50462, 14.0831, 0.4166287, 2.192102, 
    29.53002, 14.33252, 3.286679, 52.2133, 156.3645, 257.6373, 649.4648, 
    1054.655, 614.7567, 162.2067, 99.85813, 116.9508, 77.15819, 48.32669, 
    64.66377, 56.2935, 65.67332, 46.97363, 33.90272, 37.93755, 51.28942, 
    58.10233, 78.93856, 106.3503, 116.9305, 149.4504, 180.898, 213.7403, 
    292.1611, 291.1207, 281.1519, 252.0287, 285.7556, 316.2794, 374.6313, 
    325.8148, 322.2468, 325.9581, 276.3282, 228.0858, 195.2241, 187.3171, 
    175.7014, 163.5601, 151.0618, 141.3108, 129.977, 114.84, 86.42167, 
    68.05943, 63.20282, 64.60545, 60.11647, 42.99261, 50.01132, 55.99592, 
    74.10268, 81.50942, 73.58952, 83.45282, 127.7083, 226.8334,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 2.984597, 0.01858864, 0, 0.0009470581, 16.01784, 
    87.35822, 173.5935, 488.2748, 759.5725, 523.7241, 141.7197, 113.1382, 
    159.5228, 147.7596, 115.4366, 107.1132, 102.7932, 85.72213, 66.42902, 
    30.98574, 37.11678, 45.43555, 64.23547, 99.53561, 129.9766, 138.2153, 
    142.8759, 176.7178, 267.0287, 349.3065, 417.0574, 373.9982, 391.8378, 
    306.8354, 254.5319, 312.5648, 296.5179, 377.6109, 330.0472, 242.8435, 
    164.2536, 149.3302, 147.9863, 144.5899, 139.069, 133.0572, 122.3601, 
    110.4266, 95.19322, 77.43336, 63.58871, 58.07784, 51.05425, 36.38617, 
    36.80247, 46.6338, 42.84441, 35.56261, 47.46378, 56.36189, 58.939, 
    105.9327, 189.9787,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 5.923116, 0, 0, 0, 0, 0, 6.078897, 54.77836, 77.55535, 
    204.2334, 410.9161, 330.8391, 185.1925, 194.0988, 249.267, 253.3829, 
    177.0466, 158.8476, 113.1643, 101.53, 68.00449, 31.76886, 36.63785, 
    58.77195, 90.80497, 133.0862, 161.9473, 164.7115, 165.2141, 201.0824, 
    279.0718, 359.1356, 398.5262, 459.7346, 501.9608, 511.8822, 352.2849, 
    246.1968, 246.5588, 279.2735, 323.1726, 191.8587, 143.4464, 112.1324, 
    117.9595, 116.5617, 114.9787, 113.5484, 107.3903, 97.09441, 84.3097, 
    70.09772, 57.50354, 51.82816, 43.33216, 40.77794, 45.42603, 66.79871, 
    45.82823, 21.87241, 20.00079, 29.68418, 34.1625, 55.23173, 131.1202,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.007114115, 12.30466, 48.17017, 
    51.3419, 136.4395, 140.1926, 152.5834, 214.4402, 290.774, 334.6097, 
    242.1319, 179.8538, 138.1877, 94.74007, 53.06939, 31.48326, 46.89961, 
    89.87615, 131.2574, 140.4565, 168.6543, 171.5402, 207.168, 234.0502, 
    297.8369, 300.6861, 321.7401, 399.447, 557.8159, 602.8211, 392.1693, 
    231.2913, 117.9363, 190.2211, 228.4644, 181.8213, 100.4968, 90.92713, 
    91.9957, 95.57886, 98.97549, 93.66434, 91.03915, 82.98544, 72.89633, 
    60.49364, 58.69539, 60.83919, 60.2387, 64.67129, 64.97378, 60.37475, 
    50.22374, 26.93556, 10.59541, 21.63067, 16.65605, 21.7373, 41.34349,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5.366938, 28.12142, 64.29294, 
    128.7759, 176.1391, 224.7735, 297.6988, 326.8529, 254.3473, 185.0925, 
    128.5998, 87.42819, 38.13975, 29.44325, 68.62458, 118.0892, 143.8512, 
    173.974, 164.9058, 204.4256, 210.1949, 267.1867, 300.9321, 309.5306, 
    297.9662, 355.8887, 461.3635, 509.2478, 310.7938, 206.6006, 123.8932, 
    125.1484, 178.9654, 129.2888, 94.40868, 92.13621, 118.3059, 139.3436, 
    102.2285, 87.8205, 78.24416, 72.41794, 72.99378, 69.93626, 64.41702, 
    66.0837, 67.51834, 70.63937, 64.17177, 65.43086, 61.57732, 57.59845, 
    48.39719, 66.22498, 19.65588, 7.979198, 7.954746,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1979136, 16.10868, 94.42965, 
    187.4814, 245.3877, 271.5805, 257.391, 297.2609, 210.7862, 164.771, 
    95.62947, 56.90887, 40.72773, 52.8884, 92.41105, 126.1473, 166.0383, 
    207.8445, 272.0114, 271.0105, 294.9529, 248.3746, 307.0643, 316.8501, 
    327.4612, 325.9547, 386.9184, 403.7983, 311.1118, 240.8184, 164.2083, 
    103.1077, 117.4106, 99.13666, 106.3574, 154.6648, 260.3508, 285.6964, 
    234.8461, 154.5512, 112.9279, 100.7134, 123.8555, 127.3378, 90.11683, 
    76.42348, 68.03311, 66.51344, 75.3875, 112.4858, 142.2936, 124.5137, 
    93.33791, 99.31126, 54.70262, 4.06266, 0.262289,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.04155033, 10.73219, 79.11258, 
    190.445, 274.9487, 342.6148, 355.8712, 312.3603, 292.6754, 221.7762, 
    115.474, 47.77611, 50.80471, 84.23752, 95.56871, 148.4016, 177.4802, 
    241.8285, 273.5516, 339.5761, 337.356, 326.2194, 277.1494, 336.4698, 
    352.6033, 363.4337, 382.938, 416.9631, 325.3823, 303.8384, 203.988, 
    116.0254, 110.5155, 121.6094, 106.5421, 137.3756, 210.812, 317.8851, 
    344.7708, 323.2015, 252.112, 193.5985, 213.3652, 191.4196, 156.1301, 
    106.2765, 104.4049, 72.89532, 100.3581, 157.0007, 215.9135, 191.733, 
    119.1055, 115.4301, 99.49779, 31.93542, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.542466, 22.26523, 77.77408, 
    140.4331, 240.0608, 343.6068, 376.1221, 378.217, 372.9897, 356.2578, 
    217.9453, 48.16224, 56.58264, 94.03797, 155.6086, 206.1189, 244.8234, 
    262.5258, 267.4071, 294.3894, 384.4132, 383.2951, 330.3748, 318.6039, 
    351.7903, 366.8914, 400.56, 447.5571, 438.7595, 508.2295, 383.2372, 
    246.7716, 200.7712, 148.0255, 184.6252, 228.8072, 293.0768, 384.8521, 
    451.6723, 470.1341, 383.5, 297.7384, 261.2184, 257.7826, 233.8021, 
    230.1151, 168.3038, 140.5308, 159.7929, 141.3796, 184.5563, 169.6956, 
    127.2488, 153.812, 157.5335, 129.1637, 8.482048 ;

 land_mask =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0.2418439, 0, 0.1507849, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0.9672335, 0.7867691, 0.8897236, 0.7868192, 0.4295904, 0.103123, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 0.8583792, 0.24312, 0.02330228, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 0.7519304, 0.3075978, 0.05466554, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 0.7495267, 0.07681742, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.8367906, 0.08314215, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.341669, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9609066, 0.3417271, 0.0006489863, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.6232235, 0.1494775, 0.0620707, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.8576373, 0.4441393, 
    0.02198116, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9266944, 0.7165388, 0.8939224, 
    0.5627504, 0.03366798, 0.3162485, 0.02661187, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9785867, 0.3546079, 
    0.001069293, 0.5276027, 0.6956339, 0.8771922, 0.3122943, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.6351135, 0.1552348, 
    0.2120383, 0.6413907, 0.72313, 0.05286491, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.4744368, 
    0.01789349, 0.362444, 0.7183179, 0.6351389, 0.2321099, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.537541, 
    0.02737221, 0.1637618, 0.5896915, 0.6713976, 0.06366118, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.5861796, 
    0.0982726, 0.02536981, 0.1802837, 0.5701141, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.8579165, 
    0.275193, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.91327, 
    0.2402546, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.918274, 0.5621569, 0.0209811, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.588654, 0.3020536, 0.30206, 0.2020797, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 0.9413478, 0.1002747, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 0.6651581, 0.001533675, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 0.3886248, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 0.6325621, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 0.995119, 0.2749188, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 0.6972129, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.9737231, 0.9926948, 1, 1, 1, 1, 0.8642177, 0.08541915, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9564105, 
    0.4497338, 0.407091, 0.4070948, 0.4070986, 0.4071023, 0.2621634, 
    0.3688191, 0.6872182, 0.9677767, 1, 1, 1, 0.4953253, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.2941011, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.2652708, 0.8491837, 1, 1, 0.4804461, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.648157, 0.03258629, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0.4520298, 1, 1, 0.3871183, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9116583, 0.07233045, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1828122, 1, 1, 0.1171441, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.553419, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.08816408, 1, 1, 0.7507677, 0.04885805, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.6228713, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.3365233, 1, 1, 1, 0.5879625, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9385124, 0.1065637, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0.2791502, 0.6271809, 1, 1, 1, 0.9890413, 
    0.2517519, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1216078, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.6900454, 0.06213602, 
    0, 0, 0, 0, 0, 0, 0, 0.1037045, 0.7385923, 0.9886956, 1, 1, 1, 1, 1, 
    0.4103255, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.908018, 0.1728964, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.3633319, 1, 1, 1, 1, 1, 1, 1, 0.7623217, 
    0.0008263012, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.6658352, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.4360288, 0.957324, 0.635229, 0.4226641, 0.2175488, 
    0.3202175, 0.8472205, 1, 0.9694546, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.5564398, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.2841633, 0.1100108, 0, 0, 0, 0, 0.8772225, 1, 0.9926439, 
    0.7188581, 0.01636519, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.6282753, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.9419357, 1, 1, 1, 0.5849457, 0.315834, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9848972, 0.2503584, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01595704, 0.995867, 1, 1, 1, 1, 
    0.9787351, 0.2506236, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.6914676, 0.02198116, 0, 
    0, 0, 0, 0, 0, 0.08334821, 0.1012918, 0, 0, 0, 0, 0, 0.005334743, 
    0.7088248, 1, 1, 1, 0.8540698, 0.9996781, 0.6620048, 0.03839629, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9575872, 0.6579381, 
    0.3669165, 0, 0, 0, 0, 0, 0.5810857, 0.3034903, 0, 0, 0, 0, 0, 0, 
    0.07322878, 0.3065482, 0.1025856, 0.1025909, 0.06481452, 0.2606909, 
    0.8556811, 0.4936866, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9884753, 0.8030674, 
    0.2831464, 0, 0, 0, 0.4692461, 0.05008297, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.2312002, 0.6806778, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.8807496, 0.4964221, 0.118718, 
    0.2605629, 0.7617009, 1, 1, 0.9638987, 0.2762473, 0, 0.01970084, 
    0.866532, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.03466008, 0.9590737, 
    0.3642623, 0, 0, 0, 0, 0, 0, 0, 0.03183588, 0.3728453, 0.1801692, 
    0.07776905, 0.3728562, 0.2684634, 0.07811955, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.825218, 0.1281082, 0, 0, 0, 
    0.05450449, 0.1359098, 0.6320257, 0.6364659, 0.07199212, 0, 0.07605698, 
    0.7873569, 0.08185559, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.5112837, 
    0.5608108, 0.3629351, 0, 0, 0, 0, 0, 0, 0.3923621, 0.8759633, 1, 
    0.9305333, 0.6235623, 1, 0.9620325, 0.6514717, 0.1631414, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.7229308, 0.07197631, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.8089566, 0.1385804, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.718082, 0.0345762, 0, 0, 0, 0, 0, 0, 0.3329219, 0.987651, 1, 1, 1, 1, 
    1, 1, 1, 0.9168873, 0.5666844, 0.05440859, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.8832299, 0.1472945, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.4424467, 0.1988707, 0.007988392, 0.4272325, 0.7964597, 0.1058136, 0, 
    0.1016413, 0.03233812, 0, 0, 0, 0, 0, 0, 0, 0, 0.4837731, 0.6387944, 
    0.2020133, 0, 0, 0, 0.0193575, 0.5679138, 0.9483995, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 0.8473101, 0.6221716, 0.1199134, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9533704, 0.1238984, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.1078062, 4.039702e-05, 0.02094627, 0.7635151, 0.6279824, 0, 
    0.4214649, 0.03240846, 0, 0, 0, 0, 0, 0, 0, 0, 0.1298708, 0.9593522, 
    0.8726715, 0.6254805, 0.6615382, 0.6156211, 0.7938948, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 0.8723933, 0.576844, 0.1146775, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  1, 1, 1, 0.9439595, 0.8502378, 0.4763551, 0.4259781, 0.7869197, 0.754113, 
    0.2165837, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.483312, 
    0.5854645, 0, 0.1202012, 0, 0, 0, 0, 0, 0, 0, 0, 0.01637845, 0.6564068, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.859898, 0.7360823, 0.2172089, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 0.6529251, 0.507857, 0.3280367, 0.03502538, 0, 0.1547292, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1886325, 0.4330523, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.4363211, 0.7168808, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.8921524, 0.3981088, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0,
  1, 0.9714789, 0.9004541, 0.4634776, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0.05552825, 0.120399, 0.03792001, 0.00843242, 0, 
    0, 0, 0, 0, 0, 0.07417351, 0.8822758, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.8686383, 0.1390514, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.01985216, 0.09956025, 0.09957455,
  0.9850286, 0.5513424, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.01466178, 0.4497637, 0.01945193, 0, 0, 0, 0, 0, 0, 
    0.2087137, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 0.7150637, 0.00703513, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01038911, 0.03078478, 0.5223621, 
    0.5656272, 0.5656678, 0.6186966, 1, 0.975225,
  0.5147771, 0.2509983, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.01205661, 0.5400833, 0.6323332, 0, 0, 0, 0, 0, 0, 
    0.0640404, 0.8329736, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.5314379, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.06310866, 0.6251156, 1, 1, 1, 1, 1, 
    1, 1,
  0.04331701, 0.004251128, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.7602282, 0.9885215, 0.1360401, 0, 0, 0, 0, 0, 
    0.5068112, 0.1770562, 0.9897748, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9330676, 0.3697935, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.2310756, 0.410401, 0.4104408, 
    0.4104811, 0.4105217, 0.4105628, 0.6770073, 0.9558303, 1, 1, 1, 1, 1, 1, 
    1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.003479148, 0.9392874, 0.5581517, 0.007009166, 0, 0, 0, 0, 0, 0.1731326, 
    0.4696587, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9879944, 0.3274225, 0.317915, 
    0.008586753, 0.1531166, 0.007366235, 0.3192428, 0.3195822, 0.3196146, 
    0.3196478, 0.3314601, 0.8600246, 0.8667862, 0.9326418, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.01336217, 0.6549731, 0.145487, 0, 0, 0, 0, 0, 0, 0.1268012, 0.9062009, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.7842681, 0.8845835, 0.7709545, 0.9917373, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.4637389, 0.1322377, 0, 0, 0, 0, 0, 0, 0.03724731, 0.7512087, 
    0.9969589, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.03823176, 0.9980064, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.1325942, 0.07740931, 0, 0, 0, 0, 0, 0, 0, 0.1540521, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.3038891, 0.04776999, 0, 0, 0, 0, 0, 0, 0, 0.1829891, 0.9730953, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.03913443, 0.0341659, 0, 0, 0, 0, 0, 0, 0, 0, 0.009582857, 0.9771051, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.1451908, 0.07445376, 0, 0, 0, 0, 0, 0, 0, 0, 0.3511962, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0.3498454, 0.9953002, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0.2403926, 0.9019648, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.005788924, 0.01535262, 0, 0, 0, 0, 0, 0.1437764, 0.2917262, 
    0.9888229, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.1149602, 0.1676279, 0, 0, 0, 0, 0, 0.2839805, 0.2067913, 
    0.6178907, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1299978, 0.9375334, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.5485037, 0.9940798, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.4170257, 0.986974, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.8614578, 0.9180768, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0009119348, 0.393558, 0.9921986, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 0.9273752, 0.1889167, 0.7825502, 0.8380716,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0002601096, 0.8132703, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 0.6767043, 0.05085213, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.04240416, 0.8030222, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 0.8947946, 0.0665093,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.2244188, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.5003253 ;

 zsurf =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01534718, 
    0.004565009, 0.008999515, 0.009599131, 0.0008479413, 0, 0, 0.0007195598, 
    0.004574103, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.7068716, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.003399682, 
    0.0147934, 0.002706561, 0, 0, 0, 0.004826599, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.004755895, 
    0.00314351, 0.002793752, 0, 0, 0, 0.006179405, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.006290677, 
    0.007201957, 0, 0.01463142, 0.003162183, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.008779748, 0, 0, 0, 
    0.00300725, 0.002690252, 0.005241457, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 1.506357, 3.305288, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.007343553, 0, 0.009825814, 0.01535672, 0.006712195, 0, 0, 0.005644962, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19.68891, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.008339305, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.00178691, 18.51452, 0.01244308, 0, 0, 0, 
    0, 0.009080717, 0, 0, 0, 0, 0.006611669, 0.003060021, 0.008406991, 0, 
    0.005074322, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01017599, 
    0, 0, 0, 0.004030156, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.003469607, 0, 0, 0, 0, 0, 0.002995649, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.004560474, 0, 0, 0.01124365, 0.003597797, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.01154227, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.2431989, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.001374771, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.06463672, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.1425494, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  33.14798, 0, 34.79201, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.0004971988, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  668.3605, 750.8135, 625.5392, 386.1679, 158.3386, 2.453814, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1070.732, 1178.2, 1004.681, 772.6516, 403.6846, 150.0447, 26.30301, 
    1.64736, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1507.715, 1421.274, 1144.302, 833.4024, 441.414, 72.99273, 109.9673, 
    184.5779, 220.3756, 0.00647221, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1551.811, 1623.509, 1564.146, 1482.56, 1154.821, 803.4989, 487.0388, 
    202.9149, 268.4435, 226.8269, 46.07853, 0.3954178, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0,
  1557.897, 1671.874, 1696.626, 1635.232, 1700.021, 1734.235, 1559.076, 
    995.3284, 449.7531, 276.2559, 565.8065, 21.12218, 0.8193069, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1468.874, 1600.571, 1614.583, 1414.91, 1396.924, 1757.31, 2173.984, 
    2018.616, 1396.95, 1025.211, 762.0422, 232.5291, 8.014444, 1.140886, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0,
  1326.019, 1541.283, 1555.617, 1480.098, 1514.677, 1689.735, 1982.568, 
    2007.651, 1670.599, 1186.88, 1048.513, 684.1181, 117.3529, 0.1669138, 0, 
    0, 0, 14.15248, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1146.4, 1447.466, 1700.664, 1654.412, 1747.869, 2042.93, 1975.362, 
    1731.381, 1260.238, 1003.032, 874.1664, 965.1847, 711.4643, 390.3766, 
    173.5833, 3.412067, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1373.781, 1329.12, 1740.19, 1867.481, 1919.821, 2046.155, 2020.59, 
    1730.883, 1388.832, 990.3948, 863.0721, 733.3089, 488.1863, 444.3896, 
    642.3708, 630.8365, 208.2363, 11.2473, 0.03753853, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1914.861, 1386.722, 1730.161, 1876.041, 1894.845, 2047.599, 1965.026, 
    1787.49, 1283.865, 1007.386, 831.1433, 589.1078, 291.1984, 130.3001, 
    245.2175, 308.7728, 423.5323, 287.8249, 17.96172, 32.98395, 0.1041703, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.1970985, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  2061.196, 1476.068, 1648.332, 1574.314, 1569.191, 1744.371, 1828.933, 
    1790.968, 1558.644, 1149.688, 1213.996, 906.5831, 504.1509, 233.0578, 
    183.2224, 38.9668, 0.0118664, 233.6236, 272.1967, 144.2618, 56.46022, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  1840.156, 1504.441, 1582.167, 1490.926, 1402.836, 1518.827, 1694.572, 
    2058.519, 1824.339, 1671.718, 1643.01, 1482.167, 815.0604, 396.3656, 
    379.8361, 318.8223, 100.745, 65.86816, 107.3457, 244.7698, 250.1199, 
    15.35586, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0,
  1837.63, 1728.632, 1902.097, 1719.298, 1875.763, 1918.201, 2012.239, 
    2196.799, 2065.854, 1799.648, 1839.158, 1689.026, 1220.946, 556.4898, 
    653.7017, 762.9083, 615.2339, 393.6399, 83.12075, 4.564439, 169.0518, 
    231.0936, 86.59752, 8.810427, 0, 0, 0, 0, 0.004199471, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  2287.553, 2375.422, 2227.182, 2205.671, 2448.729, 2173.713, 2069.91, 
    1804.564, 1718.86, 1645.912, 1760.087, 1774.775, 1588.443, 1158.239, 
    1042.855, 1238.964, 1055.679, 720.4163, 300.8953, 74.61289, 2.083953, 
    10.21264, 134.772, 93.68505, 9.525565, 0, 0, 0, 0.06281511, 3.428892, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  2614.957, 2546.323, 2390.928, 2148.965, 2257.577, 2052.22, 1766.787, 
    1770.134, 1673.074, 1765.732, 1825.648, 1895.919, 1992.829, 1695.072, 
    1362.996, 1422.211, 1302.389, 1040.16, 627.5578, 400.1667, 51.56722, 
    2.257818, 0.1849899, 56.72547, 250.1037, 1.460486, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.967957, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1897.78, 2076.201, 2129.073, 2115.72, 2166.538, 1872.045, 2072.919, 
    1904.649, 2256.727, 1803.393, 1983.677, 2108.663, 2195.764, 2050.119, 
    1605.954, 1432.204, 1511.048, 1487.268, 1426.227, 1196.583, 721.2061, 
    185.3391, 24.12744, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0004704067, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.2958491, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1716.921, 1748.802, 1939.11, 2058.646, 2214.479, 2215.264, 2299.508, 
    2683.908, 2679.552, 2308.606, 2102.935, 2086.155, 2177.915, 2051.186, 
    1598.307, 1383.17, 1438.509, 1773.132, 2076.03, 2118.625, 1700.985, 
    1170.254, 459.9845, 48.66238, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1594.9, 1717.709, 1846.341, 2183, 2416.479, 2646.638, 2920.714, 2901.701, 
    3107.744, 2624.682, 2306.014, 2028.034, 1806.9, 1723.413, 1505.019, 
    1253.708, 1291.276, 1617.983, 1898.304, 2037.906, 2075.454, 2108.36, 
    1570.701, 841.1761, 129.8114, 0.2389687, 3.660637, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1414.581, 1499.586, 1735.549, 1988.982, 2430.141, 2544.231, 2714.589, 
    2826.258, 2566.761, 2620.082, 2419.738, 2052.477, 1891.764, 1767.929, 
    1617.863, 1432.407, 1338.126, 1367.179, 1424.379, 1473.549, 1661.907, 
    2049.929, 2230.574, 1919.274, 1373.336, 316.5095, 39.45748, 94.61289, 
    39.49365, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    7.207365e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1235.553, 1437.662, 1381.895, 1611.005, 1679.951, 1728.312, 1922.424, 
    1964.016, 1953.016, 2112.162, 2098.977, 1710.801, 1526.079, 1414.803, 
    1368.911, 1237.472, 1292.035, 1341.555, 1204.039, 1329.621, 1429.259, 
    1572.953, 1800.086, 2189.089, 2119.821, 1455.417, 1083.626, 1022.557, 
    862.4561, 51.87525, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1174.93, 1228.427, 1291.553, 1290.888, 1424, 1351.69, 1468.16, 1589.555, 
    1427.788, 1689.11, 1630.9, 1414.054, 1334.024, 1248.547, 1122.594, 
    1033.518, 1091.201, 1192.766, 1168.232, 1309.946, 1314.83, 1245.706, 
    1400.043, 1858.552, 2194.833, 2118.342, 1668, 1707.535, 1364.425, 
    595.4224, 15.76594, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  823.5144, 966.8268, 1033.309, 1192.71, 1210.489, 1193.993, 1280.92, 
    1308.805, 1209.215, 1289.174, 1294.622, 1176.932, 1193.732, 1146.91, 
    1025.355, 875.7115, 882.8735, 978.463, 1033.714, 1232.486, 1255.239, 
    1216.565, 1342.363, 1716.272, 2074.805, 2120.552, 2071.005, 1786.363, 
    1785.419, 844.6271, 169.2518, 0.001837272, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  661.3832, 741.7489, 952.168, 1073.759, 1053.268, 1013.894, 1031.548, 
    1062.557, 1014.31, 1013.214, 1007.304, 1006.718, 987.2679, 929.3942, 
    846.1819, 807.7843, 729.1191, 717.0919, 644.5469, 733.0809, 815.4983, 
    1055.672, 1469.535, 1941.911, 2045.901, 2101.024, 2062.683, 2086.129, 
    1883.878, 989.241, 529.9884, 1.092551, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0,
  574.1776, 618.1168, 795.5441, 907.0357, 894.5935, 851.0385, 820.7712, 
    843.4498, 837.6264, 813.8089, 821.1804, 790.303, 694.8225, 637.4512, 
    626.2227, 661.035, 688.275, 597.9715, 427.0944, 299.6628, 342.4961, 
    676.9834, 1214.729, 1706.491, 1881.969, 1649.495, 1733.168, 2044.59, 
    2105.82, 1415.646, 915.3256, 166.6185, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0,
  503.9159, 538.9011, 631.793, 737.8944, 750.1324, 703.1216, 655.9878, 
    654.8143, 672.593, 642.7423, 621.7355, 602.098, 473.79, 425.5311, 
    461.755, 530.6566, 568.3069, 558.3639, 330.7892, 179.9599, 143.326, 
    168.8803, 392.449, 875.6781, 1042.997, 940.2807, 1005.778, 1682.482, 
    2467.645, 1832.106, 1341.977, 441.4869, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0,
  453.9662, 441.7195, 504.0019, 592.8539, 608.1069, 578.1291, 526.2635, 
    513.4938, 532.1535, 479.4901, 447.4254, 444.3315, 379.7191, 325.8571, 
    347.1577, 396.39, 397.7914, 382.2119, 225.9507, 114.7197, 95.74188, 
    70.67721, 57.3841, 157.933, 314.682, 123.271, 156.6136, 1009.174, 
    2106.859, 2219.086, 1513.035, 924.8544, 29.27477, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  503.6515, 465.5753, 433.9768, 478.4191, 482.0991, 473.893, 436.3061, 
    425.1155, 431.4804, 382.6123, 325.8517, 340.3661, 314.822, 260.5178, 
    239.2539, 233.0164, 209.3085, 185.2675, 99.46118, 35.69082, 15.04999, 
    5.81494, 7.321244, 7.285094, 10.49513, 6.034019, 12.30279, 178.9217, 
    1494.86, 1747.576, 1843.446, 1614.362, 380.1558, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  438.2668, 471.7402, 408.1164, 400.8929, 380.3304, 374.7529, 382.5601, 
    372.2382, 382.916, 320.6809, 264.4974, 252.2818, 258.8326, 194.5873, 
    162.8055, 141.8769, 114.3217, 85.31949, 39.80796, 4.830305, 0, 0, 0, 0, 
    0, 0, 0, 0.02132653, 176.2921, 430.069, 932.7458, 1392.24, 747.5593, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  375.052, 414.3507, 415.5859, 381.3595, 361.0887, 329.3397, 313.1617, 
    313.8601, 298.01, 280.3281, 250.9803, 220.6591, 244.4896, 157.4741, 
    126.7682, 118.9209, 91.80339, 46.5208, 11.15798, 0.09899135, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 50.89595, 153.9082, 606.8809, 122.0387, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0,
  304.4448, 364.8189, 357.5074, 352.7218, 337.0601, 318.3467, 277.0119, 
    265.5412, 282.2703, 328.1339, 341.168, 288.7758, 254.3146, 138.1611, 
    97.54157, 97.74657, 73.76514, 23.01658, 0.5496842, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 3.476873, 75.94135, 449.1298, 34.83492, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  306.857, 361.5244, 342.5269, 300.4066, 292.6741, 274.3279, 251.7741, 
    245.3346, 294.167, 380.9618, 372.6419, 271.2439, 204.3829, 99.51021, 
    69.604, 73.45421, 50.67704, 12.05578, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3.512501, 149.8454, 851.515, 526.5105, 5.040119, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  319.7339, 346.4661, 325.2934, 268.1579, 235.2851, 243.1511, 224.0061, 
    242.3429, 319.4263, 334.612, 274.955, 164.2817, 109.9028, 55.26638, 
    47.65622, 41.80495, 35.97699, 2.775469, 0.03288275, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 6.357764, 280.3884, 1031.42, 1222.137, 606.0325, 0.7514994, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.07952388, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  294.8905, 319.0948, 294.4915, 238.6062, 212.2333, 193.6535, 202.8654, 
    221.7048, 288.9077, 248.9493, 137.382, 84.58096, 51.21586, 40.6296, 
    44.39739, 63.04242, 40.62316, 8.783824, 0.268134, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.7404718, 15.12963, 65.80754, 738.6376, 1257.209, 1292.93, 64.7064, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13.92286, 118.2891, 0.07517834, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  313.3622, 298.425, 277.4745, 233.6075, 198.1856, 187.4898, 173.2009, 
    175.6373, 200.6465, 144.9214, 80.57291, 77.81576, 66.51388, 73.39558, 
    92.76784, 95.03912, 61.3536, 3.831983, 0.1158118, 0, 0, 0, 0, 0, 0, 0, 
    0.6463583, 18.92656, 71.69862, 132.442, 95.90388, 289.954, 763.129, 
    1148.201, 229.1096, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.065996, 
    17.50426, 2.459143, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  289.323, 276.3043, 265.5132, 220.7219, 216.1242, 195.0884, 181.3391, 
    143.4675, 147.2648, 111.0426, 110.6656, 125.9561, 122.3719, 105.6208, 
    113.7486, 98.84241, 43.68995, 0.9661562, 0.02680171, 0, 0, 0, 0, 0, 0, 0, 
    3.878528, 38.69389, 97.16181, 132.8956, 207.0652, 216.3446, 424.0393, 
    918.3037, 351.0448, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6.011113, 
    0.1137814, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  230.5823, 241.4872, 225.9881, 214.9098, 207.3458, 206.6044, 173.4783, 
    138.0395, 130.4559, 142.9235, 167.6159, 175.7432, 143.494, 103.3232, 
    73.60364, 63.91725, 27.10206, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10.20466, 
    20.16096, 25.27402, 21.63544, 14.64767, 43.60937, 331.3476, 893.1275, 
    454.1429, 1.288543, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  191.6571, 178.5321, 189.9285, 201.3738, 214.7888, 215.5745, 179.5497, 
    147.2228, 153.1658, 179.6961, 230.3224, 239.8835, 194.1318, 137.8888, 
    87.66043, 69.8594, 27.32165, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6.084438, 
    6.930506, 0.584422, 0.003764597, 0.003457344, 0.4655042, 543.0778, 
    932.6347, 615.3885, 85.28525, 0.2777186, 0, 0, 0, 0, 0, 0.422377, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0,
  231.2289, 207.4846, 224.9596, 237.2916, 248.9516, 252.8323, 212.7034, 
    195.5234, 197.4957, 263.0653, 303.2209, 280.5213, 264.7434, 194.2222, 
    116.7919, 78.11273, 25.05218, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    4.827813, 526.7432, 777.7427, 639.5916, 362.6419, 79.72997, 29.67748, 
    0.912546, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  278.9553, 267.2621, 269.6895, 261.4806, 287.7636, 281.252, 243.8186, 
    240.3938, 298.7545, 342.4502, 399.08, 363.9893, 266.6101, 221.5975, 
    126.7727, 76.75681, 26.75876, 0.9402217, 0, 0, 0, 0, 0, 0, 0, 0.3805751, 
    0, 0, 0, 0, 0, 3.231741, 309.7996, 351.9758, 387.7886, 218.6437, 153.275, 
    263.9878, 54.07672, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  241.8856, 246.4237, 245.6055, 259.1919, 286.3187, 285.9484, 254.3894, 
    280.3928, 369.3888, 439.415, 618.7897, 387.4653, 291.7344, 174.3447, 
    113.5729, 67.22175, 24.12755, 0, 0, 0, 0, 0, 0, 0, 20.0383, 16.96434, 0, 
    0, 0, 0, 0.003687347, 0.00572379, 52.21835, 70.8857, 55.61906, 70.92522, 
    123.4313, 420.684, 636.3296, 6.528507, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  202.4083, 219.8558, 207.086, 261.2129, 295.0167, 264.0109, 249.5903, 
    352.6951, 497.0891, 679.3617, 595.9517, 404.6982, 150.7021, 114.5868, 
    78.8996, 54.99938, 26.96955, 5.426031, 1.965392, 0.1738949, 0, 0, 0, 0, 
    39.73782, 6.958992, 0, 0, 0, 0, 0, 0.0001729098, 1.584328, 6.905681, 
    0.7596173, 0.490705, 0, 84.19572, 863.5649, 289.1957, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  210.9862, 176.5489, 218.8383, 299.7639, 293.6812, 247.376, 300.3907, 
    490.8528, 720.3207, 577.838, 503.2361, 148.1991, 107.7899, 63.81637, 
    42.55847, 31.07135, 27.5754, 28.17957, 28.8343, 16.63614, 2.660592, 0, 
    0.01031376, 0.9608897, 33.86351, 0.509288, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.05132846, 0, 0, 160.5816, 333.4066, 8.909275, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  247.1366, 214.9977, 272.471, 323.8452, 298.5703, 362.521, 537.7053, 
    668.5198, 624.8367, 453.5524, 165.6625, 102.4959, 57.48196, 21.7608, 
    4.573749, 1.787246, 5.738702, 13.79587, 21.61514, 15.3555, 7.805641, 
    1.753023, 0.05135195, 1.186182, 39.27137, 0.8040789, 0, 0.01927231, 
    0.09756799, 0, 0, 0, 0, 0, 0.1619276, 0, 0, 0, 9.406398, 314.6326, 
    92.01137, 0, 0, 0.001729056, 0, 0, 0, 0, 0.6381596, 31.72947, 4.45034, 
    6.862898, 161.6274, 35.41436, 10.87154, 0.005455857, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2.744836, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  229.433, 306.0153, 351.427, 376.3137, 463.0498, 627.9566, 686.7066, 
    565.6674, 405.129, 181.5926, 102.0433, 47.04384, 16.67009, 1.10613, 0, 0, 
    0, 0.09115441, 1.67472, 5.002741, 3.653378, 0.914476, 0.0004763628, 
    1.392298, 81.95518, 36.95679, 0, 0.102858, 0, 0, 0, 0, 0, 7.409501e-05, 
    0, 0, 0, 0, 55.38284, 97.32481, 47.17434, 0, 0, 0, 0, 0, 0.03468706, 
    60.15501, 130.7003, 244.7536, 135.677, 424.9022, 731.8262, 553.5016, 
    151.7469, 15.67891, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.1039039, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  298.4516, 455.0074, 496.0555, 490.0974, 549.4736, 625.2988, 487.0647, 
    277.1122, 157.1025, 104.1153, 47.97492, 9.955524, 1.711641, 0, 0, 0, 0, 
    0, 0, 0.08672119, 0.02051163, 0.0005947647, 0, 0.02029713, 58.99087, 
    18.83587, 0.0248516, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 110.5765, 3.497101, 
    0, 0, 0, 0, 0, 0.05597858, 47.99405, 655.0215, 1362.752, 1510.303, 
    1890.99, 1900.117, 1904.355, 1649.458, 1608.771, 1245.189, 378.5316, 
    4.13827, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 1.282194, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  430.407, 573.2601, 458.0574, 384.715, 322.2038, 270.0156, 169.9159, 
    89.97162, 81.54353, 47.91539, 13.97083, 0.9449826, 0, 0, 0, 0, 0, 0, 
    0.0004252571, 0.3309443, 0.03876647, 1.728635, 0.4185002, 0, 15.5728, 
    39.27885, 1.380751, 0.007368555, 55.84319, 1.191139, 0, 0, 0, 0, 0, 0, 0, 
    0, 115.976, 114.2675, 74.08803, 0, 0, 0, 0.3069585, 74.61648, 1023.105, 
    1976.442, 2391.624, 2180.577, 1604.411, 1326.77, 901.5997, 1351.656, 
    2254.224, 2631.384, 2637.751, 1822.456, 620.1605, 20.8799, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  430.7066, 471.0601, 333.3573, 224.1613, 108.1152, 65.5984, 26.94351, 
    37.64307, 24.10448, 10.83371, 1.795868, 0, 0, 0, 0, 0, 0, 0, 0, 0.421066, 
    0.211959, 0.211567, 0.4754283, 0, 1.457668, 49.35142, 77.70663, 0.225208, 
    177.6199, 27.2492, 0, 0, 0, 0, 0, 0, 0, 0, 16.10499, 144.5139, 247.1739, 
    155.9424, 68.87181, 112.7537, 548.5216, 1326.625, 1537.927, 1522.117, 
    1053.582, 538.7177, 494.4248, 237.3714, 225.9437, 723.8336, 1495.832, 
    2103.182, 2873.699, 3292.384, 3380.365, 2269.825, 515.0248, 4.337821, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0,
  431.9473, 396.6402, 222.4012, 114.462, 25.37888, 7.691118, 6.677791, 
    7.348661, 3.157577, 0.984972, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.3024256, 
    0.2389092, 0.1394803, 0.00746349, 0, 70.57438, 149.7564, 0, 80.11617, 
    0.0417327, 0, 0, 0, 0, 0, 0, 0, 0.01057512, 27.73273, 266.8832, 915.6628, 
    1100.12, 1117.166, 1315.549, 1758.784, 2041.483, 1431.61, 474.8531, 
    232.1502, 208.0247, 196.3371, 166.9769, 139.262, 189.603, 539.9, 
    636.6401, 1134.973, 2116.188, 3255.661, 3725.555, 3525.62, 2041.445, 
    414.1652, 93.96832, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  441.435, 319.8361, 136.8747, 29.58521, 4.141918, 2.825089, 0.08903898, 
    0.08046266, 0.2208437, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.3990609, 
    0.3265876, 0.0633444, 0.05431467, 84.71734, 149.596, 0, 0.04963135, 0, 0, 
    0, 0, 0, 0, 0, 27.05583, 59.55542, 2.632703, 383.2401, 1071.188, 
    1466.155, 1676.46, 1735.292, 1635.764, 1205.279, 587.2426, 204.6946, 
    192.8305, 201.6285, 192.1485, 173.3057, 135.0386, 115.5985, 154.6932, 
    207.6518, 252.7319, 408.4037, 1234.129, 2512.059, 3625.666, 3840.744, 
    2953.312, 1398.119, 200.1961, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  298.2758, 155.1034, 25.55248, 4.920603, 0.003125044, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1279996, 0.02609903, 0.3170911, 0, 23.67887, 
    68.64729, 35.86671, 72.66331, 0, 0, 0, 0, 0, 0, 27.26858, 361.5938, 
    62.6906, 207.8889, 270.3431, 466.9674, 991.8314, 1723.766, 1665.32, 
    1134.25, 697.3764, 239.1669, 204.7155, 192.0341, 177.9332, 167.6514, 
    147.1711, 124.0248, 116.1455, 138.7632, 205.803, 202.1669, 218.9659, 
    445.2673, 918.5952, 2052.283, 3110.208, 3814.63, 3245.299, 1978.916, 
    128.154, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.621783, 0, 0, 1.331606, 2.106077,
  156.3812, 18.64756, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.02620244, 0.1723592, 0.6139864, 0.7052164, 39.91206, 73.66648, 
    34.73109, 0, 0, 0, 0, 0, 0, 103.6746, 970.1916, 637.6611, 308.0594, 
    768.11, 1294.207, 1777.075, 1670.896, 1144.713, 449.2721, 228.4367, 
    250.4818, 226.3325, 198.0396, 169.848, 146.4091, 131.5473, 124.774, 
    133.6427, 162.3437, 232.3307, 229.8633, 231.2848, 277.8121, 478.211, 
    827.6024, 1960.805, 3358.45, 4059.359, 3432.779, 1310.91, 0.5703501, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11.00629, 
    172.8352, 183.9977, 46.27448, 129.1229, 178.4515, 97.62695,
  36.70903, 1.210476, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.226078, 0.04288947, 3.178066, 257.9394, 343.0803, 13.00084, 0, 
    0, 0, 0, 0, 2.137605, 96.99342, 646.0239, 147.4564, 527.7556, 1280.455, 
    1827.782, 1949.41, 1110.227, 192.4001, 183.5117, 228.3509, 244.9112, 
    227.8943, 192.5254, 159.7048, 137.4386, 124.2721, 122.957, 142.0076, 
    164.3923, 198.738, 229.3472, 259.537, 313.7084, 313.5366, 602.6287, 
    1546.649, 3188.223, 4339.325, 4235.496, 2657.681, 348.9787, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15.4312, 110.2107, 
    133.0185, 292.7062, 324.6068, 298.3218, 359.0092, 476.8519, 554.6548,
  1.995229, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.4212663, 0.04588909, 11.18899, 517.642, 542.4244, 51.31382, 0, 0, 0, 0, 
    0, 43.47145, 14.86237, 90.16446, 49.90094, 852.6797, 695.9244, 698.5693, 
    469.248, 149.1092, 136.4317, 196.3584, 211.3587, 231.4343, 214.1757, 
    171.0396, 141.9184, 127.4874, 119.4414, 115.9838, 130.7626, 159.6196, 
    192.4039, 226.2965, 268.5108, 312.2362, 358.5796, 389.9218, 1083.607, 
    2472.518, 4258.277, 4571.348, 3741.117, 2121.892, 269.5249, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 4.388186, 133.4869, 148.3846, 211.8387, 382.2953, 
    257.1787, 180.7228, 149.7092, 212.2956, 459.678, 761.8045, 1055.912, 
    1120.853, 1110.582, 1166.25, 1085.751, 1108.78,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.001913318, 33.17125, 520.3718, 399.8852, 0, 0, 0, 0, 0, 0, 0.8113799, 
    95.28371, 460.3841, 937.3494, 915.1066, 445.8253, 106.3576, 103.3282, 
    112.4795, 164.6748, 183.3819, 200.0266, 220.7052, 195.8168, 166.651, 
    121.4309, 123.9416, 113.4673, 102.3118, 125.9921, 156.5412, 179.7962, 
    206.3467, 238.4389, 260.7508, 315.1216, 328.1903, 360.6142, 1509.248, 
    3565.005, 4402.538, 4396.66, 3602.803, 2091.149, 261.0787, 82.22005, 
    0.2868135, 0, 0.5076911, 60.36261, 183.4623, 519.5708, 450.9728, 
    353.2507, 488.7053, 617.8168, 1421.896, 2045.6, 2299.798, 2328.442, 
    2164.863, 1835.325, 1553.868, 1649.168, 1826.316, 1985.27, 1961.338, 
    1556.79, 1371.403, 1288.084, 1040.601, 1072.717,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5.771062, 165.8212, 28.28846, 0, 0, 0, 0, 0, 0.1610673, 17.69787, 
    260.4066, 714.0234, 586.6948, 462.326, 79.98116, 88.8905, 101.472, 
    127.5234, 151.2906, 172.9191, 187.4914, 183.702, 173.0886, 139.7318, 
    124.8896, 118.3931, 105.5773, 109.4129, 131.1672, 156.9932, 163.0083, 
    184.8383, 204.416, 225.2426, 266.9706, 316.145, 224.5979, 381.9278, 
    2492.509, 3806.261, 4259.841, 4400.584, 3759.828, 2950.103, 2123.126, 
    1457.011, 1071.604, 1158.814, 1261.4, 1360.847, 1651.959, 2091.039, 
    2134.101, 2298.518, 2832.512, 3516.553, 3862.269, 3539.123, 3228.904, 
    3070.49, 3133.28, 3088.744, 2907.435, 2507.032, 2134.26, 1858.328, 
    1274.926, 962.0797, 842.9384, 710.9687, 939.0226,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 51.69876, 6.425387, 0, 0, 0, 0, 0, 0, 2.873953, 169.8395, 449.1624, 
    300.1902, 62.32654, 69.31486, 78.20786, 85.0916, 97.69564, 127.4337, 
    145.2199, 162.7987, 148.36, 126.3364, 126.9805, 112.7666, 113.0274, 
    97.65716, 107.4775, 138.243, 148.1546, 151.6598, 170.6716, 190.0256, 
    201.0505, 226.6755, 261.319, 232.2254, 219.3973, 932.7808, 2511.412, 
    3070.967, 3937.193, 4288.645, 4117.858, 3970.56, 3654.04, 3348.081, 
    3098.408, 2970.42, 2560.729, 2923.75, 3655.134, 3966.941, 4254.809, 
    4391.425, 4123.873, 3285.485, 2428.365, 1895.18, 1763.043, 1610.22, 
    1446.99, 1407.953, 1387.499, 1476.249, 1487.882, 1047.58, 652.7329, 
    528.4442, 542.4118, 917.0056,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.3669669, 0.3634669, 0, 0, 0, 0, 0, 0, 0.6933007, 13.2217, 484.2191, 
    144.2932, 49.07107, 47.2271, 55.1874, 111.1454, 210.9041, 104.5796, 
    116.9778, 131.3689, 115.879, 101.3334, 98.76527, 97.77927, 91.92683, 
    82.82296, 102.0775, 115.0132, 128.6879, 136.6141, 155.6852, 166.7384, 
    172.6179, 192.5376, 207.4939, 206.3573, 175.2231, 245.1321, 792.022, 
    1577.401, 2693.881, 3723.349, 4046.354, 3911.702, 3846.095, 3873.51, 
    4067.074, 4060.027, 3885.769, 3648.284, 4000.79, 4255.121, 4298.765, 
    3941.536, 2986.297, 2167.081, 1555.988, 1086.933, 981.1671, 671.5908, 
    517.9108, 560.5896, 604.6505, 737.5284, 838.4316, 663.5747, 487.8661, 
    405.7701, 432.4994, 598.6184,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 87.07624, 9.664433, 0, 0, 0, 0, 0, 0, 0.1396964, 165.1147, 498.7843, 
    209.5764, 50.07817, 49.66368, 196.0763, 442.8151, 358.6526, 227.8948, 
    104.9866, 105.646, 125.2638, 109.2299, 82.44156, 78.38992, 73.12806, 
    72.46248, 85.68304, 100.9489, 111.212, 121.0391, 131.6541, 139.9958, 
    153.3166, 166.8747, 176.9339, 177.9256, 166.0943, 164.8257, 217.7268, 
    390.218, 1575.724, 3050.704, 3828.212, 3839.21, 3919.247, 3790.678, 
    3970.27, 4419.288, 4398.239, 4177.742, 4184.263, 4184.499, 4041.16, 
    3409.468, 2121.299, 1508.151, 989.2469, 766.4855, 749.4873, 491.5999, 
    500.2154, 587.9318, 432.9168, 407.4583, 403.593, 373.3047, 314.6314, 
    310.2964, 287.6699, 288.7629,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 137.5109, 1.268968, 0, 0, 0, 0, 0, 0, 0.1147682, 82.57735, 311.5683, 
    151.4449, 78.04676, 128.0494, 376.5229, 522.9591, 427.1115, 256.4601, 
    112.6585, 142.7851, 266.511, 196.9078, 88.25249, 66.20465, 58.85111, 
    66.82548, 83.11908, 91.31876, 101.4318, 105.2445, 110.9949, 121.9766, 
    145.8439, 152.8409, 158.7673, 160.5151, 158.0549, 151.2477, 147.5351, 
    168.9152, 567.9518, 1848.487, 3247.352, 3623.287, 3933.537, 4026.396, 
    3815.863, 3989.005, 4117.667, 4075.111, 3740.598, 3347.181, 3151.984, 
    2783.441, 1733.658, 1189.891, 689.3563, 352.485, 479.9682, 518.3051, 
    654.5156, 843.5643, 637.5115, 436.4144, 356.3743, 315.6976, 287.2369, 
    264.154, 245.379, 203.1721,
  0, 0, 0, 0, 0, 0, 0, 0, 0.0005155665, 0.00535053, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 5.954806, 0.008552877, 0, 0, 0, 0, 0, 0, 0, 
    1.392343, 147.5822, 117.1248, 79.08617, 161.021, 478.1805, 672.9123, 
    747.8989, 659.3046, 435.462, 300.6021, 411.5335, 261.7856, 93.77441, 
    56.53286, 59.12653, 61.15051, 76.3445, 85.60712, 87.65303, 86.02962, 
    90.52665, 104.9385, 125.5316, 141.8028, 161.3927, 151.9469, 148.933, 
    141.536, 144.3197, 149.6154, 172.0073, 623.9898, 1684.723, 2641.521, 
    3090.655, 3319.659, 3217.01, 3316.014, 3452.869, 3067.782, 2450.786, 
    1764.937, 1428.371, 1315.265, 759.3845, 608.1971, 375.0185, 229.107, 
    391.8174, 639.2117, 819.7453, 915.3849, 607.8117, 379.9553, 305.7845, 
    306.8441, 298.1168, 286.4967, 240.3828, 184.6151,
  0, 0, 0, 0, 0, 0, 0, 0, 0.121945, 0.03938331, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.3118506, 3.291815, 0.01598853, 0, 0, 0, 0, 0, 0.1340173, 
    4.044582, 143.5697, 233.638, 191.9344, 118.6989, 147.4646, 285.2692, 
    535.5562, 720.2246, 908.1365, 672.2578, 505.0814, 365.3874, 130.3261, 
    44.65852, 61.89712, 58.099, 59.19082, 61.83461, 73.12101, 69.1452, 
    71.91867, 79.77286, 88.05507, 108.2875, 147.0296, 195.7139, 207.4643, 
    157.7728, 145.7407, 144.7948, 163.3843, 160.5329, 192.4493, 810.9302, 
    1566.056, 2149.559, 2256.098, 2102.709, 1810.442, 1541.477, 1113.111, 
    754.5137, 622.1283, 649.4427, 513.0068, 210.115, 259.1717, 228.6151, 
    216.1971, 473.4304, 783.3362, 789.3256, 686.4561, 419.5589, 249.4682, 
    205.099, 202.2573, 216.5917, 217.1671, 199.7617, 132.155,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.005494107, 0.4346767, 0, 0, 0, 0, 0, 0, 0, 9.391527, 298.571, 237.2993, 
    140.6926, 155.2257, 256.6727, 406.4414, 433.8806, 600.3461, 683.2579, 
    620.795, 483.5708, 265.2493, 69.42221, 44.01501, 51.81279, 60.87005, 
    53.39784, 52.44471, 56.40654, 59.58292, 67.88076, 74.34882, 81.33792, 
    95.65347, 148.0806, 236.6955, 255.9585, 205.559, 151.0034, 159.6844, 
    176.646, 199.4624, 204.3659, 270.1312, 848.1915, 1003.153, 1148.617, 
    1003.102, 887.6286, 594.8246, 321.8112, 230.0089, 347.2778, 260.032, 
    255.0762, 190.1423, 159.5509, 136.5862, 182.9312, 271.9562, 310.1284, 
    283.9276, 277.2419, 213.3407, 155.9381, 136.6259, 129.9663, 124.8657, 
    144.5141, 150.6962, 106.1049,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.2010026, 5.480222, 1.905644, 0, 0, 0, 0, 0, 0, 10.41574, 79.70645, 
    33.17719, 101.7773, 211.8761, 328.2486, 519.1068, 687.5656, 568.6201, 
    426.9638, 407.4171, 258.6449, 133.8155, 46.44923, 40.82528, 43.58858, 
    52.29549, 51.97647, 43.10914, 47.15418, 57.30152, 61.27217, 67.14295, 
    78.3484, 97.84009, 141.1024, 209.3585, 245.7221, 223.8985, 178.6274, 
    164.8928, 205.0671, 272.722, 329.3512, 281.3043, 329.6042, 396.7708, 
    453.139, 536.9029, 418.7523, 345.6891, 235.4872, 214.9491, 197.1605, 
    217.0889, 210.202, 187.8262, 155.8819, 114.6811, 108.0696, 103.5813, 
    75.537, 103.2833, 131.8954, 130.8562, 121.067, 118.0025, 105.5169, 
    96.54052, 119.8245, 176.6302, 195.5793,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 1.086443, 9.708963, 25.8066, 0, 0, 0, 0.6762983, 7.368328, 15.26273, 
    7.240432, 15.79535, 109.3353, 221.0537, 269.0515, 704.3265, 939.6818, 
    701.0948, 330.6563, 190.7539, 178.3714, 105.7215, 59.61247, 39.14966, 
    45.20544, 46.21466, 48.67001, 35.86091, 46.08049, 52.98456, 62.92745, 
    69.35141, 85.43824, 110.8834, 142.6441, 180.2906, 238.7265, 252.6595, 
    239.7324, 184.5832, 228.8213, 276.7168, 392.7193, 388.6469, 296.1601, 
    280.3641, 341.4388, 353.615, 317.2159, 244.4351, 223.8407, 201.6992, 
    183.6967, 176.9333, 172.614, 165.7017, 145.3332, 110.9088, 80.85966, 
    70.93066, 76.48385, 91.80798, 97.15785, 91.67457, 100.7875, 107.6938, 
    96.9532, 86.08794, 101.3551, 185.22, 281.0552,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 2.485921, 26.4163, 34.1476, 13.50462, 14.0831, 0.4166287, 2.192102, 
    29.53002, 14.33252, 3.286679, 52.2133, 156.3645, 257.6373, 649.4648, 
    1054.655, 614.7567, 162.2067, 99.85813, 116.9508, 77.15819, 48.32669, 
    64.66377, 56.2935, 65.67332, 46.97363, 33.90272, 37.93755, 51.28942, 
    58.10233, 78.93856, 106.3503, 116.9305, 149.4504, 180.898, 213.7403, 
    292.1611, 291.1207, 281.1519, 252.0287, 285.7556, 316.2794, 374.6313, 
    325.8148, 322.2468, 325.9581, 276.3282, 228.0858, 195.2241, 187.3171, 
    175.7014, 163.5601, 151.0618, 141.3108, 129.977, 114.84, 86.42167, 
    68.05943, 63.20282, 64.60545, 60.11647, 42.99261, 50.01132, 55.99592, 
    74.10268, 81.50942, 73.58952, 83.45282, 127.7083, 226.8334,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 2.984597, 0.01858864, 0, 0.0009470581, 16.01784, 
    87.35822, 173.5935, 488.2748, 759.5725, 523.7241, 141.7197, 113.1382, 
    159.5228, 147.7596, 115.4366, 107.1132, 102.7932, 85.72213, 66.42902, 
    30.98574, 37.11678, 45.43555, 64.23547, 99.53561, 129.9766, 138.2153, 
    142.8759, 176.7178, 267.0287, 349.3065, 417.0574, 373.9982, 391.8378, 
    306.8354, 254.5319, 312.5648, 296.5179, 377.6109, 330.0472, 242.8435, 
    164.2536, 149.3302, 147.9863, 144.5899, 139.069, 133.0572, 122.3601, 
    110.4266, 95.19322, 77.43336, 63.58871, 58.07784, 51.05425, 36.38617, 
    36.80247, 46.6338, 42.84441, 35.56261, 47.46378, 56.36189, 58.939, 
    105.9327, 189.9787,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 5.923116, 0, 0, 0, 0, 0, 6.078897, 54.77836, 77.55535, 
    204.2334, 410.9161, 330.8391, 185.1925, 194.0988, 249.267, 253.3829, 
    177.0466, 158.8476, 113.1643, 101.53, 68.00449, 31.76886, 36.63785, 
    58.77195, 90.80497, 133.0862, 161.9473, 164.7115, 165.2141, 201.0824, 
    279.0718, 359.1356, 398.5262, 459.7346, 501.9608, 511.8822, 352.2849, 
    246.1968, 246.5588, 279.2735, 323.1726, 191.8587, 143.4464, 112.1324, 
    117.9595, 116.5617, 114.9787, 113.5484, 107.3903, 97.09441, 84.3097, 
    70.09772, 57.50354, 51.82816, 43.33216, 40.77794, 45.42603, 66.79871, 
    45.82823, 21.87241, 20.00079, 29.68418, 34.1625, 55.23173, 131.1202,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.007114115, 12.30466, 48.17017, 
    51.3419, 136.4395, 140.1926, 152.5834, 214.4402, 290.774, 334.6097, 
    242.1319, 179.8538, 138.1877, 94.74007, 53.06939, 31.48326, 46.89961, 
    89.87615, 131.2574, 140.4565, 168.6543, 171.5402, 207.168, 234.0502, 
    297.8369, 300.6861, 321.7401, 399.447, 557.8159, 602.8211, 392.1693, 
    231.2913, 117.9363, 190.2211, 228.4644, 181.8213, 100.4968, 90.92713, 
    91.9957, 95.57886, 98.97549, 93.66434, 91.03915, 82.98544, 72.89633, 
    60.49364, 58.69539, 60.83919, 60.2387, 64.67129, 64.97378, 60.37475, 
    50.22374, 26.93556, 10.59541, 21.63067, 16.65605, 21.7373, 41.34349,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5.366938, 28.12142, 64.29294, 
    128.7759, 176.1391, 224.7735, 297.6988, 326.8529, 254.3473, 185.0925, 
    128.5998, 87.42819, 38.13975, 29.44325, 68.62458, 118.0892, 143.8512, 
    173.974, 164.9058, 204.4256, 210.1949, 267.1867, 300.9321, 309.5306, 
    297.9662, 355.8887, 461.3635, 509.2478, 310.7938, 206.6006, 123.8932, 
    125.1484, 178.9654, 129.2888, 94.40868, 92.13621, 118.3059, 139.3436, 
    102.2285, 87.8205, 78.24416, 72.41794, 72.99378, 69.93626, 64.41702, 
    66.0837, 67.51834, 70.63937, 64.17177, 65.43086, 61.57732, 57.59845, 
    48.39719, 66.22498, 19.65588, 7.979198, 7.954746,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1979136, 16.10868, 94.42965, 
    187.4814, 245.3877, 271.5805, 257.391, 297.2609, 210.7862, 164.771, 
    95.62947, 56.90887, 40.72773, 52.8884, 92.41105, 126.1473, 166.0383, 
    207.8445, 272.0114, 271.0105, 294.9529, 248.3746, 307.0643, 316.8501, 
    327.4612, 325.9547, 386.9184, 403.7983, 311.1118, 240.8184, 164.2083, 
    103.1077, 117.4106, 99.13666, 106.3574, 154.6648, 260.3508, 285.6964, 
    234.8461, 154.5512, 112.9279, 100.7134, 123.8555, 127.3378, 90.11683, 
    76.42348, 68.03311, 66.51344, 75.3875, 112.4858, 142.2936, 124.5137, 
    93.33791, 99.31126, 54.70262, 4.06266, 0.262289,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.04155033, 10.73219, 79.11258, 
    190.445, 274.9487, 342.6148, 355.8712, 312.3603, 292.6754, 221.7762, 
    115.474, 47.77611, 50.80471, 84.23752, 95.56871, 148.4016, 177.4802, 
    241.8285, 273.5516, 339.5761, 337.356, 326.2194, 277.1494, 336.4698, 
    352.6033, 363.4337, 382.938, 416.9631, 325.3823, 303.8384, 203.988, 
    116.0254, 110.5155, 121.6094, 106.5421, 137.3756, 210.812, 317.8851, 
    344.7708, 323.2015, 252.112, 193.5985, 213.3652, 191.4196, 156.1301, 
    106.2765, 104.4049, 72.89532, 100.3581, 157.0007, 215.9135, 191.733, 
    119.1055, 115.4301, 99.49779, 31.93542, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.542466, 22.26523, 77.77408, 
    140.4331, 240.0608, 343.6068, 376.1221, 378.217, 372.9897, 356.2578, 
    217.9453, 48.16224, 56.58264, 94.03797, 155.6086, 206.1189, 244.8234, 
    262.5258, 267.4071, 294.3894, 384.4132, 383.2951, 330.3748, 318.6039, 
    351.7903, 366.8914, 400.56, 447.5571, 438.7595, 508.2295, 383.2372, 
    246.7716, 200.7712, 148.0255, 184.6252, 228.8072, 293.0768, 384.8521, 
    451.6723, 470.1341, 383.5, 297.7384, 261.2184, 257.7826, 233.8021, 
    230.1151, 168.3038, 140.5308, 159.7929, 141.3796, 184.5563, 169.6956, 
    127.2488, 153.812, 157.5335, 129.1637, 8.482048 ;
}
