netcdf atmos.1980-1981.alb_sfc.08 {
dimensions:
	time = UNLIMITED ; // (1 currently)
	lat = 18 ;
	lon = 29 ;
	bnds = 2 ;
variables:
	float alb_sfc(time, lat, lon) ;
		alb_sfc:long_name = "Surface Albedo for  Flux" ;
		alb_sfc:units = "percent" ;
		alb_sfc:_FillValue = 1.e+20f ;
		alb_sfc:missing_value = 1.e+20f ;
		alb_sfc:cell_measures = "area: area" ;
		alb_sfc:interp_method = "conserve_order1" ;
		alb_sfc:cell_methods = "time: mean within months time: mean over years" ;
		alb_sfc:time_avg_info = "average_T1,average_T2,average_DT" ;
	double average_DT(time) ;
		average_DT:long_name = "Length of average period" ;
		average_DT:units = "days" ;
	double average_T1(time) ;
		average_T1:long_name = "Start time for average period" ;
		average_T1:units = "days since 1979-01-01 00:00:00" ;
	double average_T2(time) ;
		average_T2:long_name = "End time for average period" ;
		average_T2:units = "days since 1979-01-01 00:00:00" ;
	double climatology_bounds(time, bnds) ;
	double lat(lat) ;
		lat:standard_name = "latitude" ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_N" ;
		lat:axis = "Y" ;
		lat:bounds = "lat_bnds" ;
	double lat_bnds(lat, bnds) ;
	double lon(lon) ;
		lon:standard_name = "longitude" ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_E" ;
		lon:axis = "X" ;
		lon:bounds = "lon_bnds" ;
	double lon_bnds(lon, bnds) ;
	double time(time) ;
		time:standard_name = "time" ;
		time:long_name = "time" ;
		time:climatology = "climatology_bounds" ;
		time:units = "days since 1979-01-01 00:00:00" ;
		time:calendar = "standard" ;
		time:axis = "T" ;

// global attributes:
		:CDI = "Climate Data Interface version 2.4.4 (https://mpimet.mpg.de/cdi)" ;
		:Conventions = "CF-1.6" ;
		:title = "c96L65_am5f9d8r0_amip" ;
		:associated_files = "area: 19800101.grid_spec.nc" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
		:code_release_version = "2024.05" ;
		:git_hash = "5d306c05d9fe755cab04eedc8fd3de0d3c8355a0" ;
		:creationtime = "Mon Aug 25 14:09:46 2025" ;
		:hostname = "pp050" ;
		:history = "Mon Aug 25 13:32:20 2025: ncks -d lat,,,10 -d lon,,,10 atmos.1980-1981.alb_sfc.08.nc reduced/atmos.1980-1981.alb_sfc.08.nc\n",
			"Mon Aug 25 14:40:07 2025: cdo -O -s -select,month=8 merged_output.nc monthly_nc_files/all_years.8.nc\n",
			"Mon Aug 25 14:40:01 2025: cdo -O -s -mergetime /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/shards/ts/regrid-xy/180_288.conserve_order2/atmos_month/P1M/P1Y/atmos_month.198001-198012.alb_sfc.nc /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/shards/ts/regrid-xy/180_288.conserve_order2/atmos_month/P1M/P1Y/atmos_month.198101-198112.alb_sfc.nc merged_output.nc\n",
			"Mon Aug 25 14:12:17 2025: cdo --history splitname 19800101.atmos_month.nc /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/cycle/19800101T0000Z/split/regrid-xy/180_288.conserve_order2/19800101.atmos_month.\n",
			"fregrid --debug --standard_dimension --input_mosaic C96_mosaic.nc --input_dir /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/cycle/19800101T0000Z/history/native --input_file 19800101.atmos_month --associated_file_dir /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/cycle/19800101T0000Z/history/native --interp_method conserve_order2 --remap_file fregrid_remap_file_288_by_180.nc --nlon 288 --nlat 180 --scalar_field (**please see the field list in this file**) --output_file 19800101.atmos_month.nc" ;
		:CDO = "Climate Data Operators version 2.4.4 (https://mpimet.mpg.de/cdo)" ;
		:comment = "FMS time averaging, version 3.0, precision=double" ;
		:NCO = "netCDF Operators version 5.2.4 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco, Citation = 10.1016/j.envsoft.2008.03.004)" ;
data:

 alb_sfc =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  2.366829, 2.46821, 2.420455, 2.091436, 2.318314, 2.258152, 2.254859, 
    2.254442, 2.172514, 2.196928, 2.416126, 2.159431, 2.213321, 2.410579, 
    2.483516, 2.609395, 2.625607, 2.691821, 2.562482, 2.419828, 2.586178, 
    2.560362, 2.476865, 2.379706, 2.279095, 2.655873, 2.718772, 2.558059, 
    2.42342,
  25.26284, 25.40875, 26.33274, 24.51161, 22.20685, 22.18373, 24.37224, 
    22.17222, 22.20707, 22.29963, 22.28218, 22.31068, 22.52548, 26.29648, 
    26.42618, 26.35486, 26.30699, 26.29595, 17.9051, 25.5841, 25.76107, 
    25.69589, 26.08877, 24.44001, 26.51733, 26.71969, 26.57114, 26.51045, 
    26.38241,
  33.14256, 33.68362, 3.382408, 3.699799, 3.754351, 3.920091, 33.46571, 
    16.3848, 4.289661, 3.978464, 3.672228, 3.673528, 3.072951, 3.179226, 
    3.213058, 3.270795, 2.977889, 3.123615, 3.436459, 3.739113, 4.256887, 
    4.241986, 3.989887, 4.199984, 16.36665, 27.20821, 32.29028, 33.11361, 
    33.53513,
  3.979927, 4.074976, 3.824885, 3.784202, 3.522146, 3.511045, 3.82536, 
    3.82773, 4.013837, 4.116347, 3.87122, 3.814723, 3.76345, 3.81753, 
    3.560913, 3.765203, 3.68861, 3.656616, 3.821159, 3.981951, 3.862482, 
    3.992827, 3.935484, 9.452635, 4.332763, 3.862219, 3.761817, 3.643336, 
    3.714016,
  3.64515, 3.809299, 3.98416, 3.698995, 3.731, 3.722822, 3.842741, 3.923366, 
    3.768137, 4.083189, 3.927318, 4.021428, 4.274255, 4.035739, 12.57354, 
    3.883534, 3.955111, 3.791033, 3.916451, 3.807699, 3.764191, 3.688033, 
    3.707568, 10.63035, 4.367794, 3.850884, 3.689569, 3.668735, 3.554564,
  3.777102, 3.787005, 12.33903, 3.964925, 3.874869, 3.983664, 3.853177, 
    3.918142, 3.810855, 4.22885, 9.023102, 13.51037, 10.21618, 4.054742, 
    4.108144, 3.831689, 3.785079, 3.489669, 3.698431, 3.721709, 3.863267, 
    3.754475, 3.9168, 4.648613, 8.456511, 3.673849, 3.553813, 3.759812, 
    3.68798,
  3.310161, 9.526138, 9.832544, 3.866919, 3.756557, 3.794958, 3.828189, 
    3.798339, 3.495016, 4.33229, 11.55002, 11.36397, 3.857469, 3.617673, 
    3.575799, 3.655135, 3.71266, 3.566099, 4.080117, 3.689199, 3.793124, 
    3.456768, 3.247229, 3.715207, 9.128654, 9.076441, 3.687849, 4.0109, 
    3.366214,
  3.15832, 6.050251, 9.47431, 9.011673, 3.563254, 3.669701, 3.246144, 
    3.398107, 3.488654, 3.511295, 4.732032, 3.604498, 4.104648, 3.384106, 
    3.649719, 3.467798, 3.75199, 3.937099, 3.822816, 3.705732, 3.803702, 
    3.266157, 3.314707, 9.046949, 8.646479, 9.061268, 3.906875, 3.687926, 
    3.377157,
  3.128197, 8.488458, 8.390132, 9.987049, 3.437728, 3.172434, 3.156907, 
    3.163639, 8.529546, 8.177944, 3.144166, 3.199996, 3.235384, 3.410739, 
    3.483009, 3.562577, 3.572412, 3.723848, 3.611713, 3.616317, 3.504658, 
    3.280179, 3.251914, 8.595877, 8.728022, 3.450162, 3.497264, 3.332274, 
    3.209054,
  9.62315, 9.905354, 9.594234, 9.318546, 14.89939, 3.189229, 5.053913, 
    3.02511, 3.312397, 3.219826, 4.230791, 3.135295, 3.349174, 3.377048, 
    3.187453, 3.368365, 3.284541, 3.262901, 3.249452, 3.26811, 3.152399, 
    3.246192, 8.818924, 7.323259, 3.330193, 3.120418, 2.980527, 3.124054, 
    8.483294,
  18.12294, 20.94926, 23.17325, 3.104602, 23.13115, 3.10534, 10.03437, 
    3.134645, 8.911091, 3.164966, 3.309695, 3.296278, 3.186119, 3.305102, 
    3.375503, 3.575206, 3.566499, 3.886263, 3.29626, 3.427864, 3.305232, 
    6.19355, 3.378288, 4.134084, 3.297482, 3.282988, 3.328471, 3.054445, 
    23.90358,
  24.51614, 20.68941, 21.28876, 19.93844, 13.01668, 15.05026, 12.14788, 
    9.776079, 7.008596, 10.49477, 3.567756, 3.523222, 3.617994, 3.62758, 
    3.535968, 3.906259, 3.80383, 4.023231, 3.668118, 3.893957, 12.33089, 
    11.91847, 9.170935, 3.365723, 3.608935, 3.6438, 4.017727, 3.605088, 
    11.20376,
  6.687468, 4.255378, 6.383416, 10.62898, 2.14467, 15.72688, 9.012815, 
    15.84152, 13.60104, 11.22608, 7.412081, 3.815983, 3.693043, 3.613549, 
    3.712026, 3.624846, 3.627609, 3.855302, 3.80417, 12.69293, 11.58579, 
    13.90503, 12.98967, 4.430345, 3.708153, 3.770747, 3.876454, 3.9554, 
    5.308846,
  6.207911, 12.4712, 13.82163, 14.53812, 13.83655, 12.70392, 8.41202, 
    11.28601, 7.695023, 7.102299, 7.089316, 6.866447, 4.037688, 3.784142, 
    3.734831, 3.674707, 3.901035, 3.949027, 4.112491, 9.485298, 10.97815, 
    10.04877, 7.115485, 6.904938, 5.387272, 4.077386, 4.059889, 4.139397, 
    4.116015,
  4.624712, 7.563159, 8.738003, 7.290542, 7.856249, 7.619391, 7.665995, 
    7.783946, 7.82598, 7.782948, 7.665679, 11.50543, 11.85026, 6.964451, 
    4.608799, 4.65749, 9.877812, 15.28456, 11.15907, 7.799496, 7.025727, 
    11.7302, 4.831911, 11.54305, 4.298043, 8.846851, 4.207454, 4.301073, 
    4.345144,
  4.978373, 5.632957, 8.798571, 5.421516, 5.032849, 6.019876, 14.08095, 
    13.13807, 13.95054, 13.91935, 10.33824, 10.03661, 13.68164, 7.90123, 
    20.92571, 5.096689, 10.5175, 10.55944, 6.932899, 8.581902, 23.50345, 
    20.08471, 19.06182, 29.11825, 5.551883, 52.46976, 56.56561, 8.951762, 
    4.95751,
  50.91398, 10.84881, 33.86969, 29.24585, 26.64746, 25.15069, 49.78511, 
    41.03575, 47.57872, 60.8899, 61.05832, 60.72473, 60.90753, 60.94188, 
    61.2774, 61.69684, 61.78271, 61.88842, 61.69769, 60.90642, 60.77221, 
    51.87119, 51.75109, 58.98893, 70.78397, 70.80962, 74.80889, 60.36003, 
    42.8019 ;

 average_DT = 730 ;

 average_T1 = 228.5 ;

 average_T2 = 958.5 ;

 climatology_bounds =
  228.5, 958.5 ;

 lat = -89.5, -79.5, -69.5, -59.5, -49.5, -39.5, -29.5, -19.5, -9.5, 0.5, 
    10.5, 20.5, 30.5, 40.5, 50.5, 60.5, 70.5, 80.5 ;

 lat_bnds =
  -90, -89,
  -80, -79,
  -70, -69,
  -60, -59,
  -50, -49,
  -40, -39,
  -30, -29,
  -20, -19,
  -10, -9,
  0, 1,
  10, 11,
  20, 21,
  30, 31,
  40, 41,
  50, 51,
  60, 61,
  70, 71,
  80, 81 ;

 lon = 0.625, 13.125, 25.625, 38.125, 50.625, 63.125, 75.625, 88.125, 
    100.625, 113.125, 125.625, 138.125, 150.625, 163.125, 175.625, 188.125, 
    200.625, 213.125, 225.625, 238.125, 250.625, 263.125, 275.625, 288.125, 
    300.625, 313.125, 325.625, 338.125, 350.625 ;

 lon_bnds =
  0, 1.25,
  12.5, 13.75,
  25, 26.25,
  37.5, 38.75,
  50, 51.25,
  62.5, 63.75,
  75, 76.25,
  87.5, 88.75,
  100, 101.25,
  112.5, 113.75,
  125, 126.25,
  137.5, 138.75,
  150, 151.25,
  162.5, 163.75,
  175, 176.25,
  187.5, 188.75,
  200, 201.25,
  212.5, 213.75,
  225, 226.25,
  237.5, 238.75,
  250, 251.25,
  262.5, 263.75,
  275, 276.25,
  287.5, 288.75,
  300, 301.25,
  312.5, 313.75,
  325, 326.25,
  337.5, 338.75,
  350, 351.25 ;

 time = 0 ;
}
