netcdf \20030101.atmos_static_cmip.tile2 {
dimensions:
	grid_xt = 96 ;
	grid_yt = 96 ;
	time = UNLIMITED ; // (1 currently)
variables:
	double grid_xt(grid_xt) ;
		grid_xt:units = "degrees_E" ;
		grid_xt:long_name = "T-cell longitude" ;
		grid_xt:axis = "X" ;
	double grid_yt(grid_yt) ;
		grid_yt:units = "degrees_N" ;
		grid_yt:long_name = "T-cell latitude" ;
		grid_yt:axis = "Y" ;
	double time(time) ;
		time:units = "days since 1870-01-01 00:00:00" ;
		time:long_name = "time" ;
		time:axis = "T" ;
		time:calendar_type = "JULIAN" ;
		time:calendar = "julian" ;
	float orog(grid_yt, grid_xt) ;
		orog:_FillValue = 1.e+20f ;
		orog:missing_value = 1.e+20f ;
		orog:units = "m" ;
		orog:long_name = "Surface Altitude" ;
		orog:cell_methods = "time: point" ;
		orog:cell_measures = "area: area" ;
		orog:standard_name = "surface_altitude" ;
		orog:interp_method = "conserve_order1" ;

// global attributes:
		:title = "ESM4_longamip_D1_am4p2_proto7b_whiteCapsAlbedo_salt_SIS2" ;
		:associated_files = "area: 20030101.grid_spec.nc" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
data:

 grid_xt = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19, 
    20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 37, 
    38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 54, 55, 
    56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 72, 73, 
    74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 90, 91, 
    92, 93, 94, 95, 96 ;

 grid_yt = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19, 
    20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 37, 
    38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 54, 55, 
    56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 72, 73, 
    74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 90, 91, 
    92, 93, 94, 95, 96 ;

 time = 0 ;

 orog =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.007482118, 
    4.885016, 6.027729, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4.712759, 58.8956, 
    114.3027, 105.147, 66.36284,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6.754428, 58.17822, 103.8941, 
    76.19964, 51.16923, 83.5846, 145.4227, 210.3575, 222.043, 166.9021, 
    138.0394,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12.60223, 150.9446, 238.0754, 281.3481, 
    288.7326, 300.3335, 276.3248, 277.1753, 296.433, 282.2253, 207.1847, 
    170.1954,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6.971491, 107.903, 253.5528, 311.8893, 
    314.664, 349.46, 376.1395, 363.9048, 328.7521, 316.8185, 308.9201, 
    249.6144, 213.1554,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1077713, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5.728832, 54.67075, 280.7457, 
    309.0462, 322.4052, 368.6298, 412.7725, 423.5071, 379.2067, 346.22, 
    351.7698, 329.3646, 274.3772,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2.078801, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17.70223, 257.5212, 295.4054, 
    313.6127, 373.5954, 422.1055, 435.1128, 393.682, 374.0881, 409.6835, 
    409.2048, 354.9377,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26.2593, 246.0138, 296.1431, 348.5571, 
    410.7598, 429.6357, 435.3861, 395.7879, 402.5177, 442.4218, 430.7854, 
    398.5805,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 113.7163, 268.1346, 336.5029, 392.1589, 
    444.2632, 443.9155, 420.9473, 421.8472, 452.1077, 471.5658, 444.4251, 
    418.9319,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5.859579, 200.0244, 305.7336, 330.6553, 
    391.9315, 444.2378, 439.8025, 441.541, 463.3921, 503.8092, 497.416, 
    462.6526, 441.0611,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14.25746, 228.6333, 312.2241, 361.2495, 
    416.0756, 482.3185, 484.5522, 484.6867, 507.3547, 509.7314, 483.8749, 
    461.7263, 442.7195,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0.007934935, 91.5881, 260.8788, 351.2304, 
    404.0062, 456.2148, 509.2211, 528.7908, 527.3947, 511.4882, 494.72, 
    462.9256, 467.0975, 450.041,
  7.299402, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8.026843, 190.214, 291.695, 351.6114, 
    434.4432, 470.4533, 537.1084, 567.7097, 561.1059, 537.2833, 494.2285, 
    457.0371, 454.9888, 443.677,
  46.47058, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 32.85493, 192.2326, 276.3241, 346.8046, 
    419.9743, 473.221, 539.5166, 587.4988, 579.1885, 551.3723, 502.3163, 
    438.6668, 426.6781, 416.2831,
  56.36044, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.2935236, 29.53243, 141.496, 253.5633, 
    345.4431, 426.5362, 485.1349, 548.7592, 600.852, 588.0337, 535.9756, 
    460.5315, 394.231, 382.3351, 380.9086,
  39.45049, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 32.83228, 53.73461, 1.585332, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3.041326, 10.00888, 
    106.9153, 227.8007, 348.7626, 445.4996, 478.5939, 575.4977, 600.4197, 
    570.2203, 506.0541, 415.3415, 330.4285, 332.2667, 343.1945,
  13.59347, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26.08635, 195.4105, 256.4257, 146.537, 
    55.481, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.186994, 
    18.06586, 130.0469, 253.3653, 363.8199, 394.896, 513.6748, 590.4353, 
    558.9642, 518.7917, 454.3615, 363.8717, 303.3865, 300.713, 321.3069,
  0.9656757, 0, 0, 0, 0, 0, 0.03586638, 0, 0, 0, 49.68565, 326.9774, 
    455.3936, 576.6316, 425.3625, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.01508173, 21.43529, 144.3786, 255.7441, 319.1965, 459.2542, 
    569.7118, 604.0175, 513.782, 425.8328, 371.0454, 316.678, 281.3964, 
    295.9887, 312.7417,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 188.9793, 461.0893, 744.1964, 857.3239, 
    577.0432, 10.22077, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    28.41998, 89.48728, 170.1808, 341.458, 487.3284, 552.6357, 471.7288, 
    351.3307, 336.5912, 295.8323, 257.3056, 256.7657, 275.5327, 266.8901,
  14.46666, 0, 0, 0, 0, 0, 0, 0, 0, 0, 98.10371, 430.0524, 658.2639, 
    869.6558, 593.5727, 27.91763, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 28.79319, 27.47902, 102.3828, 250.1567, 353.9292, 297.6356, 
    194.349, 196.082, 204.2073, 194.9052, 184.4335, 186.8029, 202.2491, 
    201.6232,
  63.77672, 3.367655, 0, 0, 0, 0, 0, 0, 0, 0, 20.47009, 226.3262, 481.9063, 
    847.3206, 850.9589, 97.98926, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 5.864242, 1.030459, 11.5586, 92.8717, 81.6533, 37.3248, 
    45.25832, 55.12968, 71.40536, 80.22321, 109.8221, 156.4528, 158.7244, 
    139.6773,
  92.77831, 10.55024, 0.7231424, 0, 0, 0, 0, 0, 0, 0, 0.06683189, 88.24445, 
    325.958, 897.7953, 1142.866, 334.1817, 0.2153307, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.6444512, 1.022004, 0.2444094, 0, 
    0.1744056, 0, 0, 11.61093, 95.71937, 140.5593, 109.8717, 89.47809,
  148.8612, 111.2776, 10.43683, 0.2487843, 0, 0, 0, 0, 0, 0, 0, 26.9947, 
    302.4542, 900.6857, 1410.459, 722.3347, 26.92253, 0, 0, 0, 0, 0, 0, 
    0.2948902, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.04675792, 32.30137, 73.17574, 45.04506, 113.3446,
  356.8611, 272.9169, 144.0292, 36.66886, 4.051232, 0, 0, 0, 0, 0, 
    0.00622688, 95.44665, 402.4702, 1000.551, 1468.909, 1068.681, 138.7007, 
    0, 0, 0, 0, 0, 0, 224.4563, 0.7204035, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 40.79513, 46.98636, 44.90553, 135.4555,
  607.5697, 617.0065, 415.9779, 222.5245, 82.16385, 13.76159, 0, 0, 0, 0, 
    0.7036354, 167.195, 549.0036, 865.797, 1297.997, 1084.883, 386.271, 0, 0, 
    0, 0, 0, 0, 0, 0, 38.47579, 1.349345, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.05735796, 3.489815, 17.0652, 91.46315,
  805.8144, 689.3148, 665.8074, 521.1199, 295.9792, 99.36646, 9.087084, 0, 0, 
    0.005802704, 0.3102686, 111.6922, 363.4742, 565.2116, 806.0615, 1016.094, 
    629.3563, 16.26268, 0, 0, 0, 0, 0, 0, 0, 0, 0.02296036, 0, 0, 0, 0, 
    1.214581, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.002000303, 0.005462797, 
    18.32721,
  760.7727, 661.396, 709.6733, 604.6326, 464.2514, 283.1679, 79.76301, 
    0.1074248, 0, 0, 0, 17.74922, 148.9407, 173.6682, 402.7549, 729.6694, 
    723.2713, 46.89246, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1074003,
  860.9228, 736.6833, 628.5461, 564.9741, 466.655, 335.0508, 169.4657, 
    9.562907, 0, 0, 0, 0, 7.39888, 15.74615, 103.3149, 461.4926, 652.2623, 
    214.472, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, -0.0001159482, 0, 0,
  954.5076, 825.0037, 642.887, 541.5004, 467.5988, 374.7963, 167.8485, 
    1.774008, 0, 0, 0, 0, 0, 0.3348222, 19.11695, 171.6814, 741.9515, 
    374.4197, 25.98872, 0, 0, 0, 0.0003252521, 0, 0, 0, 0, 0.001458651, 
    7.516816e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  858.3884, 673.0359, 533.1504, 448.0885, 424.8119, 345.4697, 166.7318, 0, 0, 
    0, 0, 0, 0, 0, 0.567318, 193.9483, 883.2621, 655.3737, 12.50792, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.0002288724, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.005102882, 0, 0,
  765.3333, 667.6134, 488.7987, 363.019, 313.4333, 341.2213, 122.4717, 0, 0, 
    0, 0, 0, 5.00687, 0, 0, 60.76902, 616.8209, 406.96, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  892.0968, 795.8924, 625.4323, 432.2025, 321.9835, 331.9277, 130.2014, 
    0.004251794, 0, 0, 57.24534, 20.8572, 0.7291545, 0, 0, 0, 119.2905, 
    99.81622, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 13.85986, 0.004370535, 0,
  1001.771, 792.1298, 674.5222, 541.9408, 384.3335, 350.6531, 103.3347, 
    0.1868827, 0, 0, 18.48727, 0, 0, 0, 0, 0, 9.2637, 4.286283, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.02841037, 
    1.063279, 1.850597, 3.574715, 3.295839, 153.8647, 199.7177,
  1318.781, 598.8708, 526.7117, 510.9486, 354.2004, 223.6784, 15.55483, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.01238247, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10.38296, 174.51, 148.3694, 0, 0, 0, 
    148.5062, 285.8834,
  1220.16, 848.2032, 380.6071, 390.465, 259.5177, 95.94141, 0, 0, 0, 0, 0, 0, 
    0, 0.01723676, 0.0002739781, 0.009286015, 0, 0, 0, 0.006633122, 0, 0, 0, 
    0, 0.003201818, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001933358, 
    0, 0, 0, 0, 0, 0, 0, 0, 2.528343, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.01048129, 0, 35.29255, 81.26061, 161.3701, 172.8166, 125.7769, 
    60.08969, 51.96622, 164.8291,
  1338.663, 964.2402, 591.19, 291.6062, 139.8224, 33.77381, 0.002896692, 0, 
    0, 0, 0, 0, 0, 0.09759907, 0, 0, 0, 0, 0.003041361, 0, 0, 0, 0, 0, 
    0.003417519, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2.214117, 10.05566, 31.4626, 
    198.6635, 257.3435, 200.3842, 110.9841, 79.73378, 263.6654, 36.78745, 
    1.378057, 31.15954, 8.130059, 1.005422,
  1026.086, 1045.23, 716.394, 366.1234, 142.9799, 30.33171, 0.4619157, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10.88786, 
    115.5257, 170.2808, 339.2503, 395.8933, 151.5352, 149.8366, 27.3561, 
    4.022614, 20.95062, 0, 0, 3.260029, 1.872875, 0.0508271, 0, 0, 0,
  974.4459, 1067.982, 927.8552, 494.0284, 130.0466, 22.65291, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.899872, 139.8198, 
    115.3161, 168.5896, 352.7554, 266.0829, 177.1721, 131.6926, 43.10759, 
    1.240668, 4.394837, 0.006916575, 0.0003986534, 0.0104446, 0.0172614, 0, 
    2.609623, 0, 0.001365404, 0.09803439, 0.2262536, 0.004817449,
  1204.486, 1237.256, 1141.603, 688.0075, 263.0531, 10.36784, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001947393, 0, 0, 0, 0.01043915, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01680503, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.04407993, 32.09272, 400.8964, 597.5397, 333.6716, 124.2354, 104.7639, 
    67.59129, 23.81756, 3.731113, 1.087241, 0, 0, 0, 0, 0, 0, 4.881635, 
    10.31701, 0, 6.561506, 40.6811, 3.38201, 0.01358287,
  1440.196, 1303.7, 1187.572, 799.9657, 447.4943, 28.87032, 0.287935, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.008367683, 0, 0.0005597501, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.006913288, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 17.87501, 27.6564, 41.68385, 40.07766, 2.412819, 0, 0.3703949, 0, 0, 
    2.694052, 0, 0.06298108, 0, 0, 0.007401017, 0.01018163, 0.5245222, 
    314.3598, 25.13958, 10.84065, 64.80965, 69.94651, 0.2126305, 0,
  1507.507, 1338.634, 1162.16, 895.2739, 556.3425, 113.5388, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.003531589, 0, 0.3608332, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6.645804e-05, 0.008660849, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1.399279, 1.708197, 228.0259, 260.7763, 73.72216, 0.01350134, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.04154294, 0.6853305, 0.0007041242, 0, 0, 0, 222.6289, 
    19.51247, 152.801, 98.75947, 68.60026, 0, 0,
  1593.552, 1288.948, 1293.234, 1037.663, 604.3491, 220.0716, 11.92896, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3.231213, 0.1002754, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.003929192, 0.06615317, 
    326.9998, 382.6881, 215.296, 6.51867, 0, 0, 0.0005210711, 0, 0, 0, 
    0.00945402, 0, 0.04497931, 26.08819, 57.13885, 7.390703, 0, 0, 69.87069, 
    559.0273, 111.9894, 624.2891, 262.6683, 1.642632, 0, 0,
  1658.693, 1261.843, 1404.586, 1067.003, 563.8726, 182.1493, 36.27239, 
    0.3323672, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0002778716, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3.277349, 3.089526, 
    220.2578, 271.9154, 232.9942, 11.41514, 6.090748, 2.68348, 5.510962, 
    3.529593, 0, 1.621469, 5.491666, 9.77548, 7.35185, 3.514773, 53.89715, 
    161.2589, 24.12606, 0, 0.007201126, 433.8056, 1036.646, 400.0064, 
    500.544, 149.6249, 0, 0, 0,
  1645.619, 1472.14, 1404.025, 1096.18, 483.7211, 188.2313, 50.92135, 
    15.02244, 0.3012842, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9.016459, 125.5137, 
    477.9677, 315.6645, 11.36371, 6.38086, 10.82686, 9.825094, 2.584005, 
    0.8772991, 0, 14.4698, 70.73858, 64.99486, 20.69061, 17.08455, 32.61346, 
    164.0018, 34.12597, 0.002215982, 0, 41.34579, 1159.648, 903.4078, 
    550.6257, 25.76042, 12.09169, 7.678148, 124.0715,
  1967.175, 1791.275, 1808.567, 1089.094, 523.5789, 218.3327, 97.51249, 
    52.39918, 11.84871, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26.70954, 0.01252906, 
    573.1802, 456.6572, 67.73898, 16.5005, 4.31343, 5.305326, 0.0450154, 0, 
    0.8252385, 6.159415, 65.49741, 194.1909, 179.5106, 157.9093, 77.64091, 
    91.67677, 141.2131, 99.64323, 8.659935, 0, 4.571824, 614.8233, 532.0992, 
    483.2188, 457.6458, 209.052, 8.435591, 0,
  2024.533, 2181.229, 2001.106, 1283.735, 528.7686, 242.7618, 136.9167, 
    79.82225, 23.44122, 3.95113, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.004921097, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.6401625, 
    6.308005, 158.2323, 422.013, 185.8305, 17.01043, 4.866463, 8.841109, 
    0.001300426, 0, 0, 0, 11.91, 84.76138, 176.0108, 242.7657, 291.476, 
    330.5183, 200.2534, 138.5459, 34.58592, 22.24334, 0, 0, 144.1948, 0, 
    6.173299, 15.85019, 45.24471, 0.213134, 0,
  1923.579, 1771.256, 1778.076, 1070.793, 505.6136, 241.9928, 148.163, 
    76.44843, 32.30178, 17.09214, 7.496256, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01376197, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.004098975, 22.05864, 72.32189, 406.9106, 296.7709, 13.30871, 10.29677, 
    4.396094, 1.765978, 0, 0.01962267, 0.09792335, 0.3374118, 51.71622, 
    88.17578, 76.92102, 159.3824, 380.0949, 535.228, 499.3378, 330.4606, 
    165.3464, 41.27188, 2.509667, 0.02632017, 117.6165, 245.3032, 188.3384, 
    112.4978, 172.8582, 310.4585, 94.6843,
  1794.133, 1276.998, 1319.927, 847.228, 358.8172, 233.8158, 187.9514, 
    116.8452, 68.52618, 71.37233, 45.78811, 16.83432, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.009340961, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 2.670939, 25.97792, 355.1271, 272.5902, 27.50756, 10.82965, 
    10.10394, 20.80869, 2.207196, 0, 0.004632319, 0.4954259, 0, 54.69146, 
    103.1393, 87.46021, 162.231, 378.5865, 622.8563, 789.714, 748.1737, 
    514.2153, 211.2245, 106.0069, 43.93421, 0, 117.153, 217.9034, 176.2699, 
    56.00568, 72.75879, 291.925,
  1122.184, 817.0998, 942.5208, 629.3625, 367.3386, 319.362, 310.6506, 
    233.7132, 219.4219, 172.6176, 170.9612, 87.88506, 52.56012, 6.837942, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.01282556, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.003567874, 9.907857, 7.509503, 341.4931, 669.8797, 266.7873, 
    11.2073, 57.75204, 56.43156, 49.87582, 0.7429065, 0.01104457, 0.2828173, 
    0, 0.04069449, 4.1862, 0.06066301, 11.07728, 86.06728, 187.3697, 
    479.2986, 762.8614, 937.4857, 601.6578, 195.3882, 27.83612, 0.1914168, 0, 
    0, 0, 0, 0, 0, 11.51637,
  846.5782, 504.4499, 654.7703, 570.2628, 501.0254, 542.6677, 483.9015, 
    424.1021, 332.9808, 314.234, 333.5416, 253.9334, 130.1149, 111.9619, 
    7.31144, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.0009155833, 0.003754308, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.204808, 504.0269, 598.7817, 428.9163, 
    11.3934, 12.47365, 231.9589, 136.3775, 6.838151, 0, 2.634708, 3.781463, 
    0.1162148, 0.6912898, 0.01993117, 0, 0.4706172, 7.387184, 44.55817, 
    244.1146, 594.9794, 933.8558, 513.5035, 77.61767, 4.361522, 0, 0, 0, 0, 
    0, 0, 0, 0,
  681.6527, 442.5084, 578.8173, 717.4026, 922.1249, 813.6738, 759.1872, 
    525.2695, 321.9953, 302.5872, 458.9889, 403.1359, 243.0368, 181.6122, 
    107.4319, 9.799197, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.0001312634, 0.006848679, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.3214408, 335.2546, 813.2599, 438.9796, 
    1.541609, 0.004860971, 141.2879, 433.2815, 256.4115, 14.89001, 0, 0, 0, 
    0.1404909, 6.80957, 0, 0, 0, 0, 0.4797853, 35.22785, 388.0224, 854.2148, 
    528.0695, 83.28231, 2.967625, 0, 0, 0, 0, 0, 0, 0, 0,
  545.9903, 500.1561, 701.9286, 1102.757, 1219.171, 1147.172, 956.5318, 
    675.6527, 331.725, 351.9229, 475.9785, 420.0756, 313.623, 228.7287, 
    180.0209, 134.015, 0.3182439, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01651771, 0, 0, 0, 0, 0, 0, 22.53872, 
    0.65847, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 30.20723, 195.3939, 
    90.67072, 4.860431, 0, 5.169554, 264.6625, 416.897, 223.7468, 2.467426, 
    0, 0, 0, 0.01299047, 0.1073577, 0, 0, 0, 0, 0, 2.723956, 80.23975, 
    657.4532, 634.125, 285.9821, 125.6809, 2.169004, 0.1452292, 0, 0, 0, 0, 
    0, 0,
  575.7665, 549.1124, 1004.394, 1257.504, 1520.269, 1214.792, 1053.349, 
    760.7601, 506.7095, 417.5125, 432.6968, 399.7943, 364.9707, 304.9736, 
    209.8668, 138.7341, 27.90703, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0001978899, 0.02694878, 0, 0, 0, 0, 0, 
    7.94479, 361.0423, 148.2079, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3.387879, 
    0.004412269, 0, 0, 0, 1.012016, 28.95815, 159.6374, 162.7487, 6.871452, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.002113436, 123.6737, 502.31, 
    321.5427, 69.19288, 34.57666, 4.016514, 0.6476752, 0, 0, 0, 0, 0,
  771.0378, 731.9822, 1232.212, 1579.218, 1810.72, 1665.98, 1247.325, 
    891.9006, 552.7863, 534.0606, 470.0626, 487.2615, 500.9968, 399.5934, 
    301.6216, 216.2957, 101.2677, 1.366401, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7.578414, 0, 10.02934, 
    217.377, 48.73487, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.2398228, 7.076045, 0, 
    0, 0, 0.5435731, 5.565549, 79.59003, 18.13072, 1.341174, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0.07269884, 342.0459, 154.1556, 9.21379, 
    0.01240786, 0.0236598, 5.468072, 10.2199, 0.1744068, 0, 0, 1.12455,
  1005.523, 1089.269, 1428.493, 1729.941, 2157.611, 2366.877, 1791.208, 
    1172.936, 789.075, 679.2053, 769.5369, 774.6565, 661.5249, 538.7116, 
    499.1805, 452.9259, 318.8668, 107.7354, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.003257784, 0, 0, 14.33969, 
    269.4527, 18.4388, 2.629723, 63.20306, 3.818854, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.4436082, 0.4391197, 0, 0, 0, 11.42085, 94.30405, 98.075, 
    0.03083581, 0, 0, 0, 0.03971905, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9.149135e-05, 
    0, 0, 9.795963, 11.95197, 0.4926467, 0.0001121615, 0, 0.0542269, 
    0.1652767, 35.90819, 0, 61.54511, 395.5136,
  1443.506, 1620.422, 1765.2, 1789.817, 2168.043, 2356.399, 1999.072, 
    1344.355, 974.863, 966.6523, 1036.74, 970.4948, 807.8265, 729.062, 
    640.0353, 622.3807, 558.9814, 343.8018, 29.92353, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0003971517, 0.002529405, 0, 0, 
    121.7922, 429.6986, 193.016, 6.398975, 3.334329, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.2867806, 0, 0, 0, 0, 3.61325, 129.9913, 54.15724, 0, 0, 0, 
    0.1055335, 0.3423316, 0.3816859, 0.8894814, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 3.002282, 0, 0, 0, 0, 0, 91.78906, 15.18766, 64.01128, 362.9198,
  1620.956, 2030.3, 1884.991, 2049.509, 2068.68, 2175.013, 1586.164, 
    1522.586, 1346.341, 1360.391, 1342.486, 1150.649, 1009.675, 798.4236, 
    803.64, 793.613, 751.2167, 539.5749, 185.2117, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.00889502, 0.008948714, 0, 1.305878, 
    327.1373, 460.4203, 183.9435, 19.73282, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.001868226, 3.177953, 0, 0, 0, 0, 5.91536, 94.78001, 1.925256, 0, 0, 
    0.02996243, 4.757724, 2.262005, 0.8893167, 0.6945848, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 38.47111, 40.73141, 0, 0, 0, 0, 68.93193, 198.6472, 
    337.3564, 558.7494,
  1649.085, 1708.983, 1942.575, 2064.672, 2304.163, 2042.305, 1346.739, 
    1341.973, 1536.301, 1614.115, 1351.418, 1085.79, 943.1578, 900.9448, 
    952.3292, 1066.381, 834.631, 657.6016, 280.5684, 3.45371, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001200154, 0.001476862, 0, 
    152.6915, 685.7798, 660.864, 391.5136, 81.102, 0.08322787, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.1983324, 8.214144, 0, 0, 0, 0, 7.976196, 96.0976, 
    32.68804, 0, 0, 11.5986, 136.4807, 24.27074, 1.852875, 7.053572, 
    56.97015, 4.038934, 0.03956408, 0, 0, 0, 0, 0, 9.457328e-05, 0, 0, 
    0.1137195, 89.28968, 12.82965, 0, 0.000534966, 0, 0, 46.44008, 85.76493, 
    411.291,
  1466.144, 1621.266, 1631.515, 2122.453, 2175.795, 2267.993, 1097.97, 
    824.9056, 896.3997, 932.9909, 568.8134, 122.1493, 139.7222, 230.9751, 
    585.2339, 743.4264, 595.6318, 653.7233, 457.3597, 15.86434, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.980672, 440.7948, 
    848.3855, 797.6866, 593.3608, 199.7116, 8.479733, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 11.56622, 0.1151541, 0, 0, 0, 11.44357, 154.1412, 126.2073, 
    0.02027015, 0.8643358, 204.4469, 257.3035, 118.653, 15.25982, 90.17926, 
    348.3282, 451.6818, 20.03893, 0, 0, 0, 0, 0, 0.0003784416, 0, 0, 0, 
    0.3295275, 73.48798, 1.209638, 0.001240408, 0.04867897, 35.55901, 
    205.4684, 37.47905, 55.50045,
  1265.107, 1271.335, 1965.781, 1997.247, 2257.103, 2371.452, 1157.836, 
    568.8094, 507.9307, 527.9256, 61.88685, 0, 0, 0, 0, 0, 0, 0, 25.08505, 
    2.611548, 1.012719, 54.77631, 55.46979, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 56.8435, 558.8643, 753.3204, 685.9753, 529.2399, 
    221.9993, 6.638701, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6.390496, 0.1437027, 
    0, 0, 0, 5.025319, 296.0272, 133.192, 26.48146, 105.7203, 124.3082, 
    133.4471, 18.79172, 41.91351, 168.925, 502.5459, 687.1468, 145.1467, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 9.612703, 23.07717, 0.1670243, 0.3258666, 
    40.60841, 178.4189, 98.15704, 58.47993,
  935.9797, 1371.701, 1933.655, 2314.278, 2206.839, 2331.325, 1047.749, 
    519.5513, 454.4148, 405.1205, 26.92118, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 244.4359, 
    576.6982, 579.9873, 438.5885, 334.7599, 131.4858, 3.241302, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.0453538, 0.0158177, 0, 0, 0, 75.12135, 375.2448, 
    88.78672, 19.92136, 145.9868, 126.3988, 55.09162, 79.25726, 93.2966, 
    89.02313, 311.1271, 517.6355, 122.5172, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.03161435, 9.429642, 0.6056394, 0.146424, 207.0213, 126.4081, 45.91529, 
    85.9324,
  705.9424, 1077.602, 1789.276, 2157.059, 2121.644, 2145.599, 927.7297, 
    349.9645, 414.1831, 239.4039, 205.0616, 535.8789, 337.7988, 224.2843, 
    93.21812, 12.07225, 4.108486, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21.81651, 480.2482, 616.3601, 509.2854, 
    411.6318, 353.8981, 172.9756, 23.66262, 1.744636, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.001127199, 0.426254, 0.06272013, 0, 158.0811, 521.639, 
    141.0725, 99.96737, 247.5734, 203.0635, 144.6472, 146.9874, 146.9239, 
    291.5794, 505.7589, 561.468, 82.04576, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    7.754673, 7.457764, 24.7692, 42.12467, 9.055123, 4.078703, 80.82257,
  560.522, 873.38, 1472.261, 1866.38, 1992.183, 1959.356, 668.1165, 250.8919, 
    291.7672, 17.91137, 626.5022, 1631.719, 1588.758, 1237.268, 972.5966, 
    822.8162, 666.3598, 231.6238, 95.20377, 24.35091, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 93.28631, 598.2587, 574.9574, 
    508.1927, 475.7988, 445.4901, 244.6739, 75.22868, 59.67073, 26.13394, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 7.006592, 9.506021, 2.820326, 1.543359, 
    144.5288, 485.7056, 157.8752, 139.0608, 306.2983, 182.6353, 140.4857, 
    150.7803, 237.6682, 550.9364, 811.1963, 598.2958, 25.34849, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 140.1268, 241.5589, 39.90154, 11.41144, 38.09826, 
    75.28021,
  520.9725, 685.0739, 1104.142, 1548.977, 1849.273, 1977.533, 530.145, 
    203.5752, 23.72789, 27.13107, 956.7662, 2034.414, 1627.404, 1195.415, 
    1080.397, 1104.885, 1093.357, 887.1946, 732.5614, 442.7809, 42.32203, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 227.5572, 
    614.1383, 604.0764, 532.1347, 527.2681, 501.3772, 266.3045, 197.5267, 
    319.5226, 439.0925, 52.55056, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01218646, 
    68.76542, 10.88835, 49.6851, 244.7333, 434.6059, 156.4234, 331.7645, 
    396.8661, 241.47, 169.5624, 150.5604, 254.91, 544.6859, 578.8292, 
    122.1243, 0.04935317, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.776042, 
    88.48724, 86.04845, 37.06418, 36.67148, 83.62952, 1.168923,
  520.364, 623.9707, 845.1304, 1182.964, 1794.826, 1631.395, 245.3956, 
    30.59338, 0.1295522, 65.68732, 1191.472, 1929.175, 1380.801, 898.722, 
    945.2995, 1004.129, 951.7753, 889.402, 807.7346, 725.3493, 650.4291, 
    576.4832, 399.0143, 189.4995, 1.069616, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 290.6859, 650.6129, 587.6777, 538.5913, 469.5362, 
    367.0397, 239.3359, 267.2038, 520.4188, 582.6263, 354.7753, 95.80848, 0, 
    0, 0, 0, 0, 0, 0, 0, 10.50261, 205.8622, 156.8265, 367.9012, 536.3768, 
    554.2907, 339.4029, 439.8899, 418.0555, 214.6228, 185.1647, 265.1077, 
    310.9288, 294.0193, 49.32493, 0, 0, 0, 0.0004447775, 0.0008141641, 
    0.0001843075, 0, 0, 0, 0, 0, 0.00153388, 0, 9.762164, 91.66759, 151.5858, 
    43.30084, 69.43888, 56.62251, 23.58093,
  527.755, 558.0959, 777.8425, 1038.259, 1442.285, 857.6389, 34.7822, 
    0.06794915, 0.1317989, 65.86896, 1226.782, 1676.783, 1155.866, 959.6856, 
    863.8164, 851.5259, 757.8932, 699.1624, 691.1156, 647.6199, 588.8004, 
    448.2683, 337.8521, 251.0181, 128.1548, 0.6675929, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 1.583894, 274.4207, 587.1978, 539.9442, 498.1378, 
    401.8043, 324.701, 235.9535, 351.3758, 472.5636, 586.2536, 372.6698, 
    260.64, 20.91498, 0.5449734, 0, 0, 0, 0, 0, 0.1160287, 111.142, 209.0083, 
    276.4948, 646.7979, 765.1041, 724.9354, 477.4805, 577.1857, 463.0179, 
    431.689, 425.1302, 450.4791, 382.4208, 78.48548, 0, 0, 0, 0, 0, 
    0.003998051, 0.002220947, 0, 0, 0, 0, 0, 0, 0, 105.1281, 169.7474, 
    236.0875, 9.81155, 0.1445957, 0, 0,
  489.275, 506.2431, 635.707, 891.2947, 1140.819, 104.9125, 0.5735672, 
    0.0001255112, 2.393601, 199.3139, 1536.486, 1511.392, 1079.511, 820.4056, 
    728.9279, 624.3528, 521.0572, 428.4595, 417.1996, 391.4514, 321.5363, 
    234.6511, 206.3434, 187.8103, 161.0246, 103.9707, 3.567678, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 4.888042, 22.56903, 1.230958, 202.7648, 429.525, 
    412.595, 342.0215, 395.2505, 348.6987, 285.1621, 336.5508, 375.4762, 
    287.4457, 307.1478, 204.0902, 144.1289, 12.40784, 0, 0, 0, 0, 0.09297946, 
    48.31137, 410.1348, 219.7555, 321.0481, 912.0163, 957.0075, 782.5162, 
    689.6246, 672.2351, 803.3319, 900.5595, 921.7489, 653.4254, 113.7043, 0, 
    0, 14.97981, 163.9573, 16.21266, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 34.01518, 
    399.7357, 415.947, 11.40101, 0, 0, 0,
  423.9285, 419.6786, 540.4236, 810.2414, 880.0971, 25.37736, 0, 0, 43.69834, 
    958.8488, 1720.627, 1412.165, 928.663, 770.8799, 633.066, 510.455, 
    402.9467, 319.4293, 278.5269, 235.3018, 194.7553, 149.0402, 112.7481, 
    124.9141, 133.1899, 112.3536, 20.9965, 2.64545, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 2.267793, 70.71137, 122.5515, 31.54795, 87.75684, 313.0298, 326.2078, 
    392.7047, 459.9867, 517.2142, 481.4169, 442.511, 390.7699, 276.8941, 
    289.5733, 344.4179, 305.1668, 167.0574, 9.916601, 1.032431, 1.048887, 
    0.2411555, 23.19702, 397.0361, 721.8358, 320.7461, 332.2949, 979.869, 
    1030.202, 931.765, 809.9, 823.1024, 793.5685, 951.8102, 1033.525, 
    719.0648, 119.1517, 0.833892, 0, 14.80536, 271.7417, 152.8016, 
    0.00275539, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 621.5582, 558.1843, 245.3577, 
    0, 0, 0,
  389.9949, 432.4892, 525.9587, 618.4981, 485.3033, 0.03390811, 0, 1.35604, 
    605.9611, 1549.469, 1794.849, 1175.007, 871.842, 714.1773, 567.928, 
    445.1647, 359.2397, 288.548, 230.5943, 181.9214, 144.2462, 113.5117, 
    92.68795, 83.6313, 99.99515, 113.782, 90.98781, 80.63214, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 10.24857, 59.58021, 91.44401, 35.23301, 92.64501, 269.2377, 
    433.9703, 408.1391, 449.0736, 489.8803, 490.6386, 587.921, 538.6768, 
    542.0423, 504.0613, 493.4232, 387.6947, 149.3013, 21.24825, 2.08333, 
    3.27737, 3.702941, 63.49332, 591.3827, 870.5641, 260.2408, 218.9506, 
    877.173, 980.9655, 1040.86, 1143.761, 991.8488, 921.4819, 835.4803, 
    934.3461, 614.5713, 122.0434, 14.56706, 2.029026, 0, 21.34945, 37.91715, 
    4.003912, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 419.2063, 402.9444, 268.8748, 0, 
    0, 0,
  431.8418, 536.3006, 574.058, 315.8998, 41.75761, 0, 0, 59.75841, 954.189, 
    1557.024, 1298.473, 942.2996, 752.2569, 616.2059, 486.4283, 377.0709, 
    312.1561, 255.6407, 198.0654, 142.262, 116.617, 107.7247, 90.60133, 
    80.00478, 98.95425, 307.284, 343.9886, 272.9455, 6.16348, 0, 0, 0, 0, 0, 
    0, 0, 2.050448, 40.84933, 34.03916, 33.79316, 71.37947, 217.7432, 
    315.7126, 443.3457, 437.9484, 458.0936, 444.2867, 431.0873, 447.9553, 
    504.2306, 471.0587, 559.8055, 493.2112, 392.4747, 196.1293, 47.81644, 
    8.629056, 4.509862, 7.082555, 123.9592, 629.7461, 843.9626, 281.6333, 
    305.7295, 690.8347, 1054.628, 1119.722, 1335.16, 1190.468, 1065.214, 
    984.9171, 869.7607, 546.3845, 225.0289, 150.4363, 163.5934, 3.164987, 
    1.992715, 22.49724, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 167.7594, 192.5879, 
    127.9389, 0, 0, 0,
  464.4328, 710.1633, 619.1936, 47.74748, 0.006608745, 0, 1.039034, 425.7875, 
    1205.512, 1296.795, 937.6955, 818.3823, 688.7088, 615.1889, 470.3323, 
    343.0821, 270.3759, 214.7289, 163.605, 112.6529, 104.0565, 122.8048, 
    107.724, 95.03403, 378.6848, 553.5956, 557.1316, 213.1545, 0, 0, 0, 0, 0, 
    0, 0, 3.253178, 4.987194, 15.42553, 23.11442, 53.14434, 198.1807, 
    390.6396, 476.5912, 416.6757, 370.3962, 423.6606, 388.2758, 315.9665, 
    300.9809, 279.9049, 272.6179, 240.4554, 254.8682, 231.5103, 158.6761, 
    75.81209, 21.71908, 9.130775, 31.90206, 180.6022, 519.5223, 818.9929, 
    367.1069, 232.1573, 540.9075, 1020.897, 1331.289, 1515.057, 1429.161, 
    1326.372, 1300.804, 1167.494, 857.9363, 537.9557, 430.6571, 235.6319, 
    105.8424, 52.64319, 52.60298, 48.16794, 5.177803, 0.0127918, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 7.925615, 7.623189, 0, 0, 0,
  541.9563, 702.7642, 525.0195, 0.008912559, 0, 0.7958623, 220.1246, 
    1012.623, 1381.692, 1054.735, 911.1928, 865.9833, 754.9418, 683.0833, 
    507.5714, 339.2844, 241.6909, 185.5594, 133.8963, 81.90056, 93.08733, 
    116.5835, 104.0461, 220.4304, 362.2358, 272.5128, 22.4466, 0, 0, 0, 0, 0, 
    0.464163, 2.217875, 1.132218, 118.9751, 48.45937, 24.96659, 68.75862, 
    119.5871, 168.0666, 359.0999, 420.4307, 372.978, 292.5229, 326.5298, 
    261.4095, 174.0229, 145.3442, 113.1015, 90.15494, 74.61478, 49.53991, 
    51.27683, 45.57203, 19.36777, 16.3014, 20.58949, 212.4812, 371.5741, 
    567.3152, 837.6189, 773.0519, 254.7844, 402.2862, 1117.507, 1593.182, 
    1713.899, 1657.007, 1585.993, 1660.75, 1626.9, 1297.729, 1008.488, 
    628.0763, 368.5419, 180.6032, 125.0678, 198.4454, 235.6197, 149.7811, 
    32.02615, 2.138504, 0.001609906, 0, 0.0001999206, 0, 0, 0, 0, 0, 
    0.04724865, 3.110864, 0, 0, 0,
  549.2347, 686.2816, 401.375, 0, 0, 65.01826, 822.366, 1329.428, 1219.403, 
    975.2758, 969.5549, 932.9362, 803.3354, 731.2571, 572.4413, 387.7809, 
    255.709, 181.6068, 113.3861, 42.95264, 32.65179, 33.98416, 38.83173, 
    138.7656, 318.7718, 0.7992804, 0, 4.0433, 27.02569, 43.15045, 65.88136, 
    171.93, 328.6717, 326.6402, 310.495, 300.1921, 112.6526, 39.34247, 
    116.7174, 196.2544, 210.7351, 281.5956, 376.5725, 369.3636, 290.0414, 
    245.2731, 172.5113, 134.9192, 115.1656, 85.47749, 72.11951, 66.97635, 
    58.92198, 81.27972, 173.3912, 214.537, 108.2215, 198.1225, 218.5382, 
    378.2805, 263.0815, 752.1837, 870.6851, 687.0273, 413.0518, 1141.952, 
    1943.944, 2054.098, 1926.115, 1828.285, 1968.703, 1788.26, 1402.79, 
    904.152, 675.1245, 442.3218, 270.6985, 164.4036, 201.3591, 233.2095, 
    139.005, 55.39569, 31.88385, 19.8936, 0, 0, 0, 0, 0, 0, 0, 0.36459, 
    2.782869, 0, 0, 0,
  535.8906, 600.8014, 335.9744, 0, 0, 154.2405, 912.732, 1109.16, 989.4586, 
    950.7682, 958.7252, 936.9157, 774.5905, 743.4534, 586.5957, 444.2589, 
    308.8711, 197.4996, 96.48969, 12.3244, 0.1483047, 0.03790293, 0.1436228, 
    37.92851, 155.9851, 30.76747, 221.6138, 252.8131, 416.8718, 624.1976, 
    699.0229, 728.5979, 841.8627, 953.5579, 886.6041, 601.1133, 92.53477, 
    32.85394, 103.7375, 188.0701, 216.8431, 268.9015, 362.442, 393.7513, 
    334.8778, 224.5274, 158.4746, 126.387, 112.2802, 112.7532, 257.5196, 
    397.1968, 538.8138, 1240.1, 2032.906, 2200.138, 2236.536, 1966.697, 
    1706.219, 1459.807, 783.1836, 362.6883, 642.8234, 493.0027, 840.9872, 
    1130.427, 2271.913, 2496.004, 2172.94, 1901.212, 2118.338, 2085.24, 
    1574.87, 1081.068, 810.9539, 635.4389, 423.6662, 250.8699, 288.964, 
    307.7717, 284.6146, 159.4874, 139.9633, 136.567, 123.2743, 19.75318, 0, 
    0, 0, 0, 0, 0, 0.3498602, 0, 0, 0,
  617.859, 478.8044, 162.5502, 0, 0.316467, 273.1028, 967.5567, 1024.078, 
    960.9479, 962.3912, 987.4086, 923.9738, 816.1489, 736.3137, 601.2943, 
    460.8235, 324.0718, 168.9982, 49.51987, 10.05844, 0.003400783, 0, 
    0.6139406, 3.471415, 65.67765, 299.1868, 664.0464, 680.472, 861.0681, 
    1173.805, 1176.411, 882.2818, 935.2615, 1119.443, 1414.621, 875.902, 
    96.9949, 90.53958, 68.45934, 107.9565, 151.2383, 211.1697, 253.7371, 
    301.2069, 273.2981, 195.7737, 154.6178, 177.9713, 194.5825, 716.4048, 
    1805.13, 2597.123, 3127.537, 3920.587, 4658.365, 4768.674, 4483.495, 
    4462.699, 4175.957, 3900.408, 2836.106, 1404.504, 405.8325, 765.2993, 
    1341.417, 1822.338, 2584.409, 2872.491, 2385.164, 1991.338, 2122.929, 
    2156.027, 1849.882, 1308.424, 1070.509, 911.2019, 667.9567, 410.6019, 
    468.2829, 439.6035, 464.8657, 421.4958, 294.738, 311.5735, 259.9264, 
    141.5647, 14.46012, 0, 0, 0, 196.0959, 1.784637, 0, 0, 0, 0,
  589.6921, 369.2813, 29.13641, 0, 10.16494, 462.0075, 953.4734, 992.8953, 
    961.825, 980.4223, 959.9498, 878.5264, 782.0342, 714.8068, 590.7191, 
    438.146, 255.681, 89.16268, 4.204259, 2.031146, 0, 103.8879, 350.6954, 
    283.9107, 257.0193, 369.5965, 704.6323, 645.6995, 1036.557, 1464.105, 
    1060.085, 778.238, 741.6763, 1037.683, 1462.557, 1146.481, 278.6887, 
    344.5007, 247.6657, 85.39928, 122.3622, 162.2269, 193.9326, 217.9708, 
    211.0545, 208.4449, 336.8265, 831.7836, 1583.831, 2516.133, 3871.765, 
    4676.438, 4954.179, 5109.451, 5170.38, 4871.32, 4830.958, 4825.001, 
    4712.904, 4750.763, 4316.47, 2986.506, 1810.279, 1907.389, 3094.098, 
    3158.578, 3400.082, 3428.866, 3037.146, 2417.081, 2381.95, 2137.81, 
    1823.436, 1536.647, 1236.298, 1032.425, 829.5073, 612.1199, 627.1792, 
    549.0421, 514.0405, 437.2412, 523.9689, 332.4905, 376.6574, 324.6547, 
    278.9478, 18.89644, 0.006937383, 11.19048, 622.1964, 266.2146, 0, 0, 0, 0,
  418.7992, 35.6242, 0, 0.003005615, 134.9476, 670.2584, 953.2305, 938.2223, 
    913.4232, 907.8433, 847.9294, 775.7874, 707.1496, 637.6665, 506.9577, 
    328.1991, 144.9271, 21.72296, 0.001061579, 0, 193.2861, 655.1348, 
    890.2563, 1015.931, 1077.46, 1348.436, 1022.688, 766.3108, 1302.777, 
    1343.477, 1030.237, 887.298, 1036.799, 1030.548, 1415.412, 1369.234, 
    954.7562, 897.3719, 604.0056, 161.5459, 117.0032, 160.0316, 186.1864, 
    199.844, 234.4324, 490.8765, 1452.577, 2787.096, 3704.978, 4565.677, 
    5041.605, 5282.9, 5283.827, 5293.211, 5223.339, 5147.862, 5045.44, 
    5014.276, 4810.225, 4833.973, 4828.4, 4279.334, 3368.46, 3630.062, 
    4304.909, 4239.586, 3954.809, 3997.183, 3638.99, 3208.818, 2409.19, 
    1711.776, 1245.757, 1107.457, 1129.331, 956.4644, 789.5651, 568.699, 
    588.8917, 465.5713, 293.4032, 391.9729, 524.9534, 425.9501, 367.7643, 
    501.6449, 504.5149, 232.682, 5.703031, 0.4608422, 517.0116, 853.5552, 0, 
    0, 0, 0,
  208.9919, 0.07399444, 0, 86.20094, 452.0786, 852.0658, 1002.409, 962.3193, 
    888.443, 812.5153, 720.5767, 644.718, 631.5153, 512.2603, 381.4651, 
    213.2256, 41.59562, 0.2816853, 0, 124.2844, 722.3979, 1113.143, 1471.473, 
    1611.769, 2112.062, 2108.031, 1182.046, 772.6594, 1133.844, 1030.302, 
    594.0649, 781.9883, 976.3713, 996.936, 1344.194, 1913.446, 1758.966, 
    1584.213, 828.5089, 218.7474, 120.6228, 168.4115, 186.3442, 204.9695, 
    454.7095, 1957.652, 3490.757, 4445.193, 5092.852, 5200.075, 5270.465, 
    5072.342, 5013.149, 4973.931, 4979.826, 5028.506, 4968.484, 5000.479, 
    4901.846, 4918.038, 5056.896, 4726.156, 4305.746, 4395.774, 4665.846, 
    4441.66, 4191.952, 4342.861, 4170.3, 3571.407, 2256.272, 978.5087, 
    515.0765, 648.3031, 832.2507, 1023.514, 805.8867, 528.6307, 476.446, 
    414.0162, 249.9183, 179.4859, 455.012, 263.6515, 333.0435, 479.9664, 
    632.377, 499.215, 167.3804, 1.14105, 187.7418, 1096.691, 4.065651, 0, 0, 0,
  217.0772, 0.0330215, 14.08818, 507.184, 689.6525, 956.0153, 1135.08, 
    1068.822, 935.9532, 833.0918, 700.9478, 584.4554, 511.998, 405.4882, 
    298.7473, 151.3782, 10.5746, 0, 13.38639, 627.0316, 1415.375, 1796.191, 
    1776.488, 2020.439, 2216.457, 1986.079, 824.9573, 609.1418, 1088.619, 
    704.4744, 531.5552, 655.2637, 836.7814, 991.5665, 1400.434, 1907.079, 
    2138.898, 1730.733, 856.8054, 192.3337, 187.5201, 182.8071, 191.2734, 
    306.0225, 1638.453, 3471.865, 4649.002, 5009.791, 4932.093, 5040.752, 
    4961.458, 4920.357, 4891.655, 4887.036, 4862.397, 4830.989, 4769.84, 
    4764.334, 4749.213, 4840.669, 4871.838, 4824.714, 4635.75, 4551.147, 
    4447.096, 4367.069, 4249.624, 4367.218, 4152.088, 3556.254, 2167.627, 
    517.2781, 330.44, 333.8921, 615.7012, 814.1959, 880.6069, 573.7075, 
    426.0545, 368.3916, 209.4412, 130.0882, 280.0025, 206.5527, 246.2915, 
    389.107, 555.9575, 505.8926, 402.7588, 39.14849, 0.2409696, 211.2308, 
    10.10999, 0.2490215, 8.65174, 0.6303881,
  32.38083, 0, 51.82127, 560.3418, 760.4517, 1012.509, 1175.754, 1092.682, 
    990.1829, 844.8569, 664.1961, 527.9617, 436.3003, 353.342, 264.007, 
    111.6445, 0.1420982, 0, 120.9445, 1149.31, 1999.209, 1945.943, 1973.386, 
    1762.449, 1950.817, 1315.04, 577.0366, 879.3376, 1191.386, 623.9373, 
    548.0479, 722.4045, 1082.094, 1262.284, 1544.662, 2178.558, 2164.37, 
    1978.036, 1035.92, 460.3963, 275.0108, 282.9265, 595.8168, 1425.515, 
    3292.09, 4695.376, 5096.314, 4968.224, 4930.162, 4852.206, 4795.105, 
    4827.783, 4907.193, 5035.4, 4982.63, 5017.723, 4947.738, 4862.034, 
    4921.563, 4884.641, 4879.072, 4878.018, 4793.002, 4559.51, 4386.215, 
    4295.125, 4247.954, 4282.634, 4102.235, 3924.184, 2823.693, 1224.186, 
    358.0084, 332.7956, 348.9137, 678.3985, 848.0242, 821.4729, 618.2599, 
    296.2792, 78.22495, 69.06935, 236.8286, 218.569, 131.588, 226.8546, 
    405.3286, 521.6719, 575.6138, 185.445, 0.1386309, 0, 0.01035178, 0, 0, 
    0.3566946,
  0, 3.552063, 321.7133, 849.3109, 976.9869, 1078, 1041.034, 971.9257, 
    896.7177, 738.8071, 609.843, 479.6385, 370.4907, 299.6009, 196.0335, 
    43.93956, 1.847782, 58.31754, 820.1542, 1913.927, 2158.314, 2047.404, 
    1703.193, 1653.195, 1413.601, 1037.866, 736.9638, 1415.212, 1414.237, 
    810.8496, 802.1318, 1344.746, 1755.177, 1950.15, 2215.817, 2564.552, 
    2719.364, 2259.201, 1462.947, 672.4842, 476.5094, 949.2522, 1674.35, 
    3053.793, 4114.063, 4946.655, 5076.482, 5097.934, 5060.518, 5084.558, 
    5115.013, 5053.414, 5074.056, 5093.611, 5064.592, 5146.818, 5095.178, 
    5143.528, 5132.971, 5072.526, 4904.224, 4783.976, 4806.5, 4586.318, 
    4403.593, 4429.247, 4359.3, 4282.01, 4076.977, 3919.891, 3721.054, 
    2170.56, 812.0792, 348.9857, 379.0044, 509.2384, 835.6813, 1042.576, 
    981.3938, 473.188, 59.4187, 54.51209, 257.2173, 304.478, 147.0937, 
    83.89629, 318.8223, 480.2112, 706.43, 507.7156, 43.1609, 0, 0, 0, 
    0.06568222, 0,
  0, 74.23603, 787.8488, 1047.875, 1021.896, 987.5112, 943.1434, 865.201, 
    751.0483, 636.3491, 527.4158, 403.2906, 282.5342, 179.8925, 87.43723, 
    3.748239, 13.04159, 420.638, 1624.73, 2216.099, 2128.865, 1733.536, 
    1583.128, 1268.357, 1247.077, 910.689, 1149.7, 1639.568, 1381.821, 
    977.155, 1235.957, 1915.405, 2513.842, 2519.291, 2726.454, 3145.376, 
    2913.469, 2521.798, 1770.634, 1137.481, 1062.631, 1737.886, 2865.038, 
    3579.866, 4525.335, 4868.795, 5310.432, 5363.74, 5347.537, 5387.418, 
    5274.167, 5170.409, 5133.905, 5203.841, 5101.455, 5070.62, 5106.412, 
    5089.334, 5089.588, 4879.959, 4693.276, 4713.932, 4758.439, 4678.091, 
    4520.184, 4536.472, 4453.167, 4362.481, 4144.474, 3822.403, 3798.529, 
    3049.53, 1477.426, 703.8835, 612.568, 658.7606, 819.6526, 1062.141, 
    1055.71, 575.3791, 73.42055, 27.57079, 103.5562, 207.4734, 120.4412, 
    30.39635, 148.8998, 383.1422, 591.7628, 532.1869, 174.8339, 1.234607, 0, 
    0, 0, 0,
  6.758009, 487.5991, 1021.831, 1115.679, 886.489, 892.4991, 847.3696, 
    758.7397, 623.5787, 508.0063, 426.4549, 305.7114, 158.1539, 48.50787, 
    5.502139, 5.127207, 40.45427, 1082.158, 2018.84, 2095.057, 1691.412, 
    1381.58, 1191.657, 1015.282, 1019.028, 1079.314, 1296.271, 1340.825, 
    1178.45, 832.3215, 1319.656, 1844.028, 2394.739, 2776.184, 3035.285, 
    3199.43, 3069.708, 2704.726, 3048.322, 2788.972, 2680.07, 3130.915, 
    3342.005, 4203.668, 4655.496, 5272.828, 5415.704, 5200.595, 5129.409, 
    5031.954, 5205.507, 5085.389, 5081.525, 5094.905, 5042.618, 5019.026, 
    4992.753, 5047.111, 5006.662, 4865.849, 4714.873, 4635.37, 4685.44, 
    4620.996, 4597.202, 4502.657, 4462.631, 4332.861, 4098.364, 3766.416, 
    3657.072, 3297.008, 2097.184, 1253.378, 1089.461, 1061.64, 1174.932, 
    1281.606, 1266.194, 835.1642, 263.9403, 79.5519, 32.27344, 68.0872, 
    131.0868, 118.724, 164.2968, 321.6274, 409.3891, 379.2769, 350.8774, 
    57.88399, 0.000805264, 0, 0, 0,
  238.1623, 791.4998, 1109.681, 899.7229, 803.0744, 786.03, 737.5471, 
    634.7917, 498.6732, 393.5605, 324.9799, 180.8011, 45.09904, 5.052932, 
    12.10084, 59.62862, 665.7957, 1742.159, 2304.37, 1936.526, 1518.453, 
    1209.02, 957.4006, 869.3815, 823.4235, 999.6229, 1120.257, 1287.387, 
    1058.116, 943.8759, 842.4662, 1182.286, 1637.921, 2097.368, 2345.563, 
    2374.775, 1990.883, 2252.895, 3334.049, 3940.562, 4061.273, 4010.166, 
    4178.608, 4529.894, 4820.277, 4816.019, 4359.409, 3582.755, 3025.995, 
    3098.254, 3615.333, 4245.46, 4695.494, 5053.856, 5057.838, 5040.737, 
    4995.706, 4951.887, 5012.489, 4828.667, 4652.396, 4480.73, 4422.274, 
    4482.873, 4418.603, 4365.641, 4435.617, 4158.283, 3927.431, 3744.359, 
    3460.329, 3134.216, 2236.319, 1473.672, 1232.209, 1085.229, 938.4994, 
    930.7794, 780.1253, 518.0501, 171.889, 131.0825, 128.4954, 145.3723, 
    306.1799, 273.0995, 216.7841, 302.7602, 352.1556, 292.1012, 300.0482, 
    151.9467, 1.769033, 0, 0, 0,
  762.3385, 958.6488, 967.5426, 836.1221, 672.2523, 743.9036, 705.8074, 
    585.7993, 412.0986, 315.1353, 220.0953, 76.00178, 7.931051, 19.07306, 
    352.5095, 807.7217, 1467.913, 2206.177, 2116.3, 1479.32, 1129.964, 
    788.2949, 807.8799, 715.9404, 766.021, 992.697, 1301.655, 1434.707, 
    1353.936, 786.4489, 618.7448, 572.2695, 753.1136, 781.6061, 869.8459, 
    807.5753, 789.2447, 793.95, 2282.462, 3481.706, 4177.188, 4562.651, 
    4439.226, 4581.507, 3711.448, 2810.206, 2234.735, 1677.431, 1388.387, 
    1278.489, 1672.559, 2128.335, 3001.532, 3830.48, 4550.405, 4801.908, 
    4633.007, 4499.204, 4535.861, 4201.199, 3729.332, 3460.189, 3439.621, 
    3560.627, 3621.553, 3831.16, 4091.066, 3848.02, 3584.761, 3534.397, 
    3254.213, 2773.562, 2217.112, 1683.945, 1579.851, 1373.786, 1237.948, 
    1035.855, 892.402, 538.7142, 249.4172, 148.4552, 154.6931, 130.894, 
    219.8244, 191.3214, 59.69934, 129.1412, 212.872, 166.6351, 130.7894, 
    118.5202, 14.56528, 0, 0, 0,
  989.5663, 927.1322, 930.0528, 724.9628, 672.3023, 786.1067, 760.7014, 
    580.4506, 387.8854, 255.2157, 132.3959, 20.43845, 25.85789, 478.4587, 
    1034.186, 1562.984, 1919.749, 2048.771, 1455.002, 993.2492, 1055.018, 
    1015.837, 1037.239, 1008.556, 891.994, 1129.969, 1403.661, 1486.652, 
    921.8677, 453.2355, 336.5799, 424.1663, 397.4917, 279.882, 307.3911, 
    629.627, 392.5599, 732.6076, 1854.792, 3292.929, 4316.049, 4438.208, 
    4466.581, 3936.618, 2551.772, 1529.796, 1225.804, 1185.416, 1170.846, 
    1186.658, 1149.756, 1173.267, 1364.58, 2012.139, 2864.934, 3708.189, 
    4220.437, 4108.575, 3883.59, 3378.89, 2934.686, 2709.543, 2824.293, 
    3108.43, 3076.333, 3295.794, 3656.051, 3385.662, 3217.673, 3000.589, 
    2639.363, 2225.868, 2004.855, 1872.814, 1614.911, 1220.716, 921.0709, 
    856.4285, 921.3516, 950.4296, 616.0353, 308.2891, 110.1128, 48.46398, 
    55.95203, 45.66961, 26.53019, 25.74332, 58.75687, 44.34055, 7.046542, 
    9.698866, 7.823508, 0.1154567, 0, 0,
  873.5029, 932.446, 802.8636, 679.261, 728.6178, 853.7338, 757.9206, 
    581.5193, 393.3805, 206.899, 67.25694, 23.86274, 177.6185, 981.5392, 
    1598.842, 1796.156, 1947.744, 1703.935, 1375.229, 1515.294, 1642.378, 
    1676.018, 1487.45, 1227.913, 1159.733, 1323.913, 1554.071, 1138.957, 
    556.8956, 169.3183, 218.1516, 265.9337, 235.5797, 302.2885, 690.3524, 
    1159.933, 1460.098, 1501.492, 2359.936, 3452.56, 4296.354, 4520.364, 
    4153.528, 3140.282, 1694.784, 1188.321, 1116.658, 1141.684, 1149.989, 
    1137.289, 1126.685, 1111.867, 1065.968, 976.756, 1235.389, 1905.175, 
    2724.575, 3200.128, 3303.74, 2937.104, 2721.535, 2951.062, 3359.012, 
    3876.756, 3978.864, 3924.08, 3884.962, 3585.292, 3361.129, 3095.249, 
    2504.762, 2074.735, 1898.636, 1876.1, 1742.129, 1328.015, 1136.963, 
    851.3479, 765.448, 628.5696, 611.1027, 228.0393, 106.5588, 40.51612, 
    28.73609, 26.4498, 39.7077, 42.63209, 21.35075, 11.05065, 3.122396, 
    2.336835, 0.5792097, 0.1638553, 0, 0,
  546.0862, 803.7518, 720.4936, 680.9647, 811.3162, 854.0582, 728.9124, 
    554.4362, 350.1646, 161.0941, 51.3675, 48.73245, 369.3617, 1295.04, 
    1821.616, 1891.482, 1897.59, 1783.333, 1780.204, 1693.617, 841.7841, 
    444.8978, 635.6622, 896.0977, 1128.595, 1378.011, 996.2464, 523.0845, 
    123.556, 142.2115, 182.9801, 192.1028, 208.9994, 239.5104, 673.2095, 
    1674.933, 2271.34, 2666.304, 2851.325, 3098.809, 3555.89, 3740.312, 
    3572.558, 2706.249, 1709.02, 1359.368, 1286.218, 1109.896, 1039.783, 
    1053.64, 1038.432, 1022.949, 1007.573, 974.9078, 853.291, 834.8326, 
    1136.756, 1648.817, 2111.175, 2467.282, 2775.722, 3019.613, 3544.646, 
    4111.462, 4240.049, 4245.177, 4150.613, 3692.481, 3492.051, 3113.697, 
    2519.094, 1983.502, 1739.186, 1723.87, 1627.539, 1467.329, 1415.479, 
    1188.471, 862.6572, 819.2594, 613.4723, 440.3748, 103.548, 44.31029, 
    44.08937, 32.32762, 27.8348, 27.06621, 14.8008, 2.686884, 3.042891, 
    2.475014, 0.1258945, 0, 0, 0,
  287.7358, 699.6454, 753.7252, 715.9815, 790.1022, 770.7126, 621.1946, 
    429.5545, 302.6275, 146.0066, 109.7574, 238.4723, 702.8896, 1500.438, 
    1914.869, 1864.13, 1797.373, 1384.315, 1103.181, 50.18019, -29, 
    -28.77262, 25.38564, 296.886, 687.7216, 647.961, 349.3248, 83.32568, 
    112.7014, 157.216, 171.5177, 178.561, 204.0525, 312.3961, 523.767, 
    829.8365, 1039.718, 1047.279, 1355.524, 1172.16, 1411.563, 2336.885, 
    3058.305, 3226.443, 3063.086, 2861.304, 2247.198, 1404.461, 1073.007, 
    987.9013, 956.4599, 926.052, 903.3677, 896.808, 893.4102, 892.0126, 
    796.2086, 820.1337, 984.0677, 1229.673, 1469.496, 1966.5, 2469.902, 
    3181.495, 3622.321, 3652.744, 3231.653, 2652.689, 2285.655, 2040.421, 
    1670.866, 1479.306, 1414.353, 1424.594, 1447.813, 1503.411, 1473.374, 
    1250.532, 1041.187, 973.3618, 1039.013, 789.7152, 424.5931, 71.7645, 
    43.34607, 37.34945, 45.60085, 23.38318, 6.514248, 1.005424, 1.192295, 
    0.07372784, 0, 0, 0, 0,
  280.0255, 717.2288, 800.9051, 767.515, 678.3198, 625.6271, 422.783, 
    283.5512, 241.4006, 186.5598, 174.9805, 521.5108, 1183.758, 1658.958, 
    2034.699, 1761.583, 1296.187, 204.5876, -27.33, -29, -29, -28.70372, 
    31.97342, 167.3994, 247.8943, 170.875, 60.56211, 102.6041, 146.6671, 
    170.812, 176.8664, 183.8537, 244.3707, 366.5971, 502.9418, 470.5995, 
    290.3222, 581.1486, 1270.705, 1402.007, 1254.245, 1784.784, 2600.036, 
    2944.01, 3219.255, 3399.147, 3218.488, 2378.177, 1818.334, 1375.318, 
    1074.772, 1071.595, 984.6507, 961.2864, 971.7458, 1197.327, 1193.799, 
    1028.109, 963.4049, 965.5383, 1135.214, 1159.892, 1419.062, 1704.113, 
    1884.114, 1810.738, 1669.92, 1423.683, 1450.932, 1501.812, 1357.503, 
    1354.311, 1357.144, 1350.14, 1337.69, 1373.946, 1390.578, 1208.278, 
    1047.752, 1206.215, 1150.309, 1096.129, 627.1903, 92.17794, 38.86603, 
    55.03728, 97.46461, 80.68608, 19.16875, 1.530113, 0.02449018, 0, 0, 0, 0, 0,
  278.7002, 848.4108, 836.0483, 703.4719, 592.2507, 425.2289, 267.3521, 
    212.9088, 260.6262, 199.7883, 384.8431, 1051.43, 1458.136, 1718.665, 
    1860.108, 1682.248, 920.7298, -29, -29, -29, -29, -26.10924, 98.29451, 
    120.4517, 76.57224, 60.59356, 87.99368, 121.3795, 137.9679, 144.398, 
    164.9114, 216.217, 274.5612, 275.6122, 318.0442, 259.2065, 230.8655, 
    623.9655, 1918.901, 2278.465, 2228.787, 2412.379, 2568.84, 2575.392, 
    2590.898, 2936.103, 3116.961, 3308.007, 3364.986, 2819.327, 2346.359, 
    2102.324, 1968.311, 1727.268, 1581.183, 1342.206, 1030.278, 1016.645, 
    1021.907, 1084.763, 1044.676, 1257.469, 1468.743, 1774.683, 1740.715, 
    1517.49, 1302.269, 1243.797, 1198.531, 1266.439, 1397.631, 1400.947, 
    1359.057, 1343.482, 1246.818, 1367.203, 1329.797, 1222.678, 1103.928, 
    1230.625, 1299.724, 1154.313, 827.8479, 142.0308, 30.594, 63.95813, 
    176.8368, 209.5096, 94.29587, 2.645784, 0, 0, 0, 0, 0, 0,
  372.7461, 1182.848, 984.7722, 758.8289, 559.1176, 423.6849, 319.4374, 
    300.4261, 340.6555, 502.4338, 1127.504, 1562.021, 1634.167, 1688.647, 
    1848.811, 1538.005, 454.8116, -28.99981, -29, -29, -27.34004, 37.3294, 
    157.3012, 172.0072, 120.2076, 77.74836, 81.51273, 100.2689, 110.1352, 
    113.6465, 112.3892, 174.2308, 265.0841, 238.038, 208.7626, 195.9964, 
    185.5608, 428.3402, 1028.99, 1427.11, 1409.885, 1349.094, 1442.432, 
    1663.696, 1924.178, 2039.838, 2233.458, 2097.392, 2286.286, 2274.246, 
    2335.328, 2740.635, 3043.788, 3113.309, 2620.314, 1823.444, 907.4882, 
    560.1979, 721.8196, 618.8461, 714.8278, 968.9215, 1536.432, 1776.954, 
    1845.922, 1518.606, 1331.444, 1091.121, 1037.558, 1111.581, 1316.298, 
    1388.658, 1346.563, 1293.286, 1239.811, 1305.997, 1406.889, 1326.371, 
    1211.889, 1292.238, 1407.659, 1205.926, 807.7815, 109.0812, 17.7631, 
    51.74597, 188.0972, 276.9687, 185.2122, 45.17762, 0, 0, 0, 0, 0, 0,
  23.64984, 599.7591, 511.6504, 444.8416, 378.2097, 360.2961, 380.9373, 
    438.2814, 595.3414, 1348.148, 2057.229, 2197.964, 1472.968, 1671.91, 
    1237.43, 761.7867, 28.29826, -28.70648, -28.99438, -29, -24.99033, 
    18.25178, 63.3651, 174.8866, 123.8744, 57.97906, 65.55949, 76.69518, 
    97.68421, 102.3149, 131.3378, 195.444, 256.4067, 243.5822, 187.5729, 
    165.1665, 342.9257, 405.3759, 560.9412, 516.8105, 509.3314, 621.6459, 
    699.2636, 746.7856, 760.3452, 922.6527, 823.6852, 1078.508, 1096.203, 
    1233.275, 1588.237, 2370.672, 2694.676, 2629.588, 2156.679, 1783.274, 
    1690.359, 1606.746, 1283.696, 1141.156, 1217.001, 1620.093, 1467.414, 
    1503.383, 1485.695, 1331.391, 1196.225, 1032.619, 951.8022, 972.683, 
    1066.139, 1124.131, 1171.412, 1188.777, 1279.054, 1209.068, 1229.401, 
    1345.554, 1244.472, 1249.917, 1464.447, 1206.628, 878.3694, 171.7012, 
    12.43563, 7.429965, 32.89956, 78.383, 51.98663, 29.90217, 24.32074, 0, 0, 
    0, 0, 0,
  1.67216, 340.6524, 385.0545, 416.1772, 390.3365, 441.3774, 650.9087, 
    704.9575, 1160.624, 1782.02, 2326.5, 2033.687, 1439.484, 1619.828, 
    746.22, 75.66013, 201.0358, 17.39066, -28.43431, -29, -27.93392, 
    -29.96976, 155.6212, 198.6232, 113.8873, 86.04948, 76.57941, 72.31518, 
    72.27863, 74.17043, 85.37265, 140.0728, 171.7061, 157.3423, 148.0897, 
    287.3974, 366.4878, 442.8387, 367.5465, 295.4169, 339.7092, 412.319, 
    477.4836, 479.2714, 430.4697, 594.4115, 1253.493, 1810.096, 2104.204, 
    1634.684, 1001.775, 974.5079, 900.9539, 634.2441, 554.7181, 615.168, 
    911.0193, 996.5089, 1222.358, 1436.428, 1665.35, 1462.017, 1208.923, 
    960.894, 1190.559, 1318.656, 1208.269, 1155.516, 1205.878, 1180.793, 
    1165.779, 1183.944, 1099.437, 1158.785, 1276.583, 1278.646, 1152.482, 
    1210.833, 1241.654, 1143.037, 1397.42, 1334.603, 1178.972, 665.2888, 
    53.88091, 2.508959, 0.1916037, 1.167866, 4.74597, 36.34115, 73.30758, 
    20.18326, 0, 0, 0, 0.04834903 ;
}
