netcdf atmos.1980-1981.aliq.03 {
dimensions:
	time = UNLIMITED ; // (1 currently)
	pfull = 65 ;
	lat = 18 ;
	lon = 29 ;
	bnds = 2 ;
variables:
	float aliq(time, pfull, lat, lon) ;
		aliq:long_name = "Cloud fraction for large-scale liquid clouds" ;
		aliq:units = "dimensionless" ;
		aliq:_FillValue = -999.f ;
		aliq:missing_value = -999.f ;
		aliq:interp_method = "conserve_order2" ;
		aliq:cell_methods = "time: mean within months time: mean over years" ;
		aliq:time_avg_info = "average_T1,average_T2,average_DT" ;
	double average_DT(time) ;
		average_DT:long_name = "Length of average period" ;
		average_DT:units = "days" ;
	double average_T1(time) ;
		average_T1:long_name = "Start time for average period" ;
		average_T1:units = "days since 1979-01-01 00:00:00" ;
	double average_T2(time) ;
		average_T2:long_name = "End time for average period" ;
		average_T2:units = "days since 1979-01-01 00:00:00" ;
	double climatology_bounds(time, bnds) ;
	double lat(lat) ;
		lat:standard_name = "latitude" ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_N" ;
		lat:axis = "Y" ;
		lat:bounds = "lat_bnds" ;
	double lat_bnds(lat, bnds) ;
	double lon(lon) ;
		lon:standard_name = "longitude" ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_E" ;
		lon:axis = "X" ;
		lon:bounds = "lon_bnds" ;
	double lon_bnds(lon, bnds) ;
	double pfull(pfull) ;
		pfull:standard_name = "air_pressure" ;
		pfull:long_name = "ref full pressure level" ;
		pfull:units = "mb" ;
		pfull:positive = "down" ;
		pfull:axis = "Z" ;
	double time(time) ;
		time:standard_name = "time" ;
		time:long_name = "time" ;
		time:climatology = "climatology_bounds" ;
		time:units = "days since 1979-01-01 00:00:00" ;
		time:calendar = "standard" ;
		time:axis = "T" ;

// global attributes:
		:CDI = "Climate Data Interface version 2.4.4 (https://mpimet.mpg.de/cdi)" ;
		:Conventions = "CF-1.6" ;
		:title = "c96L65_am5f9d8r0_amip" ;
		:associated_files = "area: 19800101.grid_spec.nc" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
		:code_release_version = "2024.05" ;
		:git_hash = "5d306c05d9fe755cab04eedc8fd3de0d3c8355a0" ;
		:creationtime = "Mon Aug 25 14:09:46 2025" ;
		:hostname = "pp050" ;
		:history = "Mon Aug 25 13:32:17 2025: ncks -d lat,,,10 -d lon,,,10 atmos.1980-1981.aliq.03.nc reduced/atmos.1980-1981.aliq.03.nc\n",
			"Mon Aug 25 14:40:34 2025: cdo -O -s -select,month=3 merged_output.nc monthly_nc_files/all_years.3.nc\n",
			"Mon Aug 25 14:40:11 2025: cdo -O -s -mergetime /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/shards/ts/regrid-xy/180_288.conserve_order2/atmos_month/P1M/P1Y/atmos_month.198001-198012.aliq.nc /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/shards/ts/regrid-xy/180_288.conserve_order2/atmos_month/P1M/P1Y/atmos_month.198101-198112.aliq.nc merged_output.nc\n",
			"Mon Aug 25 14:12:17 2025: cdo --history splitname 19800101.atmos_month.nc /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/cycle/19800101T0000Z/split/regrid-xy/180_288.conserve_order2/19800101.atmos_month.\n",
			"fregrid --debug --standard_dimension --input_mosaic C96_mosaic.nc --input_dir /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/cycle/19800101T0000Z/history/native --input_file 19800101.atmos_month --associated_file_dir /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/cycle/19800101T0000Z/history/native --interp_method conserve_order2 --remap_file fregrid_remap_file_288_by_180.nc --nlon 288 --nlat 180 --scalar_field (**please see the field list in this file**) --output_file 19800101.atmos_month.nc" ;
		:CDO = "Climate Data Operators version 2.4.4 (https://mpimet.mpg.de/cdo)" ;
		:comment = "FMS time averaging, version 3.0, precision=double" ;
		:NCO = "netCDF Operators version 5.2.4 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco, Citation = 10.1016/j.envsoft.2008.03.004)" ;
data:

 aliq =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, -1.167678e-06, 0, 0, 0.0003133031, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, -4.656631e-06, 0, -2.518695e-06, 0, 0, 0, 0, 0, 0, 0, 0, 
    -3.582196e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 2.737362e-05, 0, -4.020207e-06, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, -3.113808e-06, 0, 0, 0.0004285027, 0.0002200207, 
    0, 0, 0, 7.049155e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 2.533713e-05, -2.140309e-05, 0, -1.284051e-05, 0, 0, 5.345536e-06, 
    -2.010083e-05, 0, 0, 0, 0, -1.601213e-05, 0, 0, -1.488963e-06, 0, 0, 0, 
    0, 0, -1.364201e-05, -1.133428e-05, -1.834142e-05, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 9.59e-05, 0, -2.814145e-05, 3.410475e-05, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0.0002316775, 0, 0, 0.0002927076, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 2.323627e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -6.274212e-06, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, -2.896362e-05, 1.511344e-05, 0, 0, 0, 0, -8.393529e-06, 0, 0, 
    0.001337847, 0.001721214, 0, -7.298218e-06, 0, 0.0001486668, 0, 0, 0, 0, 
    0, 0, 0, 0.0001228599, 0, 0, 0,
  0, 0, -5.472744e-06, -3.083461e-05, 0, -5.197423e-05, -3.869051e-06, 
    0.0006253121, 0.001372957, 0.0001191635, 0, -2.3161e-05, 0.000136254, 
    -4.661256e-05, 0.00038098, 0.00195391, 4.013481e-05, -1.48588e-05, 0, 0, 
    0, 0, 0, -3.063311e-05, -2.761629e-05, -3.533678e-05, 0, 0, 0,
  0, 0, 0, 0, 0, -8.215857e-09, -1.814469e-05, 0, -1.412435e-06, 
    0.0009400687, 0, -7.296129e-05, 2.306214e-06, 0, 0, -2.215634e-07, 
    -1.384842e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0.002031256, 0, 0, 0.0007105857, -5.84886e-05, 0, 0, 
    0, 0, 0, 0, 0, -9.14362e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.042938e-07, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 1.670728e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2.804824e-05, 
    -5.246864e-05, 0, 0, -6.354874e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, -2.857628e-05, 0, -9.224743e-05, 0.001255759, 0, 0, -1.865342e-06, 
    -1.570604e-06, -9.561207e-06, 4.010154e-06, 0, 0.002289978, 0.004081284, 
    -7.851592e-06, -3.143133e-05, -7.435925e-05, 0.0002695633, 0, 0, 0, 0, 0, 
    0, 0, 0.001077963, -8.01412e-05, 0, 0,
  0, 0, 0.0007814702, -3.632447e-05, -2.944591e-06, -8.664257e-05, 
    0.0005788244, 0.001377287, 0.003660522, 0.0009905314, 0, 0.0001923869, 
    0.0005334225, -0.000125869, 0.001301975, 0.003987439, 0.001026125, 
    7.054981e-05, 0, 0, 0, 0, 0, 0.0008543498, 0.000806942, 0.0002939894, 0, 
    0, 0,
  0, 0, -2.262858e-05, 0, 8.215343e-06, -5.5367e-08, -2.385434e-05, 0, 
    6.408382e-06, 0.003480427, 0.001899796, -7.737974e-05, -2.134437e-05, 0, 
    -2.489197e-07, -1.99616e-06, -1.859524e-05, -1.197648e-05, 0, 0, 0, 0, 0, 
    6.948861e-06, 2.095011e-05, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0.005093509, 0, 0, 0.0008247059, -0.0001689593, 
    -4.378277e-06, -1.571152e-06, 0, 0, 0, 0, 0, -4.678643e-05, 0, 0, 0, 0, 
    0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -3.55029e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.849172e-08, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, -4.444747e-06, -3.311027e-07, 0, 0, 0,
  0, 0, -2.060806e-06, 0, 0.0001589071, 0, -2.802608e-06, 0, 0, 0, 0, 0, 0, 
    0.0001084125, 0, -4.759276e-05, 5.34973e-05, 0, 0, -2.144657e-05, 0, 0, 
    0, 0, 0, 0, 0.0002966899, 0, 0,
  0, -9.433745e-05, 0, 0.0001184265, 0.006532815, 0, 0.002088617, 
    -2.432355e-05, -3.214224e-05, -1.561938e-05, 2.926885e-05, 0, 
    0.005753683, 0.005846811, 0.003302899, 9.694599e-05, -0.0002052458, 
    0.0003186326, -4.106138e-06, 0, 0, 0, 0, 0, 0.0002835745, 0.00277189, 
    -0.0001292031, 0, 0,
  0, 0.0002910466, 0.002124045, -4.144767e-05, 5.594439e-07, -0.0001234149, 
    0.001758089, 0.002183879, 0.008368081, 0.001250865, 0.0005376327, 
    0.0002194721, 0.0009340175, 2.93651e-05, 0.001616255, 0.008582564, 
    0.002572548, 0.0004626794, -7.478227e-05, 0, 0, -2.107285e-05, 0, 
    0.002412564, 0.002336607, 0.0006147879, 0, 0, 0,
  0, 0, 0.000726103, 0, 0.0005520397, 4.817934e-05, -1.124449e-05, 0, 
    0.0003458785, 0.006452392, 0.006496461, 4.157343e-05, 0.0004403571, 
    1.241249e-06, -2.490784e-06, -5.059271e-06, -4.210347e-05, -4.143526e-05, 
    0, 0, 0, 0, 0, 0.0003784031, 0.0006260682, -1.222352e-05, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0.005802408, -8.987924e-06, 3.238721e-06, 0.001027824, 
    7.856736e-05, 0.0001718682, -6.569215e-05, -1.554586e-06, 0, 0, 
    0.0002167195, -5.67811e-09, -9.491606e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -3.59747e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -2.422174e-06, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, -2.826991e-07,
  0, 0, 0, -2.406115e-06, -3.252774e-06, -6.726646e-06, -5.89108e-06, 0, 0, 
    0, 0.0002971934, 0, 0, -5.412799e-06, 0, 0, 0, 0.000134312, 0, 0, 0, 
    0.0001484687, 0, 0, 0.0003446862, 0.0006065478, 0, 0, 0,
  0, 0, -4.844525e-05, 0, 0.001203406, 4.21304e-05, 0.00208774, 0, 0, 0, 0, 
    0, -1.009017e-05, 0.002921059, 0, 0.00082016, 0.001289875, 0, 
    -3.327804e-06, 0.0001411187, 0, 0, 0, 0, -2.685391e-07, -9.867743e-06, 
    0.001296045, 0, 0,
  0, 0.0005336081, -9.886857e-07, 0.0004228373, 0.01737272, -3.907696e-06, 
    0.004629515, -0.0001910343, -8.797106e-05, -4.970852e-05, 0.0001051602, 
    -1.401351e-05, 0.01119443, 0.009836077, 0.005676211, 0.005081087, 
    0.0007353971, 0.001145407, -3.695525e-05, 0, 0, 0, 0, 0, 0.001078883, 
    0.005003283, -0.0002505376, 0, 0,
  0, 0.0008677777, 0.003236651, -3.633231e-05, 0.0001040002, -4.740139e-05, 
    0.003292782, 0.003730493, 0.01233478, 0.001939277, 0.001655188, 
    0.002287844, 0.001374723, 0.002703298, 0.002122681, 0.01532741, 
    0.00415433, 0.0007929875, 0.0001589692, 0, 0, -9.41719e-05, 0, 
    0.007287638, 0.004747198, 0.001966579, 0.0004598903, 0, 0,
  0, 0, 0.002671096, 0, 0.001786912, 0.0001207347, 5.163504e-05, 
    -2.788607e-06, 0.001468844, 0.01100031, 0.01141315, 0.0006022485, 
    0.001815352, 6.978046e-05, -8.791119e-06, 0.0002182784, 5.554343e-05, 
    -7.895064e-05, 0, 7.517839e-06, 0, -1.429521e-05, 0, 0.0005566581, 
    0.0009606777, -9.672797e-05, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0.006280792, -4.370275e-05, 1.113017e-05, 0.002255606, 
    0.0005114645, 0.0006185835, 0.0005318393, -2.279781e-05, -5.946228e-05, 
    -1.130804e-05, 0.002617112, 0.0001628825, 0.001075509, 0, -1.447451e-05, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0002230511, -4.357995e-06, 0, 0, 0, 0, 
    0, 0.001347173, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -7.11919e-07, 0, 0, 0, 0, 0, 0.0001826213, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0003269301, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, -3.868508e-05, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 9.329755e-07, 0, 0, 0, 0, 0, 0, 2.382591e-05, 0, 0, 0, 0, 0, 0, 
    0, -4.449007e-05, 0, 0, 0, 0, 0, -7.81902e-06, 0.000183311, 0, 
    -8.480972e-07,
  0, 0, 0, -2.951759e-05, 0.0002283169, -9.523358e-05, -4.110729e-05, 
    -1.141642e-05, 0, -3.946821e-05, 0.0008839407, 0.0003586087, 0, 
    0.0005271913, 0, 0, -2.787156e-05, 0.006421343, -1.316977e-05, 
    -4.094439e-05, -2.971406e-06, 0.002191383, 0, 0, 0.002252599, 
    0.003665166, 7.647708e-05, 0, 2.967878e-05,
  0, 0, -2.014323e-05, -1.613208e-07, 0.00746176, 0.0004703008, 0.009718684, 
    0, -1.960842e-05, 0, 0.0003329534, 0, -8.722347e-05, 0.007257388, 
    -3.169369e-06, 0.002967933, 0.003760973, -6.053033e-05, -7.074528e-05, 
    0.001921223, 7.455426e-05, -2.549992e-05, 0, 0, 0.0005224525, 
    -6.51443e-05, 0.007245751, 0, 0,
  0, 0.001137515, -1.955557e-05, 0.001107833, 0.03131118, 0.0002497816, 
    0.01214102, -0.0001705518, 5.717355e-05, -9.771961e-05, 0.002561143, 
    0.0004936347, 0.01581808, 0.01502424, 0.009092841, 0.01180441, 
    0.002094575, 0.002645711, -8.706627e-05, 0, 0.0001927147, 0, 0, 0, 
    0.002518085, 0.008170258, 0.002103841, 0, 0,
  0, 0.001499706, 0.008383257, -3.270737e-05, 0.0001603708, 0.0006972335, 
    0.007241655, 0.008660658, 0.01889549, 0.003103497, 0.003034333, 
    0.00711011, 0.003048287, 0.006827723, 0.003285816, 0.02762741, 
    0.006039359, 0.001428402, 0.001655768, 0, 0, 0.0005516443, 0, 0.01114685, 
    0.01052739, 0.00333384, 0.002086784, 0, 0,
  0, 0, 0.004778591, -2.197615e-06, 0.00336966, 0.0004842966, 0.0002524789, 
    -1.792387e-05, 0.002326873, 0.01806518, 0.01498458, 0.003766104, 
    0.007021625, 0.0001481695, -3.875263e-05, 0.002489626, 0.0002064635, 
    0.0007895601, 0, 4.734053e-06, 0, -1.945874e-05, 0, 0.001736916, 
    0.001751717, 0.0007983461, 1.141428e-05, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0.006859201, -0.0001511207, 0.001914583, 0.003107162, 
    0.005100723, 0.001444649, 0.002693939, -5.290814e-05, -0.0001955483, 
    -0.0001078309, 0.006570615, 0.0005017368, 0.005601861, 3.597421e-05, 
    -6.05314e-05, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, -9.644678e-08, 0, 0, 0, 0.002054133, -8.490976e-05, 0, 
    0, 0, 0, -1.63552e-05, 0.004240076, -1.355917e-07, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, -4.884766e-06, 4.037682e-06, 0.0001265064, 0, 
    7.681482e-06, 0, 0, 0, 0.003266688, 0, 0, 0, 0, -8.321401e-06, 0, 
    -2.970812e-05, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0009626649, -6.228338e-06, 0, 0, 0, 0, 
    -4.485361e-07, 0, 0, 0, 0, -3.270389e-07, 0.0001311578, -1.318132e-05, 
    7.518483e-05, -5.224295e-06, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0.002376411, -3.876292e-07, -1.234834e-05, -3.243178e-05, 
    0.000250249, 0, 0, 0.001003161, 0, 0, 0.0003949477, 0, 0, 0, 
    -9.049184e-07, 0.001004243, -4.631162e-06, 0, -4.370986e-07, 
    -5.650319e-07, -2.842386e-06, 0.000955881, 0.001191479, -1.293281e-05, 
    0.0002869404,
  0, 0, 0, 0.0004039533, 0.006049193, 0.00166972, 0.002252951, 0.001947712, 
    0, -6.491916e-05, 0.002157978, 0.0008232584, 0.0007388527, 0.001316038, 
    -3.343014e-05, -2.317913e-06, 0.004381827, 0.01470387, 0.0007461791, 
    0.00038009, 0.0002354928, 0.004364151, 0, 0, 0.005031742, 0.008476304, 
    0.005582721, -2.284507e-05, 7.441568e-05,
  0, 0, 0.0002648807, 0.0004284618, 0.01228189, 0.004289979, 0.02239899, 
    -5.860812e-05, 0.000289351, 7.590461e-09, 0.003149354, 3.812078e-07, 
    0.0006761522, 0.02154729, 0.0002793616, 0.01094254, 0.01170012, 
    0.0004871351, 0.003961833, 0.00595115, 0.001933227, -0.0001358927, 0, 0, 
    0.004631027, 0.0009886054, 0.01604441, 0, 0,
  0, 0.005362975, 0.0004336663, 0.005504713, 0.05911029, 0.0009597035, 
    0.02349789, 0.002527667, 0.002880586, -0.0001004412, 0.006387242, 
    0.003102016, 0.02217702, 0.02373777, 0.01705807, 0.0277166, 0.01102138, 
    0.0098275, -0.0002237967, 5.910527e-05, 0.001148585, 0, 0, 0.0001911879, 
    0.006141661, 0.01158884, 0.008293901, 0, 0,
  0, 0.003516169, 0.01673029, 0.0007992586, 0.0007339787, 0.003612383, 
    0.01417929, 0.01602759, 0.02482521, 0.004021013, 0.004301508, 0.01248708, 
    0.006254137, 0.02111372, 0.01141369, 0.04737603, 0.01501493, 0.01121754, 
    0.003523377, 0, 0, 0.0006850396, 0, 0.01717511, 0.02135156, 0.007154971, 
    0.004286432, 0, 0,
  0, 0.0004015239, 0.005577961, 0.0002601359, 0.004918479, 0.004520892, 
    0.003235516, -1.896033e-05, 0.004975462, 0.02816158, 0.01920253, 
    0.01370765, 0.01700273, 0.0003636238, 0.001421652, 0.005082557, 
    0.0004505926, 0.004385224, -4.839408e-07, 0.0005727172, 0, 0.0003364603, 
    0, 0.0097006, 0.005537353, 0.002186762, 7.248401e-06, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0.009118378, 0.0006196515, 0.003946732, 0.00741847, 
    0.01364816, 0.00495326, 0.007538949, -4.466863e-05, 0.0008448485, 
    0.002602537, 0.01380999, 0.004124033, 0.01044505, 0.0001917982, 
    -0.0001464507, -2.906588e-06, 0, 0, 0, -1.667726e-07, 0, -3.913357e-06,
  0, 0, 0, 0, 0, 0, 0, 0.001876102, 0, 0, 0, 0.004896624, 0.002163997, 
    -4.76928e-06, 3.360914e-05, 0, 5.675782e-06, 0.005524504, 0.007908466, 
    -2.536157e-05, 3.094156e-06, 0, 1.183984e-05, 0, 0, 0, 0, 3.314014e-06, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001546993, 0.001643825, 0.00398817, 
    -5.512329e-06, 0.0007145397, 0, 0, -4.762668e-05, 0.009843167, 
    1.796498e-06, 0, 0, -1.131625e-05, -3.456157e-05, -9.824829e-06, 
    4.431064e-05, -3.725447e-06, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, -1.392587e-07, 0.00171272, 0.001130458, 
    0.0008739323, -1.474439e-05, -3.805376e-05, -1.756785e-05, 0.000557313, 
    -2.740269e-06, 2.00783e-05, 0, 0, -6.212292e-05, 0.002922417, 
    0.0004627191, 0.0009278419, 0.000261657, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, -6.610911e-07, -3.315357e-05, 0, 0, 4.944934e-05, 0, 0, 0, 
    -2.804049e-06, 1.677682e-05, 0, 0, -3.934928e-06, 0, 0, 0, 0, 0, 
    -1.344948e-06, 0, 0, 0, 0, 0,
  0.00164603, 5.808306e-05, 0, 0.000268816, 0.006730265, -3.193883e-06, 
    -5.578045e-05, 0.00107191, 0.003079144, 0, 0.0002196334, 0.001722993, 
    1.179004e-05, 0.0003786883, 0.001379759, -4.760622e-05, 0.0005909358, 
    0.002743006, 0.003316043, 0.004044859, 0.0008390628, 0.0006780043, 
    7.901114e-05, 0.0004549231, 3.623662e-05, 0.00326152, 0.006276483, 
    0.0003452578, 0.002846448,
  0.00135794, -0.000124288, 0, 0.00119823, 0.008551953, 0.009810917, 
    0.005811653, 0.006092805, 0, 0.002112972, 0.007183305, 0.001364886, 
    0.005065574, 0.005872103, 0.0009112369, -9.996151e-05, 0.01540454, 
    0.02706327, 0.003934645, 0.007278206, 0.003705853, 0.01124886, 
    7.457408e-06, 0, 0.009240425, 0.01609119, 0.01581611, 0.0001658439, 
    0.00153223,
  0, 0, 0.002247402, 0.004162457, 0.01744811, 0.009672066, 0.04718139, 
    0.001189287, 0.004341643, 5.276413e-05, 0.00993365, -3.929918e-06, 
    0.003690798, 0.03079222, 0.007630326, 0.028984, 0.03130296, 0.005225899, 
    0.02098715, 0.008555426, 0.01072003, -9.207703e-06, 0, 0, 0.01136738, 
    0.00616846, 0.03182917, -1.227713e-05, 8.07429e-07,
  0, 0.01244602, 0.001938009, 0.01371405, 0.1010559, 0.005516652, 0.03349884, 
    0.007018284, 0.008488383, 0.0002264748, 0.01749813, 0.005731656, 
    0.02628946, 0.032231, 0.02871703, 0.05853508, 0.03397539, 0.02103134, 
    0.001249262, 0.0007313457, 0.004851398, 0, 0, 0.002009115, 0.01084412, 
    0.02268583, 0.02692208, -1.356908e-06, 0,
  0, 0.01171185, 0.03119481, 0.00737701, 0.009036839, 0.01117207, 0.02660206, 
    0.02986705, 0.04740201, 0.006376284, 0.007585667, 0.03255936, 0.01644542, 
    0.04042039, 0.03819922, 0.07284848, 0.0283211, 0.02318946, 0.005757311, 
    -3.470604e-06, -6.876142e-06, 0.001733716, -3.815398e-06, 0.05031497, 
    0.06353143, 0.01925063, 0.005234162, -2.853782e-08, 0,
  0, 0.001667301, 0.007418589, 0.0002482989, 0.01186893, 0.01141652, 
    0.0155653, 0.0004630919, 0.02009662, 0.06504433, 0.02543517, 0.02381887, 
    0.04168209, 0.01736839, 0.01564412, 0.01166746, 0.002756394, 0.01182063, 
    3.782478e-05, 0.002554154, -4.14116e-08, 0.002362449, 4.822591e-07, 
    0.02920549, 0.01274808, 0.009934024, 3.595611e-05, -3.440479e-06, 
    -1.724577e-11,
  -7.206913e-10, 0, -2.813406e-06, 0, -1.440965e-07, -1.670094e-07, 
    1.300277e-05, 0.01477135, 0.00212966, 0.005334059, 0.02021226, 
    0.03066084, 0.01358628, 0.0152162, 0.0005900695, 0.006468547, 
    0.007846328, 0.02699049, 0.01118644, 0.01465315, 0.001625095, 
    -0.0001220035, -1.365068e-05, -1.842282e-10, -6.558744e-07, 
    -2.704421e-08, -1.011482e-08, 0, -1.383374e-05,
  0, 0, 0, 1.768236e-05, 0, 1.457691e-08, 5.910768e-06, 0.00416343, 
    -1.367647e-06, 0, 0, 0.008855041, 0.005500121, 7.018932e-05, 
    0.0004700461, -7.752958e-06, 0.0004117665, 0.02112611, 0.0251416, 
    0.005970576, 0.005323808, 0.0007785294, 0.00123567, 2.974691e-08, 0, 
    -3.340107e-08, 2.234241e-05, 0.001853048, 0,
  0, 0, 0, 0, 0, 0, 0, -1.176103e-05, 0, 0.004443945, 0.006432289, 
    0.01121744, 0.0007765846, 0.002480751, -1.950855e-09, -2.080374e-05, 
    -4.925349e-05, 0.0129818, 0.001135933, -6.496571e-05, -2.492954e-05, 
    -1.931027e-05, 0.0005906087, -4.661312e-05, 0.0007428665, 0.001358567, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, -2.025368e-05, 0.002777151, 0.004079324, 
    0.002401347, 0.00131051, 0.001389527, 0.001607934, 0.004073334, 
    0.0004260068, 0.0007197127, -1.478432e-05, 0, 0.002579726, 0.00967473, 
    0.006122513, 0.005184468, 0.001189756, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -3.969525e-06, 0, 0, 0, 0, 0, 0, 
    0, 0.000100332, 0, 0, 0.001856278, -1.58369e-06, 2.976638e-05, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.587302e-05, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 6.306899e-05, 0.002698239, 0.0001669516, 0, 0, 0.001383022, 0, 
    0, -2.74972e-05, 0.0006802324, 0.005317842, 0, 0.0001633115, 
    0.0005165605, -2.959319e-05, 1.262786e-05, 1.504283e-05, 0, 
    -1.242362e-05, 0.0005337982, 0, 0, -2.957577e-05, 0, 0,
  0.005030479, 0.00214017, 0.0004423752, 0.003333448, 0.01587755, 
    0.002252442, 0.001246633, 0.002772409, 0.008039236, 0.001410546, 
    0.001586885, 0.001761217, 0.001670415, 0.003853999, 0.00417027, 
    0.0001996661, 0.003297956, 0.0100139, 0.008972941, 0.0114897, 
    0.004213332, 0.006327784, 0.006630006, 0.004285163, 0.0009231301, 
    0.01066814, 0.01940945, 0.008612425, 0.005537166,
  0.006674461, 0.001301888, 0.0001725578, 0.004108464, 0.01458572, 
    0.02629485, 0.01725284, 0.0109916, 0.0001694813, 0.008233239, 0.01446011, 
    0.005821148, 0.007809352, 0.01762916, 0.006813966, 0.002349266, 
    0.02320312, 0.04829752, 0.01730267, 0.02169849, 0.01773322, 0.02032623, 
    0.0004481671, -1.315829e-05, 0.01343586, 0.02901075, 0.03977325, 
    0.00463124, 0.0158374,
  -3.466208e-05, -7.793285e-09, 0.004862938, 0.01300847, 0.02043831, 
    0.02418784, 0.08986327, 0.008546876, 0.0143348, 0.001584557, 0.01842141, 
    0.00122421, 0.005779706, 0.04394835, 0.04184751, 0.06198717, 0.0653021, 
    0.03229626, 0.03662354, 0.02125922, 0.02422375, 0.001803703, 
    -1.239044e-05, 3.485935e-05, 0.01905345, 0.02134752, 0.06547181, 
    0.0007197757, 0.0001739453,
  -3.101697e-09, 0.03301619, 0.008003982, 0.0685287, 0.1820525, 0.04668441, 
    0.05566237, 0.01959949, 0.06665433, 0.01228144, 0.05858712, 0.01909311, 
    0.03501296, 0.08181628, 0.1347527, 0.124611, 0.07296511, 0.07134477, 
    0.005783323, 0.003199304, 0.01006648, -1.010208e-10, -0.0001066544, 
    0.0343987, 0.08125072, 0.03533743, 0.04689211, -4.51165e-05, 0,
  -1.499644e-06, 0.03626691, 0.1046437, 0.03414272, 0.06363836, 0.05329493, 
    0.08664419, 0.08662018, 0.1599836, 0.04858337, 0.02035424, 0.1580118, 
    0.1199244, 0.1781962, 0.1687032, 0.1360161, 0.1153188, 0.05972718, 
    0.02137258, -2.217394e-05, 0.0003697872, 0.005573807, 0.001582433, 
    0.1541922, 0.2668415, 0.07461026, 0.01348534, 2.554803e-05, -8.32102e-11,
  -1.24171e-06, 0.01064166, 0.03375117, 0.003154152, 0.02618154, 0.02770631, 
    0.04529752, 0.03308255, 0.06412429, 0.1421287, 0.06630985, 0.09405822, 
    0.1502567, 0.1398949, 0.1644568, 0.0832504, 0.02944787, 0.02368282, 
    0.0002103676, 0.007867056, -0.0001073624, 0.01007619, 0.0001259293, 
    0.1270873, 0.08610035, 0.05153849, 0.003278518, 5.700856e-05, 
    -5.559337e-06,
  -2.260542e-05, -6.796971e-06, 0.0008257626, 0, -1.062572e-06, 
    -1.674418e-05, 0.0005672381, 0.03829993, 0.01708648, 0.03295064, 
    0.06049852, 0.08242448, 0.08673833, 0.04558724, 0.02761876, 0.0306516, 
    0.02150874, 0.04189156, 0.02158361, 0.02091289, 0.0061386, 0.0006940301, 
    0.0007768868, 2.99962e-07, -3.656801e-06, 0.0001218282, 0.0002262015, 
    2.358049e-05, -7.439985e-05,
  -9.316022e-12, -5.09286e-08, -2.207263e-08, 2.097108e-05, 2.717891e-10, 
    8.496735e-05, 0.001861082, 0.006058302, 0.0006102927, 2.450411e-05, 
    8.805103e-06, 0.01268944, 0.0141242, 0.001826856, 0.0003067112, 
    -1.286407e-05, 0.003549556, 0.04298368, 0.06365909, 0.01533945, 
    0.02213561, 0.0107549, 0.003964613, 2.702248e-05, 0.0001322232, 
    6.180571e-06, 0.0004238581, 0.004553743, -1.445283e-05,
  0, 0, 0, 0, -1.000733e-05, 0, -2.279553e-11, -6.029914e-05, -3.554075e-05, 
    0.01597971, 0.0175768, 0.01935157, 0.00274137, 0.004012098, 5.635778e-05, 
    -8.801759e-05, 0.001529922, 0.01679858, 0.006918615, 0.0008176714, 
    -0.0001075417, 0.009326877, 0.001876527, 0.004368401, 0.005659554, 
    0.007187382, 0.0005272388, -1.986387e-09, 0,
  0, 0, 0, 0, -1.693972e-05, 0, 0, 0, 0, 3.362211e-06, 0.005407168, 
    0.005927963, 0.004669227, 0.00782266, 0.007936236, 0.005654701, 
    0.009267589, 0.004406852, 0.001724554, -4.904579e-05, 0, 0.006271049, 
    0.02224984, 0.01888607, 0.01419467, 0.01443671, -1.931445e-06, 
    -4.398732e-06, 6.444873e-06,
  0, 0, 1.950217e-05, 0, 0, 2.202826e-05, 0, 0, 0, 0, 0, 0, 0, 0, 
    -1.029979e-05, 0, 0, 0, 1.396722e-05, 7.610746e-05, 0, 0, 0.0006538208, 
    6.13554e-05, 2.639335e-05, 0.003261666, 2.069177e-05, 0.001124532, 
    6.637531e-06,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -5.090976e-06, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, -2.212517e-05, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3.843049e-05, -2.080244e-05, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0002447772, 8.804181e-06, 0, 
    0.001368471, 1.612157e-05, 0.0001078381, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  -1.137701e-05, -4.483242e-07, 0.0003024648, 0, 0.001204851, 0.007535421, 
    0.0004239776, 9.610683e-07, 0, 0.001594789, -1.86015e-05, 4.469004e-05, 
    0.002339219, 0.002741297, 0.007628886, -3.268499e-05, 0.001662159, 
    0.002598299, 0.00182578, 0.002615171, 0.001721906, 2.304471e-05, 
    0.001432368, 0.002153471, 0.001896595, -3.95321e-05, -0.0001012451, 
    2.430606e-05, 0.0002528256,
  0.01591365, 0.008694343, 0.00225182, 0.007546179, 0.03149997, 0.01177161, 
    0.002964226, 0.006482673, 0.01087469, 0.002004198, 0.005509738, 
    0.002285327, 0.004821584, 0.007018783, 0.01528196, 0.003496672, 
    0.01042533, 0.02049087, 0.02543574, 0.02810179, 0.01151029, 0.01513736, 
    0.0207966, 0.01110322, 0.002971713, 0.02669469, 0.03133792, 0.01948052, 
    0.01179682,
  0.01664595, 0.007056844, 0.001071586, 0.01342409, 0.02804888, 0.04687279, 
    0.03705992, 0.02274352, 0.0009636382, 0.01202866, 0.0221999, 0.01008279, 
    0.01155848, 0.03369378, 0.0281109, 0.03545683, 0.04650552, 0.1020327, 
    0.07932553, 0.06027405, 0.05169617, 0.04255316, 0.002928127, 
    0.0003373949, 0.02415349, 0.0426592, 0.08592196, 0.05401226, 0.03709534,
  0.004602778, 0.0002617593, 0.01403499, 0.05523254, 0.09103892, 0.1514642, 
    0.2046625, 0.07292808, 0.06073176, 0.0415315, 0.07322511, 0.04102069, 
    0.01480813, 0.07306544, 0.09815477, 0.1291068, 0.1343715, 0.1922895, 
    0.1562834, 0.05862711, 0.04480748, 0.03333662, 0.0003844977, 0.01038006, 
    0.05405541, 0.06250328, 0.2026351, 0.05649132, 0.02012933,
  6.435357e-07, 0.08072905, 0.06810077, 0.07007109, 0.2116985, 0.06841721, 
    0.06784405, 0.04506788, 0.1107939, 0.0201184, 0.1170039, 0.04035862, 
    0.03710548, 0.08207259, 0.1580331, 0.1383329, 0.1298138, 0.1301874, 
    0.08478373, 0.06897623, 0.0203491, 0.0001487051, 0.02684587, 0.03711281, 
    0.1144921, 0.1857713, 0.1409778, 0.06798235, -1.614847e-05,
  0.006031537, 0.08400492, 0.3882363, 0.1830243, 0.1079178, 0.08817931, 
    0.1138703, 0.1513029, 0.1689829, 0.06037201, 0.02792571, 0.1386204, 
    0.1020225, 0.146571, 0.1437994, 0.134844, 0.1800706, 0.09160303, 
    0.07855044, 0.04046159, 0.005332297, 0.004137087, 0.007748067, 0.3341978, 
    0.3758829, 0.310884, 0.1129615, 0.01457942, 0.0002095332,
  0.001559961, 0.1710512, 0.3480343, 0.0378709, 0.08736931, 0.08237407, 
    0.1586008, 0.1592628, 0.2307343, 0.3407616, 0.08289118, 0.1150855, 
    0.1406203, 0.1316344, 0.127079, 0.08717507, 0.02884252, 0.02928719, 
    0.001303782, 0.01919058, 0.006013183, 0.01053152, 0.03260687, 0.3290152, 
    0.2549413, 0.1667939, 0.1279241, 0.02571829, 0.0005540076,
  0.01647525, 0.001490735, 0.03049802, -2.663978e-10, -0.0001068234, 
    0.001023881, 0.01146074, 0.05783493, 0.022372, 0.03272329, 0.07065383, 
    0.07826302, 0.07073209, 0.04052529, 0.01576829, 0.03410726, 0.05408303, 
    0.1094103, 0.05723814, 0.1011138, 0.1497724, 0.02887632, 0.01738131, 
    0.0002933387, 0.0005518197, 0.01142065, 0.0006071001, 0.03046882, 
    0.009655957,
  0.0006599247, 0.0002708789, -1.384215e-05, 0.003337875, 3.673728e-07, 
    0.003973956, 0.01273424, 0.008439773, 0.004020602, 0.0095403, 
    0.005982093, 0.01412505, 0.02634391, 0.003478492, 0.005791145, 
    0.01131661, 0.02330996, 0.09443274, 0.1861835, 0.08309526, 0.1720636, 
    0.07176068, 0.008450986, 0.002379002, 0.001748363, 0.0006621775, 
    0.00671561, 0.03015645, 0.001668771,
  -1.781339e-08, -3.523183e-09, 9.20284e-06, 4.751438e-08, 1.115356e-05, 
    -2.510779e-07, 1.910705e-05, 7.121505e-05, 0.0004649823, 0.03998359, 
    0.04124127, 0.0409474, 0.01781418, 0.01923967, 0.01151688, 0.005489873, 
    0.01323437, 0.02347483, 0.01508595, 0.007096577, 0.001445202, 0.04314159, 
    0.02883847, 0.02194486, 0.01837514, 0.01443043, 0.003959636, 0.002041, 0,
  -7.463214e-07, 0, 0, 0, 0.0009166814, -1.718953e-08, 7.420331e-06, 0, 
    -1.616755e-06, 0.001659913, 0.007377033, 0.01436237, 0.01638491, 
    0.02725095, 0.02087126, 0.0194182, 0.01916199, 0.01497107, 0.00764308, 
    0.0002638294, 0, 0.0100858, 0.03426135, 0.03416449, 0.03251721, 
    0.03380499, 0.0005918849, 0.003443601, 0.0002472294,
  0, 0, 0.0001908964, 0, 0, 0.000452865, 0, 0, 0, 0, 0, 0, 0, -6.647754e-07, 
    0.0009657277, 4.776045e-06, 8.509079e-05, 0.0008013521, 0.001516682, 
    0.0004306297, 0, 0, 0.004666815, 0.001782099, 0.001505904, 0.0127877, 
    0.003945958, 0.003730104, 0.001570756,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -9.123931e-06, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.0009500925, 0.0002027233, 0.0006191827, 0.000180053,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0002984421, 0.0002642136, 
    1.369567e-05, -3.504582e-07, 0, 0, 0.000116333, 0.0001627234, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, -1.175123e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0.002541051, 
    0.001159911, 0.0006523423, 0.003029638, 0.007889527, 0.01321736, 
    0.001940412, 0.002871573, 0.0001077929, 0.0004718352, 9.51439e-05, 0, 0, 
    -9.349474e-05, 0,
  0.0007280795, 0.004011745, 0.0003631334, -5.763688e-06, 0.003516258, 
    0.008594814, 0.004202654, 0.000380201, -2.240812e-06, 0.003626738, 
    0.0002689848, 0.001119192, 0.007466704, 0.008757423, 0.01078559, 
    0.001034684, 0.004776443, 0.01334269, 0.01251479, 0.01032516, 
    0.005970792, 0.001563665, 0.005453385, 0.007480065, 0.007677763, 
    0.0004141821, 0.00193455, 0.005379904, 0.0003967605,
  0.07168794, 0.04809924, 0.01521022, 0.02368987, 0.06702576, 0.03980979, 
    0.03191157, 0.04459079, 0.0347833, 0.0282119, 0.007793886, 0.01306101, 
    0.007831659, 0.01372196, 0.03659639, 0.01743568, 0.03173549, 0.02857368, 
    0.04876664, 0.08421589, 0.07857709, 0.04843102, 0.0573664, 0.02776951, 
    0.02330951, 0.0743193, 0.0653998, 0.05177744, 0.07037315,
  0.1139236, 0.05788288, 0.05967563, 0.09470569, 0.07675526, 0.1206072, 
    0.11631, 0.0743834, 0.06000229, 0.05965822, 0.07006907, 0.06032316, 
    0.05336231, 0.09224641, 0.05614442, 0.1000293, 0.05892025, 0.1537674, 
    0.1351747, 0.1575746, 0.1495079, 0.138427, 0.05416979, 0.007260783, 
    0.05771169, 0.08707422, 0.124662, 0.1522209, 0.1043655,
  0.00402511, 0.0109084, 0.07689853, 0.06296141, 0.09577949, 0.1533959, 
    0.233635, 0.1144848, 0.08716674, 0.06629609, 0.1350782, 0.07366027, 
    0.0408718, 0.1037212, 0.08317231, 0.1310328, 0.1271377, 0.1853762, 
    0.16604, 0.1192351, 0.1447973, 0.05642028, 0.009575346, 0.01700037, 
    0.06830847, 0.07875258, 0.2298465, 0.1080599, 0.02640821,
  -1.587664e-07, 0.06930916, 0.05379299, 0.0608032, 0.1898093, 0.05300621, 
    0.06036782, 0.03306917, 0.09412794, 0.01597048, 0.107136, 0.0294689, 
    0.02894832, 0.06499857, 0.1272986, 0.1200865, 0.1110713, 0.107412, 
    0.07101699, 0.05024064, 0.07832955, 0.006930455, 0.0125488, 0.02659213, 
    0.09944607, 0.1783428, 0.1215319, 0.06334276, 1.230034e-05,
  0.000986593, 0.05508309, 0.3655728, 0.1519425, 0.0651921, 0.06170145, 
    0.0864993, 0.1106784, 0.1466454, 0.04483135, 0.02421999, 0.1102233, 
    0.07884342, 0.1176707, 0.1226766, 0.1258232, 0.1420238, 0.07499642, 
    0.07239187, 0.02357385, 0.001035232, 0.001967877, 0.005176132, 0.3042946, 
    0.3148564, 0.266684, 0.08236386, 0.005258033, 4.67161e-05,
  0.00056341, 0.1153344, 0.2365061, 0.03429711, 0.05249402, 0.06018875, 
    0.1094561, 0.1064891, 0.1841173, 0.2870597, 0.05381295, 0.08155449, 
    0.1018842, 0.09274772, 0.09402257, 0.06211719, 0.01537885, 0.02080397, 
    0.002996937, 0.01202984, 0.0009387163, 0.004309104, 0.01016588, 
    0.2396927, 0.1889735, 0.1187712, 0.08813421, 0.006603717, 0.001258892,
  0.01614983, 0.0001759687, 0.02077034, 3.64029e-05, -5.087938e-06, 
    0.002229108, 0.008448787, 0.04833645, 0.01346203, 0.01888114, 0.05045278, 
    0.05595645, 0.05954182, 0.04164725, 0.01316418, 0.03152876, 0.05001404, 
    0.1042144, 0.04516025, 0.06655071, 0.09888498, 0.01327109, 0.006070041, 
    0.0001766518, 0.0001338281, 0.008942059, -0.0001200087, 0.01114047, 
    0.01331525,
  0.0837969, 0.02941365, 0.009605657, 0.0006688841, 1.126298e-06, 
    0.006575979, 0.01104977, 0.01462797, 0.01365052, 0.01055596, 0.01752492, 
    0.01874429, 0.03180787, 0.008432579, 0.02479224, 0.01030698, 0.04557902, 
    0.0915025, 0.2010734, 0.09914428, 0.1587018, 0.07240342, 0.007515122, 
    0.0006036889, 0.007704184, 0.0208436, 0.02383932, 0.06326634, 0.1014673,
  0.001516667, -0.0003487803, 0.01742055, 9.181078e-05, 0.00201596, 
    -9.537835e-06, 0.001108743, 0.0001526941, 0.002341216, 0.09161947, 
    0.1257906, 0.1248415, 0.07254129, 0.07447075, 0.07930329, 0.02887179, 
    0.05468779, 0.06542771, 0.06073024, 0.04325702, 0.02117628, 0.1448698, 
    0.1303498, 0.141491, 0.1442145, 0.1057933, 0.03717565, 0.007174484, 
    -0.0001585821,
  0.0002615225, 0.0001281166, 3.936887e-06, 0.0002043666, 0.006891603, 
    -2.056545e-06, 6.839624e-05, -1.358035e-05, -6.440613e-06, 0.00523382, 
    0.01169944, 0.02540843, 0.04265393, 0.05048835, 0.04511556, 0.03620319, 
    0.04307512, 0.04439051, 0.02327267, 0.004748151, 0, 0.01643095, 
    0.0533479, 0.06736567, 0.07876178, 0.09033328, 0.01470552, 0.01257208, 
    0.001475749,
  0.003926467, -5.353164e-07, 0.0007746005, 0.0005423713, 0.0004430011, 
    0.0007843723, -1.087712e-06, 0, 0, 0, 0, 0, 5.530164e-05, 0.000434437, 
    0.00343941, 0.003967987, 0.002326492, 0.00374478, 0.005835083, 
    0.000446726, -2.095125e-05, -2.056685e-05, 0.007541582, 0.004233795, 
    0.006893825, 0.03249253, 0.01354481, 0.0101249, 0.007829645,
  -2.241457e-05, -2.007175e-05, 0, 5.183111e-05, 0, -8.408259e-06, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 3.363254e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.002025001, 
    0.003715467, 0.003738776, 0.0006070534,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, -5.183047e-06, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0.0002259922, 0.001206941, 
    0.0009039008, 3.183147e-05, -7.704105e-06, 0, 0, 0.0005196861, 
    0.0003236462, -9.845557e-06, 0, 0, 0, 0,
  0, 0, 0, 0, 1.739909e-07, 0.0003898744, 0.0002991136, 0, 0, -1.889935e-05, 
    -8.024661e-07, -2.858369e-05, -1.164322e-06, 0.0003442393, 0.003608285, 
    0.002747873, 0.008443761, 0.01568933, 0.02385475, 0.04153227, 0.0232064, 
    0.0200419, 0.007591906, 0.009782442, 0.001354295, 8.639624e-07, 
    0.0001554149, 0.0004489264, 0,
  0.01048416, 0.01063203, 0.006162343, 0.002848709, 0.02081525, 0.02252158, 
    0.02770789, 0.02301802, 0.004049947, 0.01660397, 0.02141031, 0.01084354, 
    0.02881584, 0.04341258, 0.05656008, 0.03433498, 0.02812187, 0.03330427, 
    0.02721534, 0.03462963, 0.02334812, 0.009709538, 0.01944623, 0.02224168, 
    0.03360343, 0.02987306, 0.01522775, 0.01767972, 0.007969759,
  0.1348865, 0.1158931, 0.1045621, 0.1426351, 0.1763792, 0.1527388, 
    0.1185251, 0.1138795, 0.1157337, 0.08185835, 0.06998471, 0.07822278, 
    0.08401917, 0.08256195, 0.08947838, 0.0576176, 0.07147656, 0.06642147, 
    0.1004714, 0.1049594, 0.1363471, 0.09739661, 0.1434985, 0.07076397, 
    0.08589274, 0.1862721, 0.1308485, 0.08871967, 0.1311595,
  0.1142906, 0.08192943, 0.06250427, 0.08013031, 0.08381258, 0.1163169, 
    0.101183, 0.08956406, 0.08322937, 0.08828835, 0.1203013, 0.1061937, 
    0.1042802, 0.1373685, 0.1155028, 0.09699561, 0.09683342, 0.1619226, 
    0.1421513, 0.153921, 0.175091, 0.1528424, 0.06410364, 0.02793116, 
    0.08411296, 0.1050099, 0.1254225, 0.1477586, 0.1049942,
  0.004427644, 0.007874617, 0.09496336, 0.05551068, 0.07392412, 0.1357802, 
    0.2125309, 0.09483041, 0.07103042, 0.07113495, 0.1519804, 0.06926512, 
    0.04260021, 0.09602451, 0.06537365, 0.1156959, 0.1107933, 0.1748927, 
    0.1426451, 0.1038018, 0.1201956, 0.07045102, 0.01016783, 0.009422378, 
    0.05235825, 0.07966177, 0.2158058, 0.07559356, 0.01971386,
  -5.999167e-06, 0.06366274, 0.04507418, 0.05079251, 0.17964, 0.05171967, 
    0.0545024, 0.02235112, 0.07866167, 0.01671302, 0.0963968, 0.02570412, 
    0.02415521, 0.05947182, 0.1158967, 0.1118679, 0.1038003, 0.08936326, 
    0.06740347, 0.02860952, 0.05534618, 0.006831059, 0.003963592, 0.01970315, 
    0.0858074, 0.1660161, 0.09944558, 0.03578481, 1.758597e-06,
  0.000104455, 0.04425925, 0.3357167, 0.1399086, 0.05026428, 0.05481919, 
    0.07791981, 0.09881298, 0.131232, 0.03803048, 0.02769656, 0.1018698, 
    0.06448902, 0.1059661, 0.1200329, 0.1342003, 0.1281057, 0.07193899, 
    0.05802774, 0.006987691, 0.0007404101, 0.000804051, 0.003564408, 
    0.2912058, 0.2904252, 0.2432198, 0.06757122, 0.002552815, 6.532577e-05,
  0.0006077523, 0.09399599, 0.182924, 0.02208499, 0.04012297, 0.05092106, 
    0.08044177, 0.06615916, 0.1545098, 0.2602183, 0.04710779, 0.05376787, 
    0.09902394, 0.0770686, 0.08178236, 0.05237731, 0.01497253, 0.0163805, 
    0.002359369, 0.005764856, 0.001622549, 0.003487456, 0.009136165, 
    0.167262, 0.1516111, 0.09497565, 0.06957651, 0.006488529, 0.0005382759,
  0.002153575, 7.756254e-06, 0.01493356, 1.027141e-05, -9.260184e-06, 
    0.00346052, 0.005636208, 0.03611235, 0.01811565, 0.02107123, 0.03910477, 
    0.04363026, 0.04819522, 0.03919202, 0.007854235, 0.03803566, 0.05380509, 
    0.09883571, 0.03442665, 0.0488273, 0.07430393, 0.01163739, 6.305064e-05, 
    1.848274e-05, 3.519951e-05, 0.01035074, 0.004255397, 0.005170352, 
    0.01541913,
  0.1007069, 0.07423279, 0.009093115, 2.879718e-05, -0.0001119314, 
    0.01035646, 0.006331997, 0.01937892, 0.01695167, 0.01731808, 0.01629434, 
    0.0224134, 0.03443685, 0.01924452, 0.03774175, 0.007357982, 0.04804486, 
    0.07025048, 0.1873631, 0.07820632, 0.1137985, 0.05726873, 0.009001099, 
    0.0001109226, 0.00586822, 0.02272387, 0.03048909, 0.07794613, 0.09439315,
  0.03365489, 0.006517488, 0.0225121, 0.01878333, 0.007807754, 0.003304311, 
    0.0173874, 0.00128672, 0.007010611, 0.180996, 0.2028847, 0.1531552, 
    0.09302214, 0.1023159, 0.1128197, 0.095858, 0.1007366, 0.10689, 0.111452, 
    0.06305374, 0.05669998, 0.13907, 0.1516235, 0.1492273, 0.1435325, 
    0.1684807, 0.1045194, 0.07603233, 0.0589916,
  0.03030415, 0.01790585, 0.004349127, 0.0008666228, 0.02423611, 0.0176587, 
    0.0002181257, 0.0001642081, 0.001279014, 0.007093366, 0.02461443, 
    0.05240978, 0.0881991, 0.09772281, 0.09697694, 0.1132281, 0.1078202, 
    0.1568363, 0.1127502, 0.0118847, 4.539792e-05, 0.02686748, 0.09830579, 
    0.112632, 0.1328755, 0.2048402, 0.142704, 0.07075023, 0.04326413,
  0.01597051, 0.0004208246, 0.005641974, 0.002333665, 0.002065735, 
    0.006739948, 0.001713386, 0, 0, 0, 0, -4.047616e-06, 0.00144106, 
    0.003621704, 0.01598026, 0.01889972, 0.0164526, 0.04030268, 0.03434411, 
    0.001578956, 0.0001811616, 0.003210234, 0.01490157, 0.01061874, 
    0.01841867, 0.08130261, 0.1134336, 0.04898294, 0.02705509,
  0.002101813, 0.0009296412, 0.0002537988, 0.001579611, 0.0006857716, 
    0.0001364205, 0, 0, 0, 0, 0, 0, 0, -9.637723e-06, -3.274445e-05, 
    0.003550143, -0.0001272159, 0.0009018076, -5.248401e-05, -2.32376e-05, 0, 
    -6.564104e-06, 0, 0, -1.247694e-05, 0.002385339, 0.01679787, 0.01231685, 
    0.006035571,
  0, 1.235544e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0001203431, 
    0.0002927113, -3.314417e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, -6.094949e-06, 
    -4.748916e-05,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.003835133, 0.006532792, 
    0.006984174, 0.007351668, 0.002501407, -0.0002311906, -3.807887e-05, 
    0.0009480326, 0.002386008, -6.408947e-05, 0, 0, 0, 0,
  0, 0, 0, 0.0001256515, -5.550134e-05, 0.001201363, 0.01447, 0, 0, 
    -2.979566e-05, -7.681157e-06, 0.0003209851, -7.63733e-05, 0.003124851, 
    0.009483585, 0.01736597, 0.02533283, 0.02504747, 0.08849312, 0.0692862, 
    0.04609215, 0.02439095, 0.009204448, 0.008671141, 0.01392613, 
    0.004828667, 0.002701223, 0.007700219, 0.003103891,
  0.06063328, 0.03331441, 0.0227114, 0.03693978, 0.06607029, 0.06375364, 
    0.06301834, 0.06932011, 0.05473739, 0.06062824, 0.04563458, 0.06529494, 
    0.1133595, 0.1312444, 0.127187, 0.1059928, 0.07583697, 0.1026973, 
    0.09004642, 0.0790179, 0.06456017, 0.05298501, 0.07420373, 0.07135845, 
    0.09560098, 0.1016385, 0.05959181, 0.04936891, 0.03104112,
  0.1586207, 0.1459594, 0.1537854, 0.1798988, 0.2081766, 0.1824516, 
    0.1521802, 0.1614489, 0.1458369, 0.1430994, 0.1569949, 0.1584863, 
    0.1492532, 0.1179279, 0.1131385, 0.07436483, 0.1131674, 0.1214026, 
    0.1300748, 0.1137543, 0.1468716, 0.1165734, 0.1725006, 0.1067818, 
    0.1198206, 0.2237436, 0.1659474, 0.1009169, 0.1493708,
  0.09294644, 0.06590959, 0.05412253, 0.06917487, 0.07749812, 0.09486489, 
    0.09011259, 0.07575537, 0.07037985, 0.08346515, 0.1081442, 0.08037484, 
    0.08872768, 0.1329277, 0.1184183, 0.07583042, 0.09637372, 0.1574057, 
    0.1204049, 0.1414512, 0.1516851, 0.1467432, 0.05692534, 0.04122526, 
    0.06670108, 0.106523, 0.1198054, 0.1370393, 0.09092905,
  0.00456196, 0.006313142, 0.07362057, 0.04882612, 0.06954795, 0.1266024, 
    0.1887505, 0.08719586, 0.0532028, 0.06527901, 0.1598054, 0.07624015, 
    0.03886441, 0.09073219, 0.04761627, 0.1101724, 0.09772973, 0.1741357, 
    0.1389208, 0.08698874, 0.09066607, 0.05217689, 0.004794604, 0.008419574, 
    0.04526626, 0.07456065, 0.202018, 0.05559291, 0.01693269,
  2.812347e-07, 0.05391398, 0.04104172, 0.03891869, 0.1714398, 0.04576868, 
    0.05752368, 0.02123114, 0.06690697, 0.008682113, 0.08636557, 0.01945937, 
    0.01972033, 0.06046923, 0.1132181, 0.1027387, 0.09497835, 0.07578267, 
    0.06410886, 0.02182428, 0.03184323, 0.01849652, 0.00429938, 0.01594123, 
    0.08680721, 0.1694925, 0.08467199, 0.008145586, 1.114269e-06,
  -9.859323e-06, 0.05225228, 0.2965827, 0.1159127, 0.04071624, 0.04065427, 
    0.06676197, 0.08354513, 0.1053964, 0.0285954, 0.02714585, 0.09083299, 
    0.05133454, 0.08604199, 0.1094804, 0.1321391, 0.10346, 0.06074068, 
    0.04544213, 0.0009766343, 0.005146931, -3.991263e-05, 0.008362299, 
    0.2464349, 0.2566323, 0.2018318, 0.054793, 0.0009498307, 6.69768e-05,
  0.0005987423, 0.07193211, 0.1373812, 0.01574681, 0.03426627, 0.04140405, 
    0.05563617, 0.05189944, 0.1191134, 0.2108977, 0.04326605, 0.04310483, 
    0.07968316, 0.05696614, 0.06525336, 0.04721317, 0.01382167, 0.008538488, 
    0.001930095, 0.003725235, 0.008630462, 0.003716017, 0.01083408, 
    0.1149693, 0.1187812, 0.07833986, 0.04555629, 0.005494955, 0.0003278013,
  2.786675e-05, 3.938213e-06, 0.01288088, 1.687187e-05, 4.289242e-05, 
    0.002907435, 0.003125736, 0.03293474, 0.01595002, 0.01791356, 0.03480261, 
    0.03784871, 0.04125306, 0.04000636, 0.003433095, 0.03506786, 0.05827422, 
    0.09373881, 0.03359825, 0.03865725, 0.05123142, 0.009599621, 
    0.0001353702, 8.356494e-06, 0.0001935952, 0.01455658, 0.009037657, 
    0.01681967, 0.01530368,
  0.06860286, 0.05494665, 0.003768619, 0.0005989416, 0.00121291, 0.008222115, 
    0.001935473, 0.01287638, 0.01568376, 0.02335477, 0.01201942, 0.02950485, 
    0.03541482, 0.02783824, 0.02623698, 0.004362239, 0.04299295, 0.04885607, 
    0.1518045, 0.05699871, 0.09128504, 0.04684428, 0.009580464, 0.0001213803, 
    0.00209955, 0.01652956, 0.0143754, 0.06092306, 0.09700049,
  0.05284783, 0.01588169, 0.02013498, 0.02756662, 0.01120471, 0.007139973, 
    0.0233442, 0.00381961, 0.01692547, 0.2047395, 0.202823, 0.1428679, 
    0.08832541, 0.1011726, 0.09364602, 0.08795851, 0.08575086, 0.09905692, 
    0.07672381, 0.04135306, 0.07911897, 0.1113308, 0.1360505, 0.1338868, 
    0.1211596, 0.1291026, 0.09267017, 0.07029402, 0.07783042,
  0.08569141, 0.0760634, 0.03769693, 0.004764885, 0.04984374, 0.05743495, 
    0.002625672, 0.02726854, 0.03552972, 0.01920673, 0.03633247, 0.08503735, 
    0.1342664, 0.1300435, 0.1484347, 0.1574075, 0.1630944, 0.2462614, 
    0.1793418, 0.09247759, 0.001416604, 0.1006809, 0.1751651, 0.153763, 
    0.1679375, 0.2605381, 0.1597671, 0.08542471, 0.1062122,
  0.1254057, 0.04624977, 0.01889708, 0.02543223, 0.01914549, 0.03005321, 
    0.005839103, 0, 0, 0.004808661, 0.0009362608, 0.001972713, 0.009668795, 
    0.02043819, 0.05888133, 0.06093072, 0.09818434, 0.09488036, 0.09392653, 
    0.01792995, 0.009675256, 0.01000626, 0.04474314, 0.03686076, 0.0467453, 
    0.1880649, 0.2387945, 0.1475771, 0.1289087,
  0.0654669, 0.004433743, 0.005444928, 0.00825166, 0.001270268, 0.001789502, 
    -4.249929e-05, 5.562397e-06, 0, 0, 0, 0, 0, 0.005861218, 0.007353849, 
    0.01983894, 0.01433758, 0.02600408, 0.0008115546, 0.005807814, 
    -3.734813e-05, 0.0006467568, 0, -1.376087e-05, 0.002397139, 0.01678885, 
    0.06688678, 0.09076089, 0.07439122,
  -2.176514e-05, 2.412364e-05, 0.000450668, 0.0001598484, 0.001388426, 
    2.386527e-05, 0, 0, 0, 8.210149e-05, 0, 0, 0.0001949206, 0.001293694, 
    2.402653e-06, 0.005752666, 0.01754049, 0.0153145, 0.01060595, 
    0.006901385, 0, 0, 0, 0, 0, 0, -1.123622e-06, 0.006916331, 0.003054579,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8.281385e-12, 0.004599987, 
    0.01863426, 0.01769297, 0.01957336, 0.0142956, 0.00913173, 0.0001247791, 
    -7.316371e-06, 0.002326517, 0.0244355, 0.0175271, -0.001457556, 
    7.293373e-05, 5.256605e-05, 0,
  0.005306933, -4.529162e-05, -0.0001678838, 0.001595042, -0.000465597, 
    0.002247809, 0.03079911, -0.0002818168, -0.0001087776, -0.0003000312, 
    -1.230686e-05, 0.0002729751, -0.0001936614, 0.07904974, 0.0631143, 
    0.04892059, 0.05316673, 0.08749551, 0.1051972, 0.08385466, 0.07592107, 
    0.08272105, 0.06127574, 0.03572965, 0.06506988, 0.0315667, 0.02546357, 
    0.01463273, 0.01118454,
  0.09694621, 0.06606396, 0.05853146, 0.07568426, 0.1025, 0.09918731, 
    0.1159354, 0.1313331, 0.138561, 0.1123396, 0.08508869, 0.1630344, 
    0.1999729, 0.2134242, 0.1795689, 0.1571016, 0.1706418, 0.1568888, 
    0.1467733, 0.1375054, 0.1198972, 0.1208462, 0.1503806, 0.1393034, 
    0.1702647, 0.1882495, 0.1362742, 0.1114132, 0.08341001,
  0.1567743, 0.1602848, 0.1787412, 0.1915521, 0.2068338, 0.1641415, 
    0.1477379, 0.1709996, 0.1615397, 0.1595916, 0.1870266, 0.1731075, 
    0.1652826, 0.1171765, 0.1204171, 0.07994041, 0.110546, 0.1366927, 
    0.1407734, 0.1346243, 0.1453472, 0.1208365, 0.1747788, 0.139667, 
    0.1153688, 0.2228532, 0.1657976, 0.1056427, 0.1415608,
  0.0907739, 0.06138659, 0.04493592, 0.06558933, 0.07241488, 0.07609097, 
    0.07752081, 0.077301, 0.05615004, 0.06748094, 0.08257552, 0.06691831, 
    0.08549202, 0.1308748, 0.1030827, 0.06889346, 0.09962996, 0.1456816, 
    0.1133661, 0.1268398, 0.1194359, 0.1269367, 0.05116897, 0.04943732, 
    0.06229793, 0.09348768, 0.1070367, 0.1290326, 0.08648188,
  0.004764622, 0.004419871, 0.05252012, 0.03692974, 0.05767874, 0.1149334, 
    0.1820471, 0.06987348, 0.04525442, 0.05624058, 0.1656282, 0.0733518, 
    0.03652048, 0.08686912, 0.03941, 0.1025246, 0.08347939, 0.1726545, 
    0.1411772, 0.07218067, 0.0784201, 0.02883565, 0.002378352, 0.001605318, 
    0.04381798, 0.07093598, 0.1895277, 0.04991051, 0.01559802,
  7.740107e-06, 0.0487853, 0.04308842, 0.02514141, 0.1651497, 0.04052523, 
    0.05816622, 0.01480892, 0.04751018, 0.006789747, 0.06907772, 0.02003253, 
    0.01862547, 0.05228421, 0.09660407, 0.1046142, 0.08523831, 0.06447305, 
    0.05299918, 0.01589759, 0.01786892, 0.01334258, 0.008560534, 0.01147163, 
    0.08434868, 0.1637661, 0.07681303, 0.002016261, 1.041436e-06,
  0.0008310903, 0.05042015, 0.264553, 0.1068817, 0.03703668, 0.02693621, 
    0.05021266, 0.06572978, 0.07881454, 0.02334846, 0.02980141, 0.06869967, 
    0.03905184, 0.06229965, 0.099503, 0.1277286, 0.0738848, 0.05070316, 
    0.02754558, 0.0004182313, 0.004571758, -0.000323542, 0.0008315392, 
    0.2012287, 0.2149112, 0.1605098, 0.04819554, 0.0006843862, 0.000114871,
  0.0008070513, 0.05143228, 0.1078306, 0.01160853, 0.03045996, 0.03260589, 
    0.03138354, 0.03831358, 0.09894164, 0.1791256, 0.04039086, 0.02983529, 
    0.06406668, 0.0386256, 0.03968283, 0.03464967, 0.01216885, 0.003226481, 
    0.001191575, 0.003386425, 0.001352694, 0.003883669, 0.02232116, 
    0.08367827, 0.08739568, 0.06018228, 0.02753496, 0.004949994, 0.0004315707,
  8.588826e-05, 1.603029e-06, 0.008396365, 0.0006650385, 0.000486159, 
    0.003397889, 0.002221045, 0.03464534, 0.01848477, 0.01717236, 0.03114686, 
    0.03087138, 0.03398485, 0.05296444, 0.002863253, 0.01715972, 0.06456985, 
    0.08346179, 0.04250649, 0.03148148, 0.03534076, 0.007587947, 
    0.0001370235, 9.704856e-06, 0.0004068611, 0.01002156, 0.007385915, 
    0.02587508, 0.01966432,
  0.04470796, 0.02785916, 0.001872074, 0.001852603, 0.003252965, 0.002677817, 
    0.001791399, 0.009829054, 0.01049916, 0.01839373, 0.01354786, 0.0236812, 
    0.03892819, 0.03770052, 0.01629697, 0.001312761, 0.03042237, 0.02627552, 
    0.1284425, 0.0444527, 0.07739106, 0.04585985, 0.01351372, 4.513727e-05, 
    0.00132009, 0.01625725, 0.01067808, 0.03781711, 0.06287302,
  0.03597382, 0.01700017, 0.01617706, 0.02157334, 0.01219191, 0.006910538, 
    0.03883607, 0.01029957, 0.03680499, 0.1893648, 0.1881445, 0.118849, 
    0.08624271, 0.08504434, 0.07742222, 0.07534632, 0.0752752, 0.08755443, 
    0.04334523, 0.03160238, 0.06128164, 0.07765325, 0.112046, 0.1081171, 
    0.08911013, 0.09797308, 0.05757471, 0.06931219, 0.05286951,
  0.07563792, 0.07963967, 0.0616753, 0.0212095, 0.1078122, 0.1167399, 
    0.01091662, 0.1455494, 0.06833906, 0.02579918, 0.07134455, 0.1412373, 
    0.1662261, 0.1508226, 0.169587, 0.161929, 0.1991959, 0.2506482, 
    0.1830666, 0.1422524, 0.02698009, 0.1548419, 0.1976835, 0.1781769, 
    0.1873532, 0.2517869, 0.1280549, 0.08005169, 0.1043416,
  0.1273873, 0.1158851, 0.1066391, 0.1001986, 0.1031599, 0.09801378, 
    0.04843841, -3.877053e-05, 0.001948489, 0.02700255, 0.01057522, 
    0.008571913, 0.02834536, 0.05963637, 0.08456045, 0.0955584, 0.1314668, 
    0.1505584, 0.1975121, 0.04389118, 0.04419826, 0.1114357, 0.1338776, 
    0.05366187, 0.09097307, 0.2210919, 0.2728212, 0.1498844, 0.1434078,
  0.1715624, 0.05766102, 0.05600208, 0.09131401, 0.0462241, 0.03906365, 
    0.02577973, 0.01712254, 0.007106631, 6.351505e-05, -1.558292e-06, 0, 
    -0.0003015106, 0.01481098, 0.03331813, 0.05327702, 0.0672675, 0.06078987, 
    0.03298357, 0.04299077, 0.01283357, 0.01969558, 0.01135832, 0.01032059, 
    0.01732784, 0.03755216, 0.1265122, 0.1733347, 0.1689256,
  0.01761081, 0.01122618, 0.003796724, 0.01386042, 0.02045363, 0.02117102, 
    0.003204429, 0.004452149, 0.002167525, 0.004982747, 0.0009389683, 
    0.003072675, 0.004782781, 0.004623839, 0.02121174, 0.02470399, 
    0.02535158, 0.02256036, 0.01520436, 0.01729922, 0.01198471, 
    -0.0001067019, 0, 0, 0.0001365351, -1.310018e-05, -4.279316e-05, 
    0.02598612, 0.02143502,
  -9.327843e-08, -6.835111e-09, 0, -2.746768e-05, 0.002708329, 0.002742766, 
    0.0004204802, -3.474138e-05, -1.292638e-05, -1.887903e-06, 1.223742e-05, 
    0.0004399603, 0.001183148, 0.001445905, 0.001094589, 0.001477518, 
    0.0005133433, -8.573651e-06, -2.104882e-07, 0, 0, 0, 0, 0, 0, 0, 0, 
    -3.302095e-08, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3.65266e-05, 0.02265222, 0.02567066, 
    0.03487975, 0.05267412, 0.02260578, 0.0243839, 0.01088518, 0.002092564, 
    0.0164221, 0.05663451, 0.05521623, 0.01739625, 0.002286829, 0.0002084909, 
    7.501278e-05,
  0.03307595, 0.0181622, 0.06312618, 0.04403005, 0.003941832, 0.01528526, 
    0.05400665, -0.001122003, -0.0008921485, -0.0004591149, -0.0002107348, 
    0.001229135, 0.03720366, 0.1609496, 0.142371, 0.1290153, 0.1353717, 
    0.1744407, 0.1522395, 0.1289864, 0.1160447, 0.1586998, 0.1092193, 
    0.1153143, 0.2075538, 0.1215153, 0.1010886, 0.1102498, 0.06887021,
  0.1514616, 0.1081726, 0.1113007, 0.1250938, 0.1559325, 0.1652458, 
    0.1725375, 0.1841218, 0.1788249, 0.1506345, 0.1419386, 0.2415863, 
    0.2553706, 0.2321196, 0.1984801, 0.1930581, 0.2014949, 0.1960167, 
    0.2036197, 0.1790558, 0.1959083, 0.1746604, 0.1929528, 0.1833448, 
    0.2007807, 0.2222675, 0.1791505, 0.1592413, 0.1426366,
  0.1488025, 0.1738044, 0.1803242, 0.1940273, 0.2097687, 0.1578671, 
    0.1457056, 0.1775438, 0.1558277, 0.1549325, 0.1870468, 0.1646806, 
    0.1687998, 0.1099676, 0.1075285, 0.0790042, 0.1125568, 0.1300728, 
    0.1402502, 0.1383147, 0.1354691, 0.126119, 0.1838119, 0.1494265, 
    0.1172294, 0.2299864, 0.1614738, 0.104699, 0.143789,
  0.09330429, 0.0647641, 0.0448021, 0.06819782, 0.06716616, 0.07041086, 
    0.07321617, 0.06403713, 0.03851667, 0.0521031, 0.07577262, 0.06267723, 
    0.0811296, 0.1338961, 0.09029979, 0.05155075, 0.08273372, 0.1340755, 
    0.1015096, 0.1200444, 0.1068042, 0.1087185, 0.05986488, 0.03154552, 
    0.04836615, 0.08381969, 0.09348453, 0.1190223, 0.09197348,
  0.004314627, 0.002940746, 0.04221971, 0.03240796, 0.04669263, 0.1134798, 
    0.1443961, 0.05717521, 0.0419318, 0.04394948, 0.1326073, 0.07418751, 
    0.04328756, 0.08163431, 0.03386516, 0.09248022, 0.06240394, 0.1539811, 
    0.1303785, 0.06899728, 0.0623508, 0.01828567, 0.001409659, 0.001774401, 
    0.04678714, 0.05365119, 0.1663412, 0.04466944, 0.01312805,
  -7.691904e-07, 0.04631524, 0.03955714, 0.01551804, 0.1491446, 0.03684904, 
    0.05431495, 0.0162151, 0.03708184, 0.01637159, 0.04912463, 0.01571092, 
    0.02085231, 0.0455157, 0.08790068, 0.1191673, 0.0743055, 0.06068455, 
    0.04284328, 0.01128548, 0.00220372, 0.001082058, 0.003438952, 0.0102932, 
    0.07280561, 0.1440438, 0.07253055, 0.0005308526, 4.38606e-07,
  8.398249e-05, 0.06521657, 0.2161307, 0.07315502, 0.03612429, 0.02133701, 
    0.0391435, 0.0550091, 0.06408695, 0.01888338, 0.0374979, 0.06375805, 
    0.03578049, 0.04730991, 0.09846652, 0.1188019, 0.05858998, 0.0513577, 
    0.01672661, 0.0002339174, 0.001596672, -0.0002051834, -2.870197e-05, 
    0.1759534, 0.1963864, 0.1263839, 0.03848811, 0.0006626156, 0.0001292797,
  0.002122905, 0.04247703, 0.08643763, 0.01148353, 0.02157631, 0.02661845, 
    0.01777727, 0.02665874, 0.08769811, 0.1666862, 0.0393401, 0.02200606, 
    0.05827083, 0.02995326, 0.02414679, 0.03126409, 0.01565645, 0.005596146, 
    0.0009053397, 0.001282852, 0.003568436, 0.002523533, 0.02051852, 
    0.06078108, 0.08071952, 0.06126592, 0.01587143, 0.004118419, 0.0005466113,
  0.0003586979, 6.837604e-07, 0.004015154, 0.001078895, 2.218018e-05, 
    0.0009370979, 0.001619029, 0.03123766, 0.01709914, 0.02437796, 0.0311261, 
    0.02847299, 0.02760751, 0.05995919, 0.002474203, 0.01122303, 0.05622952, 
    0.07754621, 0.05126664, 0.02738879, 0.02673731, 0.005782211, 
    0.0001105243, 1.102605e-05, 0.0004827026, 0.01262204, 0.007529697, 
    0.03519451, 0.01642562,
  0.02685722, 0.00922472, 0.001577003, 0.004549722, 0.004697613, 
    0.0001192389, 0.003727708, 0.007899575, 0.008351039, 0.01184854, 
    0.0149015, 0.02140671, 0.03444165, 0.03866168, 0.006439492, 0.0004499195, 
    0.02227981, 0.01943123, 0.09593007, 0.03627216, 0.0552516, 0.04173676, 
    0.01090933, 6.610609e-05, 0.000900033, 0.009615079, 0.008756237, 
    0.01950277, 0.05131162,
  0.02665278, 0.02149033, 0.01613623, 0.01353389, 0.0149807, 0.00930644, 
    0.04542106, 0.0195357, 0.09020149, 0.1748599, 0.1762436, 0.108886, 
    0.08535822, 0.08184107, 0.05697806, 0.06774549, 0.06585337, 0.05679625, 
    0.03070104, 0.02723163, 0.04197059, 0.05603011, 0.09248789, 0.08403256, 
    0.06958196, 0.06909999, 0.04018109, 0.07430315, 0.03130721,
  0.05226075, 0.07302809, 0.08411489, 0.05114272, 0.129728, 0.1346711, 
    0.03928714, 0.1878615, 0.1163528, 0.05574276, 0.1122719, 0.1438686, 
    0.1905755, 0.1557881, 0.1703731, 0.1701002, 0.1972865, 0.2350808, 
    0.1692859, 0.1465677, 0.08483729, 0.1768658, 0.1866577, 0.1757546, 
    0.1914659, 0.2359409, 0.105022, 0.06402303, 0.08717885,
  0.126637, 0.1217202, 0.162327, 0.1788574, 0.2048752, 0.1760667, 0.1317612, 
    0.003236298, 0.02972308, 0.04768981, 0.03009375, 0.03161972, 0.05639561, 
    0.09037149, 0.1351804, 0.1219938, 0.1811667, 0.1873357, 0.2127249, 
    0.1110396, 0.105117, 0.1505745, 0.1609729, 0.1014838, 0.124282, 
    0.2163726, 0.2556159, 0.1420286, 0.1350708,
  0.2153437, 0.1438056, 0.1250187, 0.174872, 0.1469592, 0.1349171, 0.1083526, 
    0.06771007, 0.01898691, 0.02355486, 0.01640986, -0.0003006453, 
    0.01296538, 0.06687213, 0.1484191, 0.08878349, 0.1040896, 0.1171435, 
    0.08264394, 0.128169, 0.05426655, 0.0696369, 0.04864497, 0.02577366, 
    0.03949982, 0.06061272, 0.1347478, 0.2178136, 0.2050021,
  0.08432428, 0.09219106, 0.06853978, 0.1045207, 0.1160838, 0.07436737, 
    0.03855187, 0.03148322, 0.02166685, 0.04189124, 0.02263867, 0.01991655, 
    0.007734728, 0.03912953, 0.08408929, 0.04336936, 0.04361563, 0.03208821, 
    0.05423098, 0.03166069, 0.02879829, 0.005129558, 5.281693e-07, 0, 
    0.02316317, 0.0001666303, -0.0001811929, 0.06199661, 0.06828551,
  0.02376886, 0.01979123, 0.0172728, 0.02688351, 0.03396032, 0.02165976, 
    0.01605738, 0.006572514, 0.002255548, 0.006138482, 0.00693457, 
    0.01093131, 0.009218844, 0.00662052, 0.01047077, 0.02020673, 0.03097262, 
    0.01892103, 0.007739849, -0.0001110811, -4.606608e-06, 0, 0, 
    -2.930009e-05, -0.0003150104, 2.176605e-05, -2.061249e-06, -0.004209334, 
    0.02330839,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001324894, 0.03411682, 0.05514182, 
    0.1176023, 0.1156135, 0.06725078, 0.04225002, 0.02912039, 0.01052666, 
    0.03499695, 0.09098172, 0.1008691, 0.0427218, 0.05464515, 0.002161348, 
    0.0004497876,
  0.0920108, 0.08943459, 0.1604631, 0.1207704, 0.01808329, 0.02946637, 
    0.09225965, 0.0007850728, 0.004980631, 0.0005085862, 0.003898251, 
    0.01029388, 0.09942284, 0.2229349, 0.1814821, 0.1913311, 0.20702, 
    0.2918957, 0.2281549, 0.1862072, 0.2103411, 0.2198118, 0.2205933, 
    0.2017749, 0.3401956, 0.2289088, 0.1859536, 0.192895, 0.1435482,
  0.2100316, 0.1651852, 0.1674445, 0.1934538, 0.2002175, 0.2292908, 
    0.2134815, 0.2365642, 0.2490188, 0.2561382, 0.1976752, 0.2786354, 
    0.2635398, 0.2435407, 0.2092125, 0.2105673, 0.1998817, 0.198871, 
    0.2572139, 0.2263719, 0.2469077, 0.2358063, 0.2437449, 0.2326658, 
    0.271783, 0.2552365, 0.2112208, 0.1752515, 0.1630151,
  0.1405289, 0.1740851, 0.1778697, 0.2004, 0.2074216, 0.1619226, 0.1418676, 
    0.1803275, 0.1557279, 0.1650154, 0.1864832, 0.1762283, 0.1843917, 
    0.110465, 0.1026071, 0.08059065, 0.1207817, 0.1268312, 0.1408666, 
    0.1534902, 0.1373684, 0.1257817, 0.1869578, 0.151405, 0.1133346, 
    0.1948009, 0.1512058, 0.1119727, 0.1353702,
  0.08046088, 0.06206427, 0.03650931, 0.06802574, 0.06346358, 0.0568677, 
    0.06705607, 0.0459557, 0.02906229, 0.0377708, 0.06545982, 0.05140949, 
    0.0841248, 0.1310019, 0.08053116, 0.0399158, 0.06983389, 0.1243367, 
    0.09619693, 0.1026425, 0.09525771, 0.1022451, 0.05653471, 0.02820462, 
    0.04401687, 0.07123101, 0.08987366, 0.1128215, 0.07771074,
  0.005376501, 0.0005785117, 0.03579383, 0.02870458, 0.04589234, 0.1093372, 
    0.1145413, 0.05497633, 0.04266557, 0.03294711, 0.1267081, 0.07626107, 
    0.0482138, 0.08709008, 0.03256777, 0.06616499, 0.0588713, 0.145411, 
    0.1119261, 0.06711631, 0.04906382, 0.02272114, 0.003532483, 0.00024888, 
    0.04486821, 0.04413871, 0.152627, 0.03949882, 0.014359,
  3.079311e-06, 0.04095091, 0.04125414, 0.01358754, 0.1408181, 0.03308249, 
    0.0549875, 0.01804596, 0.02660077, 0.01017378, 0.04356647, 0.01376515, 
    0.02527202, 0.04480038, 0.08057851, 0.1202911, 0.07513992, 0.05171067, 
    0.03781509, 0.01208015, 0.0006305173, 6.573855e-06, 0.001141755, 
    0.008896841, 0.06120135, 0.1303495, 0.07174163, 0.004759619, 1.015339e-07,
  0.001945247, 0.06399145, 0.183482, 0.05771703, 0.03181629, 0.02067969, 
    0.03630899, 0.04699787, 0.05872216, 0.01927394, 0.04710745, 0.06669975, 
    0.03013391, 0.03909757, 0.1029729, 0.1071464, 0.04283974, 0.05560784, 
    0.01409058, 0.0002535963, -6.507559e-05, -0.0001702795, 0.0002936005, 
    0.1619817, 0.1909982, 0.1066974, 0.02910932, 0.0006440503, 0.0001366293,
  0.006768571, 0.0371189, 0.07954387, 0.01177266, 0.0171747, 0.02294838, 
    0.01360588, 0.01670231, 0.06970153, 0.1827939, 0.04596793, 0.01516238, 
    0.05004755, 0.02648509, 0.02184153, 0.03071102, 0.005855141, 0.002542184, 
    0.00141022, 0.001332286, 0.01017054, 0.001089485, 0.03122045, 0.05164968, 
    0.09286164, 0.07017224, 0.01228763, 0.005785896, 0.002720973,
  0.0001146149, 7.279865e-07, 0.0009940744, 0.00237902, 7.669682e-05, 
    0.001010381, 0.001662997, 0.02808965, 0.01840311, 0.02466558, 0.03024616, 
    0.03370714, 0.02659365, 0.04748144, 0.005442508, 0.01280607, 0.04054099, 
    0.07495262, 0.05660729, 0.03502643, 0.02478327, 0.005059749, 
    0.0001460431, 1.019888e-05, 0.001120121, 0.02595347, 0.009945235, 
    0.01382449, 0.01387871,
  0.01484269, 0.000992417, 3.229338e-05, 0.008723193, 0.004798432, 
    4.590005e-05, 0.001718689, 0.007145182, 0.006282514, 0.003816079, 
    0.009168541, 0.03249735, 0.02914052, 0.02242217, 0.004082892, 
    9.692849e-05, 0.0177949, 0.007281028, 0.0862866, 0.02803156, 0.0381307, 
    0.03763522, 0.005691137, 1.702882e-05, 0.0006260647, 0.004600283, 
    0.007282855, 0.01957228, 0.03728703,
  0.02022306, 0.02045152, 0.01264977, 0.004679183, 0.02768186, 0.01384175, 
    0.04087394, 0.03432547, 0.1551887, 0.1712639, 0.1661987, 0.09430598, 
    0.0948887, 0.07638247, 0.04945947, 0.05499826, 0.05967657, 0.04947716, 
    0.03234724, 0.02360791, 0.02940196, 0.04864992, 0.08349295, 0.06167807, 
    0.06171806, 0.05078811, 0.03521231, 0.08909029, 0.01600176,
  0.033479, 0.07511922, 0.09824529, 0.09240313, 0.1195806, 0.1177346, 
    0.08751717, 0.1659772, 0.112749, 0.08785091, 0.1300133, 0.1252959, 
    0.1878705, 0.1507749, 0.1752802, 0.1726707, 0.1898017, 0.2272999, 
    0.1584586, 0.1583844, 0.1380091, 0.1727826, 0.1767253, 0.1773208, 
    0.20175, 0.2215285, 0.08807079, 0.06074682, 0.06186254,
  0.1401281, 0.1544845, 0.1772514, 0.1770927, 0.2046293, 0.196996, 0.1956336, 
    0.07158977, 0.04359983, 0.09725228, 0.04840442, 0.0714239, 0.1089527, 
    0.1806537, 0.200221, 0.1654751, 0.2133964, 0.200018, 0.2449711, 
    0.1658748, 0.178329, 0.176493, 0.1676676, 0.137216, 0.1475014, 0.2067973, 
    0.2509866, 0.1526094, 0.1413202,
  0.251482, 0.1905788, 0.160431, 0.2328306, 0.2421173, 0.1976047, 0.201129, 
    0.1333066, 0.07786909, 0.05339949, 0.03666304, 0.01466564, 0.02154625, 
    0.1275693, 0.2011075, 0.1396016, 0.1257511, 0.1703068, 0.1523474, 
    0.1849918, 0.1236592, 0.09687164, 0.1010541, 0.04668931, 0.08694768, 
    0.103215, 0.1724376, 0.230957, 0.2400086,
  0.1042995, 0.1517255, 0.1268349, 0.1849976, 0.1716055, 0.1155896, 
    0.09277639, 0.08344086, 0.06678831, 0.0906533, 0.07986742, 0.03601949, 
    0.05089133, 0.1256531, 0.1360617, 0.08744919, 0.06484096, 0.04965948, 
    0.06842506, 0.09801544, 0.06873348, 0.02172313, 0.0004448381, 
    -1.323696e-05, 0.04401817, 0.002828686, 0.001026148, 0.08541696, 0.1007483,
  0.05875399, 0.05807485, 0.0486866, 0.07313898, 0.06429915, 0.04290752, 
    0.03773463, 0.02954752, 0.01952375, 0.01684699, 0.01910119, 0.02346442, 
    0.02222082, 0.05021419, 0.06837055, 0.07841007, 0.09492172, 0.1014061, 
    0.05920765, 0.03230246, 0.005129871, 0.004807514, -3.259007e-05, 
    -0.001407421, 0.007295899, -6.422026e-05, -0.0023532, 0.02110872, 
    0.05813608,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  -0.0006345421, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0346277, 0.09112171, 
    0.1207832, 0.187608, 0.2538227, 0.1444481, 0.07395354, 0.05017072, 
    0.02426507, 0.0653253, 0.182757, 0.1952753, 0.1628995, 0.2116459, 
    0.04083172, 0.004433447,
  0.1408665, 0.194291, 0.3351669, 0.2417124, 0.03991079, 0.04616207, 
    0.1304197, 0.03062401, 0.02548557, 0.02079133, 0.01948871, 0.03638475, 
    0.1385833, 0.2729459, 0.2331248, 0.2127421, 0.2287825, 0.3096263, 
    0.2406885, 0.1973381, 0.2457877, 0.2609461, 0.2988105, 0.31972, 0.401153, 
    0.2925002, 0.2271596, 0.2334928, 0.219493,
  0.2168748, 0.2058436, 0.247874, 0.266048, 0.2510237, 0.2516078, 0.2281342, 
    0.2536471, 0.2715069, 0.2891626, 0.2438946, 0.305386, 0.2694128, 
    0.2507439, 0.2240369, 0.2182095, 0.1988173, 0.1958717, 0.3058424, 
    0.2593755, 0.2702338, 0.2400005, 0.2686809, 0.2434213, 0.2695563, 
    0.2641394, 0.2228292, 0.1870764, 0.1707946,
  0.145057, 0.194158, 0.1846267, 0.2030835, 0.2101456, 0.1506908, 0.1342012, 
    0.173332, 0.1558711, 0.1744877, 0.2067177, 0.1707122, 0.1749008, 
    0.1144595, 0.09795354, 0.07495318, 0.1303715, 0.1363899, 0.138494, 
    0.1535769, 0.129862, 0.1349618, 0.1961364, 0.1449488, 0.1057956, 
    0.1921692, 0.1647296, 0.1132072, 0.1331906,
  0.0782564, 0.06300809, 0.03427296, 0.0666472, 0.06754707, 0.0573415, 
    0.06142418, 0.03875372, 0.0255149, 0.05169594, 0.06319547, 0.05031879, 
    0.08100867, 0.1325411, 0.06437735, 0.03430608, 0.0721979, 0.1212765, 
    0.09917961, 0.08906549, 0.09527291, 0.1183573, 0.0481102, 0.01877502, 
    0.04104542, 0.0716088, 0.08259296, 0.1008276, 0.07877915,
  0.006963133, 6.542321e-05, 0.03423651, 0.02489959, 0.04478535, 0.1041969, 
    0.09013797, 0.04678636, 0.03516414, 0.0328436, 0.1174588, 0.07965693, 
    0.05263932, 0.09174821, 0.03047512, 0.05525839, 0.06450409, 0.1337205, 
    0.1086015, 0.06756332, 0.04264595, 0.02117327, 0.005357599, 0.0001175298, 
    0.04241285, 0.03682768, 0.1386391, 0.03654274, 0.01094827,
  -5.697408e-06, 0.0481242, 0.04354174, 0.01367986, 0.1384797, 0.02967577, 
    0.05766796, 0.03045003, 0.01883188, 0.004201673, 0.03510327, 0.01412207, 
    0.03070019, 0.05015821, 0.0744302, 0.12514, 0.07777157, 0.04777935, 
    0.03622181, 0.01189644, 0.0006282537, -1.250398e-07, 4.339324e-05, 
    0.006553949, 0.05357321, 0.1194868, 0.07363395, 0.005383632, 2.610921e-06,
  0.0005402928, 0.07375651, 0.182686, 0.05691887, 0.02916987, 0.02665849, 
    0.03254754, 0.04649631, 0.05870635, 0.02715242, 0.0521604, 0.06286617, 
    0.03122055, 0.03533005, 0.09596215, 0.09534639, 0.03831208, 0.05815221, 
    0.01207544, 0.0001341621, -3.995099e-05, -0.0003978635, 0.002298722, 
    0.1453727, 0.1906029, 0.1021095, 0.01751613, 0.0008681669, 8.961761e-05,
  0.01888429, 0.03685402, 0.06328069, 0.0148216, 0.01753827, 0.01773598, 
    0.01594217, 0.01148506, 0.0663709, 0.1867076, 0.03538547, 0.01580225, 
    0.04691037, 0.02309155, 0.02255639, 0.0288626, 0.008650572, 0.0006642098, 
    0.001944659, 0.01056276, 0.01154987, 0.0007885747, 0.05875136, 
    0.05200125, 0.09720967, 0.07498887, 0.01165468, 0.008841813, 0.0065002,
  0.0002073299, 1.070977e-06, 0.0020373, 0.0009699486, 0.0003134964, 
    0.00163778, 0.002355645, 0.0281346, 0.01587242, 0.01995039, 0.0290075, 
    0.03475255, 0.03156157, 0.05372647, 0.00675856, 0.009919864, 0.03167732, 
    0.07422692, 0.06475399, 0.04900962, 0.01808394, 0.005724428, 
    0.0002213104, 3.008619e-05, 0.002058703, 0.009275896, 0.0008660406, 
    0.002273367, 0.009508557,
  0.01061814, 0.001046026, 2.044132e-06, 0.006958597, 0.009951368, 
    0.001116642, 0.0003437118, 0.007363949, 0.005750007, 0.006512242, 
    0.01614294, 0.03224984, 0.02396304, 0.01806422, 0.001782401, 
    0.0001039374, 0.01813137, 0.001671736, 0.07616074, 0.01799429, 
    0.02719978, 0.03313008, 0.004184705, 2.617936e-05, 0.000693229, 
    0.006454618, 0.000769151, 0.01391068, 0.02061689,
  0.01816434, 0.01601062, 0.009116951, 0.001250079, 0.04345949, 0.01888224, 
    0.04692021, 0.05850571, 0.2069751, 0.1729717, 0.1505309, 0.08601296, 
    0.09914466, 0.0789479, 0.04094165, 0.04025877, 0.05032191, 0.04326365, 
    0.02083971, 0.02142255, 0.02111828, 0.05250977, 0.08123722, 0.05223772, 
    0.04906858, 0.04278976, 0.03349614, 0.08271751, 0.007919637,
  0.02616253, 0.06891914, 0.1012886, 0.1067611, 0.1120157, 0.09998478, 
    0.1557442, 0.1302273, 0.09354581, 0.08898163, 0.1261925, 0.1128755, 
    0.182023, 0.1498376, 0.1762683, 0.165635, 0.1790788, 0.1998697, 0.136218, 
    0.1645002, 0.1715576, 0.1716454, 0.1697011, 0.1760921, 0.2161418, 
    0.202068, 0.07065573, 0.05012651, 0.05139031,
  0.1307964, 0.17098, 0.1732314, 0.1718563, 0.1894859, 0.1854577, 0.2020338, 
    0.1272999, 0.08204843, 0.1465073, 0.09159167, 0.135461, 0.1462666, 
    0.2047076, 0.2233803, 0.1948517, 0.2497643, 0.2120825, 0.2379051, 
    0.2116948, 0.1728315, 0.1734649, 0.1831865, 0.1578852, 0.1500365, 
    0.2097137, 0.2218568, 0.1715374, 0.1421068,
  0.2697055, 0.2384415, 0.2058257, 0.276833, 0.2711541, 0.2265049, 0.2508178, 
    0.2013912, 0.1556925, 0.110217, 0.07184491, 0.04263566, 0.1053709, 
    0.2075391, 0.2808052, 0.1792164, 0.1513707, 0.2219617, 0.2072937, 
    0.2161235, 0.1363623, 0.1449574, 0.1548225, 0.08515693, 0.1305836, 
    0.1516131, 0.190475, 0.2585704, 0.2506409,
  0.1519071, 0.2052127, 0.2535793, 0.24091, 0.2523153, 0.1752065, 0.1510499, 
    0.1398702, 0.1006285, 0.1171565, 0.1025857, 0.09469216, 0.1207086, 
    0.1515189, 0.1750067, 0.1136328, 0.09597231, 0.09890369, 0.09882827, 
    0.1609989, 0.1373594, 0.07818105, 0.05421839, -0.003529765, 0.07210736, 
    0.01179075, 0.005456336, 0.1225948, 0.149528,
  0.1025499, 0.1097175, 0.08233296, 0.09692261, 0.07420685, 0.05504708, 
    0.0691771, 0.08362351, 0.07087715, 0.07696855, 0.08645581, 0.09445979, 
    0.1033306, 0.1428427, 0.1548603, 0.1636805, 0.194571, 0.1834467, 
    0.1211563, 0.07600635, 0.03853599, 0.01085603, -0.0003232079, 
    -0.0008966154, 0.02766564, 0.002313553, -0.001276595, 0.05977362, 
    0.1007559,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -9.890031e-06, -9.890031e-06, 
    -9.890031e-06, -9.890031e-06, -9.890031e-06, -9.890031e-06, 
    -9.890031e-06, -0.0003017963, -0.0003017963, -0.0003017963, 
    -0.0003017963, -0.0003017963, -0.0003017963, -0.0003017963, 0,
  0.001585037, -5.397655e-05, 0, 0, 0, -0.0001842882, 0, 0, 0, 0, 0, 
    -2.981671e-05, 8.284889e-05, 0.0977654, 0.1534277, 0.1564369, 0.2260763, 
    0.3076191, 0.2039444, 0.1467008, 0.09383849, 0.04555356, 0.1169816, 
    0.2174816, 0.2363468, 0.2660164, 0.319593, 0.1353792, 0.02075537,
  0.1952794, 0.2647949, 0.3596333, 0.3660131, 0.08895279, 0.06791423, 
    0.1470614, 0.07550903, 0.05213136, 0.06533101, 0.07046663, 0.08973266, 
    0.1543506, 0.2953053, 0.25297, 0.2402188, 0.2501259, 0.3197842, 
    0.2640792, 0.2087587, 0.2493775, 0.2755589, 0.3035268, 0.3380632, 
    0.4132547, 0.2916408, 0.2401441, 0.2478635, 0.2519168,
  0.2094043, 0.2250062, 0.2756144, 0.2761599, 0.2693617, 0.2628223, 
    0.2606136, 0.2851384, 0.298907, 0.3045605, 0.2451309, 0.3059465, 
    0.2722211, 0.2447959, 0.2044959, 0.2142152, 0.2012598, 0.2084394, 
    0.3022872, 0.2781513, 0.2768462, 0.2501638, 0.2739898, 0.2614783, 
    0.2714776, 0.2758763, 0.1977112, 0.1835877, 0.1782564,
  0.1494925, 0.2001506, 0.1911153, 0.185921, 0.1920055, 0.1495284, 0.1487549, 
    0.1594162, 0.1648042, 0.1748468, 0.2120873, 0.1942286, 0.1691732, 
    0.1101082, 0.1014034, 0.0705907, 0.1248661, 0.1367096, 0.1360998, 
    0.1441005, 0.1381867, 0.1323974, 0.1858728, 0.1364352, 0.0952734, 
    0.1764188, 0.1635345, 0.1259347, 0.1204776,
  0.0758303, 0.06637591, 0.02863494, 0.06604835, 0.06797591, 0.05216309, 
    0.05870393, 0.04463234, 0.01703523, 0.03708563, 0.06384286, 0.04214461, 
    0.07916386, 0.1282554, 0.0625848, 0.03056605, 0.07967594, 0.1330006, 
    0.09787228, 0.08547702, 0.08235346, 0.1031931, 0.05118208, 0.01807955, 
    0.04060922, 0.06624328, 0.07377532, 0.09237237, 0.08131724,
  0.007709173, 1.13653e-05, 0.0371552, 0.01805684, 0.04169728, 0.1093089, 
    0.0659752, 0.03909644, 0.02809232, 0.01982292, 0.1077773, 0.08156092, 
    0.04797775, 0.09393119, 0.02398752, 0.04515766, 0.06934569, 0.1154007, 
    0.09591928, 0.06736386, 0.04076911, 0.02108303, 0.005324531, 
    0.0004753818, 0.04896992, 0.03066776, 0.1273459, 0.03121358, 0.009563986,
  4.630904e-05, 0.04461782, 0.04582034, 0.01666448, 0.1477686, 0.02819146, 
    0.06130802, 0.03387057, 0.01788822, 0.002607259, 0.0338846, 0.01695535, 
    0.03446045, 0.06282224, 0.08781376, 0.1376772, 0.08353439, 0.04947678, 
    0.04102074, 0.009711024, 0.001285168, 3.29369e-07, 7.284206e-06, 
    0.007998126, 0.05098221, 0.1146496, 0.07171284, 0.004052422, 4.492584e-06,
  0.003231433, 0.08780155, 0.1796919, 0.07221066, 0.0322852, 0.03123486, 
    0.03559581, 0.05249609, 0.05843865, 0.03447327, 0.05348319, 0.06322519, 
    0.04008748, 0.03959789, 0.1023348, 0.07984272, 0.04553794, 0.06164526, 
    0.01533229, 0.0001773046, -4.403624e-06, 5.134032e-06, 0.005382843, 
    0.1489759, 0.2064895, 0.107246, 0.02078423, 0.0008896747, 7.489073e-05,
  0.06679169, 0.05315469, 0.06849001, 0.01529961, 0.01503112, 0.01593489, 
    0.01489554, 0.009762393, 0.06964011, 0.1885755, 0.02736891, 0.02303975, 
    0.04604571, 0.02292752, 0.02063127, 0.02901514, 0.01120985, 0.0007162922, 
    0.002058058, 0.01135324, 0.01484875, 0.002666776, 0.09524699, 0.05997673, 
    0.1295943, 0.07803687, 0.0117341, 0.01063362, 0.01110933,
  0.0003027406, 0.0005586427, 0.01749041, 0.002292892, 7.679519e-05, 
    0.002946944, 0.002275108, 0.0309122, 0.01534507, 0.02018607, 0.0354264, 
    0.03641656, 0.0368522, 0.05658015, 0.006669919, 0.02396743, 0.03272742, 
    0.08147314, 0.06609134, 0.05812056, 0.01678093, 0.007740087, 
    0.0006250226, 0.0006292541, 0.002935595, 0.000304854, 6.532627e-05, 
    1.477459e-05, 0.01013673,
  0.004268056, 0.009479347, 6.201653e-06, 0.005115324, 0.00930714, 
    4.185452e-05, 0.0004647087, 0.007368262, 0.005970874, 0.01551984, 
    0.01822597, 0.03159808, 0.01931635, 0.01354415, 0.0009149682, 
    0.0001975068, 0.01509633, 0.003085682, 0.06596414, 0.01327485, 0.0295443, 
    0.03143562, 0.004629993, 0.001452822, 0.001126864, 0.01144778, 
    0.0002060305, 0.008684073, 0.01229704,
  0.01637232, 0.007819058, 0.00536037, 0.002348002, 0.06097572, 0.02176238, 
    0.06379046, 0.09123036, 0.2345746, 0.1769174, 0.1533802, 0.09826638, 
    0.1098725, 0.07455398, 0.03558598, 0.02947719, 0.04759277, 0.03612307, 
    0.01787348, 0.0176815, 0.01436004, 0.05974489, 0.08093357, 0.04355708, 
    0.04060543, 0.04229175, 0.0390668, 0.0605551, 0.004416746,
  0.01988319, 0.06634709, 0.09832122, 0.1172118, 0.1012078, 0.08528996, 
    0.1925491, 0.09251049, 0.0779361, 0.07017021, 0.1320301, 0.1097386, 
    0.1601968, 0.1528603, 0.1763002, 0.1626569, 0.1722905, 0.170699, 
    0.1093098, 0.1544774, 0.186663, 0.1732755, 0.1682235, 0.1819639, 
    0.2178248, 0.2020076, 0.05720504, 0.0466282, 0.03574517,
  0.1167668, 0.1695883, 0.184417, 0.1623747, 0.1835869, 0.1814648, 0.1864413, 
    0.186811, 0.1243082, 0.1641794, 0.1206899, 0.1592002, 0.1556206, 
    0.206717, 0.2386637, 0.2083462, 0.2476112, 0.2181423, 0.2320247, 
    0.2072255, 0.1549428, 0.1607891, 0.2072782, 0.1804591, 0.1601681, 
    0.207956, 0.2265178, 0.1628321, 0.1286476,
  0.2616243, 0.2402333, 0.2059352, 0.2873435, 0.2914498, 0.2359537, 
    0.2743348, 0.2365215, 0.2095118, 0.1812159, 0.1018293, 0.07908136, 
    0.1619048, 0.2428405, 0.2834903, 0.1748923, 0.1651032, 0.2399881, 
    0.2653741, 0.2248861, 0.1351141, 0.1618634, 0.1762804, 0.1918872, 
    0.1779684, 0.1819564, 0.1982939, 0.256651, 0.2350199,
  0.2522566, 0.2392038, 0.3258466, 0.2373199, 0.2374249, 0.20049, 0.2058927, 
    0.2014523, 0.1539564, 0.167731, 0.155187, 0.1239336, 0.1537652, 
    0.1383211, 0.1611967, 0.1223584, 0.1321085, 0.1222548, 0.1067914, 
    0.1721569, 0.1931686, 0.09439453, 0.09930001, 0.01848072, 0.130498, 
    0.02614222, 0.01661355, 0.2183265, 0.220653,
  0.1336831, 0.1352325, 0.1166161, 0.1261609, 0.08957167, 0.07954416, 
    0.122069, 0.1672644, 0.1526489, 0.1641495, 0.1750383, 0.159083, 
    0.1630621, 0.1939332, 0.2147878, 0.2341017, 0.2509625, 0.2225164, 
    0.1657695, 0.1206193, 0.09382547, 0.08432488, 0.02992364, -0.002126332, 
    0.07425402, 0.01513149, 0.02503946, 0.08987327, 0.2130053,
  0.009743326, 0.008572483, 0.007401641, 0.006230798, 0.005059956, 
    0.003889113, 0.002718271, 0.001629701, 0.001603721, 0.001577741, 
    0.001551761, 0.001525781, 0.001499801, 0.001473821, 0.002459998, 
    0.003356234, 0.00425247, 0.005148705, 0.006044941, 0.006941176, 
    0.007837411, 0.005742474, 0.006043062, 0.006343649, 0.006644236, 
    0.006944823, 0.00724541, 0.007545997, 0.01068,
  0.0104968, 0.002003451, -4.617024e-05, 0, -1.2865e-06, -0.001355148, 
    -0.0001243053, 0, 0, 0, 0, 0.0005394376, 0.002199296, 0.163988, 
    0.2021272, 0.2003934, 0.2587158, 0.3136967, 0.2647662, 0.1904322, 
    0.152562, 0.1127949, 0.1654867, 0.232765, 0.2435434, 0.2623105, 
    0.3193565, 0.2366281, 0.06107572,
  0.2356074, 0.2770256, 0.3381353, 0.3807272, 0.1581707, 0.1050207, 
    0.1701474, 0.1273822, 0.107079, 0.110289, 0.1479517, 0.1351621, 
    0.1602576, 0.3240982, 0.259995, 0.2381783, 0.2867865, 0.3159563, 
    0.2672548, 0.2201677, 0.240473, 0.2806047, 0.3116573, 0.356892, 
    0.4372047, 0.290832, 0.2849682, 0.2588088, 0.2706107,
  0.2191628, 0.2540779, 0.2820312, 0.2889438, 0.2676708, 0.2640004, 
    0.2764718, 0.3121356, 0.3094483, 0.3027455, 0.2572258, 0.3034058, 
    0.290403, 0.2486381, 0.2184143, 0.2207212, 0.1948674, 0.2043813, 
    0.3006894, 0.2895782, 0.2810598, 0.2741773, 0.2551102, 0.2506063, 
    0.2910582, 0.2821304, 0.1945189, 0.1987925, 0.1962871,
  0.1529445, 0.1904568, 0.2042246, 0.1869166, 0.1847726, 0.1581984, 
    0.1503914, 0.1474592, 0.1524724, 0.1809932, 0.220031, 0.1862045, 
    0.1720595, 0.0982663, 0.09557994, 0.06668855, 0.1284161, 0.1459563, 
    0.1499306, 0.1389308, 0.1206198, 0.1402244, 0.1888196, 0.1354527, 
    0.09395973, 0.1542103, 0.1614753, 0.1312933, 0.1180765,
  0.06875585, 0.06225882, 0.02713197, 0.07355817, 0.06266187, 0.05371604, 
    0.05353909, 0.04218179, 0.02413876, 0.0313739, 0.06432832, 0.03751649, 
    0.07673462, 0.1330065, 0.0628376, 0.03460994, 0.08644912, 0.1320319, 
    0.09800258, 0.07324751, 0.08028334, 0.09990798, 0.04618439, 0.01728633, 
    0.04557284, 0.07007524, 0.0700876, 0.08464716, 0.07585486,
  0.008253685, 1.539048e-06, 0.04190756, 0.01360313, 0.04059701, 0.1242182, 
    0.05476251, 0.03889195, 0.02602242, 0.01230572, 0.09847911, 0.08571128, 
    0.05065875, 0.09676494, 0.0200658, 0.04167385, 0.07411689, 0.1036191, 
    0.09454743, 0.06115884, 0.04322035, 0.02173226, 0.005794113, 
    0.0006753972, 0.04787698, 0.02781814, 0.123476, 0.02816813, 0.02197317,
  8.016127e-06, 0.05098344, 0.05408739, 0.02488827, 0.1689583, 0.02643943, 
    0.07021245, 0.03491814, 0.02391909, 0.003216663, 0.03631369, 0.02342412, 
    0.03695916, 0.07423933, 0.1072838, 0.1543757, 0.09251297, 0.06265442, 
    0.04887477, 0.01182439, 0.001251963, 1.73128e-05, 4.355143e-05, 
    0.003803455, 0.06957403, 0.1178143, 0.0737731, 0.003448847, 1.065999e-06,
  0.004250939, 0.09661664, 0.2029627, 0.09142794, 0.02914554, 0.04352276, 
    0.04090412, 0.06534238, 0.07707846, 0.04601155, 0.06572013, 0.06883435, 
    0.05777546, 0.05573169, 0.1263051, 0.07208939, 0.05494205, 0.06848937, 
    0.02233053, 0.0008355819, 0.0002751699, 0.006239295, 0.002669552, 
    0.1781271, 0.2483572, 0.1376304, 0.02290731, 0.0009967985, 0.0001639308,
  0.09896629, 0.09938774, 0.09906811, 0.02010088, 0.01674781, 0.01995749, 
    0.01797058, 0.01339275, 0.08553238, 0.2110685, 0.03225428, 0.02917597, 
    0.05482963, 0.03142416, 0.02653189, 0.03199416, 0.01460048, 0.001479564, 
    0.003787155, 0.007997856, 0.01211991, 0.01933609, 0.1105386, 0.0889634, 
    0.1282752, 0.0965028, 0.01230633, 0.009678871, 0.04173274,
  0.002236739, 0.0007293779, 0.03166514, 0.03178928, 6.798958e-06, 
    0.002887162, 0.002757326, 0.03312166, 0.01582645, 0.02482674, 0.04599199, 
    0.03909788, 0.04746023, 0.06026965, 0.007193554, 0.0375162, 0.03363818, 
    0.0730713, 0.06078969, 0.05873584, 0.01943346, 0.01348052, 0.001502692, 
    0.00220751, 0.004987611, 0.0005549802, 6.287679e-05, 9.504145e-05, 
    0.0116714,
  0.001020148, 0.003787826, 0.001622778, 0.007169169, 0.005731173, 
    6.822815e-06, 0.002736319, 0.005264261, 0.006152079, 0.04213589, 
    0.008334348, 0.03335606, 0.0140802, 0.01155599, 0.0001520564, 
    0.0007642198, 0.02276232, 0.0171651, 0.05593494, 0.009287398, 0.02620881, 
    0.03828215, 0.006281232, 0.004286988, 0.001635138, 0.01631406, 
    0.001571418, 0.003607735, 0.01210933,
  0.007135781, 0.001683271, 0.007747593, 0.005745119, 0.07557514, 0.02189638, 
    0.07763939, 0.102096, 0.2366146, 0.182934, 0.1483624, 0.1024552, 
    0.1181334, 0.07067802, 0.03914739, 0.02951799, 0.04908422, 0.03287969, 
    0.01839982, 0.01259492, 0.01020083, 0.06272885, 0.07816732, 0.03245113, 
    0.03659714, 0.0450298, 0.03872463, 0.04348328, 0.007405385,
  0.01662287, 0.06112218, 0.0956293, 0.125229, 0.09155793, 0.07309517, 
    0.2016694, 0.06132447, 0.06721644, 0.0603904, 0.1361556, 0.1084148, 
    0.1436468, 0.1478446, 0.1753708, 0.1597154, 0.1667957, 0.1498615, 
    0.09952005, 0.1456408, 0.1863635, 0.1752885, 0.1553747, 0.1728942, 
    0.2049165, 0.1898463, 0.05052718, 0.04568382, 0.02794842,
  0.09102601, 0.1747021, 0.183669, 0.1540307, 0.177981, 0.1896446, 0.1748121, 
    0.2037085, 0.1533678, 0.1602129, 0.1423245, 0.1700716, 0.1569845, 
    0.2162668, 0.2520078, 0.2028975, 0.2407714, 0.227917, 0.2208401, 
    0.2034665, 0.146645, 0.1462061, 0.2093177, 0.1960396, 0.1688293, 
    0.2077799, 0.2206937, 0.1574659, 0.1105118,
  0.2724204, 0.2381989, 0.2015261, 0.2667923, 0.292468, 0.245363, 0.2702946, 
    0.234825, 0.2265263, 0.2311788, 0.1165006, 0.128561, 0.2013275, 
    0.2726785, 0.3032953, 0.1629633, 0.1679146, 0.2587456, 0.2688764, 
    0.213811, 0.1291592, 0.1479338, 0.1871219, 0.2095208, 0.2150426, 
    0.1923549, 0.187252, 0.250535, 0.2576525,
  0.256486, 0.2285135, 0.3238615, 0.2313735, 0.238455, 0.2069946, 0.2345064, 
    0.2480239, 0.1941943, 0.1859942, 0.1509842, 0.1311414, 0.15486, 
    0.1293697, 0.151994, 0.1270035, 0.1391068, 0.1299513, 0.1087962, 
    0.1636038, 0.1997761, 0.1031647, 0.1349666, 0.03412105, 0.1958307, 
    0.05096839, 0.03951286, 0.273277, 0.2001671,
  0.1332779, 0.1427612, 0.1165082, 0.1304077, 0.1107013, 0.09269065, 
    0.1529341, 0.2192657, 0.2368096, 0.2334275, 0.2226968, 0.1899679, 
    0.1579934, 0.192645, 0.2254355, 0.2320388, 0.2742421, 0.2473501, 
    0.1865327, 0.166582, 0.1365475, 0.1529808, 0.1284345, 0.03981566, 
    0.1278467, 0.03943329, 0.06148257, 0.1963317, 0.2183594,
  0.03551299, 0.03468518, 0.03385737, 0.03302956, 0.03220176, 0.03137395, 
    0.03054614, 0.02852193, 0.02813364, 0.02774536, 0.02735707, 0.02696879, 
    0.0265805, 0.02619222, 0.01806052, 0.02089036, 0.0237202, 0.02655005, 
    0.02937989, 0.03220973, 0.03503957, 0.04385772, 0.04224396, 0.04063021, 
    0.03901646, 0.03740271, 0.03578896, 0.03417521, 0.03617523,
  0.03881848, 0.01895798, 0.001156323, -3.085437e-11, -0.0004413194, 
    0.005559039, 0.003045338, -0.0002796789, 9.542025e-07, 1.786743e-05, 
    -0.000602141, 0.008101675, 0.02156232, 0.2121493, 0.1903615, 0.2028681, 
    0.2976407, 0.3310031, 0.2954578, 0.2615928, 0.2217515, 0.1790405, 
    0.1986697, 0.2522747, 0.2692164, 0.2972391, 0.3414817, 0.2533563, 
    0.1221684,
  0.2357965, 0.2872579, 0.3215876, 0.3736158, 0.2293241, 0.132177, 0.1805262, 
    0.1952583, 0.1520397, 0.1777446, 0.2142996, 0.1690156, 0.1615915, 
    0.3448191, 0.2734811, 0.249165, 0.325315, 0.3235505, 0.2954106, 
    0.2354892, 0.2618497, 0.2868521, 0.3114167, 0.3596233, 0.4587605, 
    0.2932051, 0.2949042, 0.2423086, 0.2966818,
  0.2324072, 0.2784474, 0.2894135, 0.3140879, 0.2582234, 0.2622527, 
    0.3007316, 0.3134077, 0.3120412, 0.3332469, 0.2417616, 0.3029132, 
    0.2716231, 0.2462764, 0.2144853, 0.2073518, 0.221857, 0.2232376, 
    0.3185713, 0.2711897, 0.2586032, 0.2386155, 0.2687897, 0.2588618, 
    0.2928126, 0.2727746, 0.2193541, 0.2104043, 0.2039818,
  0.1523604, 0.1968226, 0.1975242, 0.1983461, 0.1830947, 0.1461519, 
    0.1383878, 0.1551659, 0.1604576, 0.2040183, 0.2436648, 0.1898804, 
    0.1692448, 0.1147974, 0.1002921, 0.07141379, 0.1304525, 0.1500422, 
    0.1349786, 0.155353, 0.1252914, 0.1297273, 0.1920498, 0.1358915, 
    0.08978192, 0.1439396, 0.1647783, 0.1222513, 0.1263202,
  0.06923957, 0.0640161, 0.02797001, 0.06870306, 0.05389856, 0.04635467, 
    0.05371654, 0.04128572, 0.02874775, 0.03197176, 0.06098221, 0.04194525, 
    0.0805975, 0.1378047, 0.06133698, 0.03675147, 0.0962793, 0.1293434, 
    0.09894252, 0.07525979, 0.08386002, 0.09566621, 0.04430443, 0.01583228, 
    0.05189936, 0.07187443, 0.06766855, 0.08306916, 0.08187048,
  0.007578552, 8.334733e-06, 0.04221006, 0.01402026, 0.04753949, 0.1387037, 
    0.05740444, 0.05088793, 0.02004708, 0.01324137, 0.09562617, 0.07832014, 
    0.06215745, 0.09822918, 0.02735538, 0.04703162, 0.07514073, 0.09753207, 
    0.1005886, 0.05985555, 0.04654792, 0.03521515, 0.007091926, 0.0003012575, 
    0.04832233, 0.02828592, 0.1308106, 0.0282967, 0.02289564,
  0.0001334315, 0.06119445, 0.05825987, 0.03048255, 0.18826, 0.02999178, 
    0.08347158, 0.04122671, 0.02386133, 0.004267177, 0.03892914, 0.0275379, 
    0.03861316, 0.07706884, 0.1092808, 0.1612196, 0.1021787, 0.0713158, 
    0.05701824, 0.01988425, 0.003152414, 2.011856e-05, 5.541026e-05, 
    0.001781944, 0.07541756, 0.1210089, 0.0864353, 0.001969579, 1.558318e-06,
  0.0032914, 0.08668487, 0.2362326, 0.114157, 0.03359343, 0.0446403, 
    0.04385786, 0.07287624, 0.08790249, 0.05274933, 0.06853139, 0.08655411, 
    0.08729331, 0.06910004, 0.1353228, 0.09182526, 0.06535157, 0.07206466, 
    0.0204129, 0.001873043, 6.951866e-05, 0.009300303, 0.01312568, 0.2150498, 
    0.28553, 0.1769994, 0.03375177, 0.0009247321, 0.0001482415,
  0.1123821, 0.1463271, 0.1387579, 0.03562397, 0.01592217, 0.02347283, 
    0.02272467, 0.01415444, 0.09591728, 0.2462617, 0.04408101, 0.03015433, 
    0.06316651, 0.04137766, 0.03460842, 0.03634849, 0.01639152, 0.001481881, 
    0.004752186, 0.007025433, 0.009863871, 0.01738304, 0.1189684, 0.1413531, 
    0.143686, 0.103368, 0.01101901, 0.008401267, 0.01671824,
  0.01139617, 0.004016058, 0.022158, 0.1124573, 1.43844e-05, 0.002411181, 
    0.00323011, 0.04216761, 0.01852219, 0.02658908, 0.05549754, 0.04477643, 
    0.0604196, 0.06508242, 0.01294509, 0.0355104, 0.0368961, 0.07427034, 
    0.05725011, 0.06134604, 0.0243778, 0.01506254, 0.003666941, 0.002960372, 
    0.00369118, 0.0009871462, 1.559985e-06, 0.001066481, 0.03260556,
  2.090454e-05, -2.297696e-05, 0.01380585, 0.01520776, 0.001622726, 
    2.502919e-07, 0.00827309, 0.004151778, 0.01050337, 0.04374041, 
    0.003767637, 0.03877022, 0.01762572, 0.01165108, 4.089244e-05, 
    0.001661974, 0.02893498, 0.01378023, 0.04719225, 0.009883105, 0.03476411, 
    0.03917807, 0.006481107, 0.006453601, 0.003967155, 0.02800415, 
    0.003088515, 0.0006240264, 0.0002170131,
  0.0028937, 0.0003872017, 0.01103062, 0.006821463, 0.07943977, 0.01875137, 
    0.06365447, 0.1072865, 0.2233306, 0.1968168, 0.150328, 0.1039741, 
    0.1206756, 0.07801592, 0.04243411, 0.03840783, 0.04948874, 0.03472617, 
    0.02371765, 0.009287756, 0.01066971, 0.06189682, 0.07329991, 0.03048459, 
    0.03948344, 0.05600231, 0.03117149, 0.03832562, 0.005724351,
  0.01420092, 0.05891715, 0.08567934, 0.1374839, 0.08736365, 0.06121663, 
    0.2008151, 0.03967108, 0.05762564, 0.06835161, 0.1392923, 0.1082788, 
    0.1379611, 0.138621, 0.1779264, 0.1572214, 0.1688538, 0.1454823, 
    0.1003125, 0.1396367, 0.1862666, 0.1773598, 0.1603455, 0.1679535, 
    0.2037697, 0.1885199, 0.05665633, 0.03896219, 0.02738669,
  0.09023918, 0.184247, 0.1746012, 0.1730566, 0.1872015, 0.1940573, 
    0.1716539, 0.2065748, 0.1480562, 0.1738322, 0.1358664, 0.1693623, 
    0.1447191, 0.2280379, 0.2533516, 0.2128207, 0.2460995, 0.2289357, 
    0.207151, 0.1917586, 0.1376449, 0.1406215, 0.1955539, 0.2023198, 
    0.1778584, 0.2114263, 0.216413, 0.1567524, 0.1059446,
  0.2726556, 0.2416203, 0.1929134, 0.25868, 0.3134716, 0.2599079, 0.2679671, 
    0.2463754, 0.2233514, 0.2636405, 0.1247447, 0.1479865, 0.2300877, 
    0.2814443, 0.3043084, 0.1712495, 0.1636117, 0.2721338, 0.268681, 
    0.2007201, 0.1207924, 0.1528981, 0.1903142, 0.2275543, 0.2254088, 
    0.1857834, 0.1730178, 0.2458047, 0.2522465,
  0.2437289, 0.2199483, 0.3281422, 0.2376669, 0.2516099, 0.2318329, 
    0.2409302, 0.272313, 0.2327304, 0.20983, 0.1520269, 0.1511873, 0.1704088, 
    0.1201712, 0.1370877, 0.1271665, 0.1376878, 0.1364496, 0.1090247, 
    0.1648292, 0.2127597, 0.1327638, 0.1483062, 0.08439225, 0.2152664, 
    0.09615447, 0.06770756, 0.2620357, 0.1946728,
  0.1223372, 0.1364599, 0.1195914, 0.1345527, 0.1217508, 0.1053786, 
    0.1583295, 0.2352974, 0.2575274, 0.2507263, 0.2374303, 0.2195662, 
    0.1562983, 0.1698727, 0.2222832, 0.2356683, 0.2815005, 0.2259339, 
    0.1837782, 0.1671646, 0.1393608, 0.1642282, 0.1713297, 0.06951474, 
    0.1526902, 0.1036974, 0.109101, 0.194455, 0.2008385,
  0.04494985, 0.04452401, 0.04409817, 0.04367233, 0.04324649, 0.04282065, 
    0.04239481, 0.04948217, 0.05217825, 0.05487432, 0.0575704, 0.06026648, 
    0.06296256, 0.06565864, 0.06832737, 0.07043663, 0.07254589, 0.07465514, 
    0.0767644, 0.07887366, 0.08098292, 0.06834163, 0.06396213, 0.05958264, 
    0.05520315, 0.05082365, 0.04644416, 0.04206466, 0.04529052,
  0.08404982, 0.02118674, 0.01217865, -7.536334e-05, 0.0003242293, 
    0.01520038, 0.01526851, 0.006452288, 8.959186e-05, 0.0006559779, 
    0.009947496, 0.01924823, 0.06633724, 0.2202909, 0.1720043, 0.2276994, 
    0.3199354, 0.3593781, 0.3030071, 0.2956482, 0.2978824, 0.3009141, 
    0.2261061, 0.2463945, 0.267653, 0.3141418, 0.3556583, 0.27832, 0.2049894,
  0.2643746, 0.3060038, 0.3367264, 0.371575, 0.2861901, 0.1473061, 0.2153946, 
    0.2372962, 0.173373, 0.2175429, 0.2583076, 0.185724, 0.1707068, 
    0.3428807, 0.276342, 0.2802204, 0.3716968, 0.3142318, 0.248488, 
    0.2183507, 0.2380872, 0.2890573, 0.2855818, 0.383952, 0.4785015, 
    0.3085206, 0.3066535, 0.239585, 0.3202221,
  0.2442263, 0.27929, 0.3087494, 0.3363961, 0.2918183, 0.3005525, 0.3264831, 
    0.3592499, 0.3585472, 0.3291167, 0.2760705, 0.3129063, 0.2971209, 
    0.2237422, 0.226305, 0.2096089, 0.2231855, 0.2394785, 0.3043289, 
    0.2560601, 0.2655376, 0.2478863, 0.2770756, 0.2593536, 0.2996412, 
    0.294853, 0.2279901, 0.2216738, 0.2120819,
  0.1718701, 0.2099747, 0.1997719, 0.1883631, 0.1875146, 0.1512855, 0.139863, 
    0.1571007, 0.1637671, 0.1819233, 0.2305545, 0.1897276, 0.1800443, 
    0.1151028, 0.09075109, 0.09167416, 0.1358467, 0.1575294, 0.1528713, 
    0.1649326, 0.1351667, 0.1373996, 0.1861755, 0.1307351, 0.08772088, 
    0.1354603, 0.1587306, 0.1184648, 0.1315631,
  0.07714705, 0.0701641, 0.03082494, 0.06939769, 0.0561163, 0.04547646, 
    0.06082224, 0.04414693, 0.03977455, 0.03021677, 0.05727747, 0.05257984, 
    0.08723361, 0.14335, 0.07355422, 0.04639473, 0.1200027, 0.1373414, 
    0.1010151, 0.07703623, 0.0914377, 0.09035648, 0.04876156, 0.01863215, 
    0.04792944, 0.07436655, 0.07233036, 0.0843323, 0.08898478,
  0.007252962, 0.0003136148, 0.04952185, 0.01026157, 0.05650324, 0.1441932, 
    0.06875996, 0.04631944, 0.01150997, 0.01233511, 0.08974738, 0.07755515, 
    0.08842806, 0.1139184, 0.04623646, 0.04631142, 0.08334252, 0.09585322, 
    0.1068813, 0.06776926, 0.05356278, 0.04078623, 0.009108239, 0.0006528164, 
    0.05567356, 0.0334205, 0.136065, 0.03684719, 0.02104362,
  0.0003187816, 0.0709336, 0.06572711, 0.02683692, 0.1660758, 0.02822584, 
    0.09129486, 0.03262007, 0.01129147, 0.004034375, 0.03643097, 0.02970204, 
    0.04609768, 0.06807907, 0.1080375, 0.1485844, 0.1013143, 0.05355306, 
    0.05432822, 0.02221264, 0.008616443, 0.0002139463, 1.9416e-05, 
    0.0006056632, 0.06508134, 0.1539036, 0.0847833, 0.01032727, 4.319274e-06,
  0.002097235, 0.06488406, 0.2850527, 0.1154764, 0.02838494, 0.04012866, 
    0.03616719, 0.0618009, 0.07413872, 0.0484686, 0.06412855, 0.06579413, 
    0.08111154, 0.05089314, 0.1046501, 0.07984401, 0.05656742, 0.06322238, 
    0.01643296, 0.001996349, 6.641074e-05, 0.008046316, 0.006367136, 
    0.2258583, 0.2657021, 0.2066996, 0.0281795, 0.001708285, 0.000163584,
  0.0382279, 0.1492536, 0.1512654, 0.03865168, 0.01489915, 0.02429143, 
    0.01828781, 0.01350751, 0.1003737, 0.265953, 0.05771117, 0.02275426, 
    0.05220603, 0.03256932, 0.027211, 0.03283306, 0.01502657, 0.001954524, 
    0.003578637, 0.007502217, 0.01748754, 0.007274976, 0.1122244, 0.1707714, 
    0.1433583, 0.1001353, 0.01133433, 0.009955329, 0.008002914,
  0.008119639, 0.001434599, 0.007660533, 0.1790371, 8.574249e-06, 
    0.001391686, 0.004472272, 0.04293207, 0.01585898, 0.02486351, 0.05914389, 
    0.04153132, 0.05777595, 0.06072624, 0.01270462, 0.03494234, 0.03807373, 
    0.06302744, 0.04799612, 0.06044137, 0.02301302, 0.01424602, 0.006136524, 
    0.004453088, 0.003415594, 9.750459e-05, 0.0001571907, 0.001374588, 
    0.05050822,
  4.560868e-06, 6.150638e-07, 0.001274141, 0.02361424, 5.645557e-05, 
    1.052411e-07, 0.01442852, 0.005140366, 0.01702488, 0.03338049, 
    0.00186221, 0.0397137, 0.01131914, 0.008307078, 9.681901e-05, 
    0.003884223, 0.03168983, 0.007557618, 0.04487629, 0.01722131, 0.03005774, 
    0.04167894, 0.0122157, 0.01481212, 0.005814334, 0.03428309, 0.0009043356, 
    0.0008902319, 6.69723e-06,
  0.001362268, 0.001049927, 0.009437421, 0.007375539, 0.07065637, 0.01544428, 
    0.03541293, 0.112104, 0.2080623, 0.2123356, 0.1483409, 0.107688, 
    0.1142133, 0.07161238, 0.05318866, 0.04321562, 0.05756316, 0.03841847, 
    0.02458904, 0.006576379, 0.01630509, 0.05440475, 0.0599748, 0.04147781, 
    0.04653888, 0.06882419, 0.03224095, 0.02447973, 0.0009262752,
  0.01549783, 0.04821171, 0.08131891, 0.1489676, 0.08554211, 0.04927317, 
    0.2002153, 0.02477686, 0.04744473, 0.07201019, 0.1346722, 0.1100522, 
    0.1345798, 0.1424524, 0.173801, 0.1575256, 0.1611728, 0.1452326, 
    0.1026366, 0.1406974, 0.1882056, 0.171296, 0.154296, 0.1655593, 
    0.1965531, 0.1862225, 0.05439916, 0.03786452, 0.02545515,
  0.08039922, 0.1805987, 0.1739202, 0.1766541, 0.1689309, 0.1768521, 
    0.1712424, 0.2027002, 0.1318484, 0.175592, 0.1362182, 0.1655454, 
    0.1265872, 0.2239608, 0.260015, 0.2318674, 0.2424527, 0.2467529, 
    0.2061596, 0.180439, 0.1344028, 0.138778, 0.1973052, 0.2036751, 
    0.1687208, 0.2102797, 0.2161219, 0.154257, 0.09787301,
  0.26403, 0.2368135, 0.2230334, 0.2623953, 0.3046516, 0.2511033, 0.2511363, 
    0.2429624, 0.2185415, 0.2671066, 0.145335, 0.1417658, 0.24362, 0.2993316, 
    0.3178839, 0.1793396, 0.1632408, 0.2928759, 0.2637402, 0.214238, 
    0.1180434, 0.1608634, 0.2002426, 0.2870238, 0.2354776, 0.1983189, 
    0.1844909, 0.275221, 0.2656557,
  0.2576702, 0.2327573, 0.3273786, 0.2378428, 0.282945, 0.2369701, 0.2579459, 
    0.3008694, 0.2468688, 0.2144366, 0.1830937, 0.1857321, 0.1729095, 
    0.1301885, 0.1210577, 0.1280592, 0.1332621, 0.1393136, 0.1075735, 
    0.1637878, 0.2316211, 0.1405153, 0.1658943, 0.1034232, 0.2211526, 
    0.1531871, 0.1004649, 0.2528485, 0.2010076,
  0.1047061, 0.1232872, 0.1274096, 0.1439753, 0.132905, 0.1337535, 0.171305, 
    0.2423583, 0.2671849, 0.2477196, 0.2547603, 0.2368443, 0.1612338, 
    0.1551756, 0.211589, 0.2256789, 0.2623079, 0.2057492, 0.1753828, 
    0.1623894, 0.1368424, 0.1750882, 0.1618449, 0.08739997, 0.1517001, 
    0.1172483, 0.1463462, 0.1824002, 0.1895468,
  0.08553489, 0.08394194, 0.08234897, 0.08075602, 0.07916306, 0.0775701, 
    0.07597714, 0.08869432, 0.09617741, 0.1036605, 0.1111436, 0.1186267, 
    0.1261098, 0.1335929, 0.1363201, 0.135951, 0.1355819, 0.1352128, 
    0.1348438, 0.1344747, 0.1341056, 0.1261235, 0.1206025, 0.1150814, 
    0.1095603, 0.1040393, 0.09851824, 0.09299718, 0.08680926,
  0.175584, 0.03795581, 0.02152915, 0.007667809, 0.01111486, 0.03860568, 
    0.02970476, 0.01953454, 0.01192804, 0.02780454, 0.04125502, 0.06852109, 
    0.1633897, 0.2532337, 0.1827052, 0.3172728, 0.3628134, 0.383106, 
    0.2996037, 0.294618, 0.3362775, 0.3567807, 0.2411218, 0.2631939, 
    0.3396037, 0.3370414, 0.3642692, 0.3196976, 0.218766,
  0.3142314, 0.3507543, 0.3564557, 0.3962966, 0.294016, 0.146183, 0.2760863, 
    0.2568138, 0.1800884, 0.2533879, 0.2971859, 0.1985855, 0.1792725, 
    0.3635883, 0.2797257, 0.2744836, 0.3370696, 0.2835102, 0.2579387, 
    0.3149911, 0.3294802, 0.2938451, 0.3171112, 0.3563753, 0.4709632, 
    0.3349952, 0.3290668, 0.273548, 0.3254355,
  0.2654194, 0.3096395, 0.312689, 0.3526975, 0.2982243, 0.3055665, 0.3042738, 
    0.3628474, 0.3239577, 0.3543093, 0.2655396, 0.2982572, 0.3058653, 
    0.2504784, 0.2397856, 0.2137237, 0.2369729, 0.253926, 0.3103363, 
    0.280849, 0.2782733, 0.2506554, 0.2814912, 0.2775286, 0.2906689, 
    0.2887177, 0.2246259, 0.2350927, 0.2196766,
  0.1795305, 0.2194353, 0.2066761, 0.2200778, 0.1972314, 0.173386, 0.1515954, 
    0.1665615, 0.1639016, 0.1875977, 0.2506469, 0.196759, 0.1743485, 
    0.1208392, 0.09076861, 0.104219, 0.1445865, 0.1658515, 0.1523505, 
    0.1810329, 0.1387843, 0.1462565, 0.2006581, 0.1269504, 0.0849613, 
    0.1406522, 0.1616088, 0.1341207, 0.1416789,
  0.09510998, 0.07962148, 0.03553547, 0.07431623, 0.06950482, 0.05513065, 
    0.07126771, 0.05388587, 0.05358793, 0.03528408, 0.06518743, 0.04901873, 
    0.1004806, 0.1528946, 0.08704205, 0.05548803, 0.1285376, 0.1471496, 
    0.1099694, 0.09015303, 0.09596628, 0.09457013, 0.05680751, 0.02238182, 
    0.04912478, 0.07799942, 0.07553181, 0.08783752, 0.0982309,
  0.009557237, 7.479034e-05, 0.05982033, 0.01118604, 0.06300494, 0.1298025, 
    0.1004641, 0.04070022, 0.002266052, 0.008995055, 0.07373358, 0.05403098, 
    0.09726406, 0.113733, 0.04985608, 0.05561419, 0.09597477, 0.0847716, 
    0.1030959, 0.07783086, 0.05659432, 0.04935104, 0.01227053, 0.0008215868, 
    0.0592366, 0.03231312, 0.1288533, 0.04160674, 0.02065697,
  0.0003160336, 0.07183011, 0.06441704, 0.02563892, 0.1439968, 0.02807891, 
    0.08562892, 0.03101697, 0.007847724, 0.002302841, 0.03574925, 0.04203037, 
    0.05330403, 0.05848671, 0.1066286, 0.1305944, 0.08996549, 0.04013069, 
    0.05737922, 0.02967939, 0.02117405, 0.0007480264, 4.351002e-06, 
    3.92729e-05, 0.05095645, 0.172837, 0.06276669, 0.0151563, 0.0002327381,
  0.0004996742, 0.04694863, 0.3158726, 0.0781054, 0.020653, 0.03462869, 
    0.03038349, 0.05360775, 0.06414939, 0.04787514, 0.06450839, 0.0541745, 
    0.07841498, 0.03845433, 0.08252974, 0.05648244, 0.05426062, 0.05471414, 
    0.01701671, 0.002645117, 0.001946917, 0.005992705, 0.00464044, 0.1754953, 
    0.1987473, 0.1616287, 0.02187752, 0.003205056, 0.0002743668,
  0.008638632, 0.09571493, 0.08410254, 0.03946656, 0.01447987, 0.02437637, 
    0.01697107, 0.01304046, 0.0885051, 0.2313824, 0.06348077, 0.01934553, 
    0.0427894, 0.02922435, 0.02370264, 0.02904551, 0.01540258, 0.003903685, 
    0.003552433, 0.009103068, 0.0186891, 0.006089661, 0.0913524, 0.1543519, 
    0.1141436, 0.1000372, 0.01592964, 0.01297251, 0.003948394,
  0.001199541, 2.875753e-05, 0.0004543339, 0.2448473, -3.594442e-06, 
    0.001217215, 0.005920289, 0.04219181, 0.01455993, 0.0254915, 0.07046182, 
    0.04135942, 0.05435036, 0.05233691, 0.01139683, 0.03627905, 0.03502928, 
    0.0444054, 0.04416388, 0.05173824, 0.02267079, 0.01160594, 0.01299826, 
    0.007657977, 0.004140919, 0.0001462313, 4.021823e-05, 0.0002002345, 
    0.02224831,
  2.056185e-06, 5.117197e-07, 2.091826e-05, 0.02018798, 5.122299e-05, 
    5.973441e-08, 0.01079823, 0.005659416, 0.02626127, 0.02516343, 
    0.003028231, 0.0292289, 0.01163279, 0.007405043, 0.0006244997, 
    0.006358131, 0.029669, 0.002063575, 0.03940233, 0.009381208, 0.009639719, 
    0.04273947, 0.01451378, 0.02064326, 0.01001029, 0.0379553, 0.001143954, 
    2.883442e-05, 3.199099e-06,
  0.0006115723, 0.001524284, 0.01578155, 0.01023576, 0.06039413, 0.009179786, 
    0.01884894, 0.1108052, 0.1897983, 0.2157026, 0.1527134, 0.1162178, 
    0.1221961, 0.07584308, 0.07046034, 0.05447828, 0.0673857, 0.04728517, 
    0.03375816, 0.007322833, 0.02133842, 0.05271466, 0.06347584, 0.05717596, 
    0.05403992, 0.07490156, 0.02845459, 0.01124038, 9.982388e-06,
  0.01570675, 0.04219772, 0.08309753, 0.1564758, 0.07968536, 0.0379068, 
    0.197381, 0.01726436, 0.03150132, 0.0718158, 0.1298222, 0.1052963, 
    0.1359459, 0.1533909, 0.1709711, 0.1622028, 0.1480605, 0.1458618, 
    0.1142035, 0.1585381, 0.183172, 0.1620094, 0.1602288, 0.1674795, 
    0.1935703, 0.1968693, 0.05652827, 0.0383888, 0.02817059,
  0.08378179, 0.1972364, 0.1773034, 0.1885465, 0.1833625, 0.1904329, 
    0.1594708, 0.1840103, 0.1272825, 0.1693966, 0.1219001, 0.161599, 
    0.1115121, 0.225137, 0.2723421, 0.2397007, 0.2335618, 0.2389608, 0.20328, 
    0.1855966, 0.1391867, 0.1490042, 0.2120946, 0.2166569, 0.1714885, 
    0.2016956, 0.2200486, 0.1476126, 0.1047372,
  0.2714042, 0.2302588, 0.2200955, 0.2835804, 0.3635435, 0.2643572, 
    0.3011109, 0.2528998, 0.2266694, 0.2692713, 0.1549491, 0.1372815, 
    0.2452988, 0.3037596, 0.3367998, 0.1658831, 0.1661189, 0.2993317, 
    0.2685779, 0.2520116, 0.09990551, 0.183623, 0.2218728, 0.3045624, 
    0.243208, 0.2144093, 0.1978779, 0.2855505, 0.2761736,
  0.2632295, 0.2461227, 0.3309792, 0.2560004, 0.2980365, 0.2865657, 
    0.2615021, 0.3117619, 0.2866214, 0.2496952, 0.1983839, 0.1868441, 
    0.1793227, 0.1406074, 0.1126483, 0.14283, 0.1411421, 0.1466514, 
    0.1018995, 0.164737, 0.2473117, 0.1330871, 0.1802035, 0.09315654, 
    0.2280298, 0.2027183, 0.1385517, 0.2617276, 0.1973807,
  0.09940099, 0.1252833, 0.1165829, 0.1512507, 0.1373077, 0.1393831, 
    0.1672552, 0.2540234, 0.2774206, 0.2542456, 0.2376991, 0.2255572, 
    0.1724543, 0.1580078, 0.192456, 0.2468681, 0.2596244, 0.1969501, 
    0.1708339, 0.1467538, 0.1309092, 0.1680968, 0.1489473, 0.08090147, 
    0.1408942, 0.1473867, 0.1711314, 0.172276, 0.1925555,
  0.1237352, 0.1233966, 0.123058, 0.1227194, 0.1223808, 0.1220422, 0.1217036, 
    0.1441732, 0.1523292, 0.1604852, 0.1686412, 0.1767972, 0.1849532, 
    0.1931092, 0.1952063, 0.1962129, 0.1972194, 0.198226, 0.1992326, 
    0.2002392, 0.2012458, 0.1777214, 0.1688974, 0.1600734, 0.1512494, 
    0.1424254, 0.1336014, 0.1247774, 0.124006,
  0.2011472, 0.09734012, 0.02941583, 0.02693834, 0.03840627, 0.05969895, 
    0.04555135, 0.02777209, 0.02815323, 0.05289186, 0.05851324, 0.1315373, 
    0.2052315, 0.2829196, 0.2190923, 0.3028869, 0.3804907, 0.4039832, 
    0.3060136, 0.2896824, 0.3431833, 0.3754703, 0.2386652, 0.2582274, 
    0.2881321, 0.3219415, 0.3618778, 0.3550102, 0.2277309,
  0.3129985, 0.3229042, 0.3939779, 0.4167969, 0.2905139, 0.1455347, 0.259271, 
    0.2574463, 0.2012689, 0.2671249, 0.3251463, 0.2028629, 0.1804506, 
    0.3850079, 0.2884324, 0.3116232, 0.343704, 0.2984786, 0.2671646, 
    0.2988401, 0.3262267, 0.2916271, 0.3344049, 0.3966821, 0.4648578, 
    0.3615084, 0.3475217, 0.3096416, 0.3113354,
  0.2846414, 0.3334673, 0.338554, 0.3501343, 0.3209357, 0.3755513, 0.3359454, 
    0.3762758, 0.3847764, 0.3562993, 0.3077214, 0.3396148, 0.3308713, 
    0.2571568, 0.2466588, 0.2435103, 0.2418533, 0.2626112, 0.3131178, 
    0.3175234, 0.2743947, 0.2646092, 0.2845508, 0.2920996, 0.2993674, 
    0.2772914, 0.2297099, 0.2388539, 0.2673987,
  0.1981232, 0.2485212, 0.2253332, 0.2225198, 0.1957336, 0.1629133, 
    0.1672123, 0.1869918, 0.1781717, 0.19495, 0.2582921, 0.2078713, 
    0.1948682, 0.1495275, 0.1000069, 0.1221842, 0.165255, 0.1758856, 
    0.1728594, 0.2056648, 0.1529572, 0.1454338, 0.2154194, 0.1324979, 
    0.08338024, 0.1401817, 0.1797104, 0.1425842, 0.1453445,
  0.09641925, 0.08857289, 0.04118916, 0.08255094, 0.08031885, 0.0559955, 
    0.08590965, 0.06757847, 0.05402031, 0.05931412, 0.09144297, 0.05418114, 
    0.1102838, 0.1651233, 0.09610455, 0.0685009, 0.1457573, 0.1622339, 
    0.1047454, 0.08692257, 0.1014233, 0.1035375, 0.06492103, 0.02739263, 
    0.04307803, 0.08288504, 0.07394483, 0.08479307, 0.1060818,
  0.01399543, 0.0005437497, 0.05881618, 0.01307425, 0.06512192, 0.1167756, 
    0.1049809, 0.03683327, 0.0036708, 0.008600689, 0.04255448, 0.03134508, 
    0.1140564, 0.09448551, 0.04856272, 0.06218307, 0.09699075, 0.07546832, 
    0.0984292, 0.08158936, 0.05870902, 0.06312753, 0.02149828, 0.0003060806, 
    0.05980346, 0.03406023, 0.09983769, 0.03662448, 0.02345095,
  0.001381192, 0.05401857, 0.05881029, 0.02819276, 0.1296416, 0.02859325, 
    0.08443283, 0.03842674, 0.007559584, 0.00196409, 0.04538543, 0.04713427, 
    0.057826, 0.05636777, 0.1029561, 0.1159701, 0.0785365, 0.04101587, 
    0.06205464, 0.03987525, 0.03738721, 0.001245008, 1.878919e-06, 
    -1.835407e-05, 0.04713181, 0.1483482, 0.05781621, 0.02367095, 0.00218914,
  0.000242079, 0.04316146, 0.2310674, 0.061914, 0.01783031, 0.03282715, 
    0.02969734, 0.05158073, 0.05571812, 0.04810359, 0.06465955, 0.05056648, 
    0.07879142, 0.03333879, 0.06537618, 0.0488451, 0.05380192, 0.05374326, 
    0.02419808, 0.005897462, 3.046811e-05, 0.003112494, 0.0008075213, 
    0.1635885, 0.1830589, 0.1365878, 0.02192881, 0.003883855, 0.0003650086,
  0.002831884, 0.04192994, 0.03548113, 0.04546524, 0.01392482, 0.02490875, 
    0.01973727, 0.01421568, 0.07785241, 0.2123264, 0.06396845, 0.01701505, 
    0.03995375, 0.0249229, 0.02422456, 0.03122542, 0.01866231, 0.006465779, 
    0.005699634, 0.01720086, 0.01438295, 0.009249832, 0.07931693, 0.1366949, 
    0.1091117, 0.09535915, 0.02284516, 0.0128057, 0.00369961,
  0.0002248298, 5.747571e-06, -5.215754e-05, 0.2250977, -6.478244e-05, 
    0.001858841, 0.005807811, 0.04260655, 0.01305948, 0.02743416, 0.08217834, 
    0.0511362, 0.05576398, 0.05042249, 0.01218432, 0.02926905, 0.02909393, 
    0.03757566, 0.04604055, 0.05133937, 0.0285056, 0.01309748, 0.02122265, 
    0.01457935, 0.008277657, 0.0003180413, 2.343483e-06, 2.41748e-05, 
    0.007288866,
  1.527087e-06, 2.823055e-07, -1.164119e-05, 0.0102673, 5.527645e-06, 
    -2.319704e-09, 0.002056317, 0.003057086, 0.0339999, 0.01921593, 
    0.002682283, 0.02729812, 0.01628145, 0.008058202, 0.004215283, 
    0.01104157, 0.03336763, 0.001210515, 0.02639963, 0.007547374, 
    0.0004882108, 0.05759432, 0.01760377, 0.02887706, 0.01304958, 0.03558275, 
    0.00126073, 4.502407e-06, 1.214401e-06,
  0.00114579, 0.0009162828, 0.03500962, 0.0214838, 0.05171819, 0.005683476, 
    0.008284694, 0.1015802, 0.1688431, 0.2080205, 0.149396, 0.1241825, 
    0.123477, 0.07515558, 0.08763524, 0.06875245, 0.07618191, 0.07203843, 
    0.03506263, 0.01055124, 0.02574974, 0.05722976, 0.07159129, 0.06886562, 
    0.06856823, 0.07793896, 0.02811112, 0.008842199, -0.000168072,
  0.0145383, 0.04139639, 0.09198998, 0.1682304, 0.06735135, 0.03418617, 
    0.200646, 0.01359774, 0.0140396, 0.06493457, 0.1233413, 0.09977578, 
    0.1437071, 0.1700729, 0.1777548, 0.1628929, 0.1481137, 0.167278, 
    0.1198027, 0.150516, 0.1883994, 0.1501146, 0.1822567, 0.1678308, 
    0.1922135, 0.2164478, 0.06736185, 0.03911685, 0.02891998,
  0.09987111, 0.1977882, 0.1841012, 0.2001232, 0.2143732, 0.2344639, 
    0.179226, 0.1749618, 0.128125, 0.1491588, 0.1104756, 0.1545345, 
    0.1097339, 0.2476379, 0.305105, 0.2541116, 0.2519777, 0.2556979, 
    0.2006694, 0.1912132, 0.1424047, 0.1502017, 0.2229349, 0.2140335, 
    0.1618174, 0.211419, 0.2316054, 0.1443666, 0.1175992,
  0.2623291, 0.2323843, 0.2069277, 0.2879339, 0.4015166, 0.2746929, 
    0.2981295, 0.2420533, 0.2391866, 0.2735636, 0.1864148, 0.1285001, 
    0.2762157, 0.3064637, 0.3329223, 0.186452, 0.1599269, 0.2999561, 
    0.2877453, 0.2471067, 0.09103931, 0.1774662, 0.2281532, 0.3073001, 
    0.2245368, 0.2216717, 0.2185969, 0.2972505, 0.2727533,
  0.2655929, 0.2530788, 0.3573784, 0.3147438, 0.3448979, 0.2872441, 0.317369, 
    0.3370148, 0.3097527, 0.2560382, 0.2100818, 0.1825282, 0.1747538, 
    0.1337443, 0.1040738, 0.1568384, 0.1198239, 0.1403126, 0.09791987, 
    0.1630137, 0.2242942, 0.1223793, 0.1859383, 0.08523855, 0.2232331, 
    0.2930021, 0.1849138, 0.260708, 0.2123169,
  0.1314032, 0.1523883, 0.1592135, 0.167011, 0.1410776, 0.1660226, 0.1909394, 
    0.2656853, 0.2949093, 0.2464572, 0.2116161, 0.2049579, 0.1719368, 
    0.1505319, 0.1821308, 0.2271988, 0.2396228, 0.1737141, 0.161413, 
    0.1356826, 0.1302405, 0.1680266, 0.1367766, 0.06672285, 0.1228967, 
    0.1747342, 0.1735124, 0.1626776, 0.1879434,
  0.1758035, 0.1761597, 0.1765159, 0.176872, 0.1772282, 0.1775844, 0.1779406, 
    0.2077378, 0.218023, 0.2283082, 0.2385935, 0.2488787, 0.2591639, 
    0.2694491, 0.2713853, 0.2715655, 0.2717457, 0.2719259, 0.2721061, 
    0.2722862, 0.2724664, 0.2306374, 0.2198158, 0.2089942, 0.1981726, 
    0.187351, 0.1765294, 0.1657078, 0.1755185,
  0.2194188, 0.198608, 0.05135091, 0.04335243, 0.07508383, 0.08089654, 
    0.05398444, 0.03769356, 0.05527489, 0.04753926, 0.1232632, 0.1714818, 
    0.2598799, 0.2913354, 0.218505, 0.200259, 0.2937312, 0.3591788, 
    0.3228533, 0.2625172, 0.3461907, 0.3675019, 0.2422159, 0.226852, 
    0.2221414, 0.2459147, 0.3123613, 0.3500956, 0.2407478,
  0.3149187, 0.2685075, 0.3471764, 0.3821254, 0.2792026, 0.1482092, 
    0.2254231, 0.256382, 0.2282767, 0.2705992, 0.3374541, 0.2014938, 
    0.1972121, 0.3607845, 0.2893561, 0.3291375, 0.3326927, 0.3121216, 
    0.2524568, 0.266084, 0.2691339, 0.2408101, 0.2821172, 0.3774284, 
    0.4268313, 0.3272665, 0.3093223, 0.3055888, 0.2961292,
  0.2955815, 0.3439043, 0.3389616, 0.3563414, 0.3025955, 0.3275887, 
    0.3620676, 0.3909857, 0.3882548, 0.3242204, 0.3200713, 0.3412794, 
    0.3263506, 0.2611549, 0.2589535, 0.2517693, 0.269188, 0.2864855, 
    0.3359703, 0.3481215, 0.2797575, 0.271741, 0.2917267, 0.2916576, 
    0.3135032, 0.2809322, 0.2351531, 0.25086, 0.2647233,
  0.2235361, 0.2475237, 0.2370377, 0.2348827, 0.2089073, 0.1728866, 
    0.1709193, 0.2047803, 0.1945754, 0.2106561, 0.2845352, 0.2261104, 
    0.2243243, 0.1745525, 0.1162895, 0.1368267, 0.1933307, 0.2147947, 
    0.2076337, 0.230464, 0.1791149, 0.1628296, 0.2312392, 0.1434424, 
    0.0880311, 0.1402064, 0.192727, 0.1624098, 0.1644485,
  0.1038857, 0.1047288, 0.04788961, 0.09459687, 0.08890262, 0.05705971, 
    0.08440685, 0.07936645, 0.0668611, 0.08323638, 0.101541, 0.07011232, 
    0.09760968, 0.1687361, 0.1097098, 0.07777598, 0.1600664, 0.1656885, 
    0.09974481, 0.09729864, 0.1035964, 0.1151895, 0.07256973, 0.03042806, 
    0.03568099, 0.08684514, 0.07551127, 0.08233964, 0.1094566,
  0.01601182, 0.001893553, 0.05376118, 0.02270117, 0.06360468, 0.1046094, 
    0.0896062, 0.04203655, 0.006886636, 0.008473904, 0.02116669, 0.01324588, 
    0.09995775, 0.08282436, 0.05270518, 0.06447293, 0.09791967, 0.08595528, 
    0.0970283, 0.08814026, 0.06205624, 0.07958009, 0.02864666, 0.0001451888, 
    0.04536086, 0.04874382, 0.08753246, 0.03641824, 0.03095779,
  0.002631281, 0.04264603, 0.06185566, 0.02867832, 0.1274693, 0.02961496, 
    0.08114845, 0.05089826, 0.01009972, 0.002769023, 0.03138892, 0.0400724, 
    0.05970579, 0.05697548, 0.09241351, 0.1055535, 0.07179126, 0.04137834, 
    0.07164969, 0.04448365, 0.07982045, 0.005773919, -8.027887e-07, 
    5.864507e-05, 0.04907536, 0.1425036, 0.0631614, 0.05131766, 0.007727708,
  0.0007110864, 0.036148, 0.2037362, 0.05793827, 0.01923333, 0.03184226, 
    0.03034489, 0.05249256, 0.04991584, 0.05006434, 0.06798631, 0.04953918, 
    0.08185601, 0.02902071, 0.05459016, 0.0415258, 0.05351571, 0.05500514, 
    0.03235967, 0.01118776, 2.614343e-05, 0.001362149, 0.002105346, 
    0.1535182, 0.1637836, 0.1231156, 0.02865599, 0.004690989, 0.0008538367,
  0.00207493, 0.01922652, 0.02590078, 0.0432629, 0.01557027, 0.02457656, 
    0.02319637, 0.01645685, 0.08171837, 0.2124183, 0.06484693, 0.01674284, 
    0.03385352, 0.02294078, 0.02547425, 0.03349173, 0.01908983, 0.00990501, 
    0.01251241, 0.02273442, 0.02151156, 0.01777787, 0.07461123, 0.1161884, 
    0.1030352, 0.09270824, 0.02911634, 0.01480366, 0.003411956,
  4.529496e-05, 1.322697e-06, -4.652073e-05, 0.1304166, 0.0003144847, 
    0.003520088, 0.009371819, 0.03905307, 0.01209824, 0.03133768, 0.09764471, 
    0.05826848, 0.05746509, 0.05670988, 0.01836207, 0.02725331, 0.02767548, 
    0.03666957, 0.05743314, 0.05583289, 0.03653434, 0.01571268, 0.03462128, 
    0.01537531, 0.01764679, 0.0002592067, 8.951362e-07, 1.915902e-06, 
    0.001956515,
  1.10883e-06, 2.06284e-07, -3.18697e-06, 0.002979073, 6.550783e-06, 
    1.658801e-07, 0.000245811, 0.001381157, 0.02125119, 0.01303567, 
    0.003517163, 0.02247193, 0.02651923, 0.01426035, 0.01074964, 0.01778711, 
    0.03119285, 0.003944071, 0.01967933, 0.01131241, 0.000165487, 0.07118499, 
    0.01957033, 0.03286928, 0.01554889, 0.03272761, 0.003314861, 
    -8.781654e-06, 9.291105e-07,
  0.005596913, 0.003295077, 0.04822041, 0.01432835, 0.0370174, 0.001686575, 
    0.00155753, 0.09118998, 0.1372789, 0.1922732, 0.1478551, 0.1258108, 
    0.1314077, 0.07788733, 0.0979448, 0.08180705, 0.07415612, 0.09594123, 
    0.03964248, 0.01619691, 0.03594957, 0.07146294, 0.08919666, 0.06951299, 
    0.0788113, 0.07503206, 0.03813647, 0.004617812, -3.069814e-05,
  0.01248273, 0.04578933, 0.09823854, 0.1753488, 0.05534029, 0.0258271, 
    0.1977012, 0.0129807, 0.008149672, 0.05665209, 0.1160878, 0.09682813, 
    0.1536703, 0.1880025, 0.1866064, 0.1735596, 0.1632855, 0.1990357, 
    0.1495016, 0.1576664, 0.1600179, 0.1547823, 0.1984355, 0.1586733, 
    0.2176459, 0.2527956, 0.08620765, 0.05377595, 0.02306884,
  0.1144878, 0.2068944, 0.1990277, 0.1823699, 0.1974264, 0.1897902, 
    0.1829203, 0.1637218, 0.121803, 0.1211, 0.09935605, 0.1436069, 0.1045073, 
    0.2937934, 0.3221534, 0.2469337, 0.2396846, 0.2646229, 0.2011388, 
    0.187671, 0.135425, 0.1390379, 0.1818705, 0.209157, 0.1728215, 0.2485225, 
    0.248542, 0.1617704, 0.129059,
  0.2586623, 0.2397527, 0.1952046, 0.3216098, 0.3941401, 0.2875745, 
    0.2693039, 0.2499392, 0.2383959, 0.2942915, 0.2246683, 0.1241326, 
    0.2860542, 0.3276581, 0.3299965, 0.2038363, 0.1899166, 0.3027764, 
    0.3063779, 0.201103, 0.08551706, 0.1935214, 0.1954572, 0.3220464, 
    0.2222869, 0.2541671, 0.246954, 0.3134962, 0.2817814,
  0.2772883, 0.2449681, 0.3232665, 0.2846921, 0.3172002, 0.2494978, 
    0.2644059, 0.3535419, 0.3350168, 0.2824063, 0.2162309, 0.1887936, 
    0.2022457, 0.1535552, 0.1211711, 0.1653593, 0.1022409, 0.1295139, 
    0.09492444, 0.1570665, 0.2163883, 0.1129211, 0.1831661, 0.08583139, 
    0.221958, 0.3815304, 0.2392361, 0.2628781, 0.2074175,
  0.1441181, 0.1748134, 0.1763803, 0.1910951, 0.1858804, 0.1854561, 
    0.2071081, 0.2864564, 0.3037063, 0.2516683, 0.2102473, 0.198484, 
    0.1738876, 0.1608437, 0.1941895, 0.2040491, 0.2189437, 0.156523, 
    0.1616743, 0.1390931, 0.1405593, 0.1675435, 0.1329477, 0.06059342, 
    0.1066181, 0.1553321, 0.1694057, 0.1563757, 0.1867481,
  0.2000019, 0.20188, 0.2037581, 0.2056362, 0.2075144, 0.2093925, 0.2112706, 
    0.2572009, 0.269198, 0.2811951, 0.2931922, 0.3051893, 0.3171864, 
    0.3291835, 0.3313928, 0.3294345, 0.3274763, 0.325518, 0.3235597, 
    0.3216014, 0.3196431, 0.265076, 0.2531591, 0.2412421, 0.2293252, 
    0.2174083, 0.2054913, 0.1935744, 0.1984994,
  0.2253414, 0.2428953, 0.1113357, 0.05452216, 0.09104379, 0.1024737, 
    0.06248859, 0.05119386, 0.0699855, 0.1083362, 0.1717209, 0.2002429, 
    0.2877709, 0.2567691, 0.2286581, 0.1792467, 0.278313, 0.331609, 
    0.2900768, 0.2703149, 0.3681375, 0.3808447, 0.2614724, 0.2235723, 
    0.2358243, 0.221923, 0.3498942, 0.3561243, 0.2589397,
  0.2638223, 0.2511913, 0.2940743, 0.4084949, 0.280591, 0.149875, 0.2442815, 
    0.2711768, 0.2627771, 0.2768414, 0.3363611, 0.1829238, 0.2067209, 
    0.3968654, 0.3157544, 0.3198389, 0.3114324, 0.2818738, 0.2969167, 
    0.2637846, 0.2874193, 0.208765, 0.2553553, 0.3614555, 0.373989, 
    0.2994866, 0.290596, 0.2904428, 0.2726154,
  0.2744705, 0.3195738, 0.3098192, 0.3639212, 0.2766638, 0.2865124, 
    0.3591905, 0.3579031, 0.3657864, 0.3289424, 0.2950546, 0.3110721, 
    0.3180577, 0.2669723, 0.2715719, 0.2630975, 0.2863111, 0.272713, 
    0.352717, 0.3490021, 0.2917747, 0.3007022, 0.3088194, 0.2989061, 
    0.2853897, 0.2642612, 0.2414912, 0.2603483, 0.3063408,
  0.2170043, 0.2630896, 0.232554, 0.2450611, 0.2111601, 0.1787754, 0.1850189, 
    0.2091604, 0.2079951, 0.2286575, 0.2805983, 0.2409716, 0.2292196, 
    0.1822279, 0.1138384, 0.1559187, 0.2074562, 0.2583589, 0.2391668, 
    0.2392552, 0.1842064, 0.1905083, 0.2499776, 0.15806, 0.08208758, 
    0.1338769, 0.1971437, 0.1858967, 0.1840351,
  0.1084254, 0.1186604, 0.06269035, 0.1054683, 0.105732, 0.06899437, 
    0.08301574, 0.08395682, 0.09368651, 0.1012109, 0.1075532, 0.0928911, 
    0.09323488, 0.1571141, 0.118209, 0.08477653, 0.1729025, 0.1819541, 
    0.1051634, 0.09927496, 0.09224866, 0.1398872, 0.09661502, 0.03484755, 
    0.02317155, 0.08976516, 0.09119481, 0.08499189, 0.1191746,
  0.02007318, 0.005598813, 0.05321087, 0.02991175, 0.06848004, 0.09575501, 
    0.09747683, 0.03987848, 0.0133935, 0.008455355, 0.01526415, 0.001572123, 
    0.084594, 0.09982488, 0.06603049, 0.07247191, 0.1201003, 0.08891083, 
    0.09112717, 0.09717789, 0.06090026, 0.09462777, 0.03021341, 2.923301e-05, 
    0.04088519, 0.05316588, 0.08433379, 0.04591491, 0.03678264,
  0.005346361, 0.03524693, 0.06576378, 0.03223893, 0.1175365, 0.02786146, 
    0.07316484, 0.06366096, 0.01304728, 0.004566351, 0.02249636, 0.03321222, 
    0.05936336, 0.05633248, 0.08028746, 0.09626795, 0.06925143, 0.03623239, 
    0.06758788, 0.04318163, 0.0950359, 0.03524485, -5.927621e-06, 
    0.000124743, 0.05943293, 0.1410738, 0.04835925, 0.06437576, 0.0273064,
  0.001159345, 0.0219314, 0.1849107, 0.05730161, 0.02034831, 0.02755681, 
    0.03122506, 0.0499735, 0.04173738, 0.04880976, 0.07212944, 0.04890542, 
    0.08133768, 0.0266115, 0.04356173, 0.03297919, 0.04729847, 0.0482125, 
    0.03260811, 0.01884389, 0.007428586, 0.002973054, 0.005804144, 0.1441652, 
    0.1449238, 0.1113735, 0.03810634, 0.007005027, 0.003434062,
  0.001775602, 0.01435597, 0.02564804, 0.03096214, 0.01867829, 0.02645087, 
    0.02357079, 0.01789519, 0.08752918, 0.2153323, 0.05800668, 0.01738965, 
    0.03150414, 0.02226487, 0.02428651, 0.03054158, 0.02392795, 0.01379085, 
    0.0189296, 0.02290007, 0.02583482, 0.02406106, 0.06654435, 0.09500557, 
    0.1023027, 0.08309354, 0.02850478, 0.01641487, 0.003663605,
  2.686566e-05, 4.552147e-07, -1.697163e-05, 0.06410398, 0.00165136, 
    0.003912648, 0.009887982, 0.03037529, 0.009780907, 0.03421855, 
    0.09382765, 0.05877209, 0.05455369, 0.04954365, 0.02231798, 0.02766476, 
    0.02928533, 0.04070212, 0.07204855, 0.06108142, 0.03501796, 0.01634126, 
    0.04403508, 0.01815349, 0.01924061, 0.000642115, 4.344589e-07, 
    6.602564e-07, 0.0007032299,
  7.095125e-07, 7.368465e-08, -1.66736e-06, 0.0001477778, 2.539575e-06, 
    3.540684e-07, 3.489206e-05, 0.001800984, 0.009601126, 0.01347715, 
    0.00587513, 0.03003675, 0.03366588, 0.02107121, 0.01783699, 0.02531637, 
    0.03064819, 0.01517897, 0.02373079, 0.01068815, 1.737018e-05, 0.09100085, 
    0.01997229, 0.03357119, 0.02955177, 0.03541993, 0.007665281, -1.227e-05, 
    8.149322e-07,
  0.00251627, 0.007604176, 0.0476933, 0.01293661, 0.02402697, 0.0002105619, 
    -0.001332491, 0.07719232, 0.114289, 0.1735779, 0.1432389, 0.1312104, 
    0.131447, 0.08491072, 0.1114318, 0.09574311, 0.1041207, 0.09963933, 
    0.05198297, 0.02375824, 0.03011758, 0.0851451, 0.08677241, 0.08460473, 
    0.08321768, 0.08242495, 0.0432818, 0.003518174, 0.0001139018,
  0.009531068, 0.04347783, 0.09549073, 0.189909, 0.05060448, 0.0258975, 
    0.1839563, 0.01281583, 0.009368427, 0.06150651, 0.107089, 0.113282, 
    0.1841862, 0.2289093, 0.2063027, 0.1915703, 0.1810356, 0.225464, 
    0.169789, 0.1623345, 0.1554423, 0.1703856, 0.1925181, 0.1390455, 
    0.2657264, 0.2675433, 0.1108106, 0.06117243, 0.02448367,
  0.1339586, 0.2060883, 0.2045937, 0.1737519, 0.1608059, 0.1459767, 
    0.1421854, 0.1620498, 0.1212583, 0.09517795, 0.07742282, 0.1300557, 
    0.1005868, 0.346518, 0.3166028, 0.2330374, 0.2352815, 0.2632195, 
    0.2091451, 0.1815081, 0.1237038, 0.1233098, 0.1654097, 0.2110185, 
    0.1637699, 0.2814733, 0.2861351, 0.1749527, 0.1667276,
  0.2667701, 0.2306535, 0.2152377, 0.2866139, 0.334906, 0.2569439, 0.2733617, 
    0.2864227, 0.2435265, 0.3010795, 0.2383274, 0.1319487, 0.2923838, 
    0.3136902, 0.3421417, 0.1975931, 0.1640412, 0.3125356, 0.2979877, 
    0.2075837, 0.08415404, 0.1887171, 0.1978719, 0.3141509, 0.2391143, 
    0.2548966, 0.2853588, 0.322292, 0.3134225,
  0.2793517, 0.2582515, 0.302446, 0.304192, 0.2921392, 0.2559985, 0.2672613, 
    0.3659365, 0.323927, 0.3381184, 0.2488022, 0.1918912, 0.2258217, 
    0.1404207, 0.1404253, 0.1632212, 0.1077728, 0.1136452, 0.08239439, 
    0.1614506, 0.2037487, 0.1213275, 0.1838165, 0.09996325, 0.2116128, 
    0.4335575, 0.2837645, 0.2460527, 0.219282,
  0.1510258, 0.1555861, 0.1888861, 0.1968025, 0.1922056, 0.1847841, 
    0.2252681, 0.3067742, 0.3010217, 0.2574507, 0.220586, 0.1790031, 
    0.1631008, 0.1976684, 0.1964483, 0.195707, 0.213557, 0.1431067, 
    0.1626889, 0.1402866, 0.1397669, 0.1655691, 0.1337489, 0.0618888, 
    0.09408788, 0.1404563, 0.1712041, 0.1549706, 0.2024965,
  0.2324426, 0.2343893, 0.236336, 0.2382828, 0.2402295, 0.2421763, 0.244123, 
    0.2827043, 0.2946323, 0.3065604, 0.3184884, 0.3304164, 0.3423445, 
    0.3542725, 0.3578868, 0.3550076, 0.3521284, 0.3492492, 0.3463701, 
    0.3434909, 0.3406117, 0.302075, 0.2910794, 0.2800838, 0.2690883, 
    0.2580927, 0.2470971, 0.2361015, 0.2308852,
  0.2294463, 0.2775198, 0.1896412, 0.0898283, 0.1084285, 0.1047187, 
    0.06066648, 0.05522065, 0.1038611, 0.1298078, 0.2045585, 0.2120142, 
    0.3167907, 0.2145008, 0.205231, 0.2073331, 0.2748976, 0.3146324, 
    0.2883411, 0.2820736, 0.3856504, 0.3769485, 0.2762435, 0.2288222, 
    0.2566361, 0.2567551, 0.3526776, 0.366481, 0.2735286,
  0.2829266, 0.2942808, 0.3132448, 0.4114447, 0.2765585, 0.1561728, 
    0.2705556, 0.2923971, 0.2712286, 0.2832216, 0.3154923, 0.1748339, 
    0.2156649, 0.4207758, 0.4017739, 0.3799851, 0.3519888, 0.3423343, 
    0.4305845, 0.3118337, 0.3171329, 0.2189808, 0.2767243, 0.3883182, 
    0.3652894, 0.3514467, 0.3040193, 0.3035923, 0.3520226,
  0.3057439, 0.3181703, 0.285021, 0.3767179, 0.2923445, 0.301364, 0.3833643, 
    0.4257893, 0.4078791, 0.3883002, 0.299693, 0.3210722, 0.3688623, 
    0.306304, 0.313279, 0.3096843, 0.3127968, 0.3002135, 0.4147065, 
    0.3870305, 0.3078004, 0.3505644, 0.3452612, 0.3460006, 0.3085283, 
    0.2840452, 0.2838568, 0.284911, 0.3139603,
  0.259629, 0.2703268, 0.2541012, 0.2772223, 0.2396902, 0.2021538, 0.2085299, 
    0.2704172, 0.2295447, 0.2565365, 0.2969199, 0.263146, 0.2391449, 
    0.2079027, 0.1101627, 0.1793092, 0.2277324, 0.3071411, 0.2778254, 
    0.2629784, 0.2074326, 0.2185716, 0.2615727, 0.1715026, 0.07320981, 
    0.1429867, 0.2233087, 0.2235188, 0.2102037,
  0.148048, 0.1368084, 0.1125255, 0.1211893, 0.1240588, 0.1047416, 0.115867, 
    0.1225789, 0.1269346, 0.1156086, 0.1414416, 0.101022, 0.08872601, 
    0.1444785, 0.1328613, 0.1102265, 0.2070888, 0.2166123, 0.1187663, 
    0.1289087, 0.1152729, 0.1723148, 0.1273567, 0.04021202, 0.03592724, 
    0.107434, 0.1188335, 0.1033942, 0.1326687,
  0.04142145, 0.01284698, 0.04968595, 0.04554715, 0.07897326, 0.09764679, 
    0.1176761, 0.07274476, 0.03243204, 0.01061436, 0.01627024, 0.0001700928, 
    0.06742923, 0.1030863, 0.06915511, 0.08704223, 0.1298568, 0.1059341, 
    0.09646218, 0.1018222, 0.06191369, 0.1170883, 0.045579, -6.884297e-06, 
    0.03602154, 0.05191358, 0.07851258, 0.05060545, 0.06971206,
  0.01335611, 0.0267079, 0.08961299, 0.03242842, 0.1131904, 0.02690994, 
    0.07038227, 0.06911238, 0.01803925, 0.007006733, 0.01447643, 0.02774882, 
    0.05887909, 0.05005033, 0.06311242, 0.08241084, 0.06514403, 0.02951224, 
    0.063345, 0.03485443, 0.06360506, 0.1116686, 0.004410961, 0.000282714, 
    0.07473963, 0.1509759, 0.0353288, 0.04661215, 0.06617805,
  0.003542316, 0.01800523, 0.1572251, 0.06321512, 0.0198602, 0.02401147, 
    0.03102397, 0.0430728, 0.03438443, 0.04553972, 0.07382803, 0.04625798, 
    0.07098287, 0.02490022, 0.03368293, 0.02736656, 0.03982953, 0.03207402, 
    0.03169499, 0.01936779, 0.02020545, 0.009159737, 0.02332375, 0.1260625, 
    0.1356743, 0.09993234, 0.04289504, 0.01706697, 0.01105218,
  0.002172399, 0.01546132, 0.02440415, 0.02400381, 0.02040918, 0.02924837, 
    0.02108906, 0.02021341, 0.097086, 0.2248567, 0.04774919, 0.01794593, 
    0.02925359, 0.02242643, 0.02165325, 0.03051579, 0.0227662, 0.01755108, 
    0.02522455, 0.02181888, 0.02097362, 0.02377721, 0.05562083, 0.07697553, 
    0.1001383, 0.06778665, 0.02596686, 0.01790883, 0.005117574,
  7.114569e-06, 1.420508e-07, -6.13088e-06, 0.02529521, 0.009451122, 
    0.004764487, 0.01335002, 0.02350016, 0.01065131, 0.03889341, 0.09099984, 
    0.05150209, 0.04496702, 0.04669075, 0.02206159, 0.02612183, 0.03255138, 
    0.0489675, 0.09828286, 0.06416363, 0.03019317, 0.01631237, 0.04816812, 
    0.01648295, 0.02147394, 0.003144335, 6.689611e-06, 9.996463e-08, 
    0.0002717293,
  3.495759e-07, 1.702817e-08, -5.821213e-07, 0.003125675, 6.978279e-07, 
    -8.967322e-07, 8.173271e-06, 0.001021761, 0.008702742, 0.02690004, 
    0.02336493, 0.04840933, 0.03876915, 0.03275612, 0.04423238, 0.03672275, 
    0.0446755, 0.03810102, 0.04161112, 0.0131808, 8.4257e-06, 0.1154189, 
    0.02189372, 0.02844043, 0.03660852, 0.05331902, 0.02673208, 
    -1.156715e-05, 7.242187e-07,
  0.0001235752, 0.009144854, 0.03778769, 0.01020972, 0.0176692, 
    -8.097908e-05, -0.002364496, 0.05876374, 0.1023315, 0.1566322, 0.1617369, 
    0.1620766, 0.1642853, 0.1356645, 0.1475151, 0.1643715, 0.1488353, 
    0.1133955, 0.08082409, 0.04131564, 0.02685009, 0.107631, 0.08618015, 
    0.1019117, 0.1059027, 0.1016764, 0.04926313, 0.03552182, -4.01443e-05,
  0.003999981, 0.04464324, 0.08644263, 0.1938383, 0.05292796, 0.01636719, 
    0.1688407, 0.01331143, 0.00970979, 0.07481102, 0.1003939, 0.1504694, 
    0.2344876, 0.2816853, 0.2271697, 0.2172166, 0.2158296, 0.2435649, 
    0.2057849, 0.1633755, 0.1481425, 0.1786717, 0.1877996, 0.1388036, 
    0.347136, 0.2748926, 0.1230897, 0.09076259, 0.02936915,
  0.1164437, 0.243729, 0.230497, 0.2181105, 0.1594222, 0.1535601, 0.1332904, 
    0.1628541, 0.1130781, 0.08533796, 0.05907921, 0.1186763, 0.1202395, 
    0.3976201, 0.3355694, 0.2637203, 0.2741178, 0.287686, 0.2142268, 
    0.1779721, 0.1366492, 0.1374557, 0.1646969, 0.2209137, 0.1908262, 
    0.324751, 0.3112692, 0.2023237, 0.1850682,
  0.2830278, 0.2258387, 0.2461616, 0.3248792, 0.3992448, 0.2859893, 
    0.2458083, 0.2859921, 0.2511446, 0.314099, 0.257515, 0.1408468, 0.294315, 
    0.332732, 0.3735626, 0.186176, 0.1488063, 0.3121059, 0.2973891, 
    0.2065235, 0.1051686, 0.1601219, 0.2265325, 0.2875379, 0.2561452, 
    0.2490788, 0.3245293, 0.3228246, 0.3283935,
  0.2971815, 0.3117645, 0.3353991, 0.3587441, 0.3249859, 0.2780783, 
    0.2943198, 0.3673137, 0.2857407, 0.3154626, 0.2620202, 0.2025825, 
    0.238029, 0.1455865, 0.1597522, 0.1451906, 0.1519394, 0.1189574, 
    0.08007562, 0.1740606, 0.2006975, 0.1226333, 0.1904516, 0.1024621, 
    0.2080936, 0.4371046, 0.3271663, 0.2336362, 0.2507339,
  0.1624674, 0.1535785, 0.2079889, 0.2192251, 0.1890998, 0.2492143, 
    0.2524235, 0.3707324, 0.3307586, 0.2924914, 0.2229491, 0.1753865, 
    0.1607099, 0.2080389, 0.1939794, 0.2219512, 0.2197298, 0.1571221, 
    0.167322, 0.1687249, 0.1634947, 0.1719848, 0.1456445, 0.06476369, 
    0.09004084, 0.1230225, 0.1713136, 0.1677261, 0.2433811,
  0.2675211, 0.2703813, 0.2732416, 0.2761018, 0.278962, 0.2818222, 0.2846825, 
    0.2968102, 0.3076555, 0.3185008, 0.3293461, 0.3401914, 0.3510366, 
    0.3618819, 0.3860768, 0.3824309, 0.378785, 0.3751391, 0.3714932, 
    0.3678473, 0.3642014, 0.3274426, 0.3173831, 0.3073234, 0.2972638, 
    0.2872042, 0.2771446, 0.267085, 0.2652329,
  0.224357, 0.2965442, 0.2714746, 0.1267297, 0.1251268, 0.1324668, 
    0.09139448, 0.08572219, 0.1308293, 0.1369527, 0.2196556, 0.2433693, 
    0.3397485, 0.1722695, 0.1626475, 0.2058644, 0.2820445, 0.2965263, 
    0.2897637, 0.2617719, 0.400244, 0.381173, 0.2886018, 0.2624985, 
    0.2615137, 0.2611414, 0.3715408, 0.3338313, 0.2737163,
  0.2893959, 0.2717431, 0.3596904, 0.3800995, 0.2723253, 0.1631749, 
    0.2739444, 0.3134856, 0.2742844, 0.2836862, 0.2837363, 0.1689729, 
    0.2179495, 0.4093133, 0.5329515, 0.447139, 0.4689461, 0.4792512, 
    0.437838, 0.3562902, 0.3264394, 0.234177, 0.2724621, 0.3798572, 
    0.3941178, 0.4558188, 0.3473986, 0.4585366, 0.4364181,
  0.3699309, 0.3698799, 0.3393915, 0.3550729, 0.3143069, 0.3384578, 
    0.4307381, 0.4746526, 0.4990864, 0.3788105, 0.3435718, 0.3678281, 
    0.420296, 0.3296059, 0.3445285, 0.3512816, 0.3643788, 0.3876561, 
    0.4539405, 0.4016274, 0.3280036, 0.3679168, 0.3545888, 0.3530825, 
    0.367157, 0.3660647, 0.3691605, 0.3485152, 0.3283762,
  0.3221119, 0.2956651, 0.2859467, 0.3022329, 0.2680391, 0.2300662, 
    0.2160144, 0.3121733, 0.2587635, 0.2868238, 0.3513746, 0.2981514, 
    0.3076589, 0.2368905, 0.1374389, 0.2314755, 0.2894889, 0.3375514, 
    0.284954, 0.2922083, 0.2598862, 0.2342559, 0.2958658, 0.1720829, 
    0.0676226, 0.1626136, 0.2486172, 0.2615486, 0.2691286,
  0.1927505, 0.1678667, 0.1655756, 0.1545533, 0.1758783, 0.1470105, 0.132544, 
    0.1706552, 0.1750478, 0.1497959, 0.2133721, 0.1034983, 0.08573726, 
    0.1681314, 0.1669094, 0.1491478, 0.2619562, 0.2726508, 0.1592807, 
    0.1671005, 0.1763475, 0.2131779, 0.1723345, 0.0459988, 0.03569175, 
    0.1464074, 0.1411479, 0.140604, 0.1815515,
  0.08658179, 0.02076549, 0.04554042, 0.0791901, 0.09054788, 0.1040264, 
    0.136317, 0.1018205, 0.08794643, 0.03220592, 0.01550244, 0.0005311847, 
    0.0536177, 0.1089804, 0.09171624, 0.1056867, 0.1397941, 0.1273, 
    0.1177157, 0.1031764, 0.08279498, 0.1446276, 0.1008137, 2.053814e-05, 
    0.03661552, 0.06740446, 0.08465841, 0.06032481, 0.07912643,
  0.04982434, 0.02142923, 0.07950203, 0.04475912, 0.1027534, 0.02883146, 
    0.06769659, 0.07235681, 0.03980575, 0.006372335, 0.00950848, 0.02403507, 
    0.06258637, 0.04716927, 0.0541813, 0.07188446, 0.06973637, 0.02765842, 
    0.0624208, 0.03608343, 0.0502457, 0.1452219, 0.06634381, 0.0005352162, 
    0.09996716, 0.1825413, 0.04171747, 0.04125829, 0.08032244,
  0.01912499, 0.02605538, 0.1286394, 0.07515616, 0.0220493, 0.02503073, 
    0.03326964, 0.03988315, 0.03265459, 0.04352726, 0.06867921, 0.04064883, 
    0.06483963, 0.02648687, 0.02831314, 0.02637442, 0.03447554, 0.03057087, 
    0.03242594, 0.02269215, 0.01789578, 0.02315599, 0.04413453, 0.1200094, 
    0.1256773, 0.09004122, 0.05299092, 0.03679413, 0.04550082,
  0.00395163, 0.01838449, 0.02232391, 0.01683445, 0.02478274, 0.03312337, 
    0.02282398, 0.02501163, 0.1065431, 0.2074211, 0.04170731, 0.02079638, 
    0.02870543, 0.0251525, 0.02130953, 0.02991031, 0.0226005, 0.02016654, 
    0.02313754, 0.01955843, 0.01795882, 0.0252572, 0.04508262, 0.06190028, 
    0.1051025, 0.05530021, 0.02469554, 0.01984686, 0.01338142,
  1.023341e-06, 5.399266e-08, -1.920485e-06, 0.009251447, 0.01465461, 
    0.01320668, 0.01561732, 0.02039301, 0.009622667, 0.0410682, 0.0919098, 
    0.04628336, 0.03798592, 0.04200191, 0.02783728, 0.03417683, 0.03450922, 
    0.05720299, 0.1174855, 0.06767695, 0.02916447, 0.01928731, 0.0471941, 
    0.01904316, 0.03310954, 0.02130641, 0.0006586007, 9.365584e-08, 
    0.0001210437,
  1.340646e-07, 1.366166e-08, -2.08594e-08, 0.0007279245, 5.892278e-08, 
    0.0002087031, -6.696368e-06, 0.001004533, 0.009955687, 0.04569255, 
    0.06572411, 0.08647034, 0.06291751, 0.0490739, 0.08080478, 0.07344652, 
    0.07248011, 0.06221351, 0.06718335, 0.05713412, 3.045055e-06, 0.1473857, 
    0.04048087, 0.04062037, 0.07387656, 0.07185258, 0.07464131, 5.151284e-05, 
    4.727084e-07,
  5.594035e-06, 0.008753156, 0.03519544, 0.008553604, 0.01040515, 
    -3.945909e-05, -0.002551371, 0.04209141, 0.0939514, 0.147379, 0.1847276, 
    0.1739591, 0.1899464, 0.1543788, 0.2570212, 0.2165457, 0.1626882, 
    0.1943752, 0.1521356, 0.05472591, 0.03135706, 0.1360209, 0.1068181, 
    0.1642094, 0.1661158, 0.1235912, 0.05148865, 0.0822766, -0.0001257976,
  0.0009073663, 0.02665763, 0.08026364, 0.2073993, 0.06918925, 0.01172323, 
    0.1488065, 0.008943072, 0.008537185, 0.05287065, 0.09371078, 0.1425618, 
    0.2701968, 0.2661563, 0.206973, 0.2505752, 0.2773112, 0.2544441, 
    0.2513975, 0.16711, 0.1296651, 0.1900204, 0.2001778, 0.1572962, 
    0.4077749, 0.3032136, 0.1434008, 0.1273506, 0.03646298,
  0.1312541, 0.2710465, 0.2165999, 0.2104038, 0.1273188, 0.1785501, 
    0.1419287, 0.176585, 0.1074519, 0.08249224, 0.03606043, 0.1097537, 
    0.1638113, 0.411151, 0.3952269, 0.2813371, 0.3333571, 0.3141413, 
    0.2696685, 0.1842698, 0.1366895, 0.1149104, 0.1545838, 0.247517, 
    0.2296984, 0.3991639, 0.330312, 0.2530764, 0.1874518,
  0.2942938, 0.2236867, 0.2607684, 0.3580017, 0.4535069, 0.2740264, 
    0.2788426, 0.2823342, 0.2721061, 0.3134483, 0.285494, 0.1468487, 
    0.2873966, 0.3343515, 0.454108, 0.2320217, 0.1618659, 0.3172509, 
    0.2924249, 0.1823294, 0.1242992, 0.1975856, 0.2358159, 0.2790265, 
    0.3745353, 0.2512754, 0.3051766, 0.2945068, 0.301343,
  0.3245998, 0.3321263, 0.3682236, 0.4622594, 0.3089935, 0.2824373, 0.323798, 
    0.3329451, 0.2864882, 0.2892503, 0.2823169, 0.2207049, 0.2311059, 
    0.1618165, 0.1676344, 0.1153015, 0.140573, 0.1373872, 0.07769839, 
    0.1992405, 0.2071905, 0.1572628, 0.2126499, 0.1101394, 0.1882601, 
    0.4280491, 0.3521439, 0.2233769, 0.3115734,
  0.1904605, 0.1892551, 0.2447063, 0.2221814, 0.2054779, 0.2509505, 
    0.2752822, 0.3677698, 0.3312365, 0.3021226, 0.2590573, 0.2099462, 
    0.1756855, 0.2051862, 0.2283188, 0.2144467, 0.2056701, 0.1628281, 
    0.1766305, 0.2082707, 0.1779481, 0.1850305, 0.1522491, 0.06363542, 
    0.08472946, 0.105095, 0.1719213, 0.1686498, 0.2482656,
  0.2964102, 0.3004968, 0.3045833, 0.3086698, 0.3127563, 0.3168429, 
    0.3209294, 0.3167044, 0.3258309, 0.3349574, 0.344084, 0.3532105, 
    0.362337, 0.3714635, 0.3968629, 0.3920889, 0.3873149, 0.3825409, 
    0.377767, 0.372993, 0.368219, 0.3262712, 0.3178321, 0.309393, 0.300954, 
    0.2925149, 0.2840759, 0.2756368, 0.293141,
  0.209944, 0.3116236, 0.3227966, 0.169838, 0.1562999, 0.1610828, 0.1263252, 
    0.1162412, 0.1318473, 0.1445539, 0.2355117, 0.2660734, 0.350721, 
    0.1460185, 0.1618047, 0.2033714, 0.2612609, 0.2689984, 0.2327075, 
    0.2723363, 0.4180977, 0.4211271, 0.2966377, 0.251686, 0.2880039, 
    0.291381, 0.3515104, 0.2672744, 0.2668513,
  0.2873913, 0.2655544, 0.3603023, 0.3390125, 0.2694826, 0.188358, 0.2243604, 
    0.3349116, 0.2766934, 0.2925535, 0.2791416, 0.1735306, 0.2257513, 
    0.3914332, 0.4397387, 0.4310564, 0.5073636, 0.47898, 0.4112293, 
    0.3831291, 0.3621423, 0.2891789, 0.2964363, 0.3940791, 0.4173257, 
    0.4870605, 0.5336239, 0.5239895, 0.4472522,
  0.4328558, 0.3885929, 0.3466248, 0.3661546, 0.3316943, 0.4279344, 
    0.4726017, 0.5053253, 0.5259348, 0.3849184, 0.362543, 0.3914319, 
    0.4426321, 0.3978431, 0.3622878, 0.367725, 0.424193, 0.4460333, 
    0.5000443, 0.39338, 0.3609765, 0.3779854, 0.3694512, 0.3930539, 
    0.4588359, 0.4853244, 0.4562359, 0.4658762, 0.3938427,
  0.3599926, 0.3296334, 0.3151261, 0.2897105, 0.2898273, 0.2618136, 
    0.2411483, 0.3457489, 0.3033722, 0.3067158, 0.3486423, 0.2803643, 
    0.3247754, 0.2920273, 0.1819237, 0.2338848, 0.3585184, 0.3413703, 
    0.3184335, 0.3074917, 0.3074732, 0.2705937, 0.3090115, 0.1732158, 
    0.0675939, 0.2057261, 0.2914759, 0.3166209, 0.347616,
  0.2196529, 0.2789329, 0.2192444, 0.2196179, 0.2262312, 0.2050891, 
    0.1885375, 0.2921585, 0.2856012, 0.2485693, 0.2393161, 0.1256127, 
    0.09072161, 0.237237, 0.1799062, 0.188514, 0.2792381, 0.2862574, 
    0.2001052, 0.1966953, 0.2189914, 0.2732091, 0.1872028, 0.06030539, 
    0.03277809, 0.1745383, 0.1919006, 0.1671609, 0.2072669,
  0.1522372, 0.03613669, 0.04334933, 0.1265977, 0.1263544, 0.1124138, 
    0.1415699, 0.1336467, 0.2014431, 0.04133562, 0.01824146, 0.0001138151, 
    0.03843337, 0.1163935, 0.08752549, 0.1217799, 0.1574681, 0.1528807, 
    0.1484962, 0.1298112, 0.07715628, 0.153802, 0.1624197, 8.504284e-05, 
    0.0329866, 0.0815894, 0.08747806, 0.07042991, 0.08664288,
  0.1516193, 0.01544433, 0.07302082, 0.05853309, 0.09996411, 0.0381393, 
    0.07349669, 0.08195779, 0.09426403, 0.01191561, 0.005483305, 0.01857819, 
    0.07584191, 0.07200579, 0.06377311, 0.08745763, 0.06565131, 0.03290557, 
    0.07709923, 0.0473198, 0.05763385, 0.1202602, 0.2566298, 0.0004927785, 
    0.08700652, 0.177586, 0.05169804, 0.04914569, 0.08905934,
  0.06886997, 0.03718753, 0.09685756, 0.07517814, 0.03096417, 0.03132391, 
    0.04176071, 0.04318047, 0.03734034, 0.0420859, 0.07172409, 0.04145159, 
    0.06701158, 0.03349766, 0.02919838, 0.0378959, 0.03207535, 0.04422992, 
    0.05316623, 0.04369874, 0.03726591, 0.04651312, 0.07695258, 0.09936117, 
    0.09766982, 0.07408419, 0.07265526, 0.08882027, 0.09320264,
  0.008959045, 0.01668276, 0.01891019, 0.01210143, 0.04157482, 0.06293068, 
    0.04933856, 0.0390961, 0.1106866, 0.1707356, 0.03953168, 0.02579395, 
    0.032828, 0.03426596, 0.03771017, 0.03577765, 0.02368774, 0.02033085, 
    0.02585444, 0.02111137, 0.02046472, 0.02581745, 0.02551746, 0.04283581, 
    0.09163193, 0.05111134, 0.029137, 0.02622095, 0.01822119,
  -8.392837e-07, 3.270036e-08, -1.27429e-06, 0.003123912, 0.02933772, 
    0.08760011, 0.01475229, 0.03562259, 0.01126118, 0.0564627, 0.09957314, 
    0.05004797, 0.04211779, 0.04629901, 0.05333748, 0.04520056, 0.03911069, 
    0.06461401, 0.1227815, 0.07013973, 0.04471086, 0.03367995, 0.05364536, 
    0.02806471, 0.05985112, 0.1204982, 0.01366627, 1.01516e-07, 8.703186e-05,
  3.553927e-08, 7.181434e-09, -2.784431e-09, 0.0002725838, 7.245879e-09, 
    0.001164209, -5.995947e-06, 0.003321185, 0.01254473, 0.0711696, 
    0.1031452, 0.1049783, 0.08891962, 0.08315416, 0.07895449, 0.1087965, 
    0.1510301, 0.07098478, 0.2054781, 0.1105668, -9.376823e-06, 0.165415, 
    0.05434765, 0.04440295, 0.09256962, 0.08169854, 0.130078, 0.002382615, 
    2.027533e-07,
  -8.593444e-06, 0.008430769, 0.02731481, 0.01242535, 0.007355718, 
    -1.292146e-05, -0.002472871, 0.02832838, 0.09017912, 0.1575767, 
    0.1869372, 0.1745079, 0.1966307, 0.2049059, 0.2789541, 0.2675936, 
    0.2236099, 0.2478601, 0.2305783, 0.05585422, 0.02917648, 0.1689174, 
    0.1141098, 0.2155205, 0.1694658, 0.1407751, 0.08934022, 0.04813847, 
    -0.0003282583,
  -0.0003909215, 0.02587914, 0.06825428, 0.1913598, 0.05841549, 0.0119881, 
    0.1324876, 0.004183426, 0.007378646, 0.03553352, 0.09305173, 0.1387911, 
    0.2189006, 0.1938122, 0.1634561, 0.2632385, 0.2901614, 0.2942524, 
    0.2897338, 0.1611179, 0.1107174, 0.1994916, 0.2002099, 0.1778813, 
    0.3518633, 0.2957491, 0.1425198, 0.190677, 0.07177423,
  0.1339106, 0.3143429, 0.2207058, 0.2181239, 0.1695313, 0.1661891, 
    0.1692061, 0.1800585, 0.09153856, 0.06857932, 0.01893146, 0.107216, 
    0.2493192, 0.3826213, 0.2923065, 0.3018908, 0.319049, 0.3403374, 
    0.3248399, 0.1877437, 0.1240161, 0.09943866, 0.1514865, 0.2398712, 
    0.2258177, 0.4024178, 0.334186, 0.2719173, 0.1853182,
  0.2677729, 0.2126304, 0.2882811, 0.3942435, 0.5009396, 0.3061465, 
    0.2784875, 0.2615681, 0.2413146, 0.2953549, 0.2562271, 0.1402211, 
    0.2711279, 0.3140361, 0.5266562, 0.2636847, 0.2066835, 0.3102521, 
    0.283273, 0.1562499, 0.129598, 0.2099347, 0.2617623, 0.2835526, 
    0.5659955, 0.1766205, 0.1934199, 0.249627, 0.256224,
  0.3015167, 0.2593743, 0.3806188, 0.4454555, 0.2928094, 0.246199, 0.304101, 
    0.3491003, 0.3095885, 0.3005909, 0.3219754, 0.2380927, 0.2369523, 
    0.1706136, 0.2277597, 0.1571748, 0.1299808, 0.140413, 0.0910221, 
    0.2328212, 0.2331166, 0.1747466, 0.2328877, 0.1140106, 0.1829911, 
    0.4245384, 0.3608124, 0.2124711, 0.387242,
  0.193922, 0.2205289, 0.2558545, 0.2264809, 0.2439049, 0.2729374, 0.3149797, 
    0.3868907, 0.3490103, 0.3193538, 0.3062864, 0.2414469, 0.2332117, 
    0.2555005, 0.2572567, 0.2091876, 0.2266168, 0.1989322, 0.212562, 
    0.2544274, 0.2005764, 0.203533, 0.1567008, 0.06611606, 0.08958083, 
    0.1021938, 0.1711515, 0.1775856, 0.2450889,
  0.3274852, 0.3315607, 0.3356363, 0.3397118, 0.3437873, 0.3478629, 
    0.3519384, 0.3325649, 0.3407338, 0.3489026, 0.3570715, 0.3652404, 
    0.3734092, 0.3815781, 0.3980225, 0.3908198, 0.3836173, 0.3764146, 
    0.369212, 0.3620094, 0.3548068, 0.3235424, 0.3185006, 0.3134589, 
    0.3084171, 0.3033754, 0.2983336, 0.2932918, 0.3242248,
  0.2185262, 0.3240093, 0.3605029, 0.2020106, 0.1861425, 0.1751745, 
    0.1516692, 0.1535063, 0.1366937, 0.1478276, 0.2600345, 0.2834697, 
    0.3665535, 0.1065723, 0.1796844, 0.2014452, 0.2418533, 0.2564787, 
    0.1904191, 0.3003446, 0.4329477, 0.4403039, 0.3213841, 0.2146067, 
    0.2895019, 0.3303983, 0.345677, 0.2110744, 0.2792507,
  0.281405, 0.2274558, 0.3309342, 0.2599584, 0.2724403, 0.1994778, 0.182008, 
    0.3341646, 0.2998784, 0.2976424, 0.279425, 0.1812034, 0.228552, 
    0.3262493, 0.3407706, 0.4377907, 0.448272, 0.4651598, 0.3906794, 
    0.3977637, 0.4161972, 0.3269592, 0.3125719, 0.4016573, 0.4251747, 
    0.4788762, 0.5030468, 0.4509423, 0.349236,
  0.3491676, 0.3315663, 0.3004285, 0.3547704, 0.3335867, 0.4367431, 
    0.5084197, 0.4975923, 0.4886171, 0.3486108, 0.3153008, 0.3877845, 
    0.5286534, 0.4407175, 0.3652486, 0.3740821, 0.4486537, 0.4806486, 
    0.5047027, 0.3913328, 0.3880416, 0.4024226, 0.4350547, 0.4179538, 
    0.483202, 0.5098126, 0.4682868, 0.4813064, 0.4028169,
  0.3787853, 0.3568654, 0.3229872, 0.321016, 0.2920454, 0.3321736, 0.2998172, 
    0.3665673, 0.3217326, 0.3262721, 0.3497774, 0.2973771, 0.3011712, 
    0.3286293, 0.2080996, 0.2582296, 0.3498086, 0.3608229, 0.3010185, 
    0.3039693, 0.2534067, 0.270844, 0.2866134, 0.1908072, 0.05428061, 
    0.202043, 0.3248022, 0.3896578, 0.3829737,
  0.247521, 0.3072634, 0.1752287, 0.224723, 0.2573959, 0.2509665, 0.244872, 
    0.2924969, 0.3134776, 0.2558321, 0.2158556, 0.1465972, 0.1077305, 
    0.2184483, 0.20718, 0.1761161, 0.240111, 0.2503263, 0.188311, 0.1775176, 
    0.2041093, 0.2740363, 0.2119112, 0.07839947, 0.01518727, 0.1902405, 
    0.2106754, 0.2346129, 0.2486946,
  0.1815591, 0.1177859, 0.04621962, 0.1714372, 0.1302455, 0.1241776, 
    0.1395106, 0.1130573, 0.2163355, 0.06860061, 0.01697823, -1.456938e-05, 
    0.0298373, 0.08747309, 0.08544825, 0.09579564, 0.1572048, 0.1670762, 
    0.1182597, 0.1110477, 0.1201555, 0.1311128, 0.2853791, 0.0003243704, 
    0.03359757, 0.07880525, 0.1033584, 0.1007634, 0.1023612,
  0.2647289, 0.01647912, 0.05771809, 0.08893465, 0.09760292, 0.07707705, 
    0.08566395, 0.06122532, 0.1171899, 0.0309945, 0.002667923, 0.01219736, 
    0.08994333, 0.1144271, 0.05726773, 0.09852076, 0.0972813, 0.05299363, 
    0.07933614, 0.06471229, 0.07945183, 0.07414959, 0.3752844, 0.0006522418, 
    0.06896178, 0.1646703, 0.05021416, 0.1050624, 0.1025107,
  0.2563995, 0.07189298, 0.06220968, 0.05075945, 0.08189082, 0.0715082, 
    0.0457604, 0.0793347, 0.06150467, 0.1077929, 0.07247212, 0.114832, 
    0.09229581, 0.06875893, 0.07463052, 0.1121256, 0.08710283, 0.09628004, 
    0.08588761, 0.09965383, 0.1474778, 0.1452417, 0.1660182, 0.0731098, 
    0.06766731, 0.05147133, 0.09518944, 0.1123442, 0.1816254,
  0.06043904, 0.009796283, 0.01504579, 0.009724805, 0.1238927, 0.1633593, 
    0.1939684, 0.1195146, 0.07189822, 0.1340633, 0.0572893, 0.08404773, 
    0.09211659, 0.06521721, 0.06764296, 0.06311493, 0.0344397, 0.02417518, 
    0.0469021, 0.02924348, 0.02971376, 0.03292289, 0.01808387, 0.02598532, 
    0.06145663, 0.05860725, 0.04264206, 0.04378077, 0.03782579,
  -7.91269e-07, 2.574371e-08, -2.879526e-07, 0.001371352, 0.03930887, 
    0.2461935, 0.04967314, 0.1339954, 0.03079275, 0.1003098, 0.1049035, 
    0.06621459, 0.04484264, 0.04019514, 0.05571053, 0.04178537, 0.04722053, 
    0.0862246, 0.1201909, 0.08527771, 0.07050674, 0.04773323, 0.1200785, 
    0.04253798, 0.05212575, 0.1336831, 0.132432, -3.322922e-07, 8.878016e-05,
  1.757299e-08, 6.711463e-09, -5.850342e-10, 0.0001749032, 2.408717e-09, 
    0.01431362, -8.928976e-06, 0.006781464, 0.01245466, 0.1062551, 
    0.09601821, 0.1251423, 0.1160427, 0.0956399, 0.07022387, 0.0782813, 
    0.07088991, 0.05306382, 0.1785052, 0.1987171, -0.0002905884, 0.1822444, 
    0.05281964, 0.02564364, 0.04805876, 0.04730728, 0.1089477, 0.02824201, 
    6.340718e-08,
  8.632911e-07, 0.01650672, 0.02294494, 0.01356896, 0.004394282, 
    -2.635061e-06, -0.002192297, 0.01954507, 0.08107068, 0.1677906, 
    0.1861885, 0.1352742, 0.1789624, 0.182081, 0.2057312, 0.2348668, 
    0.1668511, 0.228258, 0.258041, 0.07783307, 0.0250872, 0.1877996, 
    0.1043336, 0.170161, 0.1305586, 0.1357318, 0.1904424, 0.1133864, 
    0.0004088723,
  -0.0009487511, 0.02750373, 0.05794303, 0.2066416, 0.0463131, 0.006682293, 
    0.1223472, 0.003015801, 0.007755879, 0.03353257, 0.09111479, 0.1038666, 
    0.1755179, 0.1557705, 0.1471402, 0.2223299, 0.2824259, 0.2659258, 
    0.2962243, 0.1606742, 0.1024958, 0.2283555, 0.189513, 0.1578957, 
    0.2619624, 0.2762131, 0.1778288, 0.303317, 0.1063603,
  0.2054271, 0.3144565, 0.2165241, 0.2094538, 0.1463357, 0.1763081, 
    0.1930674, 0.1864524, 0.07346888, 0.06422759, 0.01289508, 0.1050454, 
    0.259697, 0.2966795, 0.2274329, 0.2440122, 0.283602, 0.3667848, 
    0.3312833, 0.2165823, 0.1270969, 0.09676752, 0.1370867, 0.2176811, 
    0.1986853, 0.3274152, 0.3111845, 0.2370853, 0.2481503,
  0.2683241, 0.2139127, 0.2888471, 0.3981737, 0.4681846, 0.263358, 0.2908943, 
    0.2471185, 0.210311, 0.2478123, 0.2369309, 0.1341946, 0.2361576, 
    0.2899308, 0.5736114, 0.2479717, 0.2558813, 0.28369, 0.3147309, 
    0.1395485, 0.1540848, 0.192467, 0.2752644, 0.2732293, 0.5816432, 
    0.108097, 0.1367967, 0.2286391, 0.2376781,
  0.194903, 0.1858279, 0.3729806, 0.3572525, 0.3128739, 0.2577929, 0.292074, 
    0.3778888, 0.3096689, 0.3556629, 0.366253, 0.2683695, 0.2577949, 
    0.2120873, 0.2671367, 0.1548362, 0.1428773, 0.1667873, 0.1002668, 
    0.2749587, 0.2545225, 0.2198023, 0.2534692, 0.1179929, 0.1781326, 
    0.4298475, 0.3718642, 0.1820863, 0.3857968,
  0.189234, 0.2308747, 0.2746735, 0.2554157, 0.2604007, 0.3198635, 0.335346, 
    0.4054251, 0.4079714, 0.3574149, 0.3727209, 0.314642, 0.2911323, 
    0.3203984, 0.2665707, 0.2374169, 0.2818211, 0.286662, 0.2883584, 
    0.2716149, 0.2147268, 0.2096606, 0.1557127, 0.0690219, 0.09657305, 
    0.1070599, 0.1612486, 0.1865325, 0.2488261,
  0.3558976, 0.3596848, 0.3634721, 0.3672594, 0.3710466, 0.3748339, 
    0.3786211, 0.3616071, 0.3681314, 0.3746557, 0.3811799, 0.3877042, 
    0.3942285, 0.4007528, 0.4112437, 0.4035521, 0.3958606, 0.3881691, 
    0.3804775, 0.3727859, 0.3650944, 0.3315306, 0.3289106, 0.3262907, 
    0.3236707, 0.3210507, 0.3184307, 0.3158107, 0.3528678,
  0.2337757, 0.3656875, 0.3764592, 0.2289861, 0.2156318, 0.1813065, 
    0.1697707, 0.182408, 0.1479185, 0.1795532, 0.2810206, 0.3280384, 
    0.3700995, 0.07033571, 0.1472777, 0.220772, 0.2599724, 0.2428841, 
    0.1689464, 0.3003125, 0.5103142, 0.4573719, 0.3349897, 0.205017, 
    0.2539844, 0.3384259, 0.2588936, 0.1532079, 0.2842817,
  0.2373023, 0.1831007, 0.2890477, 0.1958254, 0.2511206, 0.1947011, 
    0.1325089, 0.330186, 0.3122256, 0.293404, 0.2705662, 0.1888211, 
    0.2161317, 0.228012, 0.2484611, 0.3696728, 0.424617, 0.3878906, 
    0.3560646, 0.4183123, 0.4485091, 0.3851063, 0.3411882, 0.4281865, 
    0.4068487, 0.4830621, 0.3859976, 0.3605876, 0.2521027,
  0.2963428, 0.2864463, 0.2643223, 0.3255534, 0.3323282, 0.3965859, 
    0.4550793, 0.4352943, 0.4489108, 0.296224, 0.2828521, 0.3653988, 
    0.537074, 0.4532685, 0.3585297, 0.3975317, 0.4328901, 0.4745919, 
    0.4711046, 0.40062, 0.3755429, 0.3874546, 0.4481447, 0.403992, 0.4654964, 
    0.4996148, 0.4792864, 0.4331486, 0.3708602,
  0.405878, 0.3887994, 0.3504685, 0.3209176, 0.3042068, 0.3363225, 0.3656231, 
    0.3786009, 0.328163, 0.3302958, 0.3374866, 0.3123569, 0.310992, 
    0.3120143, 0.1871933, 0.3204562, 0.3059676, 0.3508501, 0.2708823, 
    0.2854976, 0.2244359, 0.2385565, 0.2776244, 0.194899, 0.03014229, 
    0.1995903, 0.3424519, 0.3823293, 0.3989422,
  0.2980498, 0.2537839, 0.1237775, 0.2207368, 0.2473983, 0.2462024, 
    0.2893329, 0.2380922, 0.2535557, 0.1844833, 0.1606063, 0.1191796, 
    0.08309287, 0.2259467, 0.2182255, 0.1163673, 0.1899944, 0.2031451, 
    0.1730884, 0.1895723, 0.1838807, 0.2708346, 0.1891422, 0.1046745, 
    0.01467849, 0.1771965, 0.2035605, 0.2676746, 0.2372666,
  0.1320289, 0.156749, 0.03902753, 0.07188448, 0.09467078, 0.1245885, 
    0.07658086, 0.04260427, 0.1218396, 0.04314287, 0.02060521, 0.0002293494, 
    0.02351864, 0.0644035, 0.0720914, 0.05881842, 0.09656613, 0.1688545, 
    0.1150557, 0.07276678, 0.06769807, 0.06787708, 0.1474736, 0.005875408, 
    0.03936033, 0.04737242, 0.06346543, 0.0451366, 0.07171727,
  0.1692948, 0.02202959, 0.04374663, 0.04485692, 0.0783149, 0.06802015, 
    0.05891973, 0.04171579, 0.06971505, 0.03759081, 0.0009600828, 
    0.009237619, 0.06046788, 0.04899019, 0.03810016, 0.05944858, 0.06117965, 
    0.04315329, 0.05137262, 0.01651306, 0.02302893, 0.02376679, 0.1578475, 
    0.1079784, 0.05414965, 0.1622351, 0.01645409, 0.03467026, 0.05571619,
  0.2679867, 0.1359093, 0.03940729, 0.03888063, 0.0478936, 0.03961708, 
    0.02946348, 0.05840002, 0.08263849, 0.09942377, 0.04859348, 0.05069225, 
    0.04686122, 0.04479496, 0.03055776, 0.03218304, 0.03232209, 0.03166619, 
    0.02277562, 0.04632597, 0.06171367, 0.09563588, 0.14082, 0.05609057, 
    0.04659425, 0.03220012, 0.03836873, 0.03037296, 0.06894784,
  0.1207744, 0.004764657, 0.008539215, 0.01006572, 0.1037159, 0.05553695, 
    0.03468044, 0.01879889, 0.04395583, 0.106914, 0.07853343, 0.1835254, 
    0.04114938, 0.02871951, 0.02747316, 0.05423366, 0.06089225, 0.03874028, 
    0.05750805, 0.08354094, 0.1256996, 0.1499715, 0.02963219, 0.01422519, 
    0.03035582, 0.04234631, 0.03930281, 0.07230196, 0.154871,
  -2.744035e-07, 2.341712e-08, -1.303283e-07, 0.0002873799, 0.0364551, 
    0.05657493, 0.03006204, 0.05460544, 0.02625985, 0.07312618, 0.08986241, 
    0.05833494, 0.0212829, 0.01966362, 0.01446923, 0.01393028, 0.02837208, 
    0.05664119, 0.09404337, 0.06230894, 0.02888888, 0.01760012, 0.2635568, 
    0.08546282, 0.008599408, 0.03792258, 0.07516447, -7.482345e-05, 
    3.463655e-05,
  1.271461e-08, 6.203731e-09, -1.580279e-10, 0.0003278204, 1.466078e-09, 
    0.006684218, -9.562678e-06, 0.002648655, 0.008450322, 0.1619521, 
    0.1095762, 0.09459172, 0.06515472, 0.06071312, 0.04560107, 0.0248357, 
    0.03079559, 0.04581827, 0.09656952, 0.1136224, -5.297345e-06, 0.1681998, 
    0.01788579, 0.008939851, 0.01767825, 0.02811633, 0.06221006, 0.008331063, 
    4.151568e-08,
  -3.092387e-06, 0.01321005, 0.01852343, 0.01233032, 0.00391322, 
    -1.472302e-06, -0.001912915, 0.01526778, 0.06614487, 0.160215, 0.1790017, 
    0.1200454, 0.1722766, 0.1406173, 0.1754714, 0.1947323, 0.1266074, 
    0.1265389, 0.1725382, 0.05730074, 0.02227672, 0.1983903, 0.08828656, 
    0.1182125, 0.1104595, 0.1107975, 0.129811, 0.08954981, 0.001174835,
  -0.0007679136, 0.02692256, 0.0410243, 0.2004422, 0.03748837, 0.004822954, 
    0.105496, 0.0008052365, 0.007320966, 0.03457855, 0.09151088, 0.08852471, 
    0.1483092, 0.1264551, 0.1168246, 0.1810659, 0.253394, 0.2502702, 
    0.2563081, 0.1626144, 0.0949641, 0.2261249, 0.1702916, 0.1381367, 
    0.2065237, 0.2822908, 0.160561, 0.2689728, 0.09107439,
  0.2063264, 0.2829436, 0.1630206, 0.1490717, 0.1126739, 0.2238762, 
    0.1603353, 0.1692947, 0.05741981, 0.05392713, 0.00959442, 0.1065385, 
    0.2155168, 0.2316489, 0.1864634, 0.2128509, 0.2756072, 0.3345869, 
    0.2953274, 0.2395531, 0.1166807, 0.08743241, 0.1129682, 0.1903191, 
    0.1587764, 0.2503245, 0.2795645, 0.2480115, 0.266718,
  0.2559195, 0.2402347, 0.2956536, 0.4089506, 0.4731904, 0.2356064, 
    0.3091486, 0.2160247, 0.1616308, 0.1918281, 0.2022997, 0.1480602, 
    0.2177245, 0.2461327, 0.5635908, 0.2374679, 0.2198452, 0.2618384, 
    0.3270856, 0.140816, 0.1329387, 0.1571644, 0.2667949, 0.2495964, 
    0.4677213, 0.07023256, 0.1044234, 0.2154031, 0.2196681,
  0.1354616, 0.1287649, 0.3251175, 0.2759859, 0.3501003, 0.2810499, 
    0.3044405, 0.3827546, 0.2925196, 0.3735664, 0.4599688, 0.3201264, 
    0.3025668, 0.2437647, 0.2915727, 0.1917666, 0.1893133, 0.18341, 
    0.1499787, 0.3011949, 0.2940315, 0.2681672, 0.2698438, 0.1170768, 
    0.175974, 0.412383, 0.3733846, 0.1481841, 0.330509,
  0.1714968, 0.200406, 0.3343163, 0.3165575, 0.3145623, 0.4129736, 0.3997951, 
    0.4293789, 0.4264423, 0.3925322, 0.4149318, 0.3599086, 0.3417132, 
    0.3673219, 0.2984883, 0.2982084, 0.3230676, 0.3351025, 0.3296865, 
    0.309061, 0.2346846, 0.2122683, 0.153711, 0.07108648, 0.1167042, 
    0.1201023, 0.1386457, 0.1862779, 0.2659942,
  0.3889815, 0.3894192, 0.3898569, 0.3902946, 0.3907323, 0.39117, 0.3916077, 
    0.3631904, 0.3696859, 0.3761814, 0.3826769, 0.3891724, 0.3956679, 
    0.4021634, 0.4143451, 0.4083911, 0.4024372, 0.3964832, 0.3905292, 
    0.3845752, 0.3786213, 0.3584142, 0.357435, 0.3564558, 0.3554766, 
    0.3544973, 0.3535181, 0.3525389, 0.3886313,
  0.2819541, 0.4135261, 0.3907598, 0.2613956, 0.2509989, 0.1800222, 
    0.1876988, 0.208912, 0.1515888, 0.1686155, 0.2804485, 0.3548608, 
    0.3887846, 0.04324948, 0.1305899, 0.2745878, 0.2889864, 0.236313, 
    0.1607646, 0.2694505, 0.535722, 0.4802085, 0.321219, 0.1794083, 
    0.2633404, 0.3582686, 0.1702461, 0.08532062, 0.2859748,
  0.1844605, 0.1366595, 0.2656592, 0.1403116, 0.2031886, 0.1807305, 
    0.09316474, 0.2992496, 0.2932429, 0.277045, 0.250167, 0.1979779, 
    0.1918754, 0.1552092, 0.2036704, 0.3051795, 0.384338, 0.3185137, 
    0.3122066, 0.3603211, 0.4072613, 0.3764969, 0.3747107, 0.4407329, 
    0.3859468, 0.4445517, 0.327291, 0.3028969, 0.1806312,
  0.269197, 0.2488915, 0.2200171, 0.2888399, 0.3016453, 0.3606382, 0.4024129, 
    0.3792663, 0.4037684, 0.2539399, 0.2469067, 0.3464879, 0.4944203, 
    0.4276544, 0.3500932, 0.379924, 0.4209753, 0.4827657, 0.458993, 
    0.3892193, 0.3375183, 0.366978, 0.3964148, 0.3833166, 0.4635569, 
    0.4805209, 0.4495743, 0.4135205, 0.3246203,
  0.4032718, 0.386007, 0.3361487, 0.3267588, 0.3459594, 0.3548569, 0.3889933, 
    0.3671671, 0.3262939, 0.3137754, 0.2902102, 0.2776351, 0.2696893, 
    0.3209832, 0.2030281, 0.2796649, 0.2655584, 0.3102506, 0.2544556, 
    0.262755, 0.2238544, 0.2018681, 0.2479008, 0.1823907, 0.03242081, 
    0.2020081, 0.3605101, 0.3591052, 0.3865372,
  0.273182, 0.1882999, 0.08422775, 0.1855732, 0.2086505, 0.2030267, 
    0.2112276, 0.1853598, 0.1868774, 0.1158668, 0.1165932, 0.08032733, 
    0.04399904, 0.1911618, 0.2260292, 0.06629552, 0.1606739, 0.1605248, 
    0.1540751, 0.1754192, 0.1591297, 0.2398135, 0.1442286, 0.1212373, 
    0.02458544, 0.1532372, 0.2177992, 0.2230322, 0.2492467,
  0.09498989, 0.06758638, 0.03029027, 0.02627841, 0.06945954, 0.1333899, 
    0.04571118, 0.01702798, 0.03942921, 0.02293663, 0.02220301, 0.0004311582, 
    0.02009755, 0.03949325, 0.05230933, 0.03998762, 0.05982221, 0.1536935, 
    0.09711388, 0.03625813, 0.03348938, 0.04003304, 0.05514493, 0.03656313, 
    0.0383486, 0.01845663, 0.02702838, 0.01067735, 0.02596267,
  0.08459639, 0.03947861, 0.03539338, 0.007006362, 0.0440146, 0.01984296, 
    0.02641094, 0.0212408, 0.02894155, 0.005926249, 0.0003948357, 
    0.007152366, 0.01916135, 0.01647655, 0.0150876, 0.02816208, 0.02763788, 
    0.01270236, 0.01674451, 0.004554337, 0.007400704, 0.00429845, 0.04732415, 
    0.1769009, 0.041036, 0.1605343, 0.00307128, 0.009841322, 0.01926129,
  0.07691883, 0.06330753, 0.03160954, 0.02604679, 0.006972127, 0.007652927, 
    0.00966258, 0.01529866, 0.01820311, 0.01952258, 0.02345203, 0.02305137, 
    0.01816706, 0.007523356, 0.008681669, 0.01347678, 0.01365064, 0.01067218, 
    0.004734708, 0.008211015, 0.01307177, 0.02008666, 0.02600835, 0.04813736, 
    0.03442423, 0.02714643, 0.005295659, 0.007062452, 0.01996651,
  0.01424056, 0.002869486, 0.006644269, 0.01254376, 0.0321202, 0.01579081, 
    0.00907848, 0.002837684, 0.03677312, 0.08123064, 0.01909171, 0.03069365, 
    0.01276475, 0.006556889, 0.008434493, 0.01671193, 0.02554669, 0.03312271, 
    0.01847913, 0.07949106, 0.1424115, 0.1781956, 0.1468087, 0.006705318, 
    0.01632424, 0.01493049, 0.00443892, 0.007088313, 0.02036504,
  -3.625148e-08, 2.249711e-08, 4.187662e-08, 0.0001101552, 0.02171354, 
    0.01605725, 0.006562196, 0.01289075, 0.003499237, 0.01538389, 0.05369302, 
    0.01600353, 0.005991397, 0.005351174, 0.002437224, 0.003991183, 
    0.007408045, 0.02913921, 0.04570561, 0.02822944, 0.007563221, 
    0.002110975, 0.3183964, 0.09035127, 0.0008187272, 0.01140877, 0.03295369, 
    0.001562932, 8.868139e-06,
  1.113804e-08, 5.931128e-09, 4.582179e-11, 7.032926e-05, 1.204691e-09, 
    0.001710992, -1.706763e-05, 0.0003788489, 0.005729706, 0.2796991, 
    0.05210513, 0.04841548, 0.02130625, 0.01828428, 0.009797483, 0.005551771, 
    0.01228509, 0.01964981, 0.03896776, 0.06545995, 1.221464e-05, 0.1436485, 
    0.003764809, 0.002899788, 0.006325223, 0.01477567, 0.02448364, 
    0.002463844, 3.639799e-08,
  -1.04451e-05, 0.006917621, 0.01136935, 0.009621255, 0.004616073, 
    -7.479392e-06, -0.001668881, 0.01151519, 0.048127, 0.1479349, 0.1763828, 
    0.1082573, 0.1574791, 0.1120043, 0.1661455, 0.1447747, 0.09709127, 
    0.0964741, 0.09573247, 0.03445781, 0.01964444, 0.1839022, 0.07493094, 
    0.09042092, 0.07039765, 0.07552937, 0.08605149, 0.04106062, 0.001973008,
  -0.0007698745, 0.01546639, 0.02885792, 0.2003607, 0.02034324, 0.003654393, 
    0.0886748, 0.0002976098, 0.005336105, 0.02720216, 0.09406483, 0.07398476, 
    0.1225552, 0.1049751, 0.09787288, 0.1414922, 0.2103264, 0.2137378, 
    0.2038624, 0.1573797, 0.077531, 0.2181739, 0.1552445, 0.1158501, 
    0.1616241, 0.2607865, 0.1453064, 0.1788837, 0.08093343,
  0.1585485, 0.2219999, 0.1205654, 0.1095701, 0.1862514, 0.2509145, 
    0.1189167, 0.1526111, 0.04545984, 0.04231441, 0.009541974, 0.1094041, 
    0.1636692, 0.1880784, 0.1572787, 0.1827701, 0.2753046, 0.3023753, 
    0.2352393, 0.2544867, 0.09758447, 0.07463755, 0.09351896, 0.1860072, 
    0.1122061, 0.2168564, 0.2520157, 0.2254624, 0.2381466,
  0.2102102, 0.2556677, 0.297081, 0.4316945, 0.4613833, 0.2137675, 0.2623067, 
    0.1777759, 0.112144, 0.1524807, 0.1584229, 0.1535202, 0.1956907, 
    0.1992199, 0.4982352, 0.2318648, 0.2051634, 0.2384242, 0.2839594, 
    0.1618516, 0.1234582, 0.1118936, 0.2703283, 0.1858212, 0.3769968, 
    0.0472239, 0.08579526, 0.1875653, 0.1971408,
  0.09833208, 0.09369788, 0.2679637, 0.1960493, 0.3714388, 0.2758228, 
    0.3368548, 0.3648517, 0.2911344, 0.3749663, 0.5467422, 0.349572, 
    0.361084, 0.264201, 0.3077423, 0.2581947, 0.2706733, 0.1970603, 
    0.1792838, 0.3432015, 0.3039339, 0.3280501, 0.291869, 0.1232113, 
    0.1628549, 0.3867528, 0.3784801, 0.1228753, 0.2398995,
  0.1557074, 0.1993452, 0.3931611, 0.405618, 0.4001925, 0.4890005, 0.4566607, 
    0.4673497, 0.4370323, 0.4024754, 0.4319643, 0.4172944, 0.4215127, 
    0.4327222, 0.3821008, 0.3843616, 0.3703052, 0.3769876, 0.3743778, 
    0.3437168, 0.2884212, 0.2187273, 0.1605839, 0.08217137, 0.1384627, 
    0.1395445, 0.1313725, 0.2067335, 0.3056304,
  0.3155036, 0.3162057, 0.3169078, 0.3176098, 0.3183119, 0.319014, 0.3197162, 
    0.3323184, 0.339767, 0.3472155, 0.3546641, 0.3621126, 0.3695612, 
    0.3770098, 0.3706269, 0.3655427, 0.3604586, 0.3553744, 0.3502902, 
    0.345206, 0.3401218, 0.3634031, 0.3603366, 0.3572702, 0.3542037, 
    0.3511372, 0.3480707, 0.3450043, 0.3149419,
  0.344816, 0.4035065, 0.389024, 0.2622707, 0.2691538, 0.1537988, 0.1626217, 
    0.2055485, 0.1353413, 0.1261739, 0.2237383, 0.3518239, 0.4166906, 
    0.0271016, 0.1730066, 0.3159574, 0.3554208, 0.2513413, 0.1492712, 
    0.2429682, 0.5157537, 0.5206696, 0.292339, 0.1472779, 0.2603951, 
    0.3810148, 0.1191743, 0.0438836, 0.2699452,
  0.1285644, 0.0919603, 0.2096276, 0.09338492, 0.1481509, 0.1617053, 
    0.06395323, 0.2437222, 0.2599776, 0.249994, 0.2098928, 0.1980345, 
    0.1524408, 0.1014848, 0.1718016, 0.2438609, 0.3401354, 0.2661141, 
    0.2675425, 0.2874059, 0.3240328, 0.3605191, 0.3706482, 0.4512043, 
    0.3703191, 0.4213655, 0.2796828, 0.2458486, 0.1511747,
  0.2363484, 0.2145446, 0.1822391, 0.2366565, 0.2524119, 0.3082645, 
    0.3536284, 0.3204726, 0.3380816, 0.2128595, 0.2054464, 0.3063324, 
    0.4536369, 0.3774905, 0.3086233, 0.3474339, 0.3972675, 0.4585827, 
    0.4213178, 0.3433852, 0.3035299, 0.3294753, 0.3292626, 0.3371722, 
    0.4461672, 0.4861521, 0.4247859, 0.3758148, 0.2800951,
  0.3567607, 0.3425303, 0.3040001, 0.3050974, 0.3505543, 0.3490346, 
    0.3728722, 0.3344879, 0.2939281, 0.268821, 0.2323686, 0.2193773, 
    0.2412415, 0.284659, 0.194824, 0.2216772, 0.2131027, 0.2593668, 0.230863, 
    0.2434497, 0.2037643, 0.174881, 0.2043841, 0.1569696, 0.05863982, 
    0.2096286, 0.347675, 0.325442, 0.3568515,
  0.2072958, 0.1179595, 0.05565034, 0.1398254, 0.1623328, 0.1762178, 
    0.1524161, 0.1541038, 0.1322902, 0.07504358, 0.08908129, 0.04272019, 
    0.02503196, 0.1681809, 0.2161512, 0.03622879, 0.1351431, 0.142648, 
    0.1306961, 0.1602132, 0.1261605, 0.1920823, 0.09427491, 0.1193113, 
    0.02374012, 0.1065615, 0.1669539, 0.1702105, 0.1886167,
  0.0249891, 0.02496708, 0.02642056, 0.01170941, 0.04708627, 0.1078427, 
    0.0287042, 0.008159988, 0.0167117, 0.009037839, 0.01914474, 0.0004605899, 
    0.01693167, 0.03054428, 0.03571193, 0.02724827, 0.04008943, 0.1135283, 
    0.04933059, 0.01507925, 0.01280935, 0.01974244, 0.02174165, 0.03055736, 
    0.03011029, 0.007363864, 0.01281005, 0.003025193, 0.005079337,
  0.03068912, 0.05287801, 0.02516203, 0.001602605, 0.01718896, 0.004076283, 
    0.01044139, 0.008310343, 0.01067644, 0.001647641, 0.0001106394, 
    0.004481598, 0.008013455, 0.005635643, 0.005847158, 0.01275212, 
    0.0126416, 0.00138371, 0.007142199, 0.001573965, 0.002790683, 
    0.001523996, 0.01649483, 0.06674347, 0.03143062, 0.1427882, 0.001161554, 
    0.004306003, 0.007096945,
  0.02875159, 0.02099292, 0.02416423, 0.01607001, 0.00146162, 0.001629632, 
    0.004244312, 0.006906946, 0.006510464, 0.005252107, 0.0148691, 
    0.01218212, 0.004587919, 0.001448208, 0.001836416, 0.006765629, 
    0.005956003, 0.003157841, 0.0009832637, 0.003069297, 0.004695411, 
    0.006379948, 0.008234886, 0.04711512, 0.02895431, 0.0278451, 
    0.0001497628, 0.002573742, 0.006123714,
  0.003657073, 0.001344843, 0.004719581, 0.008316385, 0.01101007, 
    0.008235491, 0.00257598, 0.0009344462, 0.03800814, 0.06848779, 
    0.007766807, 0.008158084, 0.005419235, 0.0008742734, 0.001644537, 
    0.003778625, 0.005306704, 0.003481978, 0.002804744, 0.01239104, 
    0.03442489, 0.03871392, 0.1146756, 0.004840185, 0.01186225, 0.005947201, 
    0.0002181482, 0.001195854, 0.004706068,
  -5.548036e-08, 2.213707e-08, 9.138459e-08, 0.001080176, 0.009637524, 
    0.007175087, 0.0009199935, 0.005528908, 0.0006342395, 0.005148337, 
    0.02282868, 0.004775763, 0.001705027, 0.001525491, 0.0007166815, 
    0.0002514362, 0.001393869, 0.01208315, 0.01669275, 0.00932869, 
    0.001494761, 0.0004553764, 0.2420887, 0.07649927, 0.0003372119, 
    0.004640909, 0.013585, 0.0005952027, -1.321322e-05,
  1.065555e-08, 5.665507e-09, 1.991252e-10, 2.508059e-05, 1.127334e-09, 
    0.0005758117, -5.566202e-06, 0.0001457623, 0.004031721, 0.2016666, 
    0.01670345, 0.02031362, 0.005146021, 0.008170296, 0.002860827, 
    0.001672397, 0.009554736, 0.005349606, 0.01769374, 0.03833896, 
    -1.416304e-05, 0.1139037, 0.001098555, 0.0003078585, 0.00212613, 
    0.005708802, 0.01171017, 0.001178911, 3.518159e-08,
  -2.124528e-06, 0.003477818, 0.006620562, 0.006280168, 0.004048634, 
    -8.820853e-06, -0.001514693, 0.009339224, 0.03666776, 0.130583, 
    0.1785361, 0.09045742, 0.1285386, 0.07416715, 0.1372366, 0.0916654, 
    0.07042997, 0.07340898, 0.05630632, 0.03291426, 0.0170312, 0.1601551, 
    0.06404894, 0.07427564, 0.04248707, 0.04346808, 0.03334935, 0.01624834, 
    0.003616361,
  -0.0006340522, 0.009097034, 0.01863211, 0.1908663, 0.01058381, 0.001719547, 
    0.07393921, 0.000188037, 0.00392298, 0.02078214, 0.09648248, 0.06292457, 
    0.1025028, 0.08924286, 0.07554336, 0.1121654, 0.1675823, 0.1863482, 
    0.1624937, 0.1458468, 0.06270492, 0.1878176, 0.137468, 0.09901938, 
    0.1226702, 0.187109, 0.1043538, 0.1134227, 0.05593614,
  0.1004484, 0.1591921, 0.09179339, 0.09319372, 0.1729336, 0.2253142, 
    0.08472593, 0.1292114, 0.03604868, 0.03733131, 0.01006483, 0.1050062, 
    0.1696347, 0.1512424, 0.1368605, 0.1574135, 0.265258, 0.2731639, 
    0.1993945, 0.2292884, 0.08287454, 0.06041533, 0.07833174, 0.1899166, 
    0.08545247, 0.1870961, 0.2251994, 0.1589188, 0.1941001,
  0.1579978, 0.2716511, 0.2888891, 0.4286673, 0.4175045, 0.1649178, 
    0.2002859, 0.1456547, 0.08455354, 0.12193, 0.1305301, 0.1638062, 
    0.1814567, 0.1521909, 0.427641, 0.2479402, 0.1848093, 0.2149147, 
    0.2279494, 0.1654196, 0.1176894, 0.08706834, 0.2939377, 0.1642746, 
    0.3201317, 0.03086961, 0.07315441, 0.1518739, 0.1699784,
  0.07245101, 0.07407614, 0.2222223, 0.1329393, 0.3836558, 0.2627897, 
    0.3548746, 0.3179872, 0.3076223, 0.3659303, 0.5504844, 0.3515508, 
    0.4239877, 0.3116026, 0.3150037, 0.3321077, 0.3146457, 0.2095097, 
    0.1995917, 0.3678171, 0.3056517, 0.3968982, 0.3233607, 0.1412486, 
    0.151997, 0.331938, 0.3832071, 0.1032635, 0.1727746,
  0.207614, 0.2138202, 0.4765505, 0.4363345, 0.4319665, 0.5524967, 0.5113371, 
    0.5084634, 0.4868459, 0.4344181, 0.464536, 0.4591047, 0.4641508, 
    0.475829, 0.437929, 0.4593183, 0.4195549, 0.4313281, 0.4393355, 
    0.3925215, 0.3338294, 0.2183568, 0.1787227, 0.1329672, 0.1414475, 
    0.1427969, 0.1229153, 0.2300681, 0.3577555,
  0.2669948, 0.2668634, 0.2667319, 0.2666005, 0.266469, 0.2663375, 0.2662061, 
    0.2554302, 0.2678629, 0.2802956, 0.2927282, 0.3051609, 0.3175936, 
    0.3300262, 0.385896, 0.3806024, 0.3753088, 0.3700152, 0.3647216, 
    0.359428, 0.3541344, 0.3524132, 0.3454056, 0.338398, 0.3313904, 
    0.3243828, 0.3173752, 0.3103675, 0.2671,
  0.356951, 0.347257, 0.2891999, 0.2012404, 0.2631517, 0.1241804, 0.1364967, 
    0.2012479, 0.08525044, 0.08033445, 0.1409118, 0.2880643, 0.4128953, 
    0.01075303, 0.2526652, 0.3831647, 0.4850584, 0.3294025, 0.1494894, 
    0.2415811, 0.4720864, 0.5590545, 0.2513152, 0.1184436, 0.2644941, 
    0.43283, 0.09086238, 0.01817688, 0.2341649,
  0.09133691, 0.0643307, 0.1466394, 0.06022131, 0.1084019, 0.1426054, 
    0.04752123, 0.1824068, 0.2221143, 0.2054136, 0.1679817, 0.1902899, 
    0.1148367, 0.06805276, 0.1413544, 0.1799419, 0.2821648, 0.2071066, 
    0.2166947, 0.218832, 0.2578591, 0.3278732, 0.3519514, 0.4238143, 
    0.3398546, 0.3629061, 0.2290558, 0.1811804, 0.1135363,
  0.1942678, 0.1734374, 0.142655, 0.1804392, 0.2024635, 0.2519935, 0.2909427, 
    0.2550611, 0.2636727, 0.174926, 0.1705769, 0.2576891, 0.3975717, 
    0.3022908, 0.2422491, 0.2945477, 0.3399754, 0.4087615, 0.3719475, 
    0.294131, 0.2493799, 0.2626994, 0.2550547, 0.2579022, 0.39517, 0.451845, 
    0.380564, 0.3311141, 0.234546,
  0.2891582, 0.2745457, 0.2463241, 0.2574244, 0.3048387, 0.3116886, 
    0.3311576, 0.2801667, 0.2332195, 0.2026345, 0.1675867, 0.1607867, 
    0.187822, 0.2251263, 0.1830137, 0.1714547, 0.1614745, 0.1971494, 
    0.1923513, 0.2083208, 0.1680382, 0.136694, 0.1674618, 0.1244698, 
    0.07197626, 0.2065953, 0.3199571, 0.2887399, 0.3169954,
  0.149377, 0.07766943, 0.04185184, 0.1012491, 0.1221414, 0.1415193, 
    0.1257448, 0.1298462, 0.09355991, 0.04544169, 0.06052848, 0.01980099, 
    0.01688313, 0.1277322, 0.1960692, 0.02488771, 0.1103332, 0.1273433, 
    0.1163485, 0.1308627, 0.1002568, 0.13633, 0.05961746, 0.1141328, 
    0.01265681, 0.07703765, 0.0967732, 0.1104617, 0.1247611,
  0.01028759, 0.01212117, 0.02349762, 0.004995273, 0.01798383, 0.06923917, 
    0.01005959, 0.003423292, 0.009650601, 0.004221786, 0.009303235, 
    0.000188103, 0.01134927, 0.01823182, 0.02607147, 0.01602758, 0.02562926, 
    0.07854438, 0.02205129, 0.006410916, 0.005997636, 0.007681123, 0.0103671, 
    0.01670733, 0.02376106, 0.003215767, 0.006577257, 0.001430982, 0.001761696,
  0.01485315, 0.05020091, 0.01314347, 0.0006220619, 0.005234448, 0.001838871, 
    0.002536602, 0.001852661, 0.006512783, 0.0008470514, 5.270199e-05, 
    0.002164265, 0.003626222, 0.002229024, 0.00196366, 0.005519951, 
    0.005872754, 7.127141e-05, 0.002880792, 0.0005617506, 0.001008088, 
    0.0007364886, 0.007837213, 0.03413709, 0.02342996, 0.1181426, 
    0.0004401527, 0.001849661, 0.003129254,
  0.01511217, 0.008329175, 0.02143656, 0.01080654, 0.0007190171, 
    0.0007382298, 0.002304952, 0.004032397, 0.002913841, 0.002101619, 
    0.009016069, 0.006816319, 0.001257914, 0.0006507855, 0.0006019268, 
    0.003646333, 0.00238632, 0.001432628, 0.0004080586, 0.001695749, 
    0.002424087, 0.003269733, 0.004173846, 0.0492733, 0.02759075, 0.02917629, 
    -0.0004771635, 0.001315731, 0.003198804,
  0.001783252, 0.0008860649, 0.007406255, 0.005789767, 0.005241058, 
    0.004072252, 0.001162621, 0.0005033366, 0.03455827, 0.07979344, 
    0.003529194, 0.00375413, 0.003922384, 0.0003424409, 0.0005092922, 
    0.001012457, 0.001427509, 0.0005032144, 0.0005208204, 0.002990844, 
    0.00967418, 0.0133855, 0.0308421, 0.00430478, 0.0100438, 0.002272603, 
    5.579162e-05, 0.0005935216, 0.002291925,
  2.63401e-09, 2.190126e-08, 1.220009e-07, 0.0009674928, 0.005450862, 
    0.00415461, -3.799425e-05, 0.002942593, 0.0002227388, 0.001930835, 
    0.009190083, 0.001807842, 0.0002786745, 0.0003520932, 0.000366937, 
    3.021522e-05, 0.0004056686, 0.004581495, 0.006417563, 0.004247149, 
    0.0005711628, 0.0002618275, 0.1572307, 0.06265082, 0.0001959126, 
    0.002602392, 0.00689809, 0.0001788771, -6.94566e-05,
  1.046786e-08, 5.494104e-09, 3.122907e-10, 1.260276e-06, 1.088611e-09, 
    0.0002885521, -1.319927e-05, 6.149986e-05, 0.002974745, 0.07985774, 
    0.008904442, 0.01024344, 0.002265035, 0.003934556, 0.001479115, 
    0.0006818498, 0.005127331, 0.002045918, 0.008979964, 0.02330137, 
    -9.740868e-06, 0.08421794, 0.000615265, -0.0004839235, 0.001170097, 
    0.002687495, 0.006917745, 0.0007239028, 3.519156e-08,
  1.290554e-07, 0.002115034, 0.004086508, 0.003276694, 0.004375318, 
    -4.606282e-06, -0.001452942, 0.01016243, 0.02702949, 0.0970692, 
    0.1536853, 0.06800278, 0.08818293, 0.0486648, 0.09503536, 0.06692578, 
    0.05302969, 0.0536337, 0.03565913, 0.02488715, 0.01348424, 0.1321889, 
    0.05059774, 0.05482305, 0.02451915, 0.0234396, 0.01681228, 0.008864339, 
    0.003992684,
  -0.0005569599, 0.003083499, 0.01278314, 0.17441, 0.006429899, 0.001010027, 
    0.06174058, 8.323917e-05, 0.002578734, 0.01621057, 0.09556094, 
    0.04742978, 0.08625239, 0.06936386, 0.05463061, 0.08677663, 0.1238072, 
    0.1615741, 0.1223499, 0.1330242, 0.05485907, 0.1520581, 0.117338, 
    0.0841369, 0.09252837, 0.1242326, 0.0613298, 0.07493595, 0.03459672,
  0.06178274, 0.109837, 0.06187509, 0.07638399, 0.1413221, 0.1650003, 
    0.06167745, 0.1068529, 0.03168922, 0.03454034, 0.01287672, 0.09222525, 
    0.1705721, 0.1045159, 0.117389, 0.1358092, 0.2340636, 0.2176918, 
    0.1584859, 0.1956393, 0.06798211, 0.04742116, 0.06205148, 0.1771293, 
    0.06785282, 0.1595265, 0.1788993, 0.1109075, 0.1505863,
  0.1176444, 0.2660627, 0.2648315, 0.3807778, 0.3510839, 0.129411, 0.1356447, 
    0.1109247, 0.06539802, 0.09763566, 0.1031444, 0.1639991, 0.1921421, 
    0.1284504, 0.3404025, 0.2024783, 0.2006265, 0.1895208, 0.1785305, 
    0.1507692, 0.1075105, 0.06692742, 0.2690573, 0.1653507, 0.2827644, 
    0.02137055, 0.05984725, 0.1158303, 0.1243655,
  0.05505508, 0.05623415, 0.1999936, 0.09394088, 0.3355545, 0.281624, 
    0.3242509, 0.2942854, 0.2851389, 0.3534216, 0.5556152, 0.3413785, 
    0.4706474, 0.3360048, 0.3018422, 0.374271, 0.3235588, 0.2144979, 
    0.2315169, 0.3737757, 0.3057403, 0.470551, 0.3807241, 0.1754254, 
    0.1493804, 0.2727745, 0.3877205, 0.08635959, 0.1323495,
  0.3708421, 0.249412, 0.5362445, 0.4719419, 0.4960854, 0.5953893, 0.5437199, 
    0.4933313, 0.5304375, 0.4760999, 0.5143151, 0.4926243, 0.4447024, 
    0.4739361, 0.4979946, 0.5228026, 0.4576425, 0.438634, 0.4716164, 
    0.4526283, 0.4285118, 0.2145316, 0.2131677, 0.2091422, 0.1175327, 
    0.1260615, 0.112506, 0.2007802, 0.4020918,
  0.1199178, 0.1177846, 0.1156513, 0.1135181, 0.1113849, 0.1092516, 
    0.1071184, 0.09960042, 0.1177737, 0.135947, 0.1541203, 0.1722936, 
    0.1904669, 0.2086402, 0.2999954, 0.2979857, 0.295976, 0.2939662, 
    0.2919565, 0.2899467, 0.287937, 0.2686858, 0.2546555, 0.2406252, 
    0.2265948, 0.2125645, 0.1985341, 0.1845038, 0.1216244,
  0.3360108, 0.3168287, 0.1852857, 0.1075344, 0.1722946, 0.1107462, 
    0.1018745, 0.0613481, 0.02124184, 0.04383295, 0.1165776, 0.1994388, 
    0.3416706, 0.00576187, 0.3249657, 0.4520284, 0.4988592, 0.371905, 
    0.1294951, 0.2667596, 0.4546738, 0.6125655, 0.2056314, 0.09076214, 
    0.2975458, 0.467748, 0.1056661, 0.007262255, 0.1975139,
  0.06581592, 0.04549755, 0.1008371, 0.04359302, 0.07648067, 0.1173375, 
    0.03788668, 0.1434556, 0.1829815, 0.1525811, 0.1249153, 0.187318, 
    0.08658141, 0.04846954, 0.1048974, 0.1285628, 0.2150344, 0.153146, 
    0.1687187, 0.164627, 0.1969641, 0.2808942, 0.3077537, 0.3733972, 
    0.2985953, 0.2809862, 0.1670546, 0.1193895, 0.08286177,
  0.1420579, 0.1252505, 0.1059597, 0.1336586, 0.151957, 0.1961018, 0.2242764, 
    0.1905614, 0.1947576, 0.1376658, 0.1356606, 0.2014651, 0.3234784, 
    0.2348165, 0.1710947, 0.2208427, 0.2647784, 0.3491175, 0.3157328, 
    0.2471881, 0.1983744, 0.1874444, 0.1778743, 0.1791889, 0.3169759, 
    0.3794749, 0.3102115, 0.2638529, 0.1775027,
  0.2204234, 0.210254, 0.1880064, 0.1988018, 0.2524233, 0.2547997, 0.2760631, 
    0.2249543, 0.1744799, 0.1427686, 0.1081441, 0.1029184, 0.1353462, 
    0.167762, 0.1590286, 0.1291282, 0.1131564, 0.1375176, 0.1448742, 
    0.1574839, 0.1236868, 0.09048662, 0.1135017, 0.09868082, 0.06944653, 
    0.1727174, 0.2624167, 0.241275, 0.2559481,
  0.1057883, 0.04883801, 0.03013035, 0.0687307, 0.0797462, 0.1060796, 
    0.08806862, 0.08669674, 0.05957973, 0.02469932, 0.03668889, 0.01069759, 
    0.01053183, 0.08044521, 0.172074, 0.01568509, 0.07543906, 0.0888799, 
    0.08409701, 0.09063174, 0.06608966, 0.09105007, 0.03837364, 0.1022541, 
    0.005831464, 0.05199806, 0.06522089, 0.06791177, 0.08431613,
  0.006311693, 0.007648598, 0.01846296, 0.002532142, 0.006369852, 0.03430209, 
    0.003620891, 0.001550665, 0.006537484, 0.002456837, 0.004394538, 
    7.161846e-05, 0.009564204, 0.006525374, 0.01716376, 0.007541192, 
    0.01290694, 0.0519286, 0.009019773, 0.002983438, 0.002851279, 
    0.002939131, 0.006198974, 0.01045123, 0.01843414, 0.00131047, 
    0.003116969, 0.0008360825, 0.001041032,
  0.009290742, 0.04035095, 0.005527224, 0.0003925108, -0.0002517595, 
    0.001173889, 0.0009618299, 0.000767712, 0.002586325, 0.0005524945, 
    3.477677e-05, 0.0007914326, 0.001705836, 0.001151385, 0.0006553962, 
    0.002187229, 0.002616529, 4.643529e-05, 0.0008014519, 0.0001954404, 
    0.0004534978, 0.0004550796, 0.004672241, 0.02181165, 0.01563429, 
    0.09287331, 0.000200056, 0.001063631, 0.001825175,
  0.009757964, 0.003932824, 0.01971315, 0.01400306, 0.0004670491, 
    0.000465157, 0.0009878937, 0.001846439, 0.001410265, 0.0009741839, 
    0.004449309, 0.003121414, 0.0003996743, 0.0004107632, 0.0002624246, 
    0.00178692, 0.0008828384, 0.000736134, 0.0002754321, 0.001126808, 
    0.001514919, 0.002133732, 0.002641928, 0.04257404, 0.02779936, 
    0.02669369, -0.0003727153, 0.0008510358, 0.002058701,
  0.001093661, 0.0004840976, 0.005087194, 0.004297514, 0.002737441, 
    0.002204236, 0.000769588, 0.0003230874, 0.03023428, 0.08702286, 
    0.001632212, 0.00226271, 0.00182122, 0.0002094569, 0.000244582, 
    0.0004004683, 0.0007152841, 0.0002445792, 0.0002730425, 0.001549531, 
    0.004949911, 0.006825145, 0.01205141, 0.004056261, 0.007507871, 
    0.0008564052, 2.787604e-05, 0.0003890384, 0.001427527,
  5.960831e-09, 2.180151e-08, 1.159125e-07, 0.0007767954, 0.004107309, 
    0.002799219, -0.0002232376, 0.001682273, 0.0001099875, 0.001130202, 
    0.004027531, 0.0007508812, 9.169416e-05, 0.0001172713, 0.0002428006, 
    2.332175e-05, 0.0001443519, 0.001563993, 0.002894577, 0.00208667, 
    0.0002683435, 0.0001786685, 0.1143121, 0.04687707, 0.0001292024, 
    0.001717548, 0.004305414, 9.894919e-05, -0.0002039509,
  1.046571e-08, 5.390836e-09, 3.338559e-10, -1.501355e-06, 1.062342e-09, 
    0.0001851513, -3.20315e-05, 3.868463e-05, 0.002181412, 0.03058677, 
    0.005959094, 0.00436185, 0.001683391, 0.002190444, 0.0009903456, 
    0.0004180418, 0.002241271, 0.001078982, 0.005354135, 0.01228753, 
    -6.039935e-06, 0.06614369, 0.000425969, -0.0007143926, 0.0007717129, 
    0.00138775, 0.004746151, 0.0005099486, 3.522413e-08,
  -2.259025e-06, 0.001204695, 0.002480346, 0.002131499, 0.003935603, 
    -1.717266e-06, -0.001349901, 0.01679666, 0.02224527, 0.0647822, 
    0.1294233, 0.0436137, 0.05181289, 0.03130575, 0.06379022, 0.04141322, 
    0.03844467, 0.03898004, 0.02321346, 0.01744174, 0.01000737, 0.1014548, 
    0.03401651, 0.03480584, 0.01393797, 0.01288211, 0.01058356, 0.00576761, 
    0.003526694,
  -0.0005935417, 0.001547157, 0.009156439, 0.1597472, 0.003802959, 
    0.0007076219, 0.05119342, 4.730282e-05, 0.001863191, 0.01267272, 
    0.0843649, 0.03467342, 0.06845273, 0.05060841, 0.03683518, 0.06186048, 
    0.08517392, 0.1199673, 0.08226667, 0.1181193, 0.04797337, 0.1177291, 
    0.0985602, 0.07095927, 0.06900134, 0.0752419, 0.03383018, 0.04493595, 
    0.02319759,
  0.03662417, 0.07747106, 0.03971769, 0.06031028, 0.1118239, 0.1511446, 
    0.04585125, 0.09295605, 0.0339425, 0.03245955, 0.01220954, 0.07733952, 
    0.1551754, 0.07893286, 0.0987957, 0.1065921, 0.185039, 0.1657173, 
    0.1054709, 0.1742391, 0.05536941, 0.03484792, 0.04971137, 0.1497203, 
    0.05471007, 0.1390048, 0.128598, 0.0755305, 0.1062405,
  0.07923339, 0.2456856, 0.228034, 0.3252071, 0.2864891, 0.1027053, 
    0.1051698, 0.08636367, 0.05537001, 0.08103926, 0.08052093, 0.1715748, 
    0.2082532, 0.1122151, 0.2831314, 0.1621224, 0.2177487, 0.1652563, 
    0.1448617, 0.1301745, 0.09531976, 0.06186348, 0.2111685, 0.1711848, 
    0.2578108, 0.01666537, 0.04536517, 0.08325624, 0.08300766,
  0.04239596, 0.0403396, 0.1865158, 0.06548294, 0.3103672, 0.2759342, 
    0.3355342, 0.287266, 0.2602108, 0.3533751, 0.5217024, 0.3127693, 
    0.4948496, 0.3334149, 0.2758383, 0.3703964, 0.3144556, 0.1930302, 
    0.2573621, 0.3265709, 0.2641478, 0.5064628, 0.3776705, 0.2375541, 
    0.1517883, 0.2000833, 0.392068, 0.07785268, 0.1035479,
  0.4154606, 0.269589, 0.5408052, 0.4870483, 0.5221475, 0.5550868, 0.5105274, 
    0.443056, 0.4843462, 0.4796818, 0.5182236, 0.4555601, 0.4285424, 
    0.4470488, 0.4675327, 0.434522, 0.3785377, 0.3770962, 0.438242, 
    0.4270331, 0.4037549, 0.205844, 0.2411093, 0.3114711, 0.1053133, 
    0.0849436, 0.1099937, 0.2077571, 0.3640748,
  0.06396372, 0.0629687, 0.06197369, 0.06097867, 0.05998365, 0.05898863, 
    0.05799362, 0.06983283, 0.08252311, 0.09521338, 0.1079037, 0.1205939, 
    0.1332842, 0.1459745, 0.1949239, 0.1952286, 0.1955333, 0.195838, 
    0.1961427, 0.1964474, 0.1967522, 0.1777826, 0.1657827, 0.1537827, 
    0.1417827, 0.1297828, 0.1177828, 0.1057828, 0.06475973,
  0.3555908, 0.2807987, 0.1210056, 0.02272357, 0.07833562, 0.09882177, 
    0.06405025, 0.01651254, 0.008106502, 0.01856232, 0.0748438, 0.1745672, 
    0.2645457, 0.004448777, 0.3661038, 0.5086356, 0.4362582, 0.3555277, 
    0.1023166, 0.299792, 0.4281743, 0.624815, 0.1714632, 0.07876932, 
    0.2993975, 0.4914359, 0.106438, 0.005724958, 0.1698069,
  0.05189144, 0.03629725, 0.07886304, 0.03472871, 0.05878434, 0.09117928, 
    0.03299201, 0.1253593, 0.161717, 0.1285063, 0.1082007, 0.1728594, 
    0.06922552, 0.03843208, 0.07897104, 0.09844219, 0.1610998, 0.1166521, 
    0.1361968, 0.1324202, 0.157638, 0.2395839, 0.2620709, 0.3274594, 
    0.2496342, 0.2207505, 0.1253956, 0.08950274, 0.06499165,
  0.1128746, 0.09674241, 0.08269272, 0.1058077, 0.1198929, 0.1585662, 
    0.1787789, 0.1499768, 0.1525993, 0.1172276, 0.1145295, 0.1645702, 
    0.2613545, 0.1866109, 0.1265897, 0.1695159, 0.2082246, 0.3011444, 
    0.2655046, 0.1997895, 0.1462496, 0.1391487, 0.122614, 0.1289823, 
    0.2480614, 0.3061537, 0.2500758, 0.2131181, 0.1401412,
  0.1733366, 0.1661173, 0.1482216, 0.16192, 0.2057024, 0.2138917, 0.2380538, 
    0.1851327, 0.1381199, 0.1070877, 0.07583638, 0.0692422, 0.09472609, 
    0.1236592, 0.123882, 0.09750289, 0.08142728, 0.09558515, 0.1101877, 
    0.1181163, 0.09379771, 0.06580879, 0.08063176, 0.08500139, 0.06048251, 
    0.1363943, 0.2126225, 0.1970483, 0.2084708,
  0.0746792, 0.03164944, 0.02157946, 0.04242245, 0.04762141, 0.07523684, 
    0.05938205, 0.05888045, 0.03739543, 0.01553029, 0.02693797, 0.007203008, 
    0.007145943, 0.04870133, 0.1503724, 0.01090031, 0.04526587, 0.05882587, 
    0.05559553, 0.05573469, 0.03753494, 0.05868244, 0.02469378, 0.09153534, 
    0.003541413, 0.03717078, 0.03986274, 0.04260673, 0.05967043,
  0.004596888, 0.005558501, 0.0157159, 0.001652315, 0.002902547, 0.01709276, 
    0.001780014, 0.0009358595, 0.004987897, 0.001760038, 0.002527624, 
    4.641155e-05, 0.007039739, 0.002248767, 0.01224849, 0.003757566, 
    0.007510779, 0.03177131, 0.004559126, 0.001723495, 0.001385877, 
    0.001513912, 0.004463534, 0.008066095, 0.01242967, 0.0005860387, 
    0.001657283, 0.000603263, 0.0007479419,
  0.006801018, 0.03088511, 0.003309967, 0.0002929417, -0.001165866, 
    0.0008222624, 0.0005203532, 0.0004895361, 0.001642188, 0.0004112847, 
    3.041326e-05, 0.0003599231, 0.001201781, 0.0007698401, 0.0003110991, 
    0.001164289, 0.001403666, 6.104141e-05, 0.0003050187, 0.0001116762, 
    0.0002915531, 0.0003171808, 0.003286141, 0.01614862, 0.01024115, 
    0.07719173, 0.0001238752, 0.0007229958, 0.001255598,
  0.007188063, 0.002002428, 0.01777126, 0.02078093, 0.000349656, 
    0.0003380586, 0.0004293775, 0.0008895901, 0.0008536529, 0.0007270231, 
    0.002535819, 0.001539873, 0.0001403349, 0.0003023178, 0.0001742121, 
    0.0009954147, 0.0004091648, 0.0004279678, 0.0002054863, 0.0008429749, 
    0.001086956, 0.001610852, 0.001914915, 0.03292606, 0.02054911, 
    0.02179512, -0.00049505, 0.0006294078, 0.001516308,
  0.0007754524, 0.004383737, 0.003375917, 0.003310665, 0.001625221, 
    0.001358475, 0.0005749943, 0.0002343986, 0.02667809, 0.09464683, 
    0.0008174448, 0.001580251, 0.0009467074, 0.0001556904, 0.0001645004, 
    0.0002569525, 0.0004644195, 0.0001689697, 0.0001844971, 0.00102802, 
    0.003293426, 0.004608101, 0.007284231, 0.004892617, 0.005514373, 
    0.0003876972, 1.825499e-05, 0.0002903339, 0.001026933,
  5.433758e-09, 2.179234e-08, 1.186591e-07, 0.0003674293, 0.003173504, 
    0.002113034, -0.0002964921, 0.001174482, 2.298123e-05, 0.0007660675, 
    0.001998837, 0.0003764811, 4.685538e-05, 7.269534e-05, 0.0001817058, 
    2.492091e-05, 6.956233e-05, 0.0007506291, 0.001432016, 0.001056853, 
    0.0001531236, 0.0001317184, 0.07338256, 0.03159953, 9.457512e-05, 
    0.001281374, 0.0030995, 6.70267e-05, -0.0004813481,
  1.050555e-08, 5.308274e-09, 3.590099e-10, -2.825526e-06, 1.045075e-09, 
    0.0001275806, -1.738553e-05, 2.905977e-05, 0.001655016, 0.01688141, 
    0.004008218, 0.002144806, 0.001203785, 0.001330761, 0.0007539014, 
    0.0003063313, 0.00132957, 0.0007276976, 0.003930774, 0.008230646, 
    -4.836692e-06, 0.05441452, 0.0003308774, -0.0006989226, 0.0005873244, 
    0.0009103089, 0.003634865, 0.0003972675, 3.561102e-08,
  -2.71199e-06, 0.001022964, 0.001285537, 0.001423003, 0.003471384, 
    -7.661951e-07, -0.001285751, 0.03942835, 0.02205859, 0.04922466, 
    0.1023168, 0.02586972, 0.03048897, 0.01938809, 0.04123453, 0.02336898, 
    0.02799386, 0.02455288, 0.0153606, 0.01295609, 0.008577901, 0.07942422, 
    0.02442295, 0.02210896, 0.009415556, 0.008512103, 0.007824144, 
    0.004305941, 0.002685307,
  -0.0004226574, 0.001051756, 0.007098559, 0.1523172, 0.002528994, 
    0.0005301717, 0.04255146, 3.825559e-05, 0.001503403, 0.01013704, 
    0.07508101, 0.02452578, 0.05444493, 0.03769853, 0.02730535, 0.04469392, 
    0.05737737, 0.08493057, 0.05320324, 0.1037053, 0.04389942, 0.09874082, 
    0.08442998, 0.06353405, 0.05320263, 0.04705851, 0.02031848, 0.0324175, 
    0.01628636,
  0.0255245, 0.05723994, 0.02962713, 0.05527329, 0.09820051, 0.1441145, 
    0.03629852, 0.09429987, 0.04787, 0.03022141, 0.01128311, 0.06775546, 
    0.1386686, 0.06374981, 0.08517665, 0.08528568, 0.1419237, 0.1297761, 
    0.0714386, 0.1595542, 0.04684138, 0.0314019, 0.04153605, 0.1219091, 
    0.04705787, 0.1194931, 0.09605326, 0.05197953, 0.07221556,
  0.05602792, 0.2457218, 0.2103286, 0.2976454, 0.2501996, 0.08938708, 
    0.09596904, 0.07721258, 0.05206251, 0.07345275, 0.07014479, 0.2507355, 
    0.2411927, 0.1009176, 0.2480455, 0.1439904, 0.2336444, 0.1491271, 
    0.1456689, 0.1184416, 0.08862069, 0.07251632, 0.1634464, 0.1983548, 
    0.2423639, 0.01461826, 0.03554203, 0.06332972, 0.06133662,
  0.03318632, 0.03099569, 0.1929173, 0.0516598, 0.2910246, 0.243838, 
    0.366459, 0.3023307, 0.3004779, 0.3915737, 0.5037155, 0.3052458, 
    0.5164442, 0.2931547, 0.2527921, 0.3109164, 0.3229273, 0.1674159, 
    0.2618991, 0.263555, 0.2254323, 0.445781, 0.419494, 0.2647589, 0.1667746, 
    0.147921, 0.3845536, 0.07419518, 0.08574969,
  0.4299429, 0.2935258, 0.4769163, 0.4326306, 0.4508812, 0.4240757, 
    0.3617004, 0.2992074, 0.3553006, 0.3834826, 0.339314, 0.2985731, 
    0.3091938, 0.3168855, 0.3366503, 0.287598, 0.2384734, 0.2396875, 
    0.2738433, 0.2743542, 0.2658826, 0.1909537, 0.2757763, 0.4156953, 
    0.09753898, 0.04103043, 0.1125955, 0.2118717, 0.3118407,
  0.05622332, 0.05529313, 0.05436295, 0.05343276, 0.05250257, 0.05157238, 
    0.05064219, 0.04675078, 0.05649989, 0.06624901, 0.07599813, 0.08574723, 
    0.09549636, 0.1052455, 0.1466113, 0.1475283, 0.1484453, 0.1493623, 
    0.1502793, 0.1511963, 0.1521133, 0.1386401, 0.1289042, 0.1191683, 
    0.1094323, 0.09969641, 0.08996049, 0.08022456, 0.05696747,
  0.2992794, 0.2260726, 0.06605194, 0.004431335, 0.01666638, 0.05443574, 
    0.0376883, 0.004414632, 0.005555364, 0.01105713, 0.05031259, 0.1634708, 
    0.2480744, 0.004582278, 0.3742228, 0.4702267, 0.3778804, 0.335416, 
    0.09359711, 0.3062236, 0.411229, 0.6369511, 0.1673669, 0.07508811, 
    0.2854595, 0.4965265, 0.1176901, 0.01306455, 0.1559674,
  0.05614218, 0.03180083, 0.06837287, 0.03051296, 0.05158764, 0.07318798, 
    0.03308424, 0.113091, 0.1512798, 0.1184831, 0.09880356, 0.1679775, 
    0.06170399, 0.03352627, 0.06676961, 0.08383167, 0.1312598, 0.09845965, 
    0.1172613, 0.1128019, 0.1365671, 0.212366, 0.22986, 0.2976256, 0.2250376, 
    0.1916689, 0.1022313, 0.07391837, 0.05713998,
  0.09420949, 0.0806053, 0.07018426, 0.09005949, 0.1022263, 0.1367118, 
    0.1542938, 0.1257153, 0.1273582, 0.1001301, 0.09628333, 0.1412597, 
    0.2222873, 0.1519189, 0.1037147, 0.1390103, 0.1740493, 0.254319, 
    0.2220466, 0.1620461, 0.1170139, 0.1136454, 0.09419952, 0.1018234, 
    0.2007161, 0.2518998, 0.2114537, 0.1784957, 0.1176384,
  0.14467, 0.138096, 0.1213912, 0.132915, 0.1748973, 0.1796262, 0.2043333, 
    0.1567523, 0.1174935, 0.0889044, 0.05921528, 0.0507745, 0.07432275, 
    0.09723596, 0.09987228, 0.07800221, 0.062756, 0.0732034, 0.08533949, 
    0.09076869, 0.07525682, 0.05338772, 0.06239302, 0.09261371, 0.05233349, 
    0.1084691, 0.1725617, 0.1625255, 0.1758254,
  0.05442369, 0.02285215, 0.01557267, 0.02677136, 0.03095729, 0.04955685, 
    0.04055664, 0.04202963, 0.0245886, 0.01090462, 0.01827003, 0.00569622, 
    0.004916746, 0.03325998, 0.1529427, 0.00734926, 0.02819319, 0.03951798, 
    0.03935296, 0.03914123, 0.02579954, 0.03937773, 0.01719954, 0.09255376, 
    0.002632612, 0.02935343, 0.02715353, 0.03104826, 0.04433838,
  0.00374799, 0.004576411, 0.02325379, 0.001334259, 0.001917272, 0.01016266, 
    0.001122078, 0.0007309635, 0.004239497, 0.001452813, 0.001708591, 
    3.473766e-05, 0.009939089, 0.00141235, 0.007202597, 0.002338591, 
    0.004887751, 0.0198585, 0.00312022, 0.001262037, 0.0009301017, 
    0.001049375, 0.003659298, 0.006426801, 0.0278443, 0.000396926, 
    0.00117975, 0.0004936253, 0.0006127083,
  0.005612428, 0.02450821, 0.01266204, 0.0002332496, -0.00154115, 
    0.0006617435, 0.0003862545, 0.0003707267, 0.001311673, 0.0003400134, 
    0.0003736112, 0.0005813215, 0.0009677993, 0.0006223217, 0.0002281774, 
    0.0008110408, 0.0009828918, 5.773428e-05, 0.0002068354, 8.581857e-05, 
    0.0002303358, 0.0002560853, 0.002665856, 0.01326496, 0.02625198, 
    0.1146565, 9.392026e-05, 0.0005766379, 0.001003568,
  0.005901433, 0.0009733043, 0.03634221, 0.06847238, 0.0002659002, 
    0.0002730878, 0.000236397, 0.0005792117, 0.0006206056, 0.0003582471, 
    0.001787916, 0.001005016, 8.217882e-05, 0.0002481139, 0.0001372449, 
    0.0007031214, 0.0002784575, 0.000326021, 0.0001650861, 0.000699988, 
    0.0008895996, 0.001351675, 0.001565314, 0.07127926, 0.04360262, 
    0.05623103, -0.0004730945, 0.0005216992, 0.001251815,
  0.0006198853, 0.06936877, 0.007778696, 0.003426504, 0.001214598, 
    0.00103642, 0.0004763679, 0.0001905482, 0.03390963, 0.1244812, 
    0.0005563941, 0.001247799, 0.0006406757, 0.0001207453, 0.000131463, 
    0.0002047627, 0.0003621641, 0.0001413593, 0.0001492485, 0.0007968808, 
    0.002522963, 0.003508521, 0.00538444, 0.0407109, 0.03637742, 
    0.0002469065, 1.467692e-05, 0.0002405384, 0.0008300835,
  -6.249668e-08, 2.18527e-08, 1.186436e-07, 0.0005149522, 0.002949178, 
    0.001768327, -0.0005010735, 0.0008959135, -0.0002181918, 0.0006031244, 
    0.001263073, 0.0002692825, 3.511357e-05, 5.558124e-05, 0.0001542439, 
    2.530988e-05, 5.190542e-05, 0.0005003337, 0.0009584159, 0.0006454312, 
    0.000117908, 0.0001226744, 0.08531564, 0.0266815, 8.089816e-05, 
    0.001070418, 0.002532611, 5.288836e-05, -0.001729363,
  1.055511e-08, 5.272286e-09, 3.687431e-10, -1.617173e-06, 1.056201e-09, 
    0.0001095859, -1.273014e-05, 2.454875e-05, 0.005162544, 0.01164795, 
    0.002944939, 0.001517931, 0.0008923985, 0.000968394, 0.0006367691, 
    0.0002578993, 0.001023411, 0.0005789503, 0.003301727, 0.006489484, 
    -4.23601e-06, 0.04924822, 0.0002838072, -0.0008258108, 0.0004968387, 
    0.0007242839, 0.003076517, 0.0003391572, 3.600028e-08,
  -2.381594e-06, 0.0007659824, 0.0008707982, 0.001058912, 0.003538728, 
    -4.045254e-07, -0.001307081, 0.07117708, 0.03062318, 0.04479064, 
    0.07206663, 0.01699329, 0.02058035, 0.01195092, 0.02839089, 0.01529893, 
    0.01740158, 0.01376651, 0.01123385, 0.01005089, 0.008121258, 0.07291031, 
    0.02918655, 0.01533853, 0.005811132, 0.006265389, 0.006452129, 
    0.003628776, 0.002213902,
  -4.119918e-05, 0.0007248042, 0.006404092, 0.1611427, 0.001859006, 
    0.000429517, 0.04101728, 2.871256e-05, 0.001317205, 0.008558138, 
    0.07647249, 0.01934642, 0.04871196, 0.03048463, 0.02273716, 0.03551447, 
    0.04280306, 0.06296982, 0.03786063, 0.09834525, 0.04884622, 0.08703484, 
    0.07681458, 0.05434836, 0.04373565, 0.0341991, 0.01420326, 0.02421944, 
    0.01308673,
  0.02084569, 0.04636344, 0.02662221, 0.0646826, 0.09706475, 0.146279, 
    0.03238771, 0.1390018, 0.08680069, 0.03358834, 0.01053579, 0.0775525, 
    0.1377759, 0.05528532, 0.0752129, 0.07070743, 0.1157677, 0.1057389, 
    0.05283463, 0.1601166, 0.04689051, 0.03713324, 0.04439496, 0.1209891, 
    0.04484086, 0.1052448, 0.08028006, 0.03980388, 0.05568795,
  0.04425659, 0.3013195, 0.2252896, 0.3071871, 0.2504784, 0.1091816, 
    0.1036688, 0.1009551, 0.08588497, 0.1084118, 0.08566608, 0.4012459, 
    0.3047492, 0.1131713, 0.2299355, 0.1385021, 0.2899683, 0.1455756, 
    0.1971561, 0.1349829, 0.1090182, 0.1261197, 0.135259, 0.2703029, 
    0.2372359, 0.01767395, 0.03076576, 0.05314869, 0.04885459,
  0.02744376, 0.02627932, 0.2275622, 0.04462143, 0.2769918, 0.2260555, 
    0.4087166, 0.3491864, 0.4033365, 0.4505499, 0.5398802, 0.4011417, 
    0.5123858, 0.2921206, 0.2526418, 0.2700298, 0.3773685, 0.1932142, 
    0.2670909, 0.2322338, 0.2149901, 0.3837774, 0.4016982, 0.3086909, 
    0.1506566, 0.1366416, 0.3787341, 0.07691815, 0.07774681,
  0.4966288, 0.2678288, 0.4291373, 0.3457775, 0.3683421, 0.3249768, 0.283363, 
    0.2205231, 0.2893774, 0.2790202, 0.2497741, 0.226933, 0.2415142, 
    0.2324741, 0.2602611, 0.2277394, 0.1924603, 0.1903456, 0.2171841, 
    0.2266583, 0.2075349, 0.1952335, 0.3093769, 0.4467567, 0.1059647, 
    0.02905981, 0.127183, 0.2352478, 0.2674369 ;

 average_DT = 730 ;

 average_T1 = 75.5 ;

 average_T2 = 805.5 ;

 climatology_bounds =
  75.5, 805.5 ;

 lat = -89.5, -79.5, -69.5, -59.5, -49.5, -39.5, -29.5, -19.5, -9.5, 0.5, 
    10.5, 20.5, 30.5, 40.5, 50.5, 60.5, 70.5, 80.5 ;

 lat_bnds =
  -90, -89,
  -80, -79,
  -70, -69,
  -60, -59,
  -50, -49,
  -40, -39,
  -30, -29,
  -20, -19,
  -10, -9,
  0, 1,
  10, 11,
  20, 21,
  30, 31,
  40, 41,
  50, 51,
  60, 61,
  70, 71,
  80, 81 ;

 lon = 0.625, 13.125, 25.625, 38.125, 50.625, 63.125, 75.625, 88.125, 
    100.625, 113.125, 125.625, 138.125, 150.625, 163.125, 175.625, 188.125, 
    200.625, 213.125, 225.625, 238.125, 250.625, 263.125, 275.625, 288.125, 
    300.625, 313.125, 325.625, 338.125, 350.625 ;

 lon_bnds =
  0, 1.25,
  12.5, 13.75,
  25, 26.25,
  37.5, 38.75,
  50, 51.25,
  62.5, 63.75,
  75, 76.25,
  87.5, 88.75,
  100, 101.25,
  112.5, 113.75,
  125, 126.25,
  137.5, 138.75,
  150, 151.25,
  162.5, 163.75,
  175, 176.25,
  187.5, 188.75,
  200, 201.25,
  212.5, 213.75,
  225, 226.25,
  237.5, 238.75,
  250, 251.25,
  262.5, 263.75,
  275, 276.25,
  287.5, 288.75,
  300, 301.25,
  312.5, 313.75,
  325, 326.25,
  337.5, 338.75,
  350, 351.25 ;

 pfull = 0.0252729048206747, 0.0885404738757409, 0.213072411383256, 
    0.41190537807884, 0.671080828691593, 0.987471468515016, 1.36790961365676, 
    1.82562112064242, 2.38097588033244, 3.06218961364243, 3.90121721567151, 
    4.9296281825995, 6.18008131929323, 7.68875807563375, 9.49537809361575, 
    11.643153995098, 14.1786857151188, 17.1517875598959, 20.6152476986609, 
    24.6245259348741, 29.237386591333, 34.5134757786445, 40.5138467378254, 
    47.3004421634272, 54.9355325495126, 63.4811392623337, 72.9984371159701, 
    83.5471442618119, 95.1849171805989, 107.966767294215, 121.944503506415, 
    137.166169497631, 153.675572970355, 171.511834307961, 190.708985325578, 
    211.295632932361, 233.294677858721, 256.723099608772, 281.591803639405, 
    307.905555737256, 335.66293113824, 364.856338389786, 395.47216160598, 
    427.490864234311, 460.887168786725, 495.630391513078, 531.761718445649, 
    569.289185351388, 607.768705103107, 646.445374671436, 684.792067788697, 
    722.468679913451, 759.124006783627, 794.401045766566, 827.769968639223, 
    858.597822486016, 886.389109609622, 910.841030891388, 931.860653469283, 
    949.549679924174, 964.159924710431, 976.012345333387, 985.470174132691, 
    992.77226220014, 997.948601287575 ;

 time = 0 ;
}
