netcdf \00010101.atmos_daily.tile3.ts {
dimensions:
	time = UNLIMITED ; // (182 currently)
	phalf = 66 ;
	grid_xt = 15 ;
	grid_yt = 10 ;
	scalar_axis = 1 ;
	nv = 2 ;
	pfull = 65 ;
variables:
	double average_DT(time) ;
		average_DT:_FillValue = 1.e+20 ;
		average_DT:missing_value = 1.e+20 ;
		average_DT:units = "days" ;
		average_DT:long_name = "Length of average period" ;
	double average_T1(time) ;
		average_T1:_FillValue = 1.e+20 ;
		average_T1:missing_value = 1.e+20 ;
		average_T1:units = "days since 0001-01-01 00:00:00" ;
		average_T1:long_name = "Start time for average period" ;
	double average_T2(time) ;
		average_T2:_FillValue = 1.e+20 ;
		average_T2:missing_value = 1.e+20 ;
		average_T2:units = "days since 0001-01-01 00:00:00" ;
		average_T2:long_name = "End time for average period" ;
	float bk(phalf) ;
		bk:_FillValue = 1.e+20f ;
		bk:missing_value = 1.e+20f ;
		bk:long_name = "vertical coordinate sigma value" ;
		bk:cell_methods = "time: point" ;
	double grid_xt(grid_xt) ;
		grid_xt:units = "degrees_E" ;
		grid_xt:long_name = "T-cell longitude" ;
		grid_xt:axis = "X" ;
	double grid_yt(grid_yt) ;
		grid_yt:units = "degrees_N" ;
		grid_yt:long_name = "T-cell latitude" ;
		grid_yt:axis = "Y" ;
	float height10m(scalar_axis) ;
		height10m:_FillValue = 1.e+20f ;
		height10m:missing_value = 1.e+20f ;
		height10m:units = "m" ;
		height10m:long_name = "Height" ;
		height10m:cell_methods = "time: point" ;
		height10m:axis = "Z" ;
		height10m:positive = "up" ;
		height10m:standard_name = "height" ;
	float height2m(scalar_axis) ;
		height2m:_FillValue = 1.e+20f ;
		height2m:missing_value = 1.e+20f ;
		height2m:units = "m" ;
		height2m:long_name = "Height" ;
		height2m:cell_methods = "time: point" ;
		height2m:axis = "Z" ;
		height2m:positive = "up" ;
		height2m:standard_name = "height" ;
	double nv(nv) ;
		nv:long_name = "vertex number" ;
	double pfull(pfull) ;
		pfull:units = "mb" ;
		pfull:long_name = "ref full pressure level" ;
		pfull:axis = "Z" ;
		pfull:positive = "down" ;
	double phalf(phalf) ;
		phalf:units = "mb" ;
		phalf:long_name = "ref half pressure level" ;
		phalf:axis = "Z" ;
		phalf:positive = "down" ;
	float pk(phalf) ;
		pk:_FillValue = 1.e+20f ;
		pk:missing_value = 1.e+20f ;
		pk:units = "pascal" ;
		pk:long_name = "pressure part of the hybrid coordinate" ;
		pk:cell_methods = "time: point" ;
	double scalar_axis(scalar_axis) ;
		scalar_axis:long_name = "none" ;
	double time(time) ;
		time:units = "days since 0001-01-01 00:00:00" ;
		time:long_name = "time" ;
		time:axis = "T" ;
		time:calendar_type = "NOLEAP" ;
		time:calendar = "noleap" ;
		time:bounds = "time_bnds" ;
	double time_bnds(time, nv) ;
		time_bnds:long_name = "time axis boundaries" ;
	float ts(time, grid_yt, grid_xt) ;
		ts:_FillValue = 1.e+20f ;
		ts:missing_value = 1.e+20f ;
		ts:units = "K" ;
		ts:long_name = "Surface Temperature" ;
		ts:cell_methods = "time: mean" ;
		ts:cell_measures = "area: area" ;
		ts:time_avg_info = "average_T1,average_T2,average_DT" ;
		ts:standard_name = "surface_temperature" ;

// global attributes:
		:title = "cm5_c96_am5f7c1r0_b06_piC_galb_noiceinit_alb" ;
		:associated_files = "area: 00010101.grid_spec.nc" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
		:history = "Wed Apr 30 14:48:00 2025: ncks -d grid_xt,0,14 -d grid_yt,0,9 -d time,0,181 /home/cew/Code/cmip7-sprint/testfiles/input/00010101.atmos_daily.tile3.nc -O /home/cew/Code/cmip7-sprint/testfiles/00010101.atmos_daily.tile3.nc\nFri Apr 25 14:15:06 2025: ncks -x -v sphum,psl 00010101.atmos_daily.tile3.nc -o reduce/00010101.atmos_daily.tile3.nc\nFri Apr 25 13:47:12 2025: ncks -d grid_xt,35,55 -d grid_yt,30,45 00010101.atmos_daily.tile3.nc var_select/00010101.atmos_daily.tile3.nc" ;
		:NCO = "netCDF Operators version 5.1.9 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco, Citation = 10.1016/j.envsoft.2008.03.004)" ;
data:

 average_DT = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 average_T1 = 0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 
    18, 19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 
    36, 37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 
    54, 55, 56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 
    72, 73, 74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 
    90, 91, 92, 93, 94, 95, 96, 97, 98, 99, 100, 101, 102, 103, 104, 105, 
    106, 107, 108, 109, 110, 111, 112, 113, 114, 115, 116, 117, 118, 119, 
    120, 121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 
    134, 135, 136, 137, 138, 139, 140, 141, 142, 143, 144, 145, 146, 147, 
    148, 149, 150, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 
    162, 163, 164, 165, 166, 167, 168, 169, 170, 171, 172, 173, 174, 175, 
    176, 177, 178, 179, 180, 181 ;

 average_T2 = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 
    19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 
    37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 54, 
    55, 56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 72, 
    73, 74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 90, 
    91, 92, 93, 94, 95, 96, 97, 98, 99, 100, 101, 102, 103, 104, 105, 106, 
    107, 108, 109, 110, 111, 112, 113, 114, 115, 116, 117, 118, 119, 120, 
    121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 134, 
    135, 136, 137, 138, 139, 140, 141, 142, 143, 144, 145, 146, 147, 148, 
    149, 150, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 162, 
    163, 164, 165, 166, 167, 168, 169, 170, 171, 172, 173, 174, 175, 176, 
    177, 178, 179, 180, 181, 182 ;

 bk = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.00193294, 0.00749994, 0.01640714, 0.02841953, 
    0.04334756, 0.06103661, 0.0813586, 0.1042054, 0.1294836, 0.1571101, 
    0.1870091, 0.2191095, 0.2533426, 0.2896406, 0.3279357, 0.3681587, 
    0.4102391, 0.454293, 0.5001689, 0.5468886, 0.5935643, 0.6397641, 
    0.6851825, 0.729505, 0.7723162, 0.8125153, 0.8492141, 0.8817441, 
    0.909788, 0.9332725, 0.9524949, 0.9678352, 0.9798011, 0.9889621, 0.99575, 1 ;

 grid_xt = 36, 37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50 ;

 grid_yt = 31, 32, 33, 34, 35, 36, 37, 38, 39, 40 ;

 height10m = 10 ;

 height2m = 2 ;


 nv = 1, 2 ;

 pfull = 0.0252729048206747, 0.0885404738757409, 0.213072411383256, 
    0.41190537807884, 0.671080828691593, 0.987471468515016, 1.36790961365676, 
    1.82562112064242, 2.38097588033244, 3.06218961364243, 3.90121721567151, 
    4.9296281825995, 6.18008131929323, 7.68875807563375, 9.49537809361575, 
    11.643153995098, 14.1786857151188, 17.1517875598959, 20.6152476986609, 
    24.6245259348741, 29.237386591333, 34.5134757786445, 40.5138467378254, 
    47.3004421634272, 54.9355325495126, 63.4811392623337, 72.9984371159701, 
    83.5471442618119, 95.1849171805989, 107.966767294215, 121.944503506415, 
    137.166169497631, 153.675572970355, 171.511834307961, 190.708985325578, 
    211.295632932361, 233.294677858721, 256.723099608772, 281.591803639405, 
    307.905555737256, 335.66293113824, 364.856338389786, 395.47216160598, 
    427.490864234311, 460.887168786725, 495.630391513078, 531.761718445649, 
    569.289185351388, 607.768705103107, 646.445374671436, 684.792067788697, 
    722.468679913451, 759.124006783627, 794.401045766566, 827.769968639223, 
    858.597822486016, 886.389109609622, 910.841030891388, 931.860653469283, 
    949.549679924174, 964.159924710431, 976.012345333387, 985.470174132691, 
    992.77226220014, 997.948601287575 ;

 phalf = 0.01, 0.0513470268, 0.1404240036, 0.3072783852, 0.5379505539, 
    0.8245489502, 1.170559845, 1.5862843323, 2.0879000854, 2.700272522, 
    3.4550848389, 4.3841940308, 5.5185266113, 6.8925054932, 8.5440936279, 
    10.5147802734, 12.8495031738, 15.5965148926, 18.8071691895, 
    22.5356542969, 26.8386547852, 31.7749560547, 37.4049951172, 
    43.7903613281, 50.9932617188, 59.0759326172, 68.100078125, 78.1262353516, 
    89.2131933594, 101.4173632812, 114.7922466406, 129.3878501562, 
    145.2501478125, 162.4206823438, 180.9360560938, 200.8276451562, 
    222.1212074219, 244.8367185938, 268.9881007812, 294.5831945312, 
    321.6236510156, 350.1049399219, 380.0163883594, 411.3414303125, 
    444.0575547656, 478.1367280469, 513.5456339062, 550.403556875, 
    588.6019571094, 627.3470909766, 665.9273852344, 704.0097012891, 
    741.2475327734, 777.2856108203, 811.7659041211, 843.9830114648, 
    873.3803854492, 899.5263707422, 922.2501762402, 941.5376650684, 
    957.6070185254, 970.7426572876, 981.30107, 989.65107, 995.9000099865, 1000 ;

 pk = 1, 5.134703, 14.0424, 30.72784, 53.79506, 82.4549, 117.056, 158.6284, 
    208.79, 270.0273, 345.5085, 438.4194, 551.8527, 689.2505, 854.4094, 
    1051.478, 1284.95, 1559.651, 1880.717, 2253.565, 2683.865, 3177.496, 
    3740.5, 4379.036, 5099.326, 5907.593, 6810.008, 7812.624, 8921.319, 
    10141.74, 11285.93, 12188.79, 12884.3, 13400.12, 13758.85, 13979.1, 
    14076.26, 14063.13, 13950.46, 13747.31, 13461.45, 13099.54, 12667.38, 
    12170.08, 11612.19, 10997.8, 10330.65, 9611.055, 8843.304, 8045.85, 
    7236.312, 6424.557, 5606.509, 4778.059, 3944.972, 3146.775, 2416.634, 
    1778.226, 1246.215, 826.5195, 511.2139, 290.7407, 150, 68.893, 14.999, 0 ;

 scalar_axis = 0 ;


 time = 0.5, 1.5, 2.5, 3.5, 4.5, 5.5, 6.5, 7.5, 8.5, 9.5, 10.5, 11.5, 12.5, 
    13.5, 14.5, 15.5, 16.5, 17.5, 18.5, 19.5, 20.5, 21.5, 22.5, 23.5, 24.5, 
    25.5, 26.5, 27.5, 28.5, 29.5, 30.5, 31.5, 32.5, 33.5, 34.5, 35.5, 36.5, 
    37.5, 38.5, 39.5, 40.5, 41.5, 42.5, 43.5, 44.5, 45.5, 46.5, 47.5, 48.5, 
    49.5, 50.5, 51.5, 52.5, 53.5, 54.5, 55.5, 56.5, 57.5, 58.5, 59.5, 60.5, 
    61.5, 62.5, 63.5, 64.5, 65.5, 66.5, 67.5, 68.5, 69.5, 70.5, 71.5, 72.5, 
    73.5, 74.5, 75.5, 76.5, 77.5, 78.5, 79.5, 80.5, 81.5, 82.5, 83.5, 84.5, 
    85.5, 86.5, 87.5, 88.5, 89.5, 90.5, 91.5, 92.5, 93.5, 94.5, 95.5, 96.5, 
    97.5, 98.5, 99.5, 100.5, 101.5, 102.5, 103.5, 104.5, 105.5, 106.5, 107.5, 
    108.5, 109.5, 110.5, 111.5, 112.5, 113.5, 114.5, 115.5, 116.5, 117.5, 
    118.5, 119.5, 120.5, 121.5, 122.5, 123.5, 124.5, 125.5, 126.5, 127.5, 
    128.5, 129.5, 130.5, 131.5, 132.5, 133.5, 134.5, 135.5, 136.5, 137.5, 
    138.5, 139.5, 140.5, 141.5, 142.5, 143.5, 144.5, 145.5, 146.5, 147.5, 
    148.5, 149.5, 150.5, 151.5, 152.5, 153.5, 154.5, 155.5, 156.5, 157.5, 
    158.5, 159.5, 160.5, 161.5, 162.5, 163.5, 164.5, 165.5, 166.5, 167.5, 
    168.5, 169.5, 170.5, 171.5, 172.5, 173.5, 174.5, 175.5, 176.5, 177.5, 
    178.5, 179.5, 180.5, 181.5 ;

 time_bnds =
  0, 1,
  1, 2,
  2, 3,
  3, 4,
  4, 5,
  5, 6,
  6, 7,
  7, 8,
  8, 9,
  9, 10,
  10, 11,
  11, 12,
  12, 13,
  13, 14,
  14, 15,
  15, 16,
  16, 17,
  17, 18,
  18, 19,
  19, 20,
  20, 21,
  21, 22,
  22, 23,
  23, 24,
  24, 25,
  25, 26,
  26, 27,
  27, 28,
  28, 29,
  29, 30,
  30, 31,
  31, 32,
  32, 33,
  33, 34,
  34, 35,
  35, 36,
  36, 37,
  37, 38,
  38, 39,
  39, 40,
  40, 41,
  41, 42,
  42, 43,
  43, 44,
  44, 45,
  45, 46,
  46, 47,
  47, 48,
  48, 49,
  49, 50,
  50, 51,
  51, 52,
  52, 53,
  53, 54,
  54, 55,
  55, 56,
  56, 57,
  57, 58,
  58, 59,
  59, 60,
  60, 61,
  61, 62,
  62, 63,
  63, 64,
  64, 65,
  65, 66,
  66, 67,
  67, 68,
  68, 69,
  69, 70,
  70, 71,
  71, 72,
  72, 73,
  73, 74,
  74, 75,
  75, 76,
  76, 77,
  77, 78,
  78, 79,
  79, 80,
  80, 81,
  81, 82,
  82, 83,
  83, 84,
  84, 85,
  85, 86,
  86, 87,
  87, 88,
  88, 89,
  89, 90,
  90, 91,
  91, 92,
  92, 93,
  93, 94,
  94, 95,
  95, 96,
  96, 97,
  97, 98,
  98, 99,
  99, 100,
  100, 101,
  101, 102,
  102, 103,
  103, 104,
  104, 105,
  105, 106,
  106, 107,
  107, 108,
  108, 109,
  109, 110,
  110, 111,
  111, 112,
  112, 113,
  113, 114,
  114, 115,
  115, 116,
  116, 117,
  117, 118,
  118, 119,
  119, 120,
  120, 121,
  121, 122,
  122, 123,
  123, 124,
  124, 125,
  125, 126,
  126, 127,
  127, 128,
  128, 129,
  129, 130,
  130, 131,
  131, 132,
  132, 133,
  133, 134,
  134, 135,
  135, 136,
  136, 137,
  137, 138,
  138, 139,
  139, 140,
  140, 141,
  141, 142,
  142, 143,
  143, 144,
  144, 145,
  145, 146,
  146, 147,
  147, 148,
  148, 149,
  149, 150,
  150, 151,
  151, 152,
  152, 153,
  153, 154,
  154, 155,
  155, 156,
  156, 157,
  157, 158,
  158, 159,
  159, 160,
  160, 161,
  161, 162,
  162, 163,
  163, 164,
  164, 165,
  165, 166,
  166, 167,
  167, 168,
  168, 169,
  169, 170,
  170, 171,
  171, 172,
  172, 173,
  173, 174,
  174, 175,
  175, 176,
  176, 177,
  177, 178,
  178, 179,
  179, 180,
  180, 181,
  181, 182 ;

 ts =
  261.4232, 272.5475, 265.6495, 272.4573, 269.0145, 261.5891, 265.9818, 
    266.0406, 265.0528, 248.9288, 251.1606, 254.6861, 246.4969, 248.7467, 
    236.9789,
  273.9857, 274.3366, 273.8667, 273.251, 262.0461, 259.3752, 268.0388, 
    267.6493, 267.2528, 261.5524, 253.6797, 261.9098, 261.2255, 243.566, 
    237.404,
  274.549, 274.3253, 274.1998, 273.7679, 266.4384, 246.4558, 265.5848, 
    268.087, 269.0542, 265.7857, 264.2489, 264.5054, 263.9605, 262.2203, 
    252.6757,
  275.2407, 274.548, 274.3043, 273.9989, 273.6055, 266.5992, 241.8416, 
    259.9698, 270.1733, 266.5981, 265.2796, 265.0668, 264.6185, 263.4366, 
    258.1172,
  275.598, 274.8677, 274.3722, 274.0643, 273.6554, 273.1092, 268.7558, 
    240.5218, 245.7056, 254.8214, 264.954, 265.1902, 264.7043, 264.1416, 
    263.6872,
  275.8509, 275.1342, 274.492, 274.0281, 273.6563, 273.1708, 272.5679, 
    271.3146, 262.1692, 259.521, 257.3068, 265.1455, 264.8419, 264.7994, 
    264.5615,
  276.2159, 275.3926, 274.6307, 274.0139, 273.5748, 273.1279, 272.6599, 
    272.2452, 271.8737, 271.8689, 269.0397, 265.0277, 264.8685, 264.9608, 
    264.8604,
  276.4522, 275.5732, 274.7629, 274.0305, 273.4726, 273.0077, 272.5783, 
    272.2553, 271.9786, 271.9466, 270.1411, 265.6964, 265.1457, 265.4391, 
    265.4749,
  276.076, 275.4014, 274.6709, 273.9366, 273.3167, 272.8689, 272.4659, 
    272.192, 272.1202, 271.609, 270.9261, 266.1559, 265.1629, 265.1784, 
    264.4437,
  275.1428, 274.4504, 274.0824, 273.6014, 273.04, 272.6216, 272.3374, 
    271.7111, 269.3892, 261.0533, 264.7556, 266.5723, 265.1909, 265.252, 
    264.9557,
  260.9113, 272.2013, 264.2051, 272.1252, 264.4835, 258.6393, 260.5332, 
    260.2623, 259.5305, 251.6197, 253.2786, 255.6495, 252.4703, 252.1744, 
    246.4348,
  273.7076, 274.2257, 273.8093, 273.0449, 260.6055, 256.1472, 261.8936, 
    261.2067, 260.5548, 258.2043, 254.7179, 258.2436, 257.6117, 247.8571, 
    244.5694,
  274.3864, 274.1931, 274.1149, 273.6838, 265.6578, 243.3604, 261.3607, 
    262.2855, 262.1299, 260.058, 259.6718, 259.3856, 258.4526, 257.9774, 
    251.9971,
  275.0886, 274.4305, 274.1885, 273.8976, 273.556, 266.2726, 244.3935, 
    259.4481, 263.0703, 260.6169, 260.1694, 259.7016, 258.9276, 257.6768, 
    254.7654,
  275.4106, 274.7136, 274.2326, 273.9288, 273.5631, 272.934, 268.6429, 
    247.075, 247.5125, 255.497, 260.1198, 259.8994, 259.2355, 258.479, 
    258.1149,
  275.7095, 274.9878, 274.3295, 273.8784, 273.5259, 273.0885, 272.3579, 
    271.2177, 264.4097, 262.9635, 257.2044, 260.3738, 259.7642, 259.4067, 
    259.0878,
  276.0925, 275.2771, 274.483, 273.8482, 273.4282, 273.0031, 272.5526, 
    272.0751, 271.6267, 271.6322, 265.3049, 260.7178, 260.1572, 259.9277, 
    259.4501,
  276.3787, 275.4912, 274.6779, 273.9168, 273.352, 272.8666, 272.4411, 
    272.1112, 271.8094, 271.6971, 267.1726, 261.1601, 260.6808, 260.5198, 
    259.9947,
  276.0173, 275.3458, 274.6049, 273.8161, 273.1679, 272.6839, 272.3007, 
    272.0397, 271.9105, 271.4145, 268.4091, 261.677, 261.1417, 260.8136, 
    259.8739,
  275.0603, 274.3744, 273.9991, 273.4661, 272.8647, 272.4332, 272.1444, 
    271.5997, 269.7004, 263.2733, 264.592, 262.1345, 261.5235, 261.2768, 
    260.2748,
  266.9581, 272.4611, 263.8467, 271.8894, 264.7606, 259.7199, 261.139, 
    261.0038, 260.9916, 252.8575, 252.7801, 252.9339, 250.2005, 251.7315, 
    246.3572,
  273.6947, 274.1797, 273.7932, 272.927, 259.5136, 257.1024, 262.884, 
    262.2315, 262.2334, 259.1941, 254.1138, 255.872, 257.2929, 248.7141, 
    245.2556,
  274.3526, 274.1608, 274.0523, 273.6401, 266.582, 248.0284, 262.4416, 
    263.3374, 263.0574, 260.3058, 258.2545, 257.4529, 257.6061, 259.5309, 
    253.6783,
  275.0125, 274.373, 274.1254, 273.8594, 273.5971, 267.4239, 245.8319, 
    260.0533, 262.7541, 260.4036, 258.7846, 258.2536, 258.2664, 257.8349, 
    257.0465,
  275.3269, 274.6401, 274.1682, 273.8805, 273.5484, 273.0114, 269.2608, 
    247.2702, 251.175, 257.9452, 259.4659, 259.2844, 258.9626, 258.5599, 
    258.5129,
  275.6413, 274.9382, 274.2602, 273.8158, 273.4867, 273.0997, 272.5183, 
    271.2987, 265.9336, 265.646, 259.8548, 259.8284, 259.3519, 259.224, 
    258.9186,
  276.0531, 275.2315, 274.4219, 273.7866, 273.3915, 272.988, 272.5378, 
    272.0823, 271.6559, 271.479, 263.5905, 260.5712, 259.7262, 259.902, 
    259.7477,
  276.3444, 275.4417, 274.6267, 273.8831, 273.3414, 272.8773, 272.4042, 
    272.0865, 271.7866, 271.591, 264.9236, 261.0053, 260.3088, 260.7182, 
    259.5829,
  275.9795, 275.3147, 274.5796, 273.79, 273.1452, 272.6529, 272.2452, 
    271.9998, 271.8486, 271.2299, 265.9212, 261.2701, 260.9381, 260.4531, 
    258.7062,
  274.9955, 274.3195, 273.9604, 273.4071, 272.7852, 272.3469, 272.0625, 
    271.5429, 270.0785, 265.6929, 264.393, 261.4113, 261.4474, 260.308, 
    259.8017,
  268.2433, 272.5414, 266.413, 271.8187, 265.5292, 260.7764, 261.9235, 
    259.2482, 257.4232, 248.1523, 248.8481, 248.7672, 244.2604, 245.6659, 
    235.9377,
  273.5627, 274.1088, 273.7657, 272.8929, 258.7083, 256.8725, 264.2878, 
    262.0244, 259.8647, 256.2357, 250.5677, 252.3837, 254.0294, 242.0861, 
    236.8434,
  274.2689, 274.1042, 274.0269, 273.6133, 265.3709, 247.7682, 263.1978, 
    263.3817, 261.8015, 258.4598, 255.8, 253.3345, 253.3334, 256.3084, 
    249.8748,
  274.9724, 274.3317, 274.0931, 273.8428, 273.5976, 267.2036, 250.9528, 
    260.1742, 260.8491, 257.7421, 254.9741, 253.549, 253.8431, 254.812, 
    254.4188,
  275.2951, 274.616, 274.1387, 273.8532, 273.5339, 273.027, 269.6444, 
    251.7839, 252.139, 253.649, 254.3732, 254.2474, 254.99, 256.2798, 256.8486,
  275.6046, 274.9187, 274.2285, 273.7925, 273.4683, 273.1018, 272.5204, 
    271.0408, 263.5948, 262.9958, 255.6959, 255.4267, 256.0606, 256.9972, 
    256.0624,
  276.0326, 275.2077, 274.4032, 273.7736, 273.3885, 272.9814, 272.5187, 
    272.0536, 271.5334, 271.1066, 260.8328, 256.9967, 257.3243, 257.1219, 
    256.8154,
  276.3285, 275.412, 274.5975, 273.8758, 273.3459, 272.8961, 272.3749, 
    272.0553, 271.7337, 271.1598, 261.2251, 258.3658, 257.711, 257.518, 257.2,
  275.9539, 275.2995, 274.5721, 273.7888, 273.1504, 272.6853, 272.2274, 
    271.9639, 271.7912, 270.9352, 262.8768, 259.299, 258.0822, 258.2564, 
    257.5042,
  274.935, 274.2646, 273.935, 273.3792, 272.7463, 272.3162, 272.04, 271.4784, 
    270.1179, 264.9203, 261.7554, 259.5533, 259.2415, 258.597, 259.1073,
  267.4596, 272.5972, 268.3535, 271.8336, 265.3606, 262.1751, 261.6399, 
    256.3508, 254.6736, 246.9529, 244.2722, 246.7943, 241.833, 243.1037, 
    234.2209,
  273.4676, 274.0057, 273.7329, 272.7888, 262.9688, 261.3247, 260.2725, 
    257.2383, 255.5462, 253.543, 247.2299, 252.2016, 255.3134, 239.4828, 
    232.8709,
  274.2053, 274.0147, 273.9927, 273.5595, 268.4596, 255.294, 260.3916, 
    258.8813, 256.6668, 254.9126, 254.6928, 253.7459, 255.1882, 257.3857, 
    247.0334,
  274.9181, 274.2754, 274.055, 273.8246, 273.5725, 268.175, 252.2421, 
    257.2417, 257.3658, 255.7791, 254.2335, 253.9239, 255.095, 255.6094, 
    252.3885,
  275.2532, 274.5909, 274.1123, 273.8397, 273.516, 273.1097, 268.9947, 
    248.4467, 246.8338, 251.4336, 253.6988, 254.6718, 255.7691, 256.8853, 
    258.1474,
  275.56, 274.8989, 274.2181, 273.7846, 273.4538, 273.094, 272.5924, 
    270.4323, 261.851, 260.6966, 255.0816, 255.4867, 256.4041, 257.5228, 
    257.7222,
  275.9943, 275.196, 274.4126, 273.7645, 273.3781, 272.9613, 272.5406, 
    272.0344, 270.9618, 270.5199, 260.7969, 256.4236, 256.9974, 257.8633, 
    258.1747,
  276.3141, 275.4146, 274.5933, 273.8651, 273.3329, 272.8994, 272.37, 
    272.0236, 271.6773, 270.6799, 259.509, 257.1565, 257.7242, 258.3683, 
    258.352,
  275.9433, 275.3134, 274.5847, 273.7634, 273.1164, 272.7312, 272.2384, 
    271.9082, 271.7235, 270.5957, 260.6623, 257.8233, 258.2107, 258.8047, 
    258.9296,
  274.9331, 274.2496, 273.9149, 273.3295, 272.726, 272.335, 272.0378, 
    271.4134, 269.8429, 263.5536, 259.6741, 258.383, 258.7697, 259.8268, 
    261.6818,
  263.9435, 272.2047, 266.3773, 271.6471, 263.2143, 260.9157, 261.723, 
    257.9201, 255.3701, 244.3055, 240.6227, 247.4505, 243.9388, 245.6341, 
    237.3573,
  273.3396, 273.8849, 273.6863, 272.8015, 262.4869, 261.1938, 261.6315, 
    257.4351, 254.8957, 252.3257, 244.3177, 254.1342, 257.2939, 240.5549, 
    236.5019,
  274.1534, 273.9449, 273.9348, 273.4992, 268.8662, 257.4631, 259.9808, 
    257.7526, 255.0571, 255.3475, 255.1752, 255.8233, 257.6718, 258.153, 
    247.5691,
  274.8667, 274.2186, 273.9969, 273.8016, 273.5594, 268.4082, 252.6995, 
    254.7995, 255.4984, 254.9664, 254.6343, 255.5012, 256.9476, 257.287, 
    253.1065,
  275.1965, 274.5468, 274.0687, 273.8174, 273.5121, 273.1667, 268.3338, 
    246.3331, 242.5652, 248.5963, 253.6851, 255.833, 257.4677, 258.3761, 
    259.1075,
  275.502, 274.8462, 274.1916, 273.7732, 273.4538, 273.0958, 272.6004, 
    269.7813, 260.9453, 258.4045, 253.2261, 256.8468, 258.0024, 259.3187, 
    259.8003,
  275.9421, 275.1591, 274.3956, 273.7387, 273.3783, 272.9633, 272.5465, 
    271.9915, 270.2461, 269.3599, 261.2072, 257.9833, 258.5791, 259.6784, 
    260.682,
  276.2698, 275.3829, 274.5671, 273.8432, 273.344, 272.9125, 272.3591, 
    271.9674, 271.6112, 270.4501, 259.9236, 258.4246, 258.8052, 260.5119, 
    261.1411,
  275.9336, 275.3066, 274.5935, 273.7749, 273.1505, 272.7556, 272.2344, 
    271.8367, 271.6638, 270.3604, 260.4205, 258.6363, 259.6832, 261.2455, 
    261.9372,
  275.0149, 274.2575, 273.9263, 273.3412, 272.737, 272.339, 272.0338, 
    271.3848, 269.6542, 263.8236, 260.0703, 258.8664, 259.8386, 261.6104, 
    263.7567,
  261.1124, 271.8733, 264.5701, 270.7391, 257.687, 255.2397, 258.0868, 
    256.3057, 256.2793, 247.3473, 248.9675, 252.6294, 246.2282, 246.373, 
    240.419,
  273.1369, 273.7495, 273.605, 272.7885, 257.3758, 256.3075, 259.363, 
    257.1053, 256.443, 255.9084, 251.2973, 257.7324, 257.6642, 242.5402, 
    238.7871,
  274.1075, 273.884, 273.9063, 273.474, 266.3386, 253.5141, 258.2889, 
    257.5391, 256.8131, 257.5833, 257.5655, 258.5088, 259.106, 257.8298, 
    249.6864,
  274.8271, 274.1964, 273.9559, 273.7639, 273.4939, 267.7504, 253.0625, 
    252.3206, 256.235, 256.6241, 256.9484, 258.1416, 258.8394, 257.7557, 
    253.7147,
  275.146, 274.4969, 274.0324, 273.7665, 273.4544, 273.1153, 268.1027, 
    246.1869, 239.9875, 249.3446, 256.2171, 258.3426, 258.9175, 259.8886, 
    258.9174,
  275.5153, 274.7827, 274.1498, 273.7227, 273.4118, 273.0777, 272.5275, 
    270.0615, 259.7371, 257.1087, 253.2428, 258.6251, 260.1042, 260.7333, 
    259.7813,
  275.9653, 275.1094, 274.3459, 273.6947, 273.3437, 272.9526, 272.5456, 
    271.957, 270.1925, 268.6031, 262.1385, 259.0749, 260.4636, 260.9416, 
    260.596,
  276.2911, 275.3461, 274.5255, 273.8016, 273.3205, 272.9165, 272.3547, 
    271.9429, 271.555, 270.5832, 260.5206, 259.231, 260.5456, 261.6005, 
    261.3397,
  275.9615, 275.3074, 274.6109, 273.8112, 273.1952, 272.7687, 272.2258, 
    271.8155, 271.6118, 270.2993, 260.4783, 259.2056, 260.4858, 262.3375, 
    262.2982,
  275.0998, 274.2589, 273.9467, 273.388, 272.7543, 272.322, 272.0186, 
    271.4573, 270.0175, 263.6717, 260.1099, 259.4453, 260.5099, 262.3698, 
    263.1304,
  261.7363, 271.4237, 263.3221, 268.8239, 256.9417, 252.0104, 257.9299, 
    257.2326, 256.9525, 247.4311, 245.0631, 246.8502, 242.126, 243.3412, 
    237.716,
  273.0098, 273.6548, 273.5107, 272.5155, 254.5597, 249.4205, 258.5711, 
    258.3406, 257.7094, 256.1109, 248.7267, 254.0993, 254.4664, 240.2621, 
    236.7513,
  274.1129, 273.8542, 273.8855, 273.4256, 265.4718, 248.39, 256.1584, 
    258.8839, 258.6175, 258.2431, 256.9497, 256.6734, 256.3073, 255.8174, 
    249.2625,
  274.7974, 274.1876, 273.9321, 273.7369, 273.4415, 266.8122, 242.5681, 
    253.8942, 258.6292, 258.2465, 257.4656, 256.7981, 256.5521, 255.8676, 
    252.9954,
  275.1128, 274.474, 274.0123, 273.7248, 273.4187, 273.0749, 267.4781, 
    244.0155, 244.8339, 252.6437, 257.6479, 257.8631, 257.0428, 256.7134, 
    256.826,
  275.4903, 274.7397, 274.114, 273.6739, 273.3856, 273.0449, 272.429, 
    269.8653, 260.9554, 259.0914, 254.7075, 258.5045, 257.83, 258.235, 
    257.7079,
  275.9751, 275.1031, 274.3023, 273.6597, 273.3044, 272.9131, 272.4978, 
    271.8685, 269.9613, 268.0117, 261.843, 259.5562, 258.8282, 258.73, 
    258.1916,
  276.3077, 275.3453, 274.504, 273.7691, 273.285, 272.8698, 272.2964, 
    271.8938, 271.4991, 270.1426, 260.9374, 260.3817, 260.0012, 259.4552, 
    258.351,
  275.9885, 275.3087, 274.6245, 273.8289, 273.2027, 272.7344, 272.142, 
    271.7415, 271.5593, 269.5054, 260.5508, 260.5426, 260.4678, 259.9895, 
    259.1409,
  275.1982, 274.2737, 273.9579, 273.4156, 272.7361, 272.2618, 271.9321, 
    271.3716, 269.8225, 263.5882, 261.1229, 260.5834, 260.8812, 261.0603, 
    261.5252,
  263.0708, 270.7419, 261.5298, 265.5985, 256.0223, 253.1685, 254.4779, 
    253.0471, 252.969, 242.0873, 241.0491, 244.5164, 240.7443, 243.4241, 
    236.8141,
  272.8782, 273.54, 273.2657, 271.8618, 254.4479, 252.033, 256.17, 254.4057, 
    253.5008, 251.6497, 243.2083, 252.1838, 253.9379, 236.9551, 234.5235,
  274.0759, 273.799, 273.8455, 273.3594, 264.5103, 246.7874, 255.8831, 
    255.8812, 254.6382, 254.1717, 254.0794, 254.5702, 255.29, 255.3371, 
    247.4625,
  274.7646, 274.1438, 273.8929, 273.6977, 273.3279, 266.3121, 246.9043, 
    253.1799, 254.7043, 253.9121, 253.5221, 254.0724, 255.1887, 255.4147, 
    252.7348,
  275.0877, 274.4268, 273.9696, 273.6865, 273.3756, 272.9689, 267.2433, 
    246.9314, 243.9406, 248.9307, 253.6532, 254.7244, 255.7782, 256.3349, 
    256.9955,
  275.468, 274.7034, 274.072, 273.6322, 273.3365, 272.9896, 272.1694, 
    269.0132, 260.1767, 256.9154, 253.396, 255.632, 256.0714, 256.6968, 
    257.1712,
  275.9957, 275.0956, 274.2582, 273.6196, 273.2612, 272.8442, 272.4146, 
    271.655, 268.6841, 264.8691, 259.078, 256.8132, 256.3311, 257.0309, 
    257.7691,
  276.3198, 275.3277, 274.4662, 273.7328, 273.2353, 272.7945, 272.2167, 
    271.8291, 271.3987, 268.8894, 258.9529, 257.6884, 256.7748, 257.3061, 
    257.6007,
  275.993, 275.2983, 274.6071, 273.7831, 273.1396, 272.659, 272.0416, 
    271.6628, 271.4876, 268.8007, 259.3813, 258.451, 257.6712, 257.6299, 
    257.0624,
  275.2492, 274.2621, 273.9238, 273.3662, 272.6459, 272.1527, 271.8124, 
    271.2362, 269.3967, 262.8392, 261.3418, 259.9736, 258.3296, 258.3919, 
    258.1836,
  258.7344, 269.1049, 258.2493, 261.9556, 254.0632, 250.942, 254.3486, 
    254.0804, 255.3644, 248.1058, 247.487, 250.4166, 246.2, 245.6898, 239.1406,
  272.4656, 273.3843, 272.8066, 270.6246, 251.1052, 248.064, 254.774, 
    254.721, 254.4761, 254.3661, 248.7949, 254.9108, 256.253, 245.1077, 
    242.799,
  273.9827, 273.7234, 273.771, 273.2513, 262.1109, 244.6616, 252.6146, 
    254.808, 254.5642, 254.6463, 254.4886, 255.4542, 256.9922, 257.9901, 
    252.517,
  274.7054, 274.0907, 273.8301, 273.642, 273.1999, 264.5095, 245.567, 
    249.7584, 253.7267, 253.45, 253.6119, 254.6466, 256.465, 257.7623, 
    256.6761,
  275.041, 274.3675, 273.9087, 273.6406, 273.3306, 272.8951, 266.6671, 
    242.3952, 240.0457, 246.8207, 252.8125, 254.711, 256.5843, 258.0399, 
    259.662,
  275.4219, 274.6673, 274.0138, 273.5827, 273.3003, 272.9508, 272.045, 
    269.0595, 257.0401, 253.2696, 250.0012, 255.2472, 256.5043, 258.2053, 
    259.4999,
  276.0062, 275.0853, 274.2246, 273.5873, 273.2279, 272.7715, 272.3635, 
    271.5877, 268.7217, 264.4316, 258.795, 256.1262, 256.8917, 258.4243, 
    260.0999,
  276.3353, 275.3192, 274.4251, 273.7073, 273.2012, 272.7146, 272.1321, 
    271.7705, 271.2605, 268.3074, 257.8518, 256.8062, 257.2178, 258.4415, 
    259.7106,
  276.0136, 275.2884, 274.5872, 273.7401, 273.0653, 272.5688, 271.9345, 
    271.5723, 271.3958, 267.882, 257.9074, 257.4628, 256.9693, 258.4042, 
    259.3104,
  275.3009, 274.2386, 273.8794, 273.2974, 272.5501, 272.0278, 271.6898, 
    271.1641, 268.8966, 261.3301, 260.6493, 258.2077, 256.7633, 257.79, 
    259.0513,
  256.0547, 267.5735, 255.5841, 261.2415, 255.1591, 250.2682, 254.9458, 
    255.2014, 256.9654, 252.2241, 251.9227, 253.5082, 248.1113, 247.7612, 
    241.5481,
  272.0666, 273.2245, 272.7478, 269.8798, 249.7635, 247.5349, 254.8302, 
    255.5184, 256.0513, 257.2657, 254.3952, 258.3767, 258.4517, 243.4737, 
    242.8945,
  273.9179, 273.6344, 273.7255, 273.1617, 260.5818, 244.1057, 252.132, 
    255.6209, 256.7296, 257.4854, 258.4975, 259.9125, 260.458, 260.5782, 
    256.382,
  274.6455, 274.044, 273.788, 273.6263, 273.274, 264.1954, 244.4649, 
    251.0762, 255.7589, 256.9673, 258.6336, 260.0292, 260.9445, 261.266, 
    260.2172,
  274.9929, 274.3179, 273.8784, 273.6287, 273.3345, 272.9153, 267.0238, 
    244.3012, 247.6882, 253.8584, 258.83, 260.1953, 261.0816, 260.8702, 
    261.8288,
  275.3694, 274.6462, 273.9997, 273.5833, 273.2849, 272.9394, 272.0663, 
    268.8506, 256.9297, 255.2601, 257.3967, 260.3128, 260.6381, 260.7121, 
    261.4378,
  275.9828, 275.0732, 274.2289, 273.5674, 273.2015, 272.7139, 272.3181, 
    271.304, 268.0767, 264.0417, 260.4763, 261.2055, 261.7663, 260.6693, 
    261.1686,
  276.3317, 275.3253, 274.4116, 273.6974, 273.1785, 272.6189, 272.0475, 
    271.6994, 271.0421, 266.6947, 259.746, 261.0594, 261.7307, 261.064, 
    261.1573,
  276.0236, 275.2959, 274.6054, 273.7143, 272.9988, 272.4687, 271.8117, 
    271.4673, 271.1575, 265.9151, 258.6565, 260.4384, 261.1664, 261.7325, 
    261.6529,
  275.3553, 274.2736, 273.9008, 273.2834, 272.5017, 271.919, 271.5616, 
    271.0046, 268.8804, 262.5709, 258.5878, 260.2164, 260.6185, 261.581, 
    262.1179,
  254.9844, 266.7078, 256.2479, 261.7444, 256.8997, 251.0382, 256.961, 
    258.4613, 259.8134, 253.2231, 253.7732, 256.701, 253.6305, 253.5282, 
    249.7036,
  271.4563, 273.086, 272.8708, 270.2336, 254.3277, 249.2959, 256.7924, 
    258.0692, 258.6342, 258.9026, 255.5981, 259.9731, 260.6905, 250.9922, 
    251.5643,
  273.8395, 273.5293, 273.7067, 273.1008, 261.8173, 249.184, 253.0892, 
    258.1307, 258.9257, 258.9058, 258.5948, 259.636, 260.4421, 260.6278, 
    258.9453,
  274.5888, 274, 273.756, 273.6044, 273.2786, 264.463, 244.6446, 251.8942, 
    257.5504, 257.7927, 258.0379, 258.5286, 259.4493, 259.9791, 259.8974,
  274.9623, 274.2723, 273.8523, 273.6089, 273.307, 272.8636, 266.6365, 
    244.461, 249.6289, 251.0372, 256.6053, 257.6006, 258.4891, 258.8051, 
    259.7604,
  275.3355, 274.6484, 273.9874, 273.5603, 273.2319, 272.867, 271.8957, 
    267.7462, 256.429, 255.0652, 256.5939, 257.1265, 257.6491, 258.0772, 
    258.979,
  275.9623, 275.0689, 274.2415, 273.5623, 273.1661, 272.5992, 272.2316, 
    270.7809, 266.6182, 263.8119, 258.3108, 257.6032, 257.5847, 257.7484, 
    258.2825,
  276.334, 275.3205, 274.4169, 273.7029, 273.1769, 272.5452, 271.9664, 
    271.6275, 270.5271, 265.6189, 257.8878, 257.7196, 257.7774, 257.8984, 
    258.213,
  276.0262, 275.3021, 274.6427, 273.7456, 273.0204, 272.4655, 271.7491, 
    271.3806, 270.9822, 265.1923, 257.9356, 257.4417, 257.4038, 258.1793, 
    258.9951,
  275.3715, 274.2681, 273.8803, 273.2968, 272.5431, 271.9644, 271.5353, 
    271.0184, 269.1597, 261.439, 258.8222, 258.4683, 257.0549, 257.9058, 
    259.3874,
  255.3133, 265.6208, 259.5375, 262.4636, 257.5513, 252.0197, 259.1443, 
    257.6997, 257.4532, 252.3165, 252.3258, 255.4952, 254.5423, 254.8708, 
    250.6309,
  270.3796, 272.7484, 272.7814, 269.9684, 254.146, 250.6026, 256.8045, 
    259.3344, 256.7977, 256.3917, 254.5661, 257.0272, 258.3889, 252.7138, 
    251.3291,
  273.7852, 273.3992, 273.635, 272.9759, 264.7735, 252.148, 254.6519, 
    256.5119, 256.1799, 256.117, 255.9141, 257.2132, 258.5168, 259.0701, 
    257.8647,
  274.5171, 273.9458, 273.6912, 273.5402, 273.2387, 267.1989, 250.8799, 
    251.1846, 255.1062, 255.3668, 255.5533, 256.5909, 257.8994, 258.9374, 
    258.9826,
  274.8929, 274.2115, 273.7839, 273.5614, 273.2582, 272.7612, 268.1661, 
    245.0708, 245.2993, 252.5891, 256.1136, 256.2057, 256.7911, 257.7514, 
    259.3914,
  275.2686, 274.6214, 273.9446, 273.5193, 273.1681, 272.7621, 271.791, 
    267.5242, 256.7053, 253.2679, 254.829, 256.7251, 256.5588, 257.0464, 
    258.537,
  275.9199, 275.0461, 274.2226, 273.5508, 273.119, 272.5074, 272.2066, 
    270.8007, 267.2951, 262.9399, 258.9227, 258.3706, 257.3155, 256.4828, 
    257.8602,
  276.3246, 275.2837, 274.3971, 273.6827, 273.1523, 272.4875, 271.94, 
    271.6324, 270.5158, 266.3707, 261.1541, 259.8624, 258.463, 256.9846, 
    257.6781,
  276.0309, 275.3107, 274.6389, 273.6954, 272.9686, 272.441, 271.7638, 
    271.3987, 271.1348, 267.8981, 263.859, 261.4677, 259.5493, 257.9658, 
    259.2708,
  275.4294, 274.2887, 273.821, 273.2244, 272.485, 271.9181, 271.5509, 
    271.1154, 269.4875, 267.7783, 266.9395, 263.7391, 260.8296, 258.8926, 
    258.2512,
  257.8484, 262.9321, 258.2532, 258.6942, 257.5598, 256.1154, 258.4031, 
    257.8722, 254.9996, 251.904, 252.8035, 253.4739, 252.8228, 254.2226, 
    248.4757,
  269.8528, 272.3668, 272.1473, 268.2592, 255.3764, 254.4165, 258.5296, 
    259.3849, 255.8515, 253.9002, 252.8162, 256.7096, 258.0749, 251.2712, 
    250.8299,
  273.8242, 273.3284, 273.5565, 272.8175, 265.7813, 248.0203, 258.3732, 
    259.0348, 255.828, 254.8096, 255.7894, 258.8674, 259.8073, 259.1673, 
    257.6708,
  274.4552, 273.896, 273.6314, 273.4874, 273.1468, 267.6811, 253.9932, 
    254.3598, 256.5142, 255.2372, 255.9678, 259.959, 259.9866, 260.0898, 
    258.7133,
  274.8072, 274.1448, 273.7352, 273.5175, 273.2256, 272.6704, 269.0146, 
    256.439, 253.5935, 256.5647, 256.8487, 261.2872, 260.8449, 260.3583, 
    259.472,
  275.1932, 274.581, 273.908, 273.4819, 273.1196, 272.6393, 271.7257, 
    268.472, 263.8436, 260.5077, 259.1074, 262.6526, 262.6084, 261.3609, 
    260.7387,
  275.8719, 275.0561, 274.1823, 273.5023, 273.0554, 272.4315, 272.1454, 
    270.9206, 268.2538, 266.9952, 264.7383, 264.5096, 264.4232, 263.1309, 
    261.619,
  276.2607, 275.2393, 274.3685, 273.6564, 273.123, 272.4442, 271.8976, 
    271.6105, 270.5653, 267.9244, 266.7465, 266.1372, 265.6398, 264.384, 
    263.3113,
  275.9695, 275.2695, 274.6404, 273.6423, 272.8834, 272.3953, 271.7643, 
    271.3493, 271.018, 267.4733, 266.1728, 266.0613, 266.3351, 265.3022, 
    264.5887,
  275.3896, 274.2384, 273.7788, 273.1583, 272.4116, 271.8451, 271.522, 
    271.0857, 269.4509, 266.9691, 268.8282, 267.8737, 267.0375, 266.2297, 
    265.3116,
  259.8051, 262.1688, 259.4472, 258.6809, 255.6031, 253.335, 255.7259, 
    255.1952, 255.5512, 250.886, 250.8684, 254.0594, 254.0474, 256.6777, 
    249.4466,
  269.7392, 271.3168, 270.6687, 264.8833, 254.5056, 252.6844, 256.8243, 
    257.1283, 256.8672, 256.3022, 253.4411, 257.0636, 260.2488, 259.0181, 
    251.002,
  273.9132, 273.4326, 273.5182, 272.3384, 263.1278, 248.8943, 255.1485, 
    258.5269, 259.3969, 258.5767, 258.5746, 261.4783, 262.6459, 263.8695, 
    256.2332,
  274.4861, 273.9047, 273.5846, 273.4464, 272.9479, 265.5757, 249.5002, 
    254.8813, 260.7254, 262.5602, 261.5485, 263.8246, 264.4998, 264.5926, 
    259.1998,
  274.7736, 274.1234, 273.6849, 273.4635, 273.1832, 272.5741, 267.4618, 
    252.7394, 256.3778, 262.2302, 263.9773, 264.8841, 265.2112, 265.1161, 
    261.8595,
  275.1326, 274.5336, 273.8748, 273.4467, 273.0793, 272.5741, 271.5771, 
    267.6047, 263.2307, 264.8909, 264.3774, 265.602, 265.736, 265.448, 
    264.0216,
  275.8089, 275.075, 274.1571, 273.467, 273.012, 272.3793, 272.0926, 
    270.9685, 268.496, 267.795, 266.7874, 266.321, 266.1225, 265.4735, 264.829,
  276.2372, 275.2337, 274.3397, 273.6215, 273.0972, 272.3881, 271.8414, 
    271.5706, 270.3883, 265.8582, 264.7303, 265.7419, 266.5438, 266.4671, 
    265.0345,
  275.9367, 275.2625, 274.662, 273.5799, 272.7669, 272.3225, 271.7168, 
    271.231, 270.8013, 266.7975, 265.5283, 266.9633, 267.1128, 267.0129, 
    266.6698,
  275.348, 274.2106, 273.7214, 273.0666, 272.3137, 271.7346, 271.4595, 
    270.9091, 268.9311, 265.4422, 267.7896, 268.0709, 267.8289, 267.8049, 
    267.7654,
  257.7408, 260.0534, 257.1849, 257.1173, 254.1974, 251.1339, 253.6207, 
    254.5422, 256.2919, 257.2204, 256.066, 256.5437, 250.8286, 247.9422, 
    239.5541,
  269.9369, 269.9408, 269.2879, 261.4961, 253.0112, 249.7826, 254.943, 
    255.5426, 257.7307, 260.4174, 259.8125, 260.7949, 260.2144, 249.5608, 
    245.9465,
  273.9305, 273.3701, 273.456, 271.3721, 262.0311, 245.5097, 253.4762, 
    256.0917, 259.5244, 262.7686, 264.1909, 264.8886, 264.1262, 261.6875, 
    254.5158,
  274.5044, 273.8914, 273.5399, 273.4133, 272.6728, 264.6778, 247.4635, 
    253.2871, 259.1862, 264.3049, 264.6717, 265.3629, 265.506, 264.7501, 
    259.6867,
  274.7625, 274.0936, 273.6428, 273.4323, 273.1629, 272.4818, 267.0288, 
    247.6311, 253.4996, 261.8378, 264.8713, 265.419, 265.5477, 265.6792, 
    263.021,
  275.0899, 274.5039, 273.8474, 273.4293, 273.0679, 272.5971, 271.417, 
    266.8936, 259.108, 263.3022, 263.9113, 265.64, 265.5958, 263.4796, 
    265.2494,
  275.7655, 275.0854, 274.142, 273.4499, 273.005, 272.395, 272.0625, 
    270.6679, 267.8633, 265.43, 266.1409, 265.9814, 265.6881, 264.4514, 
    266.1855,
  276.2305, 275.2447, 274.3293, 273.618, 273.0891, 272.3822, 271.8036, 
    271.5392, 269.9291, 264.6161, 265.006, 265.9821, 266.2925, 266.4375, 
    266.8127,
  275.9325, 275.2645, 274.7031, 273.5467, 272.6991, 272.2752, 271.6626, 
    270.9646, 270.4804, 266.213, 262.5095, 262.3091, 265.9637, 265.8518, 
    266.869,
  275.3578, 274.2258, 273.6504, 272.9764, 272.2437, 271.6275, 271.3204, 
    270.675, 268.5437, 262.2607, 264.8125, 263.7725, 263.7009, 266.0242, 
    266.8346,
  255.4913, 258.4057, 254.9804, 256.2148, 252.7913, 249.6349, 256.9388, 
    258.9534, 261.0703, 260.2957, 260.2229, 261.9276, 260.5851, 259.0136, 
    250.4834,
  269.3956, 268.6115, 268.3885, 259.5112, 248.369, 246.7717, 254.6773, 
    258.3635, 260.6009, 262.2577, 261.1853, 263.2956, 263.89, 259.396, 
    251.0966,
  273.8749, 273.2404, 273.3706, 270.585, 260.53, 239.7695, 252.648, 255.6781, 
    259.4355, 261.8608, 262.7415, 263.7034, 264.638, 262.953, 256.0867,
  274.4667, 273.8389, 273.4886, 273.3974, 272.7339, 264.2141, 247.0208, 
    253.0855, 257.242, 261.2064, 262.3086, 263.5543, 264.6618, 263.6299, 
    258.0237,
  274.7085, 274.0462, 273.6031, 273.4174, 273.1544, 272.4672, 267.5945, 
    248.3837, 244.4841, 256.056, 261.5176, 262.288, 264.4021, 264.0652, 
    261.124,
  275.0496, 274.4895, 273.8286, 273.4103, 273.0544, 272.6043, 271.5776, 
    267.4005, 260.6358, 257.6543, 257.631, 261.8921, 263.8722, 264.2943, 
    262.3595,
  275.7498, 275.1176, 274.1256, 273.4279, 272.9846, 272.3968, 272.0557, 
    270.8692, 267.7672, 263.5724, 261.6072, 261.6573, 263.817, 264.5846, 
    263.5871,
  276.2297, 275.2646, 274.3403, 273.6097, 273.0684, 272.3772, 271.7845, 
    271.5191, 269.7391, 265.1537, 261.8109, 261.5683, 262.4059, 263.8673, 
    264.6624,
  275.9505, 275.2633, 274.7433, 273.4926, 272.6369, 272.2443, 271.6693, 
    270.8749, 270.4726, 266.8119, 262.8987, 261.5976, 260.7947, 260.8566, 
    265.2458,
  275.3916, 274.2032, 273.4849, 272.8431, 272.1842, 271.5215, 271.1727, 
    270.7617, 269.0523, 265.3802, 266.1292, 263.2765, 260.2289, 259.8576, 
    264.7091,
  256.3999, 260.2122, 257.7697, 257.7547, 254.0236, 250.4558, 255.4427, 
    256.0873, 256.7245, 249.7368, 250.5279, 250.6935, 242.5144, 239.2376, 
    232.677,
  269.8129, 269.1241, 268.978, 261.6635, 246.9639, 247.5541, 256.0057, 
    257.4374, 258.0507, 254.9801, 251.8942, 254.7084, 250.269, 235.7221, 
    231.2793,
  273.863, 273.1712, 273.3541, 270.9569, 260.4221, 245.3307, 255.5185, 
    258.5309, 259.3324, 258.0014, 256.3949, 255.8771, 251.7251, 248.3212, 
    240.5035,
  274.4283, 273.8021, 273.453, 273.3936, 272.9745, 266.2814, 252.6779, 
    258.4551, 260.2054, 259.0168, 256.7413, 256.7397, 252.9282, 249.3103, 
    245.5215,
  274.6831, 274.0278, 273.5776, 273.4177, 273.1613, 272.5593, 269.0302, 
    253.895, 256.4208, 257.1531, 257.2198, 256.2703, 254.5514, 251.0252, 
    250.2293,
  275.0233, 274.4883, 273.8141, 273.4017, 273.0447, 272.5921, 271.7986, 
    268.7964, 263.2321, 260.7208, 256.8461, 256.8776, 256.1172, 252.4184, 
    251.4064,
  275.7327, 275.1438, 274.1218, 273.4101, 272.9698, 272.3792, 272.0386, 
    271.1184, 268.4152, 264.9672, 261.5956, 258.2572, 259.0488, 254.5694, 
    252.586,
  276.2053, 275.2741, 274.3437, 273.5945, 273.0442, 272.3465, 271.7448, 
    271.487, 269.6131, 265.7553, 262.4025, 259.8885, 260.5084, 257.2082, 
    254.388,
  275.9474, 275.2489, 274.7729, 273.414, 272.5318, 272.1577, 271.5998, 
    270.6494, 270.5451, 266.502, 262.8755, 261.3647, 258.9998, 260.5729, 
    256.0471,
  275.4208, 274.1606, 273.2431, 272.6469, 272.0695, 271.2407, 270.5667, 
    270.1634, 268.4155, 264.597, 265.6621, 262.9386, 259.9089, 258.4049, 
    260.6532,
  259.765, 261.2604, 254.5857, 258.3969, 256.2451, 254.3397, 258.1888, 
    257.3545, 252.6005, 240.3658, 238.1652, 240.4409, 237.0461, 240.0196, 
    238.3978,
  270.1086, 269.5253, 268.7261, 262.0442, 253.6621, 253.9248, 260.1737, 
    260.6653, 255.9677, 249.692, 242.4517, 247.2364, 247.8545, 236.8153, 
    238.1164,
  273.7943, 273.0945, 273.3292, 270.9405, 261.7723, 252.53, 260.6912, 
    262.3778, 259.8159, 254.4771, 251.2998, 249.7056, 248.9686, 248.9385, 
    246.263,
  274.3969, 273.7846, 273.4286, 273.361, 273.0148, 268.0624, 258.457, 
    261.3614, 260.0614, 256.6569, 252.387, 250.6059, 249.6981, 249.6912, 
    249.0191,
  274.6638, 274.0318, 273.5482, 273.405, 273.1481, 272.5963, 269.6706, 
    259.8327, 257.6483, 255.683, 253.904, 251.7775, 250.2782, 250.4131, 
    251.584,
  275.0144, 274.4876, 273.8128, 273.3782, 273.0254, 272.5782, 271.8358, 
    268.4071, 260.7597, 258.2345, 255.0059, 253.4947, 251.2734, 250.733, 
    251.9906,
  275.7466, 275.1935, 274.1363, 273.3914, 272.947, 272.3426, 271.9915, 
    270.9395, 267.0555, 262.5739, 259.4057, 255.106, 252.8938, 251.694, 
    252.325,
  276.1856, 275.2856, 274.3539, 273.5707, 272.9977, 272.2794, 271.6616, 
    271.4023, 268.799, 265.0356, 260.3691, 257.2482, 255.2074, 253.1591, 
    252.9545,
  275.9142, 275.2336, 274.7815, 273.3258, 272.3955, 272.004, 271.4297, 
    270.0335, 270.3896, 267.3374, 264.0775, 261.3741, 258.7661, 256.4271, 
    252.8472,
  275.3447, 274.1028, 273.0961, 272.4668, 271.938, 270.9314, 269.786, 
    269.8009, 267.3459, 262.9824, 265.3964, 263.382, 261.3765, 258.2724, 
    255.0062,
  257.1618, 260.1322, 255.7452, 259.7032, 258.47, 258.9236, 261.5641, 
    260.6756, 256.7481, 254.0261, 251.5913, 250.4711, 244.506, 246.055, 
    243.8724,
  269.0121, 268.8453, 268.7527, 262.9405, 257.0565, 258.1103, 262.215, 
    260.795, 258.5734, 259.2452, 255.0893, 254.9616, 250.9405, 243.2707, 
    243.7855,
  273.6679, 272.9898, 273.2352, 271.3289, 264.1736, 256.7648, 261.9223, 
    261.385, 260.028, 259.3921, 259.4135, 256.497, 252.3278, 252.5511, 250.963,
  274.3492, 273.729, 273.377, 273.3178, 273.0088, 268.2652, 255.3313, 
    260.2639, 260.6092, 259.5465, 259.1792, 257.1452, 253.1092, 253.3548, 
    252.7137,
  274.6209, 273.9923, 273.4908, 273.374, 273.1312, 272.5627, 269.5948, 
    262.0695, 261.4711, 258.2891, 258.7147, 256.7664, 254.414, 253.7513, 
    254.9216,
  274.9905, 274.4518, 273.7841, 273.3468, 273.0012, 272.5346, 271.7939, 
    268.4343, 262.7001, 263.283, 260.3106, 258.8006, 255.4392, 254.0135, 
    255.3004,
  275.717, 275.2013, 274.141, 273.3602, 272.9126, 272.2973, 271.9579, 
    270.928, 268.1529, 265.0478, 263.4847, 259.8573, 256.8588, 253.8092, 
    255.0793,
  276.1672, 275.2779, 274.3417, 273.5353, 272.9347, 272.2413, 271.6227, 
    271.2839, 268.8209, 265.9385, 263.1435, 260.5706, 258.4793, 255.4518, 
    255.0401,
  275.8836, 275.2153, 274.772, 273.2664, 272.3131, 271.9322, 271.3247, 
    269.6071, 269.7917, 266.2745, 262.7999, 261.1917, 259.2701, 258.4158, 
    254.4539,
  275.2849, 274.1093, 273.1631, 272.4637, 271.9373, 270.5397, 269.1557, 
    269.4005, 268.3123, 262.6289, 263.759, 262.5549, 260.0944, 261.4789, 
    254.432,
  258.5455, 260.0048, 257.9618, 258.3116, 256.456, 256.6202, 258.1718, 
    258.7594, 258.8764, 257.8605, 257.0996, 256.5689, 254.7032, 250.6881, 
    245.2284,
  267.7038, 267.4616, 268.3911, 262.4344, 255.7056, 256.3724, 259.9209, 
    260.1223, 260.2967, 259.7435, 258.3181, 258.9698, 257.8702, 249.021, 
    243.3015,
  273.5511, 272.9118, 273.1674, 271.3489, 264.4506, 255.1225, 261.4525, 
    261.3624, 261.2821, 260.7027, 260.6651, 260.2331, 258.9054, 256.1511, 
    248.1142,
  274.2895, 273.6789, 273.3191, 273.2758, 272.9517, 267.7283, 255.4467, 
    260.7475, 261.863, 261.7559, 261.4262, 261.16, 260.1241, 257.2688, 
    250.0364,
  274.5691, 273.9396, 273.4363, 273.3292, 273.1275, 272.5593, 269.6757, 
    258.5706, 261.4299, 260.9512, 262.0744, 261.3398, 259.8461, 257.4077, 
    252.7568,
  274.9619, 274.4014, 273.7498, 273.3208, 272.9897, 272.5237, 271.8645, 
    268.9284, 264.2185, 262.4013, 261.7179, 262.1866, 260.5555, 258.1072, 
    254.1449,
  275.6987, 275.1789, 274.1142, 273.3354, 272.9136, 272.3357, 272.019, 
    271.1593, 269.0353, 265.9861, 264.47, 263.4713, 261.579, 258.0096, 254.659,
  276.202, 275.251, 274.3218, 273.5177, 272.9291, 272.3442, 271.6817, 
    271.2896, 269.445, 266.5284, 264.8203, 263.8855, 262.3618, 258.6783, 
    253.9778,
  275.9111, 275.2562, 274.7729, 273.3042, 272.3711, 272.0134, 271.4651, 
    269.7815, 269.3014, 266.9438, 265.3837, 264.8672, 262.7949, 258.6864, 
    253.2752,
  275.2826, 274.1603, 273.2781, 272.5515, 272.0021, 270.9426, 269.1411, 
    268.913, 268.5025, 266.7578, 267.8131, 266.135, 263.4007, 259.2018, 
    253.2122,
  257.2408, 259.2545, 257.7996, 257.7455, 255.5109, 255.7518, 256.7701, 
    255.9015, 255.4782, 254.3918, 254.8634, 254.8193, 254.7322, 255.4051, 
    251.251,
  266.0839, 266.3321, 267.7519, 261.9953, 254.1998, 255.8492, 258.5388, 
    257.4074, 257.1887, 256.7464, 258.168, 259.5324, 259.1149, 256.3187, 
    250.3964,
  273.5185, 272.8719, 273.1445, 271.5328, 263.2332, 258.2949, 261.029, 
    260.1366, 260.0413, 260.6573, 261.8568, 262.5756, 261.75, 260.5084, 
    252.3062,
  274.2519, 273.6601, 273.3004, 273.2778, 272.9305, 267.4917, 256.3882, 
    261.8626, 263.8237, 264.4254, 265.7059, 265.1502, 264.2549, 262.3358, 
    252.3319,
  274.5382, 273.9296, 273.4319, 273.3287, 273.1759, 272.6329, 270.1475, 
    262.4747, 263.2605, 266.809, 267.9079, 265.5099, 264.9532, 262.7173, 
    252.6517,
  274.9944, 274.3956, 273.7484, 273.3305, 273.0586, 272.638, 272.133, 
    270.4645, 268.2478, 268.3206, 266.8927, 264.536, 264.8539, 262.8098, 
    251.8761,
  275.6975, 275.1724, 274.0934, 273.3505, 272.9596, 272.4801, 272.1797, 
    271.6091, 270.6943, 268.6085, 264.7259, 264.1185, 265.0194, 261.2762, 
    251.1647,
  276.2596, 275.2292, 274.3107, 273.5246, 272.9436, 272.4702, 271.7656, 
    271.4477, 269.9432, 266.0569, 262.5257, 265.0721, 265.3208, 259.3888, 
    249.682,
  275.9636, 275.2982, 274.7947, 273.3591, 272.434, 272.0595, 271.5509, 
    270.6318, 269.4323, 266.4699, 262.5348, 265.6458, 264.1146, 256.2823, 
    246.7563,
  275.2642, 274.2906, 273.4614, 272.6441, 272.0522, 271.161, 270.0121, 
    269.2784, 268.0649, 263.283, 266.812, 266.8287, 262.2794, 253.8378, 
    247.8748,
  255.2176, 257.2505, 255.0183, 254.3205, 251.4027, 252.1358, 253.9391, 
    252.3714, 251.745, 249.4204, 250.1017, 251.9785, 252.122, 255.0968, 
    257.0967,
  263.9683, 264.6019, 264.802, 259.4423, 250.2698, 254.5575, 256.5143, 
    253.899, 253.3924, 252.5178, 252.047, 255.0724, 256.6092, 257.9641, 
    257.9482,
  273.5501, 272.668, 273.0653, 271.2196, 259.7646, 250.7071, 259.0922, 
    256.4021, 255.0151, 254.6192, 255.327, 257.0214, 259.5905, 261.2477, 
    255.9668,
  274.2795, 273.7451, 273.381, 273.3422, 272.7873, 265.0733, 252.9165, 
    257.9372, 258.2026, 257.0858, 257.6763, 259.6982, 261.215, 262.2988, 
    253.8214,
  274.5779, 273.9961, 273.558, 273.3848, 273.213, 272.6584, 268.9424, 
    254.5214, 254.8228, 259.2424, 260.9365, 261.5836, 262.4968, 262.0359, 
    254.4305,
  275.1104, 274.4443, 273.7893, 273.3686, 273.1443, 272.7885, 272.3354, 
    269.2272, 261.0244, 259.6162, 260.6879, 262.4651, 263.5399, 260.584, 
    251.8785,
  275.7755, 275.2254, 274.1018, 273.3737, 273.0326, 272.6858, 272.3557, 
    271.7706, 269.5887, 263.5669, 262.39, 263.1355, 262.8331, 257.916, 251.451,
  276.3286, 275.2251, 274.3158, 273.5371, 272.9827, 272.6343, 271.9421, 
    271.6789, 270.1666, 265.8268, 263.8296, 263.6819, 262.7558, 255.6921, 
    249.2518,
  276.0054, 275.3188, 274.8228, 273.4669, 272.5674, 272.1721, 271.7829, 
    271.1333, 270.2589, 267.7849, 265.0698, 264.5752, 261.6354, 253.4746, 
    246.7913,
  275.2088, 274.307, 273.5334, 272.7013, 272.1494, 271.5162, 271.0345, 
    270.7685, 270.2915, 268.5139, 267.4306, 265.2571, 260.4205, 252.065, 
    248.028,
  257.5839, 259.4006, 255.1185, 254.4659, 250.3105, 250.8833, 253.7178, 
    250.7767, 249.3303, 243.7212, 244.0152, 246.4687, 243.1907, 244.7571, 
    240.8385,
  263.3293, 264.3548, 262.5408, 257.2349, 249.1114, 254.1671, 255.6238, 
    251.8483, 250.8727, 248.5475, 246.6271, 249.869, 249.5187, 244.2839, 
    238.0291,
  273.4686, 271.8941, 272.2135, 269.3552, 256.0433, 248.266, 258.1459, 
    254.0362, 252.0791, 250.3408, 250.5912, 250.1963, 250.3256, 250.8261, 
    245.7233,
  274.2995, 273.7518, 273.3999, 273.3279, 271.6852, 262.1872, 249.7182, 
    256.0474, 255.2117, 252.8592, 251.8204, 251.4317, 251.669, 253.0149, 
    250.4192,
  274.559, 273.9901, 273.5477, 273.3637, 273.1767, 272.4173, 267.4933, 
    250.194, 251.0845, 255.3389, 255.8887, 254.2383, 252.949, 254.6861, 
    253.2577,
  275.1367, 274.416, 273.7405, 273.3247, 273.1206, 272.7885, 272.3514, 
    268.842, 259.1638, 256.53, 256.3115, 256.4973, 254.9452, 255.1307, 
    253.0535,
  275.8188, 275.2771, 274.0569, 273.3147, 273.0007, 272.734, 272.4352, 
    271.9037, 270.0084, 262.5981, 259.3196, 257.3875, 256.1146, 255.7249, 
    252.7049,
  276.3302, 275.2278, 274.2772, 273.455, 272.9102, 272.6602, 272.0147, 
    271.8365, 270.3573, 264.2873, 261.5746, 259.5772, 257.1716, 255.4298, 
    251.9996,
  276.0013, 275.3087, 274.8162, 273.3798, 272.4781, 272.1068, 271.7961, 
    271.3369, 269.9147, 266.7169, 263.4074, 261.3708, 257.6349, 255.9137, 
    250.0415,
  275.1629, 274.271, 273.4054, 272.3837, 272.0106, 271.1245, 269.3828, 
    269.4795, 269.6342, 268.5923, 266.7255, 263.2189, 259.2096, 256.0294, 
    251.2969,
  257.9846, 260.2383, 257.4946, 256.8639, 252.9679, 253.5941, 256.3068, 
    251.6525, 250.5468, 244.3374, 243.1411, 243.8471, 238.097, 238.2909, 
    233.1817,
  263.0524, 264.2772, 262.2477, 257.7983, 251.4593, 256.1444, 256.3396, 
    252.2338, 251.3289, 249.2435, 246.2572, 248.9768, 247.508, 235.9785, 
    231.9022,
  273.139, 270.9613, 270.6339, 265.8912, 257.5349, 250.4442, 256.7338, 
    253.1002, 251.952, 250.6457, 251.6358, 249.5214, 247.4429, 246.0038, 
    238.8611,
  274.2741, 273.7215, 273.3588, 273.1169, 270.0858, 262.3517, 250.0483, 
    253.5003, 253.089, 251.4441, 251.06, 250.2439, 248.7409, 247.9058, 
    244.3198,
  274.5521, 273.9572, 273.5092, 273.3179, 273.0782, 271.7834, 267.068, 
    248.8077, 248.2294, 251.9908, 253.1551, 252.5349, 250.4329, 250.8084, 
    249.7747,
  275.1724, 274.3629, 273.6976, 273.2752, 273.0797, 272.7534, 272.2237, 
    267.9279, 258.7344, 255.0169, 254.9373, 254.7903, 251.9631, 251.3439, 
    249.3944,
  275.822, 275.3112, 274.0594, 273.2678, 272.9647, 272.7124, 272.4189, 
    271.8678, 269.5392, 261.1646, 257.4056, 255.2584, 253.2736, 252.0195, 
    250.1723,
  276.2973, 275.2265, 274.2392, 273.4134, 272.8535, 272.637, 272.001, 
    271.8039, 269.8463, 261.7938, 257.2992, 255.5166, 254.2171, 251.9277, 
    249.5964,
  276.0026, 275.3013, 274.8289, 273.3494, 272.445, 272.0746, 271.7484, 
    271.3371, 268.8109, 261.9336, 258.0487, 256.8496, 254.838, 252.235, 
    248.7702,
  275.1239, 274.254, 273.3891, 272.4114, 271.9694, 271.0024, 268.9856, 
    268.2802, 266.3049, 261.657, 262.5665, 259.1699, 256.281, 253.3983, 
    250.6303,
  257.3974, 259.3055, 257.3921, 256.4687, 252.0229, 251.6227, 254.4621, 
    249.3326, 249.6694, 242.1081, 239.8974, 242.3671, 238.8073, 239.1202, 
    235.7393,
  263.3317, 264.0448, 263.2162, 256.9912, 250.936, 253.2241, 252.6225, 
    250.0126, 249.5572, 248.5078, 243.8342, 247.9144, 247.6811, 235.7902, 
    232.946,
  271.9964, 269.7082, 269.2904, 262.5642, 257.5266, 247.2527, 251.8458, 
    250.6836, 250.5468, 249.8687, 250.7668, 247.9116, 246.6388, 245.8637, 
    238.5804,
  274.246, 273.6585, 273.2713, 272.1198, 268.8778, 260.9869, 246.0151, 
    250.3982, 250.8472, 249.7423, 249.1476, 247.7763, 246.9193, 246.4116, 
    244.3435,
  274.5376, 273.9007, 273.4701, 273.2679, 272.7692, 270.64, 266.1456, 
    246.3027, 242.8291, 246.5489, 250.3294, 249.9253, 248.3321, 248.7202, 
    249.1043,
  275.1648, 274.2884, 273.6589, 273.2292, 273.0457, 272.7052, 271.7821, 
    266.9371, 258.361, 254.0828, 251.0541, 252.6142, 249.7502, 248.9411, 
    247.9025,
  275.797, 275.2505, 274.0341, 273.2294, 272.9352, 272.6911, 272.3976, 
    271.6802, 268.8371, 261.4758, 256.8692, 253.6195, 251.0448, 249.7973, 
    248.1467,
  276.3008, 275.2379, 274.21, 273.404, 272.832, 272.6361, 272.0127, 271.7712, 
    269.3201, 260.7247, 255.89, 253.2117, 252.0289, 249.7044, 247.701,
  276.0572, 275.3099, 274.8426, 273.3829, 272.4914, 272.0625, 271.75, 
    271.4413, 268.8755, 259.7021, 255.8278, 254.2458, 252.8054, 250.1986, 
    247.3439,
  275.1562, 274.2844, 273.4535, 272.5233, 272.043, 271.2617, 269.6443, 
    268.6699, 263.6026, 257.913, 259.5656, 256.199, 253.541, 251.5326, 
    249.6402,
  257.4521, 258.2274, 255.5104, 254.7123, 250.2363, 248.9707, 251.9292, 
    248.8988, 251.291, 244.469, 242.8387, 245.1734, 241.8293, 240.945, 
    237.0543,
  264.8885, 262.763, 262.1396, 254.8195, 249.2115, 248.2616, 250.1127, 
    249.3316, 249.5894, 251.0685, 245.8151, 249.1857, 250.0144, 239.0983, 
    236.0677,
  271.2649, 267.9334, 267.567, 259.0616, 256.8001, 243.297, 249.1681, 
    250.2745, 250.4766, 250.1766, 250.7491, 249.2624, 249.3917, 248.9642, 
    242.5973,
  274.1644, 273.4067, 272.972, 269.957, 267.7047, 259.6415, 243.9872, 
    249.0561, 250.2373, 249.3274, 249.0091, 248.7189, 249.0112, 249.4817, 
    248.1353,
  274.5092, 273.8067, 273.3994, 273.1853, 272.2384, 269.596, 265.9099, 
    243.4655, 239.4586, 245.3037, 249.818, 250.3722, 249.7821, 250.4848, 
    251.9268,
  275.0787, 274.214, 273.6041, 273.1562, 272.9766, 272.5529, 271.0225, 
    265.8235, 257.0087, 253.0668, 249.454, 252.0919, 250.5391, 250.4632, 
    251.2423,
  275.713, 275.0955, 273.9364, 273.1538, 272.8747, 272.6291, 272.3139, 
    271.134, 267.6054, 260.1685, 255.0851, 252.7498, 251.4361, 250.8238, 
    250.4841,
  276.2202, 275.1645, 274.1198, 273.3406, 272.765, 272.5799, 271.9516, 
    271.6836, 267.1855, 258.6861, 254.3005, 252.9212, 252.3999, 250.5809, 
    250.7149,
  276.0113, 275.2356, 274.7756, 273.3801, 272.4804, 271.9947, 271.692, 
    271.0983, 267.2644, 256.8272, 254.8345, 254.4334, 253.9112, 251.8138, 
    250.9388,
  275.1264, 274.2669, 273.5304, 272.5751, 272.0034, 271.0981, 269.2435, 
    267.8434, 259.5915, 253.5431, 257.7595, 255.6172, 254.4427, 253.6789, 
    252.1361,
  256.2746, 257.5533, 254.0743, 254.9568, 250.8271, 249.1298, 251.8147, 
    250.1349, 252.3763, 244.7259, 241.9314, 244.5828, 242.2917, 242.1575, 
    238.6417,
  265.054, 262.0869, 261.3595, 255.3523, 248.651, 247.1106, 250.8935, 
    250.9965, 251.1021, 253.0903, 247.8186, 251.8668, 253.4694, 243.2242, 
    241.2866,
  271.3152, 266.9032, 267.0373, 259.5907, 257.9151, 241.4212, 249.6796, 
    251.8373, 252.9228, 253.3464, 253.8209, 253.7143, 254.4439, 254.2383, 
    248.552,
  274.0993, 273.1487, 272.6738, 269.1543, 268.3638, 260.375, 240.7971, 
    250.9343, 253.2367, 253.4199, 253.562, 254.1458, 254.7355, 255.0873, 
    253.5862,
  274.4668, 273.7447, 273.3539, 273.1531, 272.321, 269.9882, 266.3231, 
    243.634, 245.4554, 252.5764, 254.3455, 255.4681, 255.229, 255.9684, 
    256.5717,
  274.9944, 274.1907, 273.5665, 273.1268, 272.9574, 272.4264, 270.6579, 
    265.8049, 258.7833, 257.02, 253.8152, 255.7851, 256.42, 256.5999, 257.9458,
  275.6849, 275.0205, 273.8943, 273.1256, 272.8561, 272.6041, 272.2311, 
    270.769, 266.8594, 260.3363, 256.8398, 256.088, 256.3405, 256.7915, 
    257.7694,
  276.1913, 275.1321, 274.0812, 273.3196, 272.7349, 272.5338, 271.8901, 
    271.5464, 265.468, 259.079, 256.8101, 255.6787, 255.7464, 255.9022, 
    257.4897,
  275.9829, 275.2013, 274.7446, 273.3934, 272.4686, 271.9475, 271.6088, 
    270.394, 266.1137, 258.4798, 257.7256, 256.8001, 255.1494, 255.1968, 
    256.5917,
  275.1001, 274.2632, 273.6003, 272.5879, 271.9432, 270.8187, 268.7047, 
    267.6531, 259.6153, 255.7826, 259.0283, 256.8707, 254.954, 254.2061, 
    255.8466,
  254.1161, 257.9501, 253.0348, 254.8094, 250.5652, 247.839, 250.2364, 
    249.129, 250.9357, 242.0159, 240.1481, 243.6634, 242.5377, 244.2217, 
    241.0517,
  265.1042, 262.2183, 260.5763, 255.6806, 248.6924, 246.5492, 251.4139, 
    251.1435, 250.7698, 251.0127, 245.2794, 249.9681, 251.3574, 241.6057, 
    239.0264,
  271.7818, 267.5018, 267.8704, 260.4503, 258.1057, 240.187, 251.2689, 
    254.0592, 253.8924, 253.5131, 252.8562, 251.8599, 251.6858, 251.1175, 
    245.2935,
  274.0724, 273.2577, 272.7676, 269.7541, 268.8676, 262.2003, 245.613, 
    252.815, 255.0368, 254.1364, 252.8099, 252.19, 251.8052, 252.5608, 
    250.1825,
  274.4107, 273.7129, 273.3458, 273.1797, 272.7254, 270.4934, 267.4274, 
    249.3441, 249.0307, 251.8792, 253.8612, 253.1291, 253.183, 255.3174, 
    253.3496,
  274.9336, 274.1894, 273.5632, 273.1249, 272.9749, 272.4213, 270.5567, 
    266.1417, 260.6613, 257.541, 254.3233, 256.1063, 256.3432, 255.3706, 
    253.6412,
  275.6716, 275.0376, 273.888, 273.1171, 272.8534, 272.5955, 272.1342, 
    270.6456, 266.2964, 262.1576, 260.3064, 258.0371, 257.35, 255.5912, 
    254.1984,
  276.1874, 275.1228, 274.0721, 273.3124, 272.6979, 272.5018, 271.8423, 
    271.1288, 264.438, 261.2134, 260.152, 259.9408, 259.1609, 259.412, 260.107,
  275.9585, 275.1785, 274.7184, 273.3971, 272.4479, 271.9045, 271.4261, 
    269.5452, 265.0253, 260.9955, 260.4804, 260.2276, 259.2066, 257.6466, 
    256.9321,
  275.0826, 274.2427, 273.6453, 272.5838, 271.9053, 270.2486, 268.4061, 
    267.0065, 262.0448, 259.5826, 260.3714, 257.7854, 257.1207, 256.1399, 
    257.0607,
  253.1099, 256.1921, 252.171, 254.0396, 250.2621, 249.2637, 252.8562, 
    253.4417, 255.8459, 252.224, 251.0199, 251.1218, 247.0618, 247.0502, 
    242.6216,
  263.3271, 260.6336, 258.9454, 255.0649, 248.5797, 247.366, 252.4522, 
    253.5781, 254.0506, 256.0924, 252.3246, 254.2985, 254.4421, 245.9573, 
    242.1832,
  271.4276, 266.4766, 266.817, 259.2923, 256.5161, 241.8642, 251.0937, 
    253.6473, 254.463, 255.0117, 255.2888, 254.2202, 254.3996, 252.785, 
    247.402,
  274.0431, 273.1837, 272.5995, 268.3494, 267.3824, 259.7665, 243.5015, 
    250.6545, 253.5056, 253.7616, 253.6221, 253.3419, 253.5508, 252.6574, 
    250.6391,
  274.3841, 273.6919, 273.3, 273.1218, 272.6639, 269.6481, 266.2161, 245.497, 
    243.5335, 250.6455, 254.1523, 254.4897, 254.506, 254.2551, 253.1869,
  274.9441, 274.2058, 273.5624, 273.0866, 272.9543, 272.2946, 269.9509, 
    264.8732, 259.0874, 257.1989, 253.9452, 256.0368, 255.8408, 254.6507, 
    254.0274,
  275.7346, 275.1613, 273.924, 273.109, 272.8218, 272.5489, 271.9723, 
    269.9324, 265.1796, 260.0078, 258.4264, 256.6062, 255.9302, 253.8126, 
    253.6113,
  276.249, 275.171, 274.099, 273.2876, 272.651, 272.4335, 271.7762, 270.9297, 
    263.5533, 259.6612, 258.3961, 257.4798, 257.0883, 255.6969, 254.6959,
  275.9928, 275.2042, 274.7374, 273.3633, 272.4213, 271.8487, 271.3405, 
    269.4715, 263.724, 260.2927, 259.5827, 259.312, 257.7398, 254.7487, 
    253.6403,
  275.0726, 274.2224, 273.6266, 272.4986, 271.8418, 270.0565, 268.9704, 
    267.7858, 262.6658, 260.8493, 261.3207, 259.0689, 255.3562, 253.4216, 
    254.1455,
  251.4681, 255.7788, 250.8235, 254.8812, 249.7813, 250.9408, 256.4041, 
    255.3145, 255.069, 248.6559, 248.187, 248.157, 244.3119, 242.4046, 
    238.4978,
  260.8959, 260.1083, 259.3758, 255.5512, 247.1116, 249.34, 256.1734, 
    256.0118, 255.1262, 254.5261, 247.6773, 250.6775, 250.2852, 241.0845, 
    240.1223,
  270.4635, 266.5772, 267.1268, 260.5518, 258.6562, 248.7139, 255.0821, 
    256.8192, 256.1246, 254.4206, 253.0108, 251.3809, 250.8321, 250.3852, 
    245.5341,
  273.9788, 273.1358, 272.6374, 268.8552, 267.6557, 261.8646, 249.5057, 
    253.8112, 253.0882, 252.6526, 251.3931, 250.2177, 249.8697, 249.6259, 
    249.7967,
  274.3799, 273.6537, 273.2578, 273.0742, 272.5873, 269.4557, 266.6178, 
    247.6555, 245.8061, 249.2591, 251.0592, 250.2711, 250.1853, 250.8262, 
    251.2147,
  274.9768, 274.1867, 273.5465, 273.0521, 272.9328, 272.1469, 269.5549, 
    264.6026, 259.8364, 257.2274, 251.7672, 251.4923, 250.9796, 251.0322, 
    251.4568,
  275.7752, 275.2395, 273.9755, 273.0966, 272.7901, 272.4908, 271.8429, 
    268.9964, 263.7325, 257.7569, 254.8433, 252.6791, 251.7225, 250.9346, 
    251.3348,
  276.2927, 275.2279, 274.1313, 273.246, 272.5981, 272.3619, 271.7059, 
    270.7208, 262.2509, 257.2063, 254.6604, 253.3227, 252.1593, 251.1425, 
    251.4176,
  276.0703, 275.24, 274.7689, 273.3117, 272.3831, 271.7628, 271.2152, 
    268.7807, 261.1973, 256.8266, 255.0476, 254.0198, 252.1987, 251.2677, 
    251.8877,
  275.1141, 274.2129, 273.5556, 272.3948, 271.7679, 270.033, 269.0065, 
    266.9785, 259.6298, 258.101, 257.166, 254.5811, 252.6616, 252.0983, 
    252.671,
  248.9198, 255.3319, 251.2292, 255.9121, 253.6618, 253.3477, 254.9478, 
    253.1472, 254.1902, 248.2948, 245.7835, 246.2175, 243.3771, 241.5579, 
    237.0471,
  259.5123, 259.3848, 258.7333, 256.0197, 249.0624, 250.4051, 254.1403, 
    253.078, 252.772, 253.1079, 248.7374, 250.1749, 250.8346, 240.4587, 
    238.0164,
  269.5685, 267.1025, 267.2154, 261.3081, 256.1218, 244.5208, 251.4761, 
    252.6851, 253.1365, 253.5631, 253, 250.5443, 250.566, 250.8917, 244.8284,
  273.8984, 273.1169, 272.7786, 269.5369, 267.7686, 260.3098, 243.9233, 
    249.3667, 252.0858, 252.356, 251.1642, 248.6685, 248.8862, 248.7862, 
    249.4867,
  274.3961, 273.5835, 273.192, 273.0051, 272.6305, 269.5181, 266.1531, 
    243.3089, 241.7229, 247.7632, 249.813, 248.5959, 248.8314, 249.764, 
    250.909,
  275.0541, 274.1627, 273.5388, 273.0184, 272.9129, 272.1521, 269.5251, 
    263.7668, 257.4698, 255.6619, 250.0385, 249.3747, 249.2716, 249.7533, 
    250.5287,
  275.8438, 275.2972, 274.0477, 273.077, 272.7588, 272.4412, 271.8243, 
    267.9873, 261.6664, 255.2629, 252.6296, 250.5163, 249.9587, 249.7338, 
    250.4733,
  276.3104, 275.3196, 274.1892, 273.2077, 272.5406, 272.3162, 271.6502, 
    270.795, 261.209, 254.0663, 251.8837, 250.9335, 250.3645, 249.6588, 
    250.1877,
  276.1419, 275.2851, 274.7917, 273.2291, 272.3141, 271.6714, 271.1694, 
    268.8577, 259.1045, 253.0279, 251.3775, 251.2904, 250.5268, 249.8486, 
    250.7094,
  275.152, 274.1856, 273.3727, 272.2148, 271.5926, 270.041, 269.1037, 
    266.9337, 258.2263, 253.8731, 254.4631, 252.2057, 251.2635, 251.1693, 
    251.5549,
  250.9916, 254.9588, 251.2384, 256.8748, 253.5828, 251.6057, 252.3947, 
    249.8441, 249.0851, 240.8763, 239.7119, 244.9798, 244.341, 239.6141, 
    233.8912,
  258.253, 258.3376, 258.4221, 257.1427, 249.6232, 247.341, 251.1536, 
    250.7276, 248.7654, 248.5828, 243.0863, 249.2433, 252.0812, 237.962, 
    234.0253,
  268.7014, 266.9093, 266.3731, 261.1729, 257.4292, 243.1647, 248.0502, 
    250.2701, 249.6869, 249.5782, 249.2242, 250.0524, 251.8389, 250.3592, 
    243.3525,
  273.8438, 273.0887, 272.8058, 269.9133, 267.6759, 261.1727, 242.5165, 
    248.2352, 251.0977, 249.7037, 248.0465, 247.7475, 249.1666, 250.4836, 
    248.0103,
  274.3906, 273.5419, 273.1373, 272.9281, 272.6264, 269.9988, 265.5868, 
    243.4818, 241.9013, 248.7223, 248.0305, 247.5223, 248.4883, 249.8371, 
    249.9851,
  275.0467, 274.127, 273.5189, 272.981, 272.8809, 272.1895, 269.6862, 
    263.2824, 257.5309, 256.4718, 251.145, 248.8263, 248.4202, 248.6481, 
    248.9314,
  275.8218, 275.232, 274.0206, 273.0493, 272.7299, 272.3868, 271.8955, 
    267.9938, 263.0237, 257.4594, 253.6852, 249.7434, 248.9394, 248.4084, 
    248.7997,
  276.2523, 275.2907, 274.1722, 273.1698, 272.4984, 272.2493, 271.5903, 
    271.002, 263.7486, 256.3093, 252.82, 250.3744, 249.1239, 248.1884, 248.328,
  276.1106, 275.265, 274.744, 273.1786, 272.2488, 271.5043, 271.1202, 
    269.2352, 260.7984, 254.7581, 252.7836, 251.3666, 249.6111, 248.3539, 
    248.6759,
  275.1497, 274.1418, 273.2144, 272.0735, 271.3949, 269.5202, 268.821, 
    267.3398, 259.9612, 256.3078, 256.308, 252.3901, 250.4729, 249.9325, 
    249.4377,
  256.2216, 255.8438, 253.5358, 254.5523, 252.7565, 249.1104, 248.1023, 
    247.9798, 247.9537, 239.2133, 238.2341, 242.1687, 239.3678, 237.4415, 
    231.7962,
  259.3495, 258.6533, 257.4804, 256.1133, 251.515, 246.8957, 247.9223, 
    247.7342, 246.838, 246.755, 242.0114, 248.6534, 249.663, 235.6185, 232.252,
  267.0787, 266.2352, 263.4526, 259.435, 255.3161, 242.5214, 246.9189, 
    247.5124, 247.108, 248.2099, 248.9582, 250.0945, 251.0307, 248.8377, 
    242.1992,
  273.8237, 272.7597, 272.2201, 268.1805, 264.5037, 256.4087, 241.7403, 
    245.5747, 246.8666, 247.1748, 247.2468, 248.5026, 251.2439, 249.7354, 
    246.6447,
  274.3411, 273.5347, 273.1399, 272.9276, 272.4421, 268.2218, 263.3477, 
    242.3742, 239.8401, 245.0989, 247.0635, 248.0223, 250.5528, 251.7527, 
    249.1626,
  274.9766, 274.0958, 273.492, 272.9774, 272.8546, 272.0922, 269.0747, 
    262.6012, 256.4459, 255.3415, 251.1415, 248.9799, 248.9644, 249.9489, 
    248.7636,
  275.7298, 275.0738, 273.9169, 273.0197, 272.728, 272.371, 271.9065, 
    267.516, 263.7223, 258.4695, 253.9239, 249.6044, 249.0255, 249.2159, 
    248.6393,
  276.1982, 275.1733, 274.084, 273.1797, 272.5744, 272.2977, 271.5504, 
    270.9574, 265.6963, 260.7762, 254.7693, 250.578, 249.0831, 248.088, 
    247.7999,
  276.0409, 275.2072, 274.6552, 273.3866, 272.3855, 271.4953, 270.8924, 
    268.8925, 262.5913, 261.1925, 259.0763, 254.776, 250.3772, 247.9753, 
    247.1773,
  275.12, 274.1942, 273.5717, 272.4172, 271.5469, 269.3432, 268.1049, 
    266.0171, 261.1167, 260.644, 262.4797, 259.1064, 255.1835, 251.3601, 
    248.3136,
  264.2712, 262.4092, 258.0812, 253.6475, 249.5433, 246.9764, 247.9901, 
    248.125, 248.66, 239.6874, 238.0395, 240.2962, 237.0039, 236.7011, 
    230.6905,
  265.7346, 264.0482, 260.6443, 254.4781, 248.5598, 245.5392, 246.9679, 
    247.5795, 247.5703, 246.7787, 241.8177, 246.7174, 246.5787, 234.5442, 
    231.2742,
  270.0378, 268.4935, 263.5876, 257.2388, 253.2885, 242.2089, 245.8106, 
    247.2767, 247.515, 248.4281, 248.4841, 248.4159, 248.3168, 246.7545, 
    241.2826,
  273.8704, 273.061, 271.52, 265.7963, 260.7081, 255.4077, 241.7094, 
    244.6169, 246.5392, 247.7237, 247.5567, 248.0138, 248.2952, 247.4673, 
    245.0144,
  274.325, 273.5225, 273.128, 272.7355, 270.9522, 265.9546, 262.3366, 
    242.0899, 239.7778, 244.5512, 247.4326, 248.5104, 248.5712, 248.6752, 
    247.6759,
  274.9778, 274.0892, 273.4594, 272.9564, 272.8117, 271.8737, 267.7545, 
    261.1922, 255.3836, 254.8468, 250.798, 249.7592, 248.8509, 248.7054, 
    247.486,
  275.764, 275.0428, 273.8655, 272.9903, 272.7156, 272.3963, 271.7026, 
    265.2187, 260.4065, 256.8994, 253.6048, 249.8972, 249.3965, 248.6379, 
    247.8431,
  276.2041, 275.1299, 274.0563, 273.1906, 272.6376, 272.4221, 271.6294, 
    270.4015, 262.9222, 255.6949, 252.5627, 250.2223, 249.5748, 248.1504, 
    247.6404,
  276.0355, 275.1832, 274.6097, 273.5705, 272.618, 271.6865, 271.0397, 
    268.9676, 259.5729, 255.0842, 253.29, 251.299, 249.767, 247.9862, 246.6318,
  275.1302, 274.1876, 273.7263, 272.8222, 271.9072, 269.9682, 267.9725, 
    264.0702, 257.8773, 255.9524, 258.1293, 254.9928, 252.1638, 249.5937, 
    247.5457,
  264.8376, 266.6855, 266.2374, 261.1334, 254.4167, 249.4921, 250.007, 
    248.7418, 247.2183, 238.2913, 237.6193, 239.0633, 235.6888, 235.6104, 
    231.1857,
  266.8638, 268.3983, 267.4174, 260.4619, 250.9598, 247.8916, 248.0402, 
    247.519, 246.1313, 244.8852, 240.7733, 244.7794, 244.346, 233.2941, 
    230.4253,
  271.0384, 269.8776, 268.2294, 261.2747, 254.8114, 243.3681, 246.1768, 
    247.1348, 246.7383, 246.3795, 245.9865, 245.6228, 245.4221, 244.1422, 
    239.0371,
  273.8917, 273.3023, 272.2925, 266.5638, 261.6694, 256.4609, 241.696, 
    244.52, 245.8308, 246.1315, 245.0354, 245.042, 244.8213, 244.5234, 
    243.1342,
  274.341, 273.5213, 273.1414, 272.4619, 268.6402, 264.8018, 261.6974, 
    240.8943, 237.8516, 242.8212, 244.7879, 245.4069, 245.3941, 245.5959, 
    245.6923,
  275.0287, 274.1216, 273.4573, 272.9691, 272.7603, 271.4397, 267.0188, 
    260.2139, 254.317, 254.306, 248.7426, 247.0641, 246.176, 245.8655, 
    245.4709,
  275.8333, 275.1405, 273.8792, 273.008, 272.7065, 272.395, 271.2053, 
    263.0855, 257.8555, 255.4659, 251.7533, 247.7025, 247.0538, 246.1781, 
    246.0484,
  276.2359, 275.1218, 274.0517, 273.2187, 272.6535, 272.4647, 271.7157, 
    269.3546, 260.3687, 253.4185, 250.428, 248.2521, 247.5569, 246.5829, 
    246.2887,
  276.0851, 275.226, 274.6212, 273.5784, 272.7204, 271.7506, 271.4021, 
    269.4075, 257.3737, 251.9681, 250.1451, 249.0115, 248.2686, 246.9071, 
    245.9997,
  275.1794, 274.1555, 273.6474, 272.9306, 272.0193, 270.6844, 268.1062, 
    262.9472, 254.0783, 251.9884, 254.1052, 250.5337, 249.5056, 248.4081, 
    246.6353,
  263.8649, 264.5756, 264.1212, 264.0512, 260.8704, 257.2018, 255.6522, 
    252.511, 248.7819, 239.5549, 238.5541, 239.5162, 235.3382, 235.1175, 
    231.3656,
  265.1851, 265.245, 264.8302, 264.1109, 259.8521, 254.9155, 252.9822, 
    250.1265, 247.3721, 245.4428, 241.5154, 245.0121, 244.7108, 232.2352, 
    229.1841,
  271.2666, 269.7313, 267.5161, 265.3408, 261.975, 250.8986, 249.4168, 
    248.7629, 246.7803, 246.3294, 246.107, 245.8245, 245.3283, 243.9384, 
    238.1039,
  273.867, 273.36, 272.557, 269.4612, 266.1053, 260.0972, 245.8576, 244.843, 
    245.5413, 245.392, 245.5036, 244.9079, 244.2091, 243.6959, 241.9912,
  274.4067, 273.5294, 273.1265, 272.7211, 269.0633, 265.5799, 262.9719, 
    242.564, 238.9225, 242.4482, 244.6405, 244.8008, 244.2866, 244.1396, 
    244.1299,
  275.1111, 274.1438, 273.4511, 272.9801, 272.7119, 271.0701, 267.4582, 
    261.1193, 254.5889, 253.799, 248.2499, 246.0312, 245.0869, 243.6823, 
    243.3546,
  275.9305, 275.2438, 273.9271, 273.0054, 272.7346, 272.4095, 271.037, 
    263.08, 256.7528, 255.4013, 251.3748, 246.533, 245.5281, 243.746, 243.1948,
  276.2755, 275.1885, 274.0504, 273.1809, 272.6893, 272.5022, 271.7405, 
    268.6928, 258.1267, 251.5373, 248.6592, 246.5094, 245.4748, 243.7554, 
    243.219,
  276.1713, 275.3016, 274.6462, 273.5558, 272.7823, 271.7881, 271.5359, 
    269.2523, 254.7341, 249.272, 247.3541, 246.2238, 245.4281, 243.993, 
    243.0918,
  275.277, 274.1682, 273.5616, 272.9324, 272.062, 271.104, 268.588, 260.9873, 
    250.4657, 248.7352, 250.6692, 247.0278, 246.6107, 245.5358, 244.4229,
  264.9955, 265.2259, 264.1137, 263.3201, 261.7794, 260.7383, 261.0329, 
    258.404, 255.7749, 248.2613, 244.2262, 243.0608, 236.9497, 236.0605, 
    235.226,
  267.2143, 266.0282, 264.9137, 263.5848, 261.4948, 260.1719, 259.2984, 
    257.0688, 254.0924, 250.9866, 246.2688, 247.2402, 245.7505, 233.046, 
    232.3322,
  271.8588, 269.9702, 267.8288, 264.2735, 262.334, 256.4315, 256.3895, 
    255.7337, 252.3498, 250.6424, 249.1399, 248.1996, 246.7401, 244.6214, 
    238.5482,
  273.8374, 273.3841, 272.6489, 269.5504, 266.206, 263.713, 251.0067, 
    249.4351, 249.3361, 249.0392, 248.0875, 246.4161, 245.5191, 244.1981, 
    241.7343,
  274.4969, 273.504, 273.0948, 272.8323, 268.6993, 267.2382, 264.4823, 
    245.3517, 242.3009, 245.5678, 246.6161, 245.9769, 245.2654, 244.806, 
    244.7643,
  275.2175, 274.1355, 273.4511, 272.9596, 272.6024, 270.835, 267.8789, 
    262.4724, 257.5152, 255.7381, 250.5105, 247.261, 245.8129, 244.071, 
    243.4138,
  276.0266, 275.3433, 274.004, 272.9834, 272.7181, 272.384, 270.8119, 
    264.898, 260.9588, 258.3773, 253.8029, 247.5505, 245.8867, 243.5254, 
    242.8596,
  276.3087, 275.3611, 274.0876, 273.1459, 272.6923, 272.5045, 271.7059, 
    268.8931, 260.0093, 252.8994, 250.0553, 247.1663, 245.4886, 243.119, 
    242.2569,
  276.2038, 275.3493, 274.6462, 273.5443, 272.7915, 271.7788, 271.5334, 
    269.0077, 255.1479, 249.8213, 247.6924, 246.5629, 244.8571, 243.0098, 
    241.8183,
  275.2642, 274.2666, 273.7536, 272.9352, 272.0454, 271.2556, 268.954, 
    260.0207, 249.9538, 248.5914, 250.5425, 247.1413, 245.6896, 244.2763, 
    243.1654,
  263.5825, 264.3999, 262.9669, 262.4062, 260.4833, 259.3706, 260.1083, 
    259.0638, 258.4248, 253.3089, 252.4293, 252.5663, 248.2325, 246.5484, 
    243.7915,
  267.3286, 264.9192, 263.6924, 262.0604, 259.7216, 259.0504, 259.2169, 
    258.1284, 257.5, 257.1385, 254.9183, 255.8457, 253.0741, 243.071, 240.6434,
  272.2733, 270.6076, 268.5581, 265.2131, 262.462, 257.4176, 257.9413, 
    257.3614, 255.7427, 255.8909, 256.1127, 254.7558, 252.1089, 248.9265, 
    244.0969,
  273.8353, 273.4185, 272.8547, 270.8642, 267.5674, 264.331, 253.5382, 
    252.8448, 252.295, 253.3237, 253.554, 252.5275, 250.5606, 247.6469, 
    244.6033,
  274.5991, 273.4813, 273.0566, 272.8658, 270.8212, 269.2035, 266.1864, 
    253.6379, 250.9117, 250.0441, 251.7993, 251.5095, 249.3261, 247.2984, 
    245.2198,
  275.3148, 274.1438, 273.4411, 272.9208, 272.7094, 271.5736, 268.5692, 
    264.4291, 259.9037, 259.0979, 254.2649, 251.0666, 248.7276, 245.9033, 
    243.8956,
  276.0823, 275.3646, 274.0669, 272.9529, 272.7083, 272.3662, 270.7464, 
    264.5563, 260.6283, 260.9341, 257.0399, 250.9648, 247.8986, 244.9726, 
    243.1361,
  276.2759, 275.3832, 274.0843, 273.0824, 272.6681, 272.4615, 271.5698, 
    267.9058, 259.1176, 255.0396, 252.9162, 249.1947, 247.1914, 243.8483, 
    242.6329,
  276.1533, 275.31, 274.6003, 273.4838, 272.7516, 271.6961, 271.2931, 
    267.6764, 254.9886, 250.8088, 249.3108, 247.9535, 245.6317, 243.4237, 
    242.5557,
  275.1654, 274.2593, 273.7552, 272.8694, 271.9716, 271.1754, 269.0087, 
    260.5956, 250.3057, 248.6398, 250.6495, 247.3095, 246.092, 244.2492, 
    244.4112,
  263.8031, 265.2842, 263.5369, 262.303, 259.5475, 256.9249, 257.624, 
    255.3058, 253.4595, 246.4843, 246.8529, 249.7597, 247.2273, 246.686, 
    244.7404,
  269.4368, 268.1623, 266.9151, 264.9341, 261.2884, 259.7237, 257.8944, 
    255.0329, 253.4016, 252.0505, 250.7067, 253.717, 253.0289, 245.5247, 
    244.2104,
  272.3623, 271.0725, 269.4193, 267.8227, 264.6574, 258.9158, 259.0899, 
    257.5557, 255.0888, 253.8287, 254.2215, 254.4885, 254.1036, 253.0023, 
    248.3423,
  273.8203, 273.4078, 272.9094, 271.4865, 268.7131, 265.3005, 257.2347, 
    255.3661, 254.8028, 254.869, 254.3204, 254.0276, 253.3793, 252.6512, 
    249.8041,
  274.624, 273.4536, 273.0197, 272.795, 271.4158, 270.0712, 266.4003, 
    254.8598, 252.0357, 254.8757, 254.8812, 254.593, 253.6512, 252.4273, 
    250.8394,
  275.2762, 274.093, 273.4393, 272.8941, 272.6173, 271.9505, 269.0592, 
    266.264, 263.4205, 262.8775, 258.4525, 256.1432, 254.4029, 251.202, 
    248.5834,
  276.009, 275.2168, 273.9904, 272.9178, 272.6826, 272.3512, 270.8353, 
    265.511, 263.3983, 264.068, 260.5847, 256.5061, 253.8201, 249.9697, 
    247.874,
  276.2372, 275.3018, 274.0043, 273.0042, 272.6408, 272.4206, 271.3439, 
    267.3368, 259.9227, 258.4836, 256.8915, 254.6512, 252.3237, 248.5743, 
    246.6039,
  276.1558, 275.3061, 274.5764, 273.425, 272.6686, 271.5267, 270.7758, 
    265.9448, 254.701, 253.6314, 253.486, 252.5813, 249.8839, 246.7316, 
    244.3254,
  275.1599, 274.2403, 273.6919, 272.7567, 271.8, 270.6489, 267.9908, 260.307, 
    250.7682, 249.219, 252.7812, 250.5016, 248.8779, 246.6514, 244.8548,
  267.1424, 267.9669, 265.3858, 266.6588, 264.9429, 263.1674, 263.1456, 
    261.1554, 258.0447, 249.1245, 248.8381, 252.0096, 249.1107, 248.789, 
    246.9653,
  267.4896, 265.251, 263.6689, 265.7778, 264.2351, 263.9926, 263.2695, 
    261.5181, 259.613, 254.9712, 253.2319, 255.0115, 253.2441, 245.5741, 
    245.156,
  272.221, 270.7922, 267.0637, 263.6399, 263.7311, 260.9674, 261.9909, 
    261.8249, 260.479, 258.3517, 256.8728, 255.6349, 253.0218, 251.2462, 
    247.6648,
  273.7779, 273.3471, 272.8748, 270.1732, 265.0824, 263.5508, 257.3059, 
    257.479, 257.1919, 256.7188, 255.3191, 253.265, 252.8122, 251.8867, 
    249.4706,
  274.6696, 273.4064, 272.9418, 272.7224, 270.0966, 268.7296, 265.1359, 
    249.7842, 253.9555, 254.853, 256.1656, 254.9329, 253.3023, 252.5966, 
    251.3092,
  275.3244, 274.0476, 273.3791, 272.838, 272.5544, 271.637, 268.0198, 
    264.3112, 260.7745, 261.9682, 258.6468, 256.4109, 254.6471, 252.4419, 
    250.721,
  276.0431, 275.1699, 273.946, 272.8661, 272.6189, 272.2878, 270.6479, 
    263.8739, 261.0585, 262.6249, 260.8775, 256.6653, 254.6033, 252.4144, 
    250.4467,
  276.2457, 275.3409, 274.0368, 272.9942, 272.6259, 272.3626, 270.9984, 
    265.94, 258.2297, 257.0221, 257.4212, 256.0852, 254.5398, 251.6431, 
    249.4879,
  276.2083, 275.3754, 274.6222, 273.4154, 272.6047, 271.3571, 270.5294, 
    264.9535, 254.7088, 253.1449, 255.3978, 255.2109, 253.5037, 250.1208, 
    247.0838,
  275.2138, 274.2533, 273.6327, 272.6792, 271.6836, 270.4805, 268.0692, 
    262.2862, 251.2436, 246.6118, 253.7504, 254.664, 252.854, 249.5261, 
    248.0045,
  262.1857, 263.5632, 257.3104, 262.0073, 259.6715, 259.4481, 262.0602, 
    261.5788, 260.7632, 255.9426, 255.6046, 255.4745, 252.4488, 251.924, 
    249.8085,
  263.2982, 261.2001, 259.7246, 260.2074, 257.6928, 259.5024, 261.3029, 
    260.9213, 260.7875, 258.5679, 257.1983, 257.9873, 257.4361, 250.7382, 
    248.8446,
  272.0396, 270.5219, 266.617, 263.1595, 260.2078, 257.9544, 260.8681, 
    261.2595, 260.7289, 258.3516, 258.0365, 258.0299, 256.0835, 254.7561, 
    251.3174,
  273.706, 273.3096, 272.8968, 270.9175, 267.6271, 266.1137, 261.4441, 
    259.5063, 258.9954, 257.6004, 254.9595, 254.0759, 253.9671, 253.5073, 
    252.2706,
  274.7224, 273.369, 272.9245, 272.7319, 271.5612, 270.9571, 268.831, 
    260.6085, 255.3098, 253.8217, 254.4495, 254.2315, 252.8436, 254.4976, 
    253.0728,
  275.4049, 274.06, 273.4034, 272.8716, 272.6756, 272.1504, 270.1937, 
    266.9146, 261.5025, 259.469, 255.1971, 254.6185, 253.8182, 252.7414, 
    251.4984,
  276.1184, 275.1522, 273.9608, 272.9046, 272.668, 272.3263, 271.3326, 
    265.7506, 262.3054, 261.8685, 255.8277, 252.5963, 253.648, 253.0656, 
    251.39,
  276.2591, 275.3644, 274.0893, 273.0665, 272.6857, 272.3806, 271.0129, 
    266.9547, 261.26, 257.8759, 252.4971, 250.5327, 252.7698, 251.8198, 
    250.353,
  276.2415, 275.3969, 274.6282, 273.4016, 272.5833, 271.1956, 270.4702, 
    265.5824, 259.4849, 255.3893, 250.6094, 250.4415, 251.4694, 250.5604, 
    248.6974,
  275.2505, 274.2539, 273.6232, 272.6347, 271.5634, 270.155, 267.5437, 
    261.975, 256.8417, 249.8201, 248.0475, 250.7348, 251.7596, 250.44, 
    249.3105,
  258.4344, 260.9731, 257.2294, 260.4416, 259.7751, 260.0849, 261.7463, 
    261.1169, 261.334, 260.0338, 261.1302, 261.9497, 260.5061, 259.0499, 
    254.7351,
  262.2694, 263.4084, 262.0828, 261.5349, 260.1939, 261.5663, 261.8733, 
    261.069, 260.5547, 260.3381, 261.4746, 262.8926, 261.9741, 256.0568, 
    253.4842,
  271.8927, 270.835, 268.9024, 265.9787, 262.0673, 257.4507, 261.7218, 
    261.7706, 260.7203, 258.9812, 260.5033, 261.4428, 259.9645, 258.1269, 
    254.513,
  273.652, 273.376, 272.9453, 271.8251, 266.8979, 260.5696, 255.3078, 
    257.6251, 258.5, 257.0389, 257.6931, 258.0309, 257.7903, 257.6828, 256.103,
  274.7381, 273.3647, 272.954, 272.7441, 271.8675, 270.2811, 261.6538, 
    254.0173, 254.7205, 253.8758, 254.8311, 255.2373, 256.17, 257.851, 
    257.3705,
  275.3899, 274.0854, 273.4175, 272.855, 272.6898, 272.1112, 267.9173, 
    263.7554, 259.8426, 257.746, 252.8675, 255.5897, 257.4579, 257.7432, 
    254.8511,
  276.1306, 275.1176, 273.8907, 272.8391, 272.6297, 272.2529, 271.0593, 
    263.7872, 260.0479, 258.0887, 253.4827, 252.7997, 256.3466, 253.9359, 
    252.0447,
  276.2624, 275.3151, 274.0388, 273.0327, 272.6656, 272.3394, 270.6542, 
    266.2478, 259.4254, 256.1223, 251.6298, 251.0361, 250.0601, 249.4072, 
    248.4128,
  276.2375, 275.3737, 274.599, 273.3581, 272.5342, 271.1265, 270.3139, 
    265.976, 258.5338, 253.4728, 250.9926, 248.723, 248.3202, 247.5968, 
    247.4788,
  275.2787, 274.2278, 273.4866, 272.4801, 271.5398, 270.2581, 268.1623, 
    263.8378, 258.6569, 252.456, 248.2429, 248.7706, 247.8689, 247.8456, 
    247.5572,
  259.7058, 261.1056, 257.6552, 258.4177, 256.6455, 257.4155, 259.9093, 
    257.7872, 256.2256, 250.515, 252.9295, 255.707, 252.831, 251.6681, 
    247.7207,
  264.9595, 262.088, 258.8499, 258.6729, 255.6329, 258.9966, 260.4536, 
    259.1279, 257.493, 253.325, 252.6293, 255.7331, 254.5401, 247.491, 244.846,
  271.8166, 269.8803, 267.4335, 264.0962, 259.7693, 256.2852, 262.9379, 
    261.3481, 260.0744, 254.4971, 254.9585, 255.2066, 254.4194, 252.9465, 
    248.9747,
  273.6327, 273.3631, 272.9474, 271.623, 267.6553, 263.5656, 261.6033, 
    260.8553, 260.8186, 256.374, 253.9565, 256.0721, 254.8823, 252.445, 
    250.7816,
  274.7569, 273.3445, 272.9324, 272.7119, 272.0568, 271.1628, 267.9552, 
    261.8599, 260.2993, 258.4151, 254.4944, 255.7552, 254.8231, 253.5162, 
    256.3385,
  275.3894, 274.1261, 273.4017, 272.8449, 272.675, 272.2033, 270.7759, 
    268.4927, 266.8408, 263.631, 255.0236, 256.1459, 253.5707, 252.0308, 
    249.6893,
  276.153, 275.1748, 273.8932, 272.8134, 272.6456, 272.2764, 271.6909, 
    269.7314, 268.2711, 266.0963, 259.1581, 254.0547, 254.1403, 248.7711, 
    247.1146,
  276.279, 275.3289, 274.0587, 273.0063, 272.702, 272.3687, 271.2124, 
    270.3751, 268.7959, 266.8877, 262.062, 255.4505, 252.973, 250.8143, 245.61,
  276.2724, 275.404, 274.6096, 273.3022, 272.5128, 271.2377, 271.1745, 
    270.0761, 269.0455, 267.4041, 263.4937, 257.7619, 253.5397, 248.6838, 
    245.7953,
  275.3858, 274.2307, 273.2744, 272.2604, 271.4167, 270.1598, 270.1835, 
    269.6389, 269.3486, 267.7412, 264.9632, 260.0364, 255.1981, 250.6978, 
    247.614,
  260.9863, 262.0452, 263.2642, 266.5576, 265.7618, 265.8605, 266.7978, 
    264.6841, 258.6557, 244.744, 248.8865, 251.6571, 247.3335, 244.3564, 
    242.5595,
  263.595, 264.3477, 266.6391, 266.852, 265.2227, 266.2051, 266.7898, 
    263.9554, 262.2278, 253.2445, 247.3214, 253.2531, 252.5754, 241.5202, 
    239.4204,
  271.359, 270.061, 270.0178, 268.2882, 265.8099, 263.278, 266.666, 265.7747, 
    265.673, 260.6617, 254.9426, 253.2158, 252.502, 253.4588, 249.4222,
  273.5819, 273.3376, 272.98, 271.7115, 269.2344, 267.087, 263.3783, 260.826, 
    266.4007, 264.6834, 259.5202, 255.3742, 251.2305, 251.3448, 253.1336,
  274.7737, 273.3474, 272.9063, 272.665, 272.0522, 271.2673, 268.3827, 
    263.4547, 264.4885, 266.3118, 262.734, 259.9228, 253.3173, 250.21, 
    251.9469,
  275.432, 274.2046, 273.4082, 272.8088, 272.6144, 272.1255, 270.6111, 
    268.6709, 267.2524, 267.6553, 264.9007, 263.0606, 258.7032, 252.9309, 
    249.8867,
  276.2002, 275.255, 274.0056, 272.8334, 272.6253, 272.2354, 271.6659, 
    269.3645, 268.3967, 267.3821, 266.9257, 263.8937, 261.5626, 256.2022, 
    250.999,
  276.3054, 275.3981, 274.188, 273.0528, 272.7045, 272.3165, 271.1436, 
    270.1968, 268.6414, 267.1378, 267.1686, 264.747, 262.9213, 258.9468, 
    253.635,
  276.3152, 275.466, 274.6428, 273.1729, 272.4177, 271.3076, 271.0369, 
    269.9436, 268.874, 268.1526, 267.6236, 265.1062, 263.9045, 260.9231, 
    255.9344,
  275.5091, 274.2908, 273.1305, 272.1653, 271.5407, 270.7185, 269.3578, 
    267.8631, 268.9192, 267.3148, 267.593, 266.3282, 264.1617, 261.5593, 
    258.1965,
  265.5417, 265.4822, 264.6469, 264.7645, 264.4337, 264.3524, 265.0551, 
    262.9978, 261.6739, 251.9585, 247.3303, 249.1224, 241.347, 242.0529, 
    241.3186,
  266.8918, 266.3261, 265.6113, 264.0049, 262.3565, 263.8398, 262.5971, 
    264.3973, 263.5671, 261.3013, 253.8942, 253.5723, 252.6275, 246.198, 
    242.8944,
  270.8498, 268.9745, 268.4733, 266.3998, 264.3658, 259.0244, 264.7567, 
    264.6234, 264.4154, 263.4218, 261.7052, 259.6595, 257.1063, 255.339, 
    250.5651,
  273.5719, 273.2484, 272.9484, 271.1633, 268.0238, 265.1742, 262.3501, 
    260.4583, 261.4829, 261.6714, 262.1048, 261.8765, 260.9571, 258.9045, 
    257.0824,
  274.7731, 273.3401, 272.871, 272.6008, 271.9781, 271.1168, 268.2034, 
    263.1129, 263.2772, 262.8518, 264.2169, 264.4014, 263.5137, 261.5324, 
    259.5701,
  275.4534, 274.2699, 273.4118, 272.7578, 272.565, 272.0803, 270.7373, 
    268.8297, 268.2267, 267.2323, 267.0002, 265.1614, 265.2484, 264.0807, 
    262.1324,
  276.2383, 275.3224, 274.0752, 272.8417, 272.6178, 272.2448, 271.7803, 
    270.1337, 269.4219, 268.5459, 267.5476, 266.1848, 265.8065, 265.2248, 
    264.0784,
  276.3238, 275.437, 274.2599, 273.1117, 272.7306, 272.3671, 271.4263, 
    271.0301, 270.3116, 269.7208, 269.3173, 267.3823, 266.7105, 266.16, 
    264.6792,
  276.2864, 275.4757, 274.6458, 273.188, 272.4611, 271.5988, 271.5252, 
    271.2316, 270.878, 270.442, 269.9639, 269.0146, 268.1187, 266.1773, 
    264.9194,
  275.4557, 274.3524, 273.5168, 272.3551, 271.7944, 271.4575, 271.4531, 
    270.9008, 271.2465, 270.7271, 270.57, 269.8804, 269.0902, 267.3554, 
    264.7454,
  266.2019, 263.4551, 259.8967, 257.9187, 254.3646, 254.9731, 257.5441, 
    258.0667, 258.8882, 257.9193, 259.4132, 260.1769, 259.3808, 258.9901, 
    259.9278,
  266.4654, 264.0808, 261.0669, 257.8975, 253.6301, 254.6518, 259.3762, 
    259.5687, 259.9939, 259.6373, 260.2663, 262.6188, 263.416, 262.0981, 
    261.5356,
  270.0049, 266.7931, 265.1737, 260.9676, 256.8026, 251.021, 259.209, 
    259.8879, 261.9698, 262.6302, 263.6709, 265.3318, 266.2931, 266.1531, 
    265.4285,
  273.5241, 273.0314, 272.7849, 270.1512, 264.8652, 259.46, 258.7143, 
    261.7816, 265.3589, 266.7007, 267.5973, 268.3289, 267.8181, 267.016, 
    266.085,
  274.7281, 273.3, 272.8342, 272.559, 272.0383, 271.0736, 268.2714, 265.0007, 
    266.4371, 268.1554, 269.8581, 269.3293, 267.917, 266.8658, 266.187,
  275.41, 274.2622, 273.3911, 272.7339, 272.5928, 272.1649, 271.4304, 
    269.5733, 270.1509, 270.5824, 270.3494, 268.2851, 267.0772, 266.325, 
    265.4037,
  276.2063, 275.2868, 274.0099, 272.8233, 272.6158, 272.3272, 271.9939, 
    271.3703, 271.5391, 270.9609, 268.3848, 266.7185, 265.8391, 264.9578, 
    264.2464,
  276.3009, 275.3725, 274.1819, 273.0979, 272.7378, 272.5067, 271.8294, 
    271.5897, 271.4664, 268.6506, 266.2915, 264.8777, 264.3805, 263.3425, 
    263.1761,
  276.226, 275.4112, 274.5942, 273.2854, 272.5484, 271.8077, 271.8352, 
    271.613, 269.4336, 267.0228, 265.4129, 263.2037, 262.2, 261.584, 261.7984,
  275.3311, 274.2928, 273.7339, 272.648, 271.9489, 271.7436, 271.5464, 
    268.4556, 266.6268, 262.6353, 264.5779, 262.0088, 260.7061, 260.2259, 
    260.1727,
  266.3993, 264.8229, 262.4151, 259.9966, 256.153, 254.4873, 256.1296, 
    252.8419, 251.5787, 249.7008, 251.9059, 255.6396, 257.6511, 259.7136, 
    256.879,
  267.5602, 266.8361, 263.6435, 260.4395, 255.8454, 254.9569, 256.748, 
    253.8224, 253.4495, 252.624, 254.2252, 258.9751, 261.2792, 257.8906, 
    254.7111,
  270.5204, 268.4767, 267.2751, 263.8799, 258.508, 254.4162, 258.8419, 
    257.946, 257.1099, 256.2344, 258.0056, 260.7807, 261.1384, 258.5388, 
    255.1245,
  273.5143, 273.0942, 272.782, 270.6721, 265.863, 259.8291, 256.4024, 
    257.2772, 258.5237, 258.5493, 261.1462, 262.3574, 260.6917, 259.1396, 
    256.3559,
  274.6588, 273.2776, 272.8321, 272.5482, 272.022, 270.6782, 265.8167, 
    259.1491, 257.7156, 263.2297, 266.0291, 263.7159, 261.8839, 260.6471, 
    259.106,
  275.326, 274.2516, 273.3813, 272.7247, 272.5802, 272.1651, 271.4685, 
    267.5372, 265.2751, 266.7055, 267.0455, 264.8725, 263.5034, 261.5472, 
    258.9412,
  276.1107, 275.2331, 273.9805, 272.8108, 272.6063, 272.3226, 272.0306, 
    270.7838, 268.6712, 268.3344, 267.3353, 265.2457, 263.4985, 261.2653, 
    258.4838,
  276.2505, 275.3093, 274.1365, 273.0864, 272.7051, 272.5425, 271.8624, 
    271.1024, 268.9734, 268.1652, 267.2315, 264.8053, 263.0564, 260.3278, 
    258.1669,
  276.1819, 275.382, 274.5517, 273.2547, 272.5038, 271.7691, 271.4991, 
    270.4236, 269.3712, 268.9623, 268.14, 264.9631, 262.5455, 259.6313, 
    257.8102,
  275.3102, 274.2921, 273.7039, 272.3697, 271.2725, 270.8069, 270.2346, 
    269.3723, 269.4732, 267.6749, 268.1039, 264.4904, 261.4473, 258.6849, 
    256.5536,
  267.2129, 266.4179, 266.3036, 266.3236, 264.761, 263.5384, 263.1969, 
    259.9304, 256.9395, 250.5798, 249.7067, 251.5012, 248.9693, 247.6992, 
    246.303,
  266.9453, 266.8938, 266.7766, 266.4668, 264.8014, 263.5108, 263.9352, 
    260.4788, 257.9661, 255.7283, 254.0449, 254.9085, 253.7298, 249.2047, 
    249.0615,
  270.9435, 269.5103, 268.6579, 267.6676, 266.2557, 262.1836, 264.6854, 
    263.1667, 258.6942, 257.8922, 258.057, 257.9426, 257.4608, 258.2432, 
    257.3627,
  273.5515, 273.2763, 272.8959, 271.5415, 269.2726, 265.6631, 262.1785, 
    262.2612, 261.1139, 260.687, 260.8093, 260.4912, 261.3536, 260.1084, 
    256.9872,
  274.5965, 273.2674, 272.8303, 272.5389, 272.0511, 271.101, 268.0919, 
    261.5843, 261.7336, 263.4556, 264.8994, 263.8416, 262.6569, 258.5551, 
    257.0297,
  275.2921, 274.2962, 273.3766, 272.7104, 272.5596, 272.1391, 271.5977, 
    269.4355, 266.737, 265.6916, 266.932, 265.336, 260.8862, 257.6148, 
    256.3272,
  276.0676, 275.2208, 273.9787, 272.7985, 272.5878, 272.2915, 272.0157, 
    270.8759, 266.318, 267.2131, 265.7785, 261.515, 257.9507, 256.1929, 
    254.9878,
  276.2493, 275.2842, 274.1346, 273.0748, 272.6664, 272.5336, 271.8361, 
    271.0826, 268.5772, 266.6296, 261.4157, 257.4402, 255.7207, 254.058, 
    253.3753,
  276.1764, 275.3983, 274.5351, 273.1638, 272.4228, 271.7492, 271.3893, 
    270.6244, 268.5959, 265.8481, 263.1521, 256.2294, 253.8288, 252.4151, 
    252.138,
  275.3494, 274.2855, 273.5663, 272.1728, 271.0564, 270.4362, 269.7793, 
    267.9533, 265.9419, 260.6219, 262.2389, 255.8159, 252.5187, 251.137, 
    250.2212,
  262.8116, 263.7238, 263.5239, 266.1033, 265.8125, 267.4249, 268.3117, 
    268.0323, 266.8921, 263.9668, 261.3156, 260.0544, 256.2135, 253.7088, 
    249.8924,
  264.7351, 265.0204, 267.162, 268.6396, 267.9943, 269.3922, 269.869, 
    268.8982, 267.2636, 263.9164, 262.7429, 261.8089, 259.7289, 253.9366, 
    251.9368,
  270.9826, 269.8822, 269.9982, 270.8331, 270.4888, 269.6832, 270.0133, 
    269.3829, 267.2505, 264.7677, 264.0781, 262.8909, 261.853, 260.557, 
    257.5813,
  273.5363, 273.3615, 272.9518, 272.1184, 271.9132, 271.4777, 269.7739, 
    268.7077, 266.9694, 265.6714, 264.1934, 263.3131, 263.3385, 262.3562, 
    260.9053,
  274.5902, 273.3163, 272.8701, 272.57, 272.1448, 271.8206, 271.2935, 
    267.836, 266.7484, 265.9029, 266.8708, 266.4944, 265.3385, 263.6912, 
    262.0641,
  275.3409, 274.3767, 273.4104, 272.7408, 272.5854, 272.1484, 271.7305, 
    270.6253, 269.6273, 268.6986, 267.7667, 267.2269, 266.1969, 264.4545, 
    261.5033,
  276.0729, 275.2582, 274.0258, 272.8474, 272.6298, 272.3105, 272.0412, 
    271.2921, 268.3111, 267.1225, 266.311, 266.8275, 265.0633, 262.7144, 
    257.6987,
  276.2778, 275.3125, 274.1872, 273.1209, 272.6943, 272.56, 271.8442, 
    271.3427, 269.3281, 268.3778, 267.9535, 266.2452, 264.2059, 258.5146, 
    253.6002,
  276.1947, 275.4501, 274.5703, 273.1221, 272.4275, 271.7879, 271.6434, 
    270.7175, 269.5258, 269.1759, 268.848, 264.6074, 258.74, 253.177, 251.7335,
  275.3944, 274.3257, 273.5646, 272.3135, 271.6842, 271.115, 270.2506, 
    269.4171, 269.8113, 268.0223, 266.8225, 259.7879, 253.1116, 249.9035, 
    248.0187,
  259.617, 261.6701, 261.6107, 263.0143, 262.7346, 264.7657, 266.5186, 
    266.7595, 265.798, 265.0623, 264.5154, 265.0399, 263.615, 264.5858, 
    263.6672,
  263.7336, 263.8291, 263.4698, 263.0299, 263.3061, 267.0608, 267.1713, 
    266.0974, 265.534, 264.3478, 264.3748, 264.8581, 265.3761, 265.4543, 
    265.2933,
  271.1048, 269.2915, 268.0737, 266.0732, 267.8657, 266.5052, 268.9042, 
    266.4183, 265.3549, 264.8282, 265.6929, 266.6711, 268.4174, 268.3392, 
    267.3625,
  273.4943, 273.3468, 272.9321, 271.6769, 269.6162, 269.8442, 268.3898, 
    267.8751, 267.0023, 266.6609, 267.658, 268.9568, 269.277, 268.867, 
    265.9005,
  274.5499, 273.3209, 272.846, 272.5464, 272.1554, 271.5721, 270.7778, 
    267.7699, 267.7715, 269.2151, 270.2438, 269.9932, 269.7901, 268.9272, 
    265.4212,
  275.3075, 274.335, 273.383, 272.7162, 272.5805, 272.1526, 271.7642, 
    270.8733, 270.1254, 270.5622, 270.054, 269.8269, 269.7856, 268.3693, 
    262.8107,
  276.0091, 275.23, 274.0327, 272.8455, 272.6339, 272.3208, 272.0685, 
    271.5686, 270.5842, 269.5874, 269.2609, 269.4967, 269.6941, 266.2338, 
    259.1068,
  276.2553, 275.3116, 274.1872, 273.1247, 272.6977, 272.5955, 271.8853, 
    271.5477, 270.5142, 269.5946, 269.1627, 270.0543, 268.5354, 261.1888, 
    254.0797,
  276.1785, 275.4548, 274.582, 273.1174, 272.4399, 271.8055, 271.7159, 
    271.027, 270.2369, 270.0018, 270.5858, 269.8649, 264.4836, 254.758, 
    250.7329,
  275.3685, 274.3427, 273.612, 272.3361, 271.7043, 271.3492, 270.6894, 
    269.6766, 269.7783, 269.4792, 270.5466, 267.5731, 257.4786, 250.6939, 
    247.3719,
  258.4252, 260.031, 259.2716, 259.615, 257.2449, 257.3978, 260.6736, 
    260.7722, 262.5562, 263.235, 264.0945, 264.9583, 264.7411, 265.1204, 
    265.3149,
  263.2697, 262.9278, 260.8537, 259.3682, 258.0883, 262.9023, 264.9879, 
    264.3543, 265.3988, 265.6366, 265.8434, 266.0692, 265.2705, 265.0094, 
    266.2041,
  271.6316, 269.8479, 267.6798, 265.4147, 266.7875, 265.343, 268.2636, 
    267.6609, 266.8917, 266.172, 265.3649, 265.5666, 266.7293, 268.3651, 
    269.1781,
  273.5672, 273.3848, 272.9128, 272.0577, 269.8145, 268.2768, 266.6955, 
    269.1433, 267.2819, 264.6721, 265.9717, 267.3679, 268.8501, 269.6667, 
    269.4095,
  274.4646, 273.2972, 272.8665, 272.5358, 272.2183, 271.2994, 270.1184, 
    266.3055, 266.9165, 268.241, 269.7182, 269.3956, 269.9538, 269.928, 
    269.2636,
  275.2054, 274.2393, 273.3726, 272.7032, 272.5961, 272.1695, 271.7753, 
    270.6137, 269.5846, 270.0434, 270.3066, 270.2265, 270.1563, 270.0305, 
    268.2637,
  275.9168, 275.1581, 273.9846, 272.8251, 272.6231, 272.3247, 272.0775, 
    271.6254, 271.0108, 270.6276, 270.5758, 270.4575, 270.2506, 269.756, 
    266.062,
  276.2155, 275.2754, 274.1617, 273.1299, 272.6911, 272.6228, 271.9098, 
    271.6327, 271.2587, 270.8666, 270.6863, 270.5782, 270.3973, 268.6475, 
    264.1252,
  276.1247, 275.4267, 274.5904, 273.1517, 272.4518, 271.8257, 271.7972, 
    271.5036, 271.3151, 271.2498, 271.2787, 270.742, 270.0799, 267.0079, 
    261.7885,
  275.2435, 274.3284, 273.6839, 272.4246, 271.8298, 271.6006, 271.3786, 
    271.1015, 271.3025, 271.5259, 271.402, 270.8646, 269.0205, 265.0959, 
    259.4162,
  257.5888, 259.249, 258.6602, 259.5597, 257.4293, 257.5934, 258.9878, 
    257.3445, 257.7643, 257.8221, 259.6331, 260.3739, 260.8979, 262.1771, 
    262.7328,
  263.003, 261.355, 259.1487, 258.0856, 255.8516, 260.89, 262.8879, 261.4229, 
    261.0563, 261.4636, 262.2603, 263.2755, 263.8958, 263.5149, 264.3643,
  272.0959, 270.6219, 267.6503, 264.2244, 260.5131, 260.5348, 267.2551, 
    265.2237, 264.1271, 263.8455, 263.8938, 264.6171, 265.3148, 265.8885, 
    266.3225,
  273.6465, 273.4414, 272.9228, 272.3669, 268.9817, 264.5754, 263.5533, 
    268.1522, 267.1821, 266.1211, 265.4735, 264.8074, 265.9664, 266.4769, 
    266.7333,
  274.3867, 273.3031, 272.9027, 272.56, 272.2984, 271.0958, 269.2155, 
    264.7191, 265.6899, 266.723, 268.381, 265.9598, 266.2354, 267.2864, 
    266.4668,
  275.1317, 274.1917, 273.3565, 272.7092, 272.6118, 272.1967, 271.77, 
    269.9078, 267.3834, 267.9051, 268.062, 266.7773, 266.9095, 267.6568, 
    268.0326,
  275.8184, 275.0723, 273.9062, 272.7942, 272.5995, 272.3145, 272.0641, 
    271.6178, 270.1506, 268.0752, 267.6865, 267.412, 268.019, 268.2186, 
    268.5048,
  276.1429, 275.1862, 274.0844, 273.0858, 272.6561, 272.6176, 271.8957, 
    271.6, 270.5037, 268.6958, 268.0318, 267.7694, 267.7599, 267.8638, 
    268.5667,
  276.0309, 275.336, 274.5472, 273.2074, 272.4568, 271.8196, 271.7946, 
    271.3665, 270.2293, 269.7611, 270.05, 268.5174, 268.6187, 268.6992, 
    268.6146,
  275.0351, 274.1876, 273.6457, 272.469, 271.3294, 270.8208, 270.5136, 
    270.366, 270.5427, 270.418, 270.8947, 270.3648, 269.7429, 269.3161, 
    268.9783,
  257.0275, 258.5514, 258.3503, 259.259, 255.6421, 256.0599, 257.1558, 
    254.5353, 252.4643, 252.0817, 252.9886, 253.4942, 252.2196, 251.8752, 
    251.4125,
  262.1255, 259.1576, 257.566, 256.2385, 254.1121, 259.2172, 260.8375, 
    257.0621, 254.3383, 253.3211, 254.0905, 255.0885, 254.3876, 252.3958, 
    253.3374,
  272.3159, 270.1377, 266.5883, 261.3094, 255.0662, 253.5243, 265.3074, 
    261.4197, 258.0418, 255.3024, 256.1754, 256.3998, 255.5538, 255.6169, 
    256.1923,
  273.6753, 273.4559, 272.9145, 272.3814, 267.5505, 259.4362, 257.2731, 
    265.8293, 263.6035, 260.6438, 259.4542, 260.1441, 260.2647, 260.9674, 
    261.1835,
  274.3521, 273.2971, 272.8977, 272.552, 272.3235, 270.1896, 266.0356, 
    260.2221, 261.281, 263.6058, 265.4756, 264.2286, 263.8584, 263.9111, 
    263.8571,
  275.1205, 274.1603, 273.3127, 272.6843, 272.5912, 272.2212, 271.7672, 
    269.5705, 263.9951, 264.2016, 264.8233, 265.9051, 265.9119, 265.8243, 
    265.6363,
  275.7404, 274.9904, 273.8264, 272.7334, 272.5503, 272.2773, 272.0437, 
    271.6192, 270.1424, 266.6673, 267.1958, 267.15, 266.9965, 266.7928, 
    266.4106,
  276.0725, 275.0794, 273.957, 272.9725, 272.5621, 272.5634, 271.8296, 
    271.5604, 269.8047, 264.8181, 265.9496, 266.0219, 266.5884, 266.7796, 
    266.6035,
  275.9512, 275.2238, 274.426, 273.0844, 272.3155, 271.6818, 271.6352, 
    270.6942, 267.557, 266.058, 268.524, 266.6438, 266.5421, 266.1188, 
    266.0224,
  274.8577, 273.7884, 273.189, 271.87, 269.8705, 267.3199, 263.3215, 
    260.2935, 263.9553, 264.7719, 267.8375, 267.3782, 265.3396, 265.6891, 
    266.1124,
  259.4874, 260.3489, 260.0607, 260.6207, 258.1136, 258.5215, 259.4492, 
    256.8496, 255.2615, 253.5978, 253.1339, 254.1424, 251.9299, 251.2668, 
    249.3127,
  264.7248, 261.2207, 259.3977, 258.1694, 255.9321, 260.6499, 261.5324, 
    258.4799, 255.8772, 255.0491, 255.4855, 256.032, 254.2177, 250.5154, 
    249.41,
  272.4667, 270.4749, 268.138, 262.7576, 257.7968, 255.8427, 264.501, 
    261.0665, 258.1753, 255.5597, 257.062, 255.9462, 254.6749, 252.8855, 
    251.1701,
  273.6537, 273.4246, 272.8888, 272.3383, 268.2645, 259.7957, 256.8864, 
    264.7908, 262.5665, 259.186, 257.9304, 257.5959, 255.7485, 255.1727, 
    253.3602,
  274.3622, 273.2783, 272.8531, 272.4986, 272.2487, 270.1461, 264.6422, 
    257.5705, 257.4815, 261.8367, 263.127, 260.0357, 257.8585, 255.9205, 
    254.2217,
  275.1409, 274.105, 273.2689, 272.6026, 272.5196, 272.1566, 271.6476, 
    268.0887, 262.0287, 259.6765, 261.6192, 262.3015, 262.5296, 262.2085, 
    261.5618,
  275.698, 274.9491, 273.7824, 272.6652, 272.5047, 272.2097, 271.9857, 
    271.5054, 269.9667, 266.1613, 264.7666, 264.5708, 264.0037, 263.5516, 
    263.4481,
  276.0386, 275.052, 273.8991, 272.8975, 272.4805, 272.4989, 271.7092, 
    271.3397, 268.252, 257.5721, 255.6352, 255.2609, 254.7744, 255.546, 
    255.9279,
  275.934, 275.1852, 274.4012, 273.0115, 272.2, 271.4745, 271.109, 269.5703, 
    264.6599, 261.1567, 264.9253, 255.1681, 253.7155, 253.0368, 253.9736,
  274.8053, 273.6943, 273.0626, 271.4397, 269.6807, 266.937, 261.257, 
    256.1098, 256.5564, 254.3773, 259.8407, 255.1988, 254.2038, 254.1245, 
    254.6224,
  259.5141, 261.1654, 260.3459, 261.2226, 258.3525, 259.1678, 260.1729, 
    258.8778, 257.5536, 255.5845, 255.6648, 256.19, 255.2811, 254.5789, 
    254.0363,
  266.2959, 264.1576, 261.4086, 259.7472, 256.5803, 261.6212, 262.9001, 
    259.8714, 258.1398, 257.2781, 257.8931, 257.9286, 256.5502, 253.8343, 
    253.7548,
  272.4223, 270.8537, 269.3261, 264.7105, 259.261, 257.2164, 265.0692, 
    262.4646, 260.332, 258.4662, 259.1959, 258.3904, 257.0011, 256.2332, 
    254.9445,
  273.6013, 273.3645, 272.8461, 272.1501, 268.0407, 260.9975, 257.7769, 
    265.1198, 263.6368, 260.6077, 260.5152, 259.7986, 258.459, 257.4841, 
    256.2206,
  274.4149, 273.2639, 272.8206, 272.4537, 272.1214, 269.8008, 265.3878, 
    259.2801, 260.284, 261.6211, 263.3521, 261.1851, 259.941, 258.5201, 
    257.692,
  275.1878, 274.0824, 273.2814, 272.547, 272.4554, 272.0885, 271.4568, 
    267.9007, 262.8261, 259.4322, 259.3258, 259.6316, 259.3914, 259.4344, 
    259.1372,
  275.7049, 274.961, 273.7905, 272.6389, 272.4855, 272.1635, 271.9305, 
    271.2973, 268.5481, 263.746, 261.4055, 260.8976, 261.3166, 260.4219, 
    258.4448,
  276.0548, 275.0782, 273.8936, 272.8578, 272.4012, 272.4135, 271.5116, 
    270.8107, 265.8189, 257.0833, 255.9784, 255.7599, 255.5085, 255.414, 
    254.4553,
  275.9485, 275.1709, 274.3975, 272.9061, 271.9755, 270.6125, 269.6284, 
    266.6776, 260.9843, 257.6153, 261.037, 251.4124, 251.9077, 250.9417, 
    250.0473,
  274.632, 273.3607, 272.6549, 270.164, 266.9894, 262.7599, 257.1188, 
    254.2197, 254.1043, 250.0492, 254.0388, 248.9429, 248.4425, 247.8214, 
    249.9206,
  260.796, 262.1544, 261.339, 261.3478, 258.1153, 257.1975, 259.3176, 
    257.425, 256.2739, 252.904, 254.3954, 255.1884, 252.9041, 251.3217, 
    250.406,
  266.4415, 264.3941, 262.2983, 259.9831, 258.5806, 262.2366, 262.5268, 
    258.3563, 255.8292, 254.1635, 255.9089, 257.3057, 255.8261, 251.7323, 
    251.7868,
  272.4471, 271.0953, 269.3868, 264.4872, 259.996, 257.3217, 264.6871, 
    261.4247, 258.3856, 254.4494, 256.9997, 256.9497, 255.4738, 254.8703, 
    253.2303,
  273.5941, 273.324, 272.8766, 271.9834, 268.0404, 261.2384, 258.039, 
    264.0443, 261.5656, 258.0464, 257.4809, 257.0085, 255.6166, 255.978, 
    255.1336,
  274.4369, 273.2235, 272.7759, 272.4095, 272.0542, 269.2909, 263.8752, 
    258.4258, 258.6143, 260.5052, 261.3456, 259.229, 257.4156, 256.4163, 
    255.4666,
  275.1595, 274.0287, 273.2364, 272.4724, 272.3992, 272.0071, 271.1864, 
    266.8506, 261.7724, 260.2104, 260.009, 259.4098, 258.5063, 257.5388, 
    256.2419,
  275.6602, 274.8771, 273.7101, 272.5669, 272.4286, 272.1033, 271.841, 
    270.6686, 266.4048, 261.8921, 260.0746, 259.0655, 258.9893, 258.2548, 
    257.6782,
  276.0289, 275.0295, 273.812, 272.7524, 272.2843, 272.2841, 270.9515, 
    269.4313, 260.9182, 255.7156, 255.9309, 256.4408, 256.9569, 256.6931, 
    256.4802,
  275.9472, 275.1302, 274.3533, 272.8402, 271.6504, 269.5731, 267.7792, 
    263.7655, 258.727, 255.7405, 257.1746, 251.2243, 250.9033, 251.2355, 
    252.024,
  274.7241, 273.4572, 272.4626, 269.4321, 266.0283, 261.0604, 256.0958, 
    253.3719, 252.2496, 248.136, 249.9594, 246.4073, 245.8501, 246.269, 
    248.3954,
  263.4989, 263.3398, 261.8231, 262.0274, 257.8688, 257.768, 258.7488, 
    256.4366, 255.8676, 252.6535, 253.2039, 253.7838, 249.4416, 248.0734, 
    245.8754,
  267.0827, 265.2071, 262.6913, 261.4232, 258.1365, 262.2015, 262.1362, 
    257.9399, 255.8908, 255.0891, 255.3784, 256.7192, 254.3219, 248.5182, 
    247.119,
  272.451, 270.9428, 268.8775, 263.3363, 261.0733, 258.4611, 264.5856, 
    261.3639, 258.0557, 255.0207, 257.904, 257.5777, 254.8938, 253.3579, 
    250.2575,
  273.5721, 273.2602, 272.8488, 271.4796, 267.2533, 262.3413, 258.5616, 
    263.2534, 261.552, 257.9155, 257.1779, 257.2753, 256.2173, 255.1175, 
    253.2411,
  274.4532, 273.1983, 272.7422, 272.3593, 271.8151, 268.1916, 264.1394, 
    258.3539, 255.9982, 259.3603, 260.9657, 258.2466, 257.5142, 256.5136, 
    254.437,
  275.1302, 273.9904, 273.1782, 272.4166, 272.3326, 271.9218, 270.5302, 
    265.0579, 257.7693, 255.862, 257.7806, 259.0048, 257.4879, 256.7572, 
    255.048,
  275.6414, 274.8176, 273.6585, 272.5386, 272.4031, 272.0599, 271.7022, 
    269.0381, 261.4911, 257.058, 257.2979, 256.6916, 257.0245, 256.4543, 
    255.8543,
  276.0158, 275.0313, 273.826, 272.7086, 272.2079, 272.1991, 270.4782, 
    268.2808, 258.4894, 252.9574, 252.0259, 254.1499, 256.9509, 256.2738, 
    255.87,
  275.9268, 275.0923, 274.3467, 272.751, 271.4554, 269.2531, 267.6261, 
    263.0736, 257.4825, 253.4946, 252.7164, 250.3784, 253.2791, 256.0321, 
    255.667,
  274.6565, 273.2935, 272.0197, 267.4762, 263.4888, 259.2328, 256.3286, 
    254.0592, 250.5184, 245.1722, 246.7389, 246.3779, 249.8736, 254.8152, 
    255.6954,
  266.3373, 266.6425, 265.4037, 264.2509, 260.6729, 259.5548, 260.6503, 
    257.1045, 257.9081, 255.2384, 255.9423, 256.2124, 252.0522, 249.1591, 
    245.8963,
  267.6804, 266.0492, 264.7731, 263.1618, 260.0432, 262.8686, 262.5864, 
    258.7665, 257.8704, 258.2169, 257.9663, 258.9186, 256.5894, 250.0502, 
    246.9382,
  272.5032, 270.5911, 267.9276, 263.9613, 260.9688, 257.9801, 263.8073, 
    261.2767, 258.46, 256.3954, 260.5186, 259.8492, 257.3042, 254.9141, 
    251.2141,
  273.5465, 273.2479, 272.8142, 270.6438, 264.8434, 260.1135, 256.3771, 
    261.8282, 260.6446, 257.8536, 257.6528, 257.7697, 257.5439, 256.4236, 
    254.116,
  274.4283, 273.152, 272.7228, 272.3288, 271.5332, 266.6365, 261.261, 
    256.9066, 257.0092, 258.378, 259.4753, 257.3059, 256.701, 257.0841, 
    255.8604,
  275.035, 273.9162, 273.1339, 272.3675, 272.2874, 271.85, 269.7927, 
    263.5756, 257.7074, 256.2779, 256.4518, 258.0962, 256.7837, 255.6284, 
    254.8566,
  275.5836, 274.743, 273.6097, 272.5254, 272.3928, 272.052, 271.638, 
    269.2792, 262.3379, 258.3854, 254.7232, 252.61, 253.5411, 253.7796, 
    253.8195,
  275.9731, 274.9892, 273.7829, 272.6283, 272.1349, 272.1322, 270.4541, 
    268.8469, 261.652, 255.8991, 252.0229, 250.4379, 248.7828, 248.5379, 
    249.281,
  275.8317, 274.9607, 274.2412, 272.6729, 269.8435, 266.8328, 267.0011, 
    265.2455, 261.0796, 256.8586, 252.3722, 248.3927, 246.4949, 245.0852, 
    245.5809,
  274.4431, 273.0766, 271.6979, 264.4708, 258.8762, 254.5939, 255.3477, 
    258.2135, 256.2619, 251.9028, 248.3932, 245.6276, 243.7844, 243.8903, 
    245.026,
  259.6546, 264.9276, 264.2466, 265.5115, 264.1454, 264.2561, 264.4707, 
    261.4751, 259.446, 255.9729, 254.1493, 252.4697, 247.8217, 247.4662, 
    247.7153,
  264.8755, 263.8149, 263.9841, 263.7193, 261.7851, 265.3572, 265.6127, 
    262.0249, 259.9664, 257.5606, 256.4327, 256.7001, 253.0992, 245.4035, 
    246.8122,
  272.469, 269.9156, 266.3132, 263.6126, 262.8212, 262.0798, 265.5292, 
    262.9896, 260.275, 258.5355, 259.9726, 258.1978, 252.7228, 250.5692, 
    248.3544,
  273.5057, 273.1756, 272.7606, 269.967, 265.6669, 262.8953, 260.6978, 
    262.5699, 260.7898, 258.136, 258.0731, 257.9555, 254.1638, 251.6912, 
    250.392,
  274.409, 273.0872, 272.6934, 272.2938, 271.1168, 266.7941, 262.5673, 
    256.7285, 255.7958, 257.4186, 257.4048, 256.8331, 255.4982, 254.0803, 
    250.6472,
  274.9618, 273.8338, 273.0737, 272.3082, 272.2294, 271.7341, 269.3999, 
    263.884, 259.5428, 258.0414, 256.6685, 256.7931, 257.0326, 256.5155, 
    252.1673,
  275.5247, 274.6684, 273.5151, 272.4604, 272.3508, 271.9934, 271.4946, 
    269.6836, 263.1716, 260.1623, 257.2824, 256.0438, 256.1754, 257.0407, 
    255.7919,
  275.9181, 274.8673, 273.6506, 272.5306, 272.0869, 271.8896, 269.5124, 268, 
    260.2725, 257.3715, 258.1045, 256.7015, 255.955, 255.922, 256.1066,
  275.7473, 274.8805, 274.1679, 272.6003, 267.7961, 264.0921, 262.4177, 
    259.2763, 255.2571, 254.4377, 259.0869, 257.6639, 255.9386, 254.9637, 
    254.1311,
  274.3489, 272.8357, 271.1656, 263.102, 256.7216, 252.5395, 251.4574, 
    252.7435, 252.1, 251.2443, 257.1728, 256.6649, 255.3224, 254.421, 254.3555,
  259.0945, 261.7176, 258.9331, 262.3412, 261.8521, 262.5234, 262.6436, 
    260.2773, 257.3482, 257.041, 256.6996, 257.4236, 256.8247, 256.4772, 
    255.4115,
  265.2934, 263.4417, 261.0409, 259.8875, 260.6419, 263.1209, 263.1836, 
    261.7594, 259.2524, 258.7539, 259.0265, 260.3337, 259.308, 254.7429, 
    254.2553,
  272.4167, 269.8807, 265.8751, 261.4167, 259.0481, 257.2587, 263.5735, 
    263.1762, 262.0529, 260.0014, 261.5132, 260.3712, 258.5004, 257.4, 
    254.1973,
  273.4343, 273.1357, 272.7513, 269.899, 263.7296, 261.4178, 259.0708, 
    263.3231, 262.9146, 260.6553, 260.218, 260.1214, 258.2664, 256.8474, 
    254.6212,
  274.3583, 273.0148, 272.653, 272.2453, 270.728, 266.1226, 263.6588, 
    259.9963, 259.432, 259.8407, 260.5202, 259.2833, 257.3143, 255.7999, 
    253.2124,
  274.9075, 273.7422, 272.9986, 272.2528, 272.1962, 271.5849, 269.2563, 
    265.2867, 262.5337, 261.9067, 261.0812, 259.9161, 257.447, 254.9089, 
    252.6388,
  275.4474, 274.6067, 273.422, 272.3856, 272.3193, 271.9774, 271.3371, 
    269.2808, 264.934, 263.2789, 261.3665, 258.8653, 256.4193, 253.6407, 
    251.3281,
  275.9022, 274.809, 273.5488, 272.4389, 272.015, 271.5105, 269.048, 
    267.7071, 262.5303, 261.208, 259.9829, 258.2953, 255.9328, 253.0441, 
    250.7436,
  275.7697, 274.8874, 274.1478, 272.3553, 265.9788, 262.7239, 260.7225, 
    258.1875, 258.263, 259.1595, 259.0065, 257.4693, 254.0737, 252.5938, 
    250.7098,
  274.4087, 272.7931, 270.7038, 262.239, 254.8331, 251.3761, 250.83, 
    253.1998, 252.335, 251.7654, 256.6029, 255.243, 253.5665, 252.1842, 
    251.9873,
  260.9606, 262.8603, 258.3127, 261.6676, 260.7036, 259.9873, 261.2365, 
    258.9669, 257.36, 255.2707, 255.8925, 258.5995, 258.1948, 257.9652, 
    256.757,
  264.6526, 260.6516, 260.0658, 259.1856, 259.3103, 260.9724, 261.3217, 
    258.7744, 256.3209, 257.9471, 257.7755, 260.0176, 260.4053, 256.2386, 
    255.4127,
  272.3986, 269.658, 263.5257, 258.1619, 259.087, 254.0184, 260.8974, 
    259.729, 258.052, 258.4626, 260.1295, 259.1953, 257.9809, 258.2353, 
    256.4302,
  273.4419, 273.1059, 272.6872, 269.0225, 260.6221, 258.9212, 255.6619, 
    259.0991, 259.149, 258.627, 258.8623, 258.8174, 257.1274, 256.8612, 
    257.5804,
  274.2583, 272.9374, 272.5954, 272.1971, 270.053, 263.7521, 261.378, 
    252.5448, 254.0732, 257.8159, 258.8599, 258.3541, 257.197, 256.9545, 
    257.3455,
  274.8955, 273.6689, 272.9213, 272.1703, 272.1243, 271.3398, 267.7314, 
    263.1039, 260.5124, 260.1078, 260.486, 259.4975, 257.8861, 256.3441, 
    255.7797,
  275.4387, 274.586, 273.3499, 272.3192, 272.2856, 271.944, 271.0313, 
    268.408, 262.9805, 261.9948, 260.7957, 259.0431, 257.1534, 256.3462, 
    256.4766,
  275.9161, 274.84, 273.504, 272.3657, 271.9363, 271.21, 269.6521, 267.5331, 
    262.0314, 259.8676, 258.1794, 259.0099, 257.7666, 256.2876, 256.603,
  275.8079, 274.8988, 274.1242, 271.8025, 264.4283, 262.6924, 262.5566, 
    261.9547, 260.2159, 259.2316, 257.8687, 258.8469, 257.8843, 256.7358, 
    255.6939,
  274.3128, 272.4663, 270.0839, 260.8147, 253.5571, 251.5975, 253.5323, 
    258.6498, 257.4313, 256.3954, 258.2589, 259.132, 258.1289, 257.4677, 
    255.5081,
  261.2717, 264.5676, 260.6876, 263.2983, 261.8976, 260.7939, 261.8486, 
    260.5477, 260.0972, 255.8938, 255.7107, 257.2783, 254.4798, 253.1226, 
    251.6639,
  265.7742, 263.8473, 263.278, 262.4718, 260.2881, 260.3821, 261.6, 259.564, 
    257.4244, 258.5975, 256.6797, 259.2792, 259.5356, 252.0677, 251.0388,
  272.5482, 269.6129, 265.8564, 262.913, 259.6905, 254.0734, 259.6464, 
    258.2969, 256.9793, 257.9147, 259.2509, 257.6773, 257.57, 258.4203, 
    254.245,
  273.5387, 273.2374, 272.7584, 269.6805, 261.6739, 258.382, 249.8297, 
    255.6758, 256.8596, 256.8397, 256.7679, 256.9963, 256.5424, 257.267, 
    257.715,
  274.1925, 272.911, 272.5804, 272.1921, 269.5605, 262.3202, 259.7466, 
    250.2382, 251.6672, 254.6542, 255.8534, 256.7717, 256.6819, 257.3284, 
    257.799,
  274.889, 273.6796, 272.873, 272.1162, 272.0984, 271.0356, 265.657, 
    261.7879, 259.9172, 260.7445, 259.1383, 258.0194, 257.2548, 255.7809, 
    254.5856,
  275.4377, 274.5333, 273.3108, 272.2846, 272.2694, 271.901, 270.8713, 
    266.8925, 262.7972, 263.0443, 260.9611, 258.4757, 256.9581, 254.8793, 
    251.9201,
  275.8897, 274.824, 273.4521, 272.3115, 271.9436, 271.1049, 269.8938, 
    267.1785, 261.3029, 259.9351, 258.1941, 257.3925, 255.4134, 251.7253, 
    249.5168,
  275.7778, 274.8695, 274.0464, 270.7808, 265.4904, 265.4991, 264.756, 
    262.5588, 260.1392, 258.0334, 256.2738, 255.2406, 252.5972, 250.9111, 
    250.2373,
  273.88, 271.6243, 268.8763, 260.8651, 258.1988, 259.6879, 260.439, 
    261.2766, 257.7355, 255.9399, 254.9156, 253.7023, 252.683, 251.2689, 
    251.8006,
  262.5247, 265.3215, 264.0033, 263.6715, 261.1655, 262.3289, 261.5924, 
    258.8268, 258.0913, 255.6035, 257.1654, 257.8587, 255.9759, 253.9682, 
    251.5872,
  267.9325, 265.1882, 262.283, 258.512, 255.204, 260.4875, 261.8193, 
    259.2246, 257.3886, 258.3657, 257.3211, 259.3318, 259.3208, 252.621, 
    250.6082,
  272.6463, 269.7642, 264.2969, 258.0283, 255.9374, 256.6867, 260.8687, 
    258.7915, 258.0287, 258.3514, 258.318, 258.0706, 257.5064, 256.8036, 
    252.7099,
  273.6204, 273.316, 272.8128, 268.3945, 260.1014, 260.2931, 255.1379, 
    257.1521, 257.6877, 256.8416, 256.6536, 256.4699, 255.9438, 258.0504, 
    257.324,
  274.1849, 272.9116, 272.553, 272.1347, 267.8576, 262.1682, 261.7852, 
    252.0535, 252.7283, 252.8775, 255.1835, 255.6422, 255.978, 257.1462, 
    258.4099,
  274.8694, 273.6807, 272.8124, 272.072, 272.0358, 269.9138, 262.9032, 
    260.7653, 259.2113, 259.101, 256.2122, 256.3201, 256.4484, 256.4096, 
    256.2154,
  275.3845, 274.4982, 273.2769, 272.2395, 272.2294, 271.7175, 270.1694, 
    264.5754, 260.8708, 261.9622, 259.7814, 256.2812, 255.6936, 254.463, 
    253.5089,
  275.8536, 274.7817, 273.4017, 272.1639, 272.0915, 270.8967, 269.6075, 
    266.0023, 258.5046, 256.8418, 256.0322, 254.9635, 252.9176, 252.2755, 
    250.8825,
  275.7164, 274.8325, 273.9695, 270.1853, 266.1866, 265.6422, 264.1836, 
    260.7319, 256.8492, 253.3286, 251.732, 253.5362, 252.4417, 250.5995, 
    249.5925,
  272.9717, 270.6259, 268.4306, 262.2444, 258.8739, 257.6407, 257.7254, 
    259.5548, 254.9359, 251.2984, 249.935, 251.6096, 250.7295, 248.5688, 
    249.015,
  259.0594, 260.4117, 256.5064, 259.3853, 255.6192, 255.2365, 257.9043, 
    257.3987, 256.7132, 249.1468, 249.985, 258.6036, 257.0949, 255.3027, 
    258.5386,
  265.8105, 260.4805, 258.4048, 257.0361, 255.6887, 257.7407, 259.4408, 
    257.2072, 252.19, 258.4021, 254.4046, 261.0996, 260.9005, 255.0895, 
    255.2845,
  272.4719, 268.3197, 262.7958, 259.9695, 260.6637, 255.7227, 257.11, 
    255.4373, 254.5572, 256.2429, 258.8556, 259.094, 259.6381, 258.973, 
    256.574,
  273.678, 273.329, 272.6145, 267.1205, 261.2271, 260.644, 251.2829, 
    251.5423, 253.8609, 254.4169, 255.328, 256.6206, 257.6886, 258.6017, 
    258.343,
  274.1769, 272.8907, 272.5331, 271.8012, 265.3416, 262.2036, 261.7845, 
    245.2659, 250.6481, 253.75, 255.0135, 255.5452, 256.0429, 258.6951, 
    258.7129,
  274.847, 273.6166, 272.7477, 272.0458, 271.7437, 268.1479, 262.1685, 
    261.3177, 257.2503, 259.4851, 256.3829, 256.3642, 257.2078, 257.1763, 
    255.9777,
  275.3337, 274.4773, 273.251, 272.1839, 272.187, 271.4533, 269.4818, 
    262.5121, 260.2741, 260.1836, 257.0792, 255.895, 256.1493, 255.8867, 
    254.5617,
  275.8365, 274.7977, 273.3876, 272.1609, 272.2885, 271.0657, 269.7089, 
    265.1411, 257.8497, 255.8587, 254.188, 254.4342, 253.1372, 252.8829, 
    251.042,
  275.7376, 274.8404, 274.0199, 270.6672, 266.7466, 265.8002, 264.3968, 
    258.6823, 254.2146, 250.8972, 249.2766, 250.0955, 249.9244, 249.9766, 
    250.39,
  273.1393, 271.4408, 269.3667, 261.9268, 258.8546, 255.3834, 255.6484, 
    256.2596, 251.246, 247.2048, 247.6308, 249.9058, 250.3784, 249.8964, 
    251.3905,
  258.9599, 260.0194, 256.5262, 256.9224, 253.9537, 253.6313, 256.356, 
    256.8848, 257.4827, 256.0832, 256.148, 260.0696, 259.2657, 258.1195, 
    256.4995,
  264.9008, 261.3712, 258.7211, 256.75, 254.0102, 252.5405, 254.9353, 
    254.8919, 255.3674, 258.742, 256.8945, 260.5026, 260.9635, 256.7428, 
    255.0182,
  272.05, 267.0549, 261.3986, 257.7141, 257.156, 247.5238, 254.4672, 
    255.5285, 255.8209, 255.0048, 257.6074, 257.9246, 259.3516, 259.4714, 
    257.6481,
  273.642, 273.286, 272.1061, 265.8249, 259.8408, 258.3354, 247.1387, 
    248.1539, 251.1411, 252.5932, 253.7141, 256.8236, 256.3668, 257.6071, 
    258.7881,
  274.2054, 272.8127, 272.4681, 271.2745, 263.9833, 262.1783, 262.4992, 
    249.6394, 250.7398, 250.6826, 252.4495, 253.1317, 255.0602, 256.5207, 
    258.2218,
  274.9118, 273.6019, 272.7146, 271.9808, 271.4387, 267.4413, 260.7271, 
    262.0122, 256.6493, 257.5114, 251.5296, 254.9934, 254.683, 256.3849, 
    256.2454,
  275.4428, 274.5507, 273.3087, 272.1409, 272.1616, 271.3582, 268.914, 
    261.1883, 257.4868, 255.5284, 252.6996, 254.758, 255.3109, 256.8565, 
    255.893,
  275.8838, 274.9374, 273.4919, 272.1892, 272.3526, 271.3571, 269.5038, 
    263.1196, 253.7773, 251.5656, 250.5007, 253.8295, 256.6502, 256.7982, 
    254.4882,
  275.8409, 274.9171, 274.0556, 270.9475, 267.0159, 264.7074, 263.0365, 
    256.8624, 252.2203, 250.3148, 248.7681, 249.6612, 253.8672, 254.7075, 
    254.2638,
  273.6508, 271.8488, 269.6584, 260.2981, 257.9695, 252.3379, 251.9772, 
    252.8453, 250.8786, 248.6201, 245.886, 248.3718, 248.5586, 252.0001, 
    252.7183,
  257.1446, 259.8371, 256.472, 258.1072, 256.7612, 255.3257, 255.8961, 
    255.3389, 257.2112, 257.0406, 257.7213, 258.4482, 255.4362, 253.9836, 
    255.2035,
  262.6311, 259.3404, 258.0506, 256.59, 255.8876, 252.231, 255.9941, 
    255.0231, 256.2417, 258.4708, 258.4205, 260.4415, 258.996, 252.8269, 
    252.5828,
  271.9044, 266.2172, 260.8501, 256.4602, 255.3535, 250.1969, 255.7203, 
    255.0676, 255.6481, 257.5635, 259.2833, 260.4654, 259.0002, 257.7046, 
    254.9254,
  273.5775, 273.2525, 272.1338, 265.6521, 258.9377, 259.4004, 253.2591, 
    252.1529, 254.9308, 256.4738, 258.3133, 259.1388, 258.0907, 256.905, 
    257.2379,
  274.2552, 272.7465, 272.4361, 271.1952, 262.9105, 261.9305, 260.9454, 
    250.2016, 251.4174, 255.7072, 256.7426, 256.7979, 256.755, 256.5886, 
    257.7593,
  275.0107, 273.6719, 272.7164, 271.9538, 271.4179, 267.495, 260.3697, 
    259.3002, 256.954, 257.1604, 255.5405, 255.8947, 255.19, 254.8338, 
    255.6999,
  275.6084, 274.6599, 273.3994, 272.0979, 272.1537, 271.4995, 268.7219, 
    260.5423, 256.8301, 255.1909, 255.3875, 255.2905, 254.2491, 254.1177, 
    253.7637,
  275.9572, 275.0901, 273.6525, 272.1901, 272.404, 271.4424, 269.0344, 
    262.2911, 254.5494, 254.0838, 253.8384, 254.7876, 254.1602, 253.5144, 
    252.8084,
  275.9471, 275.0639, 274.0921, 271.2745, 267.3645, 264.0931, 261.2242, 
    255.3647, 252.6819, 252.4753, 251.4452, 251.6873, 253.7288, 252.5448, 
    253.6608,
  274.2874, 272.6759, 270.9753, 263.2744, 259.2817, 256.0779, 254.7262, 
    253.5685, 249.8499, 250.1688, 246.6412, 248.9318, 248.9178, 250.7645, 
    252.7841,
  256.4814, 259.0824, 258.8637, 259.3612, 258.7901, 257.1351, 257.6859, 
    256.9637, 257.5657, 254.8968, 251.9905, 252.1908, 251.8174, 253.3633, 
    254.6246,
  262.6754, 259.5424, 258.9857, 258.2303, 258.0347, 255.9005, 258.4064, 
    257.5533, 257.0442, 257.7173, 254.8237, 255.8172, 257.079, 253.6592, 
    253.7438,
  272.1181, 266.4084, 262.6973, 260.0224, 260.4764, 256.9932, 259.537, 
    257.6502, 256.931, 257.7569, 256.9421, 255.7321, 256.2546, 258.6968, 
    257.5111,
  273.5425, 273.2211, 272.3739, 267.8637, 263.79, 263.2154, 253.5292, 
    255.966, 257.2495, 257.2685, 257.5031, 256.1235, 255.321, 256.8092, 
    259.2628,
  274.2444, 272.6998, 272.4279, 271.693, 265.7359, 262.1342, 260.6368, 
    249.4179, 250.5785, 256.0619, 256.0281, 254.8234, 254.7785, 256.6601, 
    259.1776,
  274.9966, 273.7105, 272.6857, 271.954, 271.5196, 266.9668, 260.524, 
    259.6876, 257.4058, 257.6918, 254.9334, 254.1119, 254.4414, 257.824, 
    257.983,
  275.6129, 274.6842, 273.4223, 272.0561, 272.1027, 271.4176, 268.1345, 
    260.813, 257.9145, 256.2324, 254.8945, 253.776, 254.6176, 257.274, 
    257.3297,
  275.9547, 275.1259, 273.7426, 272.2003, 272.3894, 271.1861, 268.015, 
    260.0216, 256.0698, 254.5016, 253.1042, 252.701, 256.0143, 256.6788, 
    255.0426,
  275.9288, 275.1532, 274.104, 270.8204, 265.0641, 262.6425, 259.7726, 
    255.8024, 254.3739, 252.8994, 252.371, 253.3189, 254.8789, 255.2393, 
    254.2823,
  274.2549, 272.6413, 270.5107, 259.5549, 256.2605, 254.2355, 253.5109, 
    254.2597, 251.6226, 249.9514, 249.2967, 251.5032, 252.3875, 251.7078, 
    251.8233,
  259.8631, 259.602, 258.4859, 256.981, 255.1913, 254.8802, 256.0842, 
    254.4879, 254.2674, 252.8407, 253.3438, 254.9569, 254.5797, 254.4415, 
    252.0469,
  263.8566, 260.6142, 259.3263, 257.3401, 255.6616, 256.2578, 257.2292, 
    255.8933, 255.5175, 257.1531, 256.5771, 257.6141, 259.4334, 253.0672, 
    249.8941,
  272.3206, 266.0375, 262.1095, 258.7659, 257.8625, 253.4015, 257.288, 
    257.3012, 256.8036, 259.0737, 257.9599, 255.8654, 258.6742, 259.5486, 
    253.9097,
  273.4812, 273.1827, 272.3833, 267.7995, 260.8354, 260.1324, 252.3211, 
    255.2179, 257.2099, 256.7222, 254.533, 252.8897, 257.0544, 256.7781, 
    255.0688,
  274.2465, 272.6699, 272.4097, 271.7752, 264.0296, 261.1687, 262.4978, 
    251.405, 251.5724, 249.5391, 249.1008, 253.4269, 256.0222, 256.0371, 
    255.8701,
  274.993, 273.6976, 272.5882, 271.8618, 271.0445, 266.5657, 261.524, 
    260.7713, 256.5405, 255.3032, 250.9687, 255.3428, 255.2436, 254.7302, 
    253.5748,
  275.5454, 274.6288, 273.3394, 271.9743, 272.043, 271.2237, 266.5217, 
    259.2718, 256.3603, 255.3078, 255.3063, 254.1115, 253.2457, 251.0795, 
    249.7432,
  275.8632, 274.9762, 273.5842, 272.2313, 272.255, 270.872, 267.7474, 
    259.6271, 255.1342, 253.8901, 253.3951, 252.6469, 251.0128, 249.2363, 
    247.0558,
  275.7563, 274.9614, 273.9787, 270.161, 266.1605, 263.9921, 260.8808, 
    256.7937, 253.7067, 252.7358, 252.3033, 252.1562, 251.0187, 250.0936, 
    249.964,
  273.9895, 272.5174, 268.8995, 258.4139, 257.166, 255.2672, 254.8063, 
    256.4702, 253.2797, 251.9247, 251.1666, 251.9891, 252.3035, 250.0768, 
    251.2854,
  260.5865, 261.4242, 259.8529, 259.0652, 255.7873, 254.3885, 255.6098, 
    252.9617, 251.0067, 244.9999, 245.461, 247.6796, 245.1874, 245.865, 
    245.3301,
  263.9491, 262.6833, 261.0201, 259.0295, 256.2479, 256.4225, 256.0026, 
    253.5887, 251.9271, 251.2301, 249.7422, 252.8901, 253.4716, 248.3926, 
    248.1439,
  272.2503, 266.8392, 262.1855, 259.8428, 258.2526, 253.2572, 255.3209, 
    253.6996, 251.8295, 252.8725, 253.6181, 254.3464, 256.2003, 257.9372, 
    256.4128,
  273.3944, 273.1481, 271.8246, 266.1934, 259.6409, 259.5916, 251.039, 
    250.9521, 250.7959, 250.7762, 253.1276, 254.5056, 256.8004, 257.717, 
    257.6982,
  274.2358, 272.6151, 272.3757, 271.5047, 261.8523, 259.7968, 260.5553, 
    246.8982, 244.5823, 246.5923, 247.9577, 252.0274, 254.9527, 255.4305, 
    255.6064,
  274.9578, 273.5982, 272.5143, 271.704, 269.4482, 264.4995, 259.2184, 
    260.4949, 254.5621, 255.5688, 248.7714, 251.8553, 252.5246, 251.9902, 
    252.8714,
  275.4601, 274.5579, 273.2831, 271.9399, 272.0033, 270.9772, 264.5993, 
    258.6888, 254.0675, 252.968, 251.8916, 251.0802, 250.2119, 248.8351, 
    249.5666,
  275.8039, 274.8903, 273.5141, 272.2777, 272.2301, 270.8215, 267.5418, 
    257.9006, 252.8826, 250.1703, 248.5898, 248.5047, 247.5258, 246.0618, 
    247.0848,
  275.6418, 274.8291, 273.9008, 271.2233, 268.3838, 265.7605, 260.8128, 
    254.1147, 250.5007, 247.278, 246.4794, 246.5153, 245.8995, 245.7696, 
    245.6443,
  274.1826, 272.9869, 268.9546, 259.1511, 256.8239, 255.0137, 252.9646, 
    253.8003, 248.813, 243.114, 242.3684, 245.9263, 245.792, 245.4556, 
    246.0951,
  259.1696, 261.4662, 261.0815, 260.4169, 256.8549, 255.6836, 256.9158, 
    254.0131, 250.6825, 244.6628, 243.9519, 245.1392, 241.6819, 242.8457, 
    241.4035,
  261.3535, 261.1794, 261.1136, 259.4754, 255.4894, 255.8396, 256.2176, 
    253.1357, 249.1865, 248.5485, 245.8464, 250.5472, 250.8295, 245.1293, 
    245.4049,
  272.0183, 265.3487, 261.3056, 259.0875, 258.1468, 252.0065, 254.501, 
    251.8907, 248.4331, 249.2781, 250.5135, 251.3488, 253.3715, 255.2322, 
    253.9019,
  273.3377, 273.0671, 271.0493, 264.3133, 259.8882, 259.478, 247.7511, 
    248.4393, 247.2389, 246.8423, 249.7892, 251.864, 254.2399, 256.3497, 
    255.948,
  274.2337, 272.5775, 272.3442, 271.0133, 260.7134, 259.6979, 260.4322, 
    245.0948, 240.3021, 245.533, 246.5, 249.6616, 253.8384, 254.113, 254.8605,
  274.9122, 273.4661, 272.4675, 271.3942, 267.8546, 262.6721, 258.631, 
    259.9866, 252.6227, 250.7954, 245.7722, 249.6659, 251.32, 251.0645, 
    251.3873,
  275.3685, 274.4726, 273.2278, 271.8915, 271.9428, 270.5418, 263.0861, 
    256.1115, 251.3916, 249.6348, 249.3356, 249.0358, 248.8915, 247.2036, 
    249.0522,
  275.7612, 274.8595, 273.5012, 272.2733, 272.2286, 270.8979, 267.3734, 
    258.8097, 251.1186, 248.7982, 248.3058, 247.8905, 247.6025, 246.6543, 
    248.1839,
  275.6089, 274.7833, 273.8626, 271.7433, 269.8098, 266.9825, 262.041, 
    253.3018, 249.3477, 246.6534, 245.8897, 246.667, 246.5597, 247.4449, 
    247.5611,
  274.2987, 273.1945, 269.0548, 259.9994, 257.5954, 254.8839, 254.85, 
    251.7941, 247.7038, 241.8185, 240.4769, 244.8396, 245.0281, 244.8661, 
    245.8154,
  259.6088, 260.9905, 259.6631, 257.8233, 255.611, 252.1186, 257.6465, 
    257.0772, 255.9929, 251.918, 250.8458, 250.7971, 246.7553, 245.083, 
    241.0278,
  262.6853, 258.0966, 258.6836, 257.1794, 250.9131, 253.916, 256.8338, 
    255.7285, 254.4804, 254.1733, 251.0314, 251.5514, 250.1384, 240.8517, 
    241.1037,
  271.6891, 264.9216, 259.5443, 256.8665, 256.338, 249.7398, 253.5977, 
    253.4476, 252.7958, 252.8168, 251.4341, 249.6924, 249.8046, 250.6667, 
    250.1256,
  273.2829, 273.0212, 270.635, 262.7473, 258.1106, 259.2571, 246.6338, 
    249.453, 249.2251, 246.7339, 248.4753, 249.1982, 251.0084, 252.8573, 
    253.9211,
  274.2401, 272.5414, 272.2993, 270.0197, 257.627, 259.2943, 259.9664, 
    243.0191, 237.6842, 242.4251, 246.5981, 248.7687, 251.1508, 252.266, 
    254.6588,
  274.936, 273.362, 272.4206, 270.8512, 266.031, 259.8691, 258.0673, 259.646, 
    251.7865, 249.5233, 245.7467, 247.5714, 249.7271, 250.5896, 253.2414,
  275.3643, 274.4428, 273.2061, 271.8224, 271.86, 269.8387, 261.5082, 
    255.4035, 251.1901, 249.6301, 247.9676, 247.225, 247.0747, 248.2503, 
    250.5793,
  275.7715, 274.8869, 273.5242, 272.2494, 272.2341, 270.8599, 266.8486, 
    255.7146, 250.4577, 248.4094, 247.1726, 246.8611, 246.3801, 247.2377, 
    248.9243,
  275.6484, 274.8181, 273.8485, 271.9599, 269.7841, 266.5344, 260.8394, 
    252.7945, 249.9576, 247.611, 247.0508, 247.2189, 247.5155, 247.9093, 
    248.7333,
  274.3793, 273.2914, 269.4502, 262.4212, 258.1624, 255.9212, 255.4554, 
    251.3522, 248.2344, 243.4877, 244.3643, 247.0987, 247.5022, 246.981, 
    248.0615,
  260.4787, 261.7389, 259.4434, 255.556, 251.5312, 250.2576, 254.183, 
    254.7769, 255.8515, 250.6791, 249.0646, 250.8064, 249.675, 245.858, 
    242.1237,
  262.486, 258.3177, 256.7177, 253.7328, 249.0538, 249.3065, 252.0676, 
    252.6048, 253.6681, 254.9178, 250.4764, 251.3992, 251.1046, 239.66, 
    236.286,
  271.0037, 263.5158, 257.1821, 254.2061, 253.5033, 243.0643, 248.4238, 
    250.2092, 251.239, 253.3275, 253.1838, 251.8484, 251.6767, 250.3146, 
    246.6385,
  273.2122, 272.8782, 270.0196, 261.8691, 255.3249, 257.3934, 240.6842, 
    247.0974, 249.6743, 250.1421, 252.5315, 252.719, 253.3748, 252.7577, 
    249.8791,
  274.2428, 272.5255, 272.2618, 268.878, 254.8212, 257.7577, 259.744, 
    240.067, 240.9039, 247.1503, 249.7, 250.9679, 252.0523, 251.7513, 251.2891,
  274.9935, 273.327, 272.3704, 270.3055, 264.8222, 258.3596, 257.4606, 
    258.9108, 252.3751, 251.1552, 248.2931, 249.9489, 250.7002, 250.2424, 
    250.4941,
  275.4125, 274.4478, 273.1986, 271.7609, 271.7667, 269.2777, 258.9603, 
    253.5866, 251.3524, 249.7925, 248.8026, 248.6323, 248.8477, 247.8548, 
    249.0576,
  275.7748, 274.9108, 273.5736, 272.2078, 272.2317, 270.7525, 265.3923, 
    253.8451, 250.2482, 248.3009, 247.8321, 247.5563, 247.5401, 248.0578, 
    249.2243,
  275.6651, 274.8554, 273.8367, 271.9459, 269.6838, 265.1043, 256.8426, 
    251.9609, 249.3303, 247.2109, 246.8884, 247.0326, 247.3419, 247.7156, 
    249.2783,
  274.4764, 273.4926, 269.2017, 260.4489, 255.0113, 252.9314, 251.9942, 
    251.6419, 248.0887, 244.5391, 244.1308, 246.8575, 246.5381, 246.1583, 
    247.4584,
  259.43, 259.0674, 255.6512, 254.7086, 250.8981, 248.1916, 250.6408, 
    250.0411, 251.0863, 244.8849, 243.8487, 246.4203, 244.926, 242.3899, 
    239.8359,
  259.941, 257.1175, 255.6418, 252.4523, 247.2508, 244.4439, 247.5073, 
    247.9252, 248.6007, 250.8872, 245.5333, 249.0529, 249.4653, 237.7634, 
    235.1716,
  269.3198, 261.1945, 255.8955, 253.5664, 251.7647, 239.8668, 244.437, 
    246.3327, 246.4212, 248.7357, 249.5554, 249.4342, 249.7957, 248.466, 
    241.947,
  273.0931, 272.5113, 269.6005, 262.3768, 256.8117, 256.6157, 238.9997, 
    244.118, 247.1406, 245.9697, 247.9007, 248.8513, 249.6482, 248.8516, 
    245.5701,
  274.1941, 272.5106, 272.258, 269.0538, 255.0724, 259.498, 259.0038, 
    238.4008, 240.2622, 244.9521, 246.4517, 247.4182, 249.461, 249.4277, 
    249.9759,
  275.006, 273.3341, 272.2811, 270.0905, 264.8024, 258.3817, 257.4925, 
    258.2664, 252.1586, 250.8656, 246.1339, 247.1986, 248.5393, 249.2088, 
    249.9837,
  275.4402, 274.4828, 273.2253, 271.7039, 271.7394, 268.6773, 258.3528, 
    254.228, 252.2166, 250.4369, 248.5505, 246.9264, 246.1739, 245.8215, 
    247.4581,
  275.7629, 274.9315, 273.6607, 272.1855, 272.2288, 270.7128, 264.3574, 
    253.9148, 251.1255, 249.2879, 247.7287, 246.4572, 244.907, 244.6938, 
    246.2852,
  275.6541, 274.8816, 273.8463, 271.9684, 269.5645, 265.0477, 256.7905, 
    252.7229, 250.2499, 246.772, 245.7189, 245.0279, 244.2809, 244.149, 
    244.7063,
  274.5017, 273.5526, 269.2547, 259.1728, 254.0471, 252.7112, 252.6865, 
    252.2477, 247.5596, 242.2125, 240.5472, 243.9599, 242.8866, 242.5169, 
    243.7603,
  258.1907, 258.8572, 256.3211, 256.3411, 254.7811, 252.9251, 253.1042, 
    252.4525, 252.678, 246.7261, 244.6268, 244.9948, 241.3746, 239.8895, 
    235.9352,
  258.5123, 257.1925, 256.2868, 254.3613, 252.0598, 247.2206, 249.7383, 
    249.7144, 249.5625, 250.1578, 243.9541, 247.0221, 247.6603, 237.2442, 
    235.5956,
  267.7568, 258.9985, 256.3255, 254.6778, 253.7638, 242.1491, 245.4062, 
    247.1383, 246.6226, 247.7644, 247.7554, 247.6464, 248.5591, 248.3302, 
    241.9048,
  272.9007, 272.2509, 268.5122, 259.7621, 256.1412, 256.1417, 239.727, 
    243.6596, 245.2052, 244.0032, 245.6695, 247.1856, 248.6483, 248.9703, 
    245.6466,
  274.1699, 272.4995, 272.2889, 268.5241, 254.555, 258.3133, 258.0126, 
    239.1371, 237.1562, 241.128, 243.9848, 246.1634, 248.4506, 248.9447, 
    249.0916,
  275.0352, 273.3286, 272.1402, 269.5504, 264.0786, 256.6103, 258.4141, 
    258.1757, 250.0672, 246.4512, 242.1488, 245.1972, 247.0725, 247.761, 
    247.9451,
  275.4847, 274.5575, 273.2603, 271.6219, 271.6607, 267.8269, 258.3606, 
    253.6946, 249.3132, 246.9578, 244.9672, 244.3293, 244.1843, 244.4803, 
    245.1619,
  275.7812, 274.9828, 273.7733, 272.2065, 272.2206, 270.5521, 263.4162, 
    252.7909, 248.5755, 245.2345, 243.6667, 242.9806, 241.9991, 242.8808, 
    245.1833,
  275.6859, 274.9523, 273.8826, 271.894, 269.4733, 265.0724, 257.09, 
    251.2084, 247.34, 243.5492, 242.6883, 242.4181, 242.4361, 243.8966, 
    245.6364,
  274.5453, 273.5621, 269.5274, 260.6513, 257.1375, 255.075, 252.8393, 
    250.2941, 245.4331, 239.503, 239.3989, 243.4092, 243.8689, 245.283, 
    247.1755,
  258.8004, 259.1078, 256.8472, 257.411, 258.3888, 256.613, 256.8646, 
    257.1333, 258.7336, 255.4659, 253.773, 254.0701, 251.723, 250.4962, 
    246.875,
  259.409, 258.6281, 257.847, 258.2368, 257.3169, 253.2266, 254.5882, 
    254.9165, 255.9276, 256.4686, 252.4887, 253.248, 252.9126, 245.2023, 
    242.5052,
  266.8798, 260.2284, 258.7259, 258.8072, 258.4747, 248.5589, 250.6363, 
    251.8451, 252.2074, 253.1056, 252.2798, 251.3003, 251.4602, 250.6313, 
    245.1383,
  272.7533, 272.4661, 267.744, 260.0857, 258.1843, 258.3276, 245.1137, 
    247.8513, 248.0655, 247.4878, 248.5539, 248.9895, 249.8479, 249.5839, 
    246.6244,
  274.1421, 272.4673, 272.3308, 266.7253, 255.8648, 256.8748, 258.3817, 
    239.6915, 236.8975, 242.1297, 244.9446, 247.5254, 248.2108, 248.2407, 
    248.6624,
  275.0616, 273.3067, 271.9774, 268.5518, 262.6186, 255.8023, 258.0801, 
    257.9146, 249.2823, 245.4091, 241.6819, 244.4211, 245.4341, 246.347, 
    246.6989,
  275.518, 274.5852, 273.2843, 271.5101, 271.4725, 267.1614, 257.7515, 
    252.0389, 247.3236, 245.9536, 244.5235, 243.2775, 243.2804, 243.9831, 
    244.1166,
  275.7961, 274.9697, 273.8119, 272.2352, 272.1394, 270.4814, 261.7361, 
    251.0146, 247.6323, 246.057, 244.7638, 244.1455, 243.0312, 242.8265, 
    244.4766,
  275.7237, 275.0088, 273.9028, 271.8769, 269.4856, 264.8893, 256.1817, 
    251.5233, 249.5602, 248.8624, 248.4287, 248.2074, 247.3742, 247.7602, 
    247.0798,
  274.6536, 273.6475, 270.3719, 263.0328, 257.5746, 254.9988, 253.5034, 
    252.9224, 251.9377, 249.9093, 251.0732, 251.8335, 250.3188, 250.0193, 
    249.4837,
  259.6781, 260.6625, 258.83, 258.9066, 260.173, 258.3745, 260.6538, 
    261.8452, 263.7401, 260.904, 260.9009, 262.8369, 261.6283, 260.2476, 
    257.3708,
  259.592, 260.7215, 260.1227, 261.8474, 260.0248, 255.4794, 256.7141, 
    259.6638, 261.6363, 262.9886, 260.1108, 262.096, 262.3113, 256.9912, 
    254.4223,
  266.4127, 262.7101, 261.3254, 262.7239, 261.6755, 252.9832, 254.2203, 
    255.1156, 257.5823, 259.7875, 260.1452, 260.1577, 260.3246, 260.0181, 
    255.7889,
  272.8208, 272.808, 268.7046, 262.2997, 261.9383, 261.7914, 250.0261, 
    252.033, 251.9096, 254.1541, 256.2878, 256.6939, 257.1088, 256.3901, 
    254.6369,
  274.121, 272.4713, 272.4021, 266.6713, 259.8199, 260.5043, 261.3893, 
    243.9802, 241.0144, 247.6457, 251.1571, 252.9212, 254.4314, 254.2656, 
    253.6877,
  275.1059, 273.3383, 271.9311, 268.6966, 262.6949, 258.39, 259.0488, 
    258.6301, 249.6194, 246.5628, 244.8225, 247.601, 250.5598, 251.2695, 
    251.3522,
  275.5497, 274.614, 273.3408, 271.5339, 271.5219, 267.657, 258.0262, 
    253.2361, 248.8948, 247.2242, 244.8407, 244.7483, 245.9493, 247.3173, 
    248.0689,
  275.7971, 274.9461, 273.8324, 272.2658, 272.0612, 270.8011, 263.165, 
    254.8827, 255.1941, 251.0238, 247.2492, 245.2798, 243.7906, 243.448, 
    247.6083,
  275.7317, 274.9977, 273.8853, 271.5831, 269.1044, 264.7765, 258.6472, 
    255.9743, 254.3759, 253.6851, 252.3282, 249.8186, 247.0997, 246.2874, 
    246.2421,
  274.7303, 273.7089, 269.5036, 262.622, 259.8992, 258.3505, 256.9821, 
    255.3775, 252.0756, 249.197, 253.3465, 253.8645, 250.7313, 249.3187, 
    248.1377,
  259.5938, 263.5518, 258.9337, 259.3853, 262.0176, 257.8409, 258.6132, 
    260.4178, 262.1269, 258.2808, 257.8349, 263.5099, 260.3489, 261.0625, 
    257.5914,
  261.1052, 262.9237, 260.3318, 261.9106, 261.3174, 255.6868, 256.492, 
    259.1756, 262.9087, 263.5103, 259.7782, 263.8396, 264.1777, 260.4861, 
    257.7878,
  267.3782, 265.3337, 261.7117, 262.8511, 262.4826, 253.5352, 254.7867, 
    255.9019, 257.5066, 260.7038, 262.4824, 262.8291, 263.4555, 263.4121, 
    259.8583,
  273.0147, 273.0616, 270.1289, 262.2192, 263.6103, 262.9471, 249.5713, 
    253.1927, 253.7963, 254.2548, 258.2271, 260.8243, 261.9709, 261.7815, 
    260.4412,
  274.1268, 272.5185, 272.6017, 266.9779, 261.6205, 263.1075, 262.3784, 
    243.3296, 243.8206, 249.031, 251.3436, 255.9242, 258.882, 260.4222, 
    260.6281,
  275.072, 273.422, 271.9735, 268.8012, 265.6946, 264.5045, 262.4502, 
    260.2638, 251.4242, 247.7519, 245.7257, 249.0498, 252.8492, 256.7229, 
    258.7005,
  275.5351, 274.6837, 273.4427, 271.5466, 271.5645, 269.1668, 262.1134, 
    257.4688, 255.6942, 251.4269, 246.4602, 245.4711, 246.9328, 249.5406, 
    254.1833,
  275.8289, 274.9994, 273.874, 272.2881, 271.9821, 270.9241, 263.6721, 
    256.9346, 256.6613, 255.4934, 252.2045, 245.2322, 243.7567, 244.7115, 
    248.5964,
  275.7318, 275.0174, 273.8571, 271.2771, 268.0079, 262.3917, 256.2407, 
    252.72, 251.7468, 250.8457, 248.8431, 249.3437, 246.7396, 244.3615, 
    244.5607,
  274.7761, 273.7292, 270.0489, 262.9868, 257.6908, 253.7775, 252.7635, 
    251.8601, 249.879, 247.709, 249.109, 248.9283, 246.471, 244.0277, 243.7136,
  260.6398, 261.2549, 259.6977, 257.6264, 257.1772, 250.1156, 251.7934, 
    255.6342, 260.2357, 260.028, 257.1023, 260.4227, 259.4512, 255.4312, 
    254.0698,
  262.1429, 261.3932, 260.3196, 261.3967, 259.019, 247.26, 250.3139, 
    251.9923, 257.0998, 259.6954, 260.3753, 264.377, 264.8841, 258.5468, 
    255.7169,
  267.4194, 263.7004, 262.2266, 262.6028, 261.934, 250.7954, 248.5342, 
    249.8963, 251.6787, 253.9176, 256.925, 259.7121, 262.4601, 263.516, 
    261.6289,
  273.008, 272.9493, 270.1448, 263.9321, 263.4439, 262.232, 248.4958, 
    249.1505, 250.3648, 249.8622, 251.6972, 255.4436, 257.7211, 258.5811, 
    258.1513,
  274.1067, 272.5584, 272.7067, 268.096, 262.8687, 263.9033, 262.7494, 
    244.3853, 241.5215, 246.7003, 247.7769, 250.2171, 253.6694, 255.7412, 
    257.377,
  275.0268, 273.4484, 271.9856, 269.5355, 265.5479, 263.2354, 263.7091, 
    262.3289, 253.7701, 248.9159, 244.1622, 246.923, 248.916, 251.5704, 
    254.4405,
  275.5017, 274.681, 273.4585, 271.5561, 271.4033, 268.7962, 262.3599, 
    258.656, 255.7488, 254.362, 247.9169, 245.4005, 245.8439, 247.0103, 
    250.1438,
  275.8221, 274.9937, 273.8809, 272.2979, 271.9348, 271.0087, 263.4387, 
    257.3928, 254.7284, 255.2172, 252.0139, 245.4328, 243.6728, 244.5862, 
    247.2084,
  275.7133, 275.0349, 273.8633, 271.5786, 269.1722, 265.153, 259.4631, 
    255.4399, 254.2249, 252.0711, 250.9737, 246.5248, 243.5224, 243.663, 
    245.3651,
  274.8387, 273.8339, 271.3484, 265.7158, 261.1992, 259.1758, 257.2859, 
    255.999, 252.5266, 251.2, 252.9408, 247.7918, 242.9536, 242.627, 243.8527,
  260.4153, 260.601, 259.5498, 260.2839, 259.2316, 252.535, 251.0961, 
    252.3159, 258.5429, 260.6726, 260.3444, 262.0056, 260.5826, 252.6794, 
    251.8049,
  265.1947, 261.2311, 261.0304, 261.6637, 260.0303, 251.1383, 250.3828, 
    250.1261, 253.2506, 257.8323, 259.9854, 263.5287, 262.9988, 258.9315, 
    254.0759,
  268.1478, 264.4604, 262.1292, 263.4637, 262.509, 253.8992, 249.5099, 
    248.7114, 249.8901, 251.7717, 253.5881, 256.4331, 258.1589, 259.7172, 
    255.7322,
  273.0378, 272.7518, 270.1215, 265.3316, 264.4427, 262.7045, 253.2398, 
    248.4379, 249.2431, 248.7281, 250.7711, 252.0187, 252.7576, 252.9495, 
    251.9332,
  274.1052, 272.6221, 272.7359, 269.2259, 264.6198, 264.2521, 263.4354, 
    255.6407, 253.5568, 246.5816, 247.2484, 249.0677, 250.5176, 250.896, 
    251.547,
  275.0144, 273.4684, 272.1119, 270.2728, 266.5842, 264.3688, 264.0709, 
    263.3047, 256.0044, 251.2623, 245.9175, 246.5076, 247.4837, 248.6922, 
    250.0664,
  275.4741, 274.6529, 273.4396, 271.5092, 271.1707, 268.9217, 263.7617, 
    260.2627, 256.6051, 252.9223, 248.8759, 246.5434, 245.2127, 245.7212, 
    248.7094,
  275.8087, 274.9757, 273.8539, 272.3075, 272.1031, 271.1729, 265.3426, 
    259.4661, 254.8416, 252.5024, 249.3709, 247.882, 243.3445, 244.3581, 
    248.4043,
  275.6962, 275.0258, 273.9124, 271.9695, 270.7615, 267.8021, 263.4123, 
    258.0514, 253.6098, 252.157, 248.7492, 248.4699, 242.5574, 243.9671, 
    247.8237,
  274.8717, 273.8909, 271.99, 268.372, 266.1717, 265.1483, 261.6178, 
    256.2777, 251.9432, 249.8121, 249.6235, 246.6727, 242.1373, 242.9602, 
    246.311,
  266.5439, 264.6774, 261.337, 260.9308, 256.513, 255.1918, 256.9372, 
    258.7992, 261.8239, 260.2247, 259.9045, 260.6326, 259.5923, 256.1285, 
    253.0727,
  266.9889, 265.159, 261.4611, 260.2429, 255.1287, 252.3137, 256.1183, 
    257.8327, 260.0284, 262.0286, 261.2427, 262.7991, 262.4353, 249.8884, 
    251.8482,
  270.0323, 267.4024, 263.9798, 263.037, 259.8144, 250.1751, 253.6763, 
    255.5292, 257.5544, 258.4493, 259.4359, 259.8552, 258.2026, 257.1497, 
    248.0327,
  273.0482, 272.6327, 270.0876, 264.6514, 262.2987, 261.6577, 250.9744, 
    253.4012, 254.3809, 255.2259, 256.186, 254.9761, 254.0509, 252.1127, 
    248.9071,
  274.128, 272.656, 272.7462, 269.0863, 262.0106, 262.8805, 262.1261, 
    249.5895, 249.0818, 250.7515, 252.4255, 252.6962, 252.1749, 250.8078, 
    250.4683,
  275.0578, 273.5025, 272.1226, 269.9714, 264.8948, 262.35, 263.021, 
    262.9366, 258.717, 254.5793, 250.1348, 249.7417, 248.7573, 248.2378, 
    249.0487,
  275.516, 274.6724, 273.427, 271.3319, 270.4788, 268.2745, 262.624, 
    261.2745, 258.175, 254.7393, 251.5823, 248.7775, 246.2613, 245.759, 
    248.3423,
  275.8459, 274.9921, 273.8447, 272.2765, 272.1154, 271.1838, 264.627, 
    259.6599, 256.1375, 253.008, 250.1934, 247.8025, 243.6658, 244.7509, 
    248.5396,
  275.7488, 275.0577, 273.9308, 272.111, 271.3296, 268.3214, 263.2994, 
    259.0208, 254.562, 251.4305, 248.8299, 245.7105, 242.6738, 244.4734, 
    247.7997,
  275.0108, 273.9426, 272.0958, 267.2232, 263.5083, 264.3096, 262.2171, 
    257.2631, 252.3113, 249.3486, 247.3087, 244.7651, 242.198, 243.7429, 
    246.9771,
  267.3691, 266.361, 265.5461, 264.2054, 258.0256, 251.0632, 254.8842, 
    256.9943, 258.8, 255.9777, 256.5318, 256.9198, 255.2807, 253.2158, 
    248.8688,
  267.837, 267.0732, 266.2478, 263.1862, 255.6834, 248.874, 252.0004, 
    255.5001, 258.419, 259.8636, 258.8098, 259.8577, 259.148, 250.9849, 
    249.1748,
  269.6921, 267.663, 266.2772, 263.5048, 259.3261, 247.1438, 250.3279, 
    254.0302, 257.9332, 260.3087, 261.0014, 260.3502, 259.6114, 258.5676, 
    253.2354,
  272.9974, 272.4644, 270.4538, 264.7583, 261.5797, 260.3322, 249.1026, 
    253.2249, 256.6364, 258.8332, 259.2859, 258.679, 257.8383, 256.3087, 
    252.6238,
  274.1426, 272.6883, 272.7962, 268.8646, 258.6025, 261.1599, 262.8043, 
    248.6703, 249.7007, 255.0258, 256.2654, 256.0794, 255.6705, 254.4866, 
    252.8358,
  275.0849, 273.5493, 272.1193, 270.0241, 260.8665, 258.0605, 262.4564, 
    262.839, 259.1288, 257.0618, 254.0331, 253.6838, 253.2978, 252.6119, 
    251.1418,
  275.5274, 274.6919, 273.406, 271.2036, 269.6307, 266.9979, 261.6427, 
    260.0454, 257.2792, 255.9866, 253.7069, 252.2474, 250.7722, 249.6792, 
    249.2866,
  275.8454, 274.9804, 273.7867, 272.2245, 272.0728, 270.8065, 261.5439, 
    257.9783, 255.1763, 253.761, 251.6278, 250.1426, 246.8863, 246.707, 
    248.2023,
  275.7414, 275.0467, 273.91, 272.046, 271.1954, 266.6958, 259.3856, 
    256.5177, 253.0379, 250.596, 248.946, 247.3875, 244.3337, 245.5576, 
    247.0123,
  275.0955, 273.9959, 272.0558, 265.1299, 259.5369, 259.7523, 257.3287, 
    254.6597, 251.1216, 247.9411, 246.2887, 246.0441, 243.1948, 244.2306, 
    246.0378,
  269.5026, 268.8225, 268.4525, 267.941, 266.9363, 264.939, 263.0189, 
    261.3358, 260.1566, 256.2009, 255.1867, 255.674, 254.4336, 254.2958, 
    251.218,
  269.4416, 269.1334, 268.6007, 267.583, 265.3025, 259.6059, 258.5428, 
    257.0888, 257.4237, 256.7875, 255.9731, 258.0602, 258.1295, 252.0875, 
    250.2323,
  270.1181, 268.8595, 267.5454, 266.503, 264.1872, 255.7367, 256.7991, 
    257.4971, 256.025, 256.1873, 257.1875, 258.0943, 258.7675, 259.1112, 
    255.3946,
  273.0111, 272.584, 270.3035, 266.0015, 264.0949, 260.9439, 251.7346, 
    254.1112, 253.1488, 254.0225, 255.9218, 257.536, 258.749, 258.7556, 
    256.1418,
  274.1392, 272.6956, 272.7742, 267.9512, 262.8317, 262.8606, 262.3989, 
    249.0466, 245.021, 252.5457, 255.3719, 257.4911, 258.5023, 258.4144, 
    256.9712,
  275.0396, 273.4754, 272.1024, 269.2672, 264.6027, 260.7212, 261.8297, 
    261.1631, 257.7299, 255.9142, 255.1288, 256.8021, 257.464, 257.2066, 
    256.4873,
  275.443, 274.5836, 273.3282, 270.9185, 269.7782, 266.0115, 259.7465, 
    258.8434, 257.1168, 256.9518, 256.4355, 256.4403, 256.1546, 255.7399, 
    255.3491,
  275.7605, 274.8918, 273.7112, 272.156, 272.0025, 269.6756, 259.3861, 
    256.9862, 255.9384, 255.5662, 255.409, 255.1291, 254.2037, 254.2401, 
    253.8466,
  275.6409, 274.9759, 273.8524, 271.9621, 270.4688, 264.7497, 257.4765, 
    255.5483, 254.1536, 253.6612, 253.3495, 253.11, 251.9488, 251.8578, 
    250.2944,
  274.9916, 273.9548, 271.4405, 261.5417, 256.1399, 257.1428, 255.8391, 
    254.2792, 252.4126, 250.8542, 250.3618, 250.8586, 249.2874, 248.3464, 
    247.9785,
  264.3358, 262.3791, 260.4057, 260.3383, 261.5548, 257.0281, 255.8687, 
    257.3257, 258.4814, 257.8019, 257.7218, 259.1094, 258.9014, 259.6219, 
    258.3502,
  264.0065, 262.346, 260.1769, 260.3132, 259.4236, 255.9386, 254.1843, 
    252.6494, 254.3076, 256.1425, 255.2288, 257.9478, 257.0878, 251.7597, 
    255.0326,
  268.2289, 262.3528, 259.8756, 260.3922, 260.7096, 252.476, 253.5418, 
    253.2438, 253.8622, 255.2157, 256.7593, 257.9617, 258.3131, 258.8868, 
    257.3067,
  272.9469, 272.4271, 268.9489, 262.6563, 262.2708, 260.6881, 249.5482, 
    251.0373, 253.2644, 254.7963, 256.2881, 258.3123, 258.6568, 259.0453, 
    257.8289,
  274.1102, 272.6678, 272.7306, 266.6061, 261.1039, 261.4104, 260.8491, 
    244.3804, 246.0229, 253.487, 256.06, 257.1478, 258.8604, 259.0278, 
    258.1323,
  275.0084, 273.4359, 272.061, 268.5543, 262.7639, 259.9985, 260.3384, 
    259.7118, 256.8571, 256.7462, 255.3529, 256.811, 257.9611, 257.879, 
    256.8889,
  275.4133, 274.54, 273.2697, 270.7678, 269.6962, 264.1729, 258.1872, 
    257.2684, 256.8877, 257.683, 257.3987, 257.2904, 257.2272, 256.9031, 
    256.5619,
  275.739, 274.8636, 273.6464, 272.0772, 271.9624, 268.0775, 256.876, 
    255.5133, 255.1342, 256.0605, 256.721, 256.9626, 256.35, 256.0801, 
    256.0102,
  275.6364, 274.96, 273.8119, 271.6809, 268.8613, 261.0751, 255.5925, 
    254.6906, 254.0922, 253.8924, 254.4501, 254.7406, 254.2417, 254.0659, 
    252.7429,
  275.0131, 273.9332, 271.0094, 260.4691, 253.9536, 253.6024, 254.0386, 
    253.8486, 252.6492, 251.027, 251.1238, 252.3503, 251.9409, 251.5846, 
    250.7054,
  267.1716, 263.2942, 259.3987, 257.3455, 256.7599, 252.7489, 252.6857, 
    252.4543, 254.868, 254.0029, 255.545, 257.0833, 256.6121, 255.2825, 
    254.4698,
  268.1913, 263.5404, 260.9297, 257.3423, 255.8974, 250.3767, 252.6434, 
    251.5736, 253.7766, 256.117, 256.025, 258.8506, 258.9989, 251.741, 
    253.5859,
  270.0583, 264.5409, 262.3533, 258.4672, 258.7979, 248.0598, 251.7263, 
    254.1367, 255.5419, 257.1696, 258.2154, 259.3288, 259.4422, 258.6344, 
    259.8053,
  272.932, 272.6781, 270.1263, 260.7535, 261.7522, 258.0241, 247.101, 
    251.5848, 255.0218, 257.3139, 258.8138, 259.3371, 259.3143, 258.938, 
    258.7901,
  274.1384, 272.6972, 272.7773, 265.9466, 259.0055, 259.056, 258.5872, 
    243.5465, 249.3925, 256.1855, 258.2049, 258.5667, 259.0164, 258.2988, 
    258.5195,
  275.037, 273.4773, 272.0882, 268.7695, 262.4637, 258.4942, 258.4707, 
    256.4102, 255.0306, 257.1088, 256.0365, 257.6021, 258.3383, 257.8684, 
    257.4309,
  275.4385, 274.5774, 273.2784, 271.0444, 270.4068, 263.9914, 256.5424, 
    253.7547, 253.5344, 254.8996, 254.7464, 255.7945, 256.3602, 256.1641, 
    256.1165,
  275.7588, 274.9169, 273.6664, 272.0618, 271.9692, 267.4458, 255.0897, 
    252.6698, 251.6754, 252.1864, 252.6291, 253.2476, 253.1422, 253.5259, 
    253.5817,
  275.6654, 274.9988, 273.8475, 271.8841, 269.5391, 260.3301, 254.4426, 
    251.9079, 250.4831, 249.4986, 249.894, 250.3921, 250.7157, 250.9065, 
    250.6274,
  275.0444, 273.9981, 272.2333, 268.946, 262.4441, 255.0748, 253.1642, 
    252.1897, 249.1738, 245.5689, 246.1705, 248.742, 248.6233, 248.9569, 
    249.7081,
  272.4455, 270.3125, 265.7239, 259.7213, 253.9937, 249.8455, 248.7894, 
    250.1204, 256.0867, 254.8494, 256.2732, 257.5027, 255.0526, 253.2183, 
    248.9969,
  272.3829, 269.9299, 265.1559, 258.0833, 252.4408, 248.6283, 249.6878, 
    250.1663, 254.0297, 255.9905, 255.8476, 259.4399, 258.9755, 250.444, 
    244.9212,
  272.0077, 269.8389, 264.9496, 259.2435, 256.74, 247.0605, 249.059, 
    251.4552, 255.0717, 256.583, 257.1792, 257.4774, 256.7822, 255.8604, 
    252.8981,
  273.008, 272.6795, 269.5547, 261.4797, 260.404, 257.0796, 245.0016, 
    250.7092, 253.6911, 256.1076, 257.3882, 257.006, 256.6591, 256.643, 
    257.4054,
  274.2119, 272.7737, 272.8297, 265.9432, 260.0587, 260.1339, 258.7277, 
    244.6128, 250.1244, 253.5623, 255.9939, 257.0775, 258.2823, 258.5537, 
    259.0059,
  275.0881, 273.5443, 272.0823, 268.4543, 262.3859, 259.1873, 259.5145, 
    256.5919, 252.6753, 255.2285, 253.7388, 255.9878, 257.2658, 257.2346, 
    257.6181,
  275.4813, 274.6636, 273.2794, 270.5536, 269.5861, 262.9922, 257.6154, 
    253.5372, 252.1793, 252.7576, 252.5227, 254.3957, 255.2343, 255.7778, 
    256.4871,
  275.7869, 274.9526, 273.7076, 272.0658, 271.9691, 266.9494, 256.194, 
    253.1174, 250.8574, 250.1529, 250.4453, 251.6504, 252.3253, 253.9848, 
    254.4858,
  275.6729, 275.0151, 273.9025, 272.2638, 270.91, 262.2312, 255.1084, 
    252.549, 250.1745, 248.8179, 249.175, 250.1351, 250.8532, 252.4242, 
    253.601,
  274.9923, 273.9767, 272.1117, 267.7691, 261.6054, 256.7401, 254.2479, 
    252.9773, 250.3322, 247.1016, 247.3678, 250.134, 251.1359, 252.5, 253.6561,
  260.9599, 257.9031, 255.2676, 254.6004, 253.4953, 252.7623, 253.9178, 
    248.7867, 251.1697, 248.1497, 249.8076, 252.8124, 251.5941, 249.4843, 
    247.1681,
  261.722, 258.1299, 256.9372, 255.0309, 253.9311, 252.1835, 254.2723, 
    250.8476, 251.2057, 250.5767, 249.6655, 253.5649, 253.9952, 245.436, 
    244.2781,
  268.6425, 260.4238, 258.58, 258.5208, 257.882, 248.4196, 252.7691, 
    253.4775, 255.3015, 253.944, 253.5725, 254.1452, 253.5882, 252.9955, 
    250.125,
  272.8957, 271.3744, 266.6506, 260.2231, 261.587, 259.681, 250.2144, 
    253.6121, 255.3785, 256.6731, 257.6458, 256.6579, 255.319, 254.6923, 
    252.6794,
  274.1315, 272.6917, 272.4397, 264.5256, 261.213, 261.373, 260.8783, 
    246.9533, 250.4477, 255.2516, 257.1027, 258.727, 259.0191, 257.8202, 
    256.4374,
  274.9734, 273.393, 271.8238, 266.9809, 262.1273, 259.7936, 259.7504, 
    258.3078, 256.0253, 256.7451, 255.3314, 256.9402, 258.2315, 258.3076, 
    257.7332,
  275.3852, 274.5092, 273.125, 270.018, 269.0494, 261.5229, 258.2785, 
    256.7127, 256.0091, 256.1512, 256.5267, 256.4804, 257.0273, 257.6273, 
    258.0382,
  275.6936, 274.8172, 273.6031, 272.0057, 271.7979, 264.8845, 257.8197, 
    256.4568, 255.4641, 255.3941, 256.2202, 257.2891, 256.5432, 257.34, 
    257.7262,
  275.5786, 274.8906, 273.8834, 272.3489, 269.9733, 261.6926, 257.9075, 
    256.5609, 255.6988, 255.3686, 255.1569, 256.869, 257.5673, 257.7591, 
    258.7493,
  274.8896, 273.9593, 272.0927, 265.5419, 260.0628, 258.836, 257.1022, 
    257.6334, 255.5409, 253.9203, 253.7389, 255.354, 257.1969, 258.2813, 
    259.1978,
  260.6612, 259.5373, 259.8752, 259.5754, 254.0597, 250.5457, 250.7972, 
    250.3324, 250.8753, 245.8155, 245.5979, 249.4847, 250.2693, 250.6588, 
    250.3581,
  261.2411, 258.5789, 259.7155, 259.0103, 255.3057, 250.5965, 251.9609, 
    250.7394, 252.251, 249.9273, 246.2463, 250.9682, 254.6788, 246.9767, 
    247.6035,
  268.6479, 261.9407, 260.0821, 260.4779, 259.7817, 248.6604, 251.5799, 
    252.5113, 254.0201, 253.5255, 251.8744, 251.7866, 253.2551, 255.1533, 
    253.0041,
  272.8059, 271.686, 267.4766, 261.5757, 261.7722, 259.2473, 248.9751, 
    251.4926, 253.855, 253.6722, 254.8825, 253.2098, 252.5109, 254.4255, 
    253.6125,
  274.0961, 272.6627, 272.0824, 264.1687, 260.8606, 260.1237, 259.4547, 
    245.3231, 248.5216, 251.9686, 253.0046, 253.6294, 253.0698, 253.3279, 
    254.3201,
  274.9075, 273.3331, 271.5778, 266.7773, 263.068, 259.1603, 258.1293, 
    256.1891, 255.1426, 255.4307, 250.1993, 253.2074, 254.6785, 253.0503, 
    253.1036,
  275.3388, 274.443, 272.9879, 269.8426, 269.0577, 260.5249, 257.2573, 
    254.5074, 254.7758, 256.5207, 254.4164, 253.5552, 252.4124, 252.1367, 
    252.2051,
  275.639, 274.7419, 273.5096, 271.9862, 271.2229, 262.3202, 256.7672, 
    253.6895, 252.4698, 254.4166, 256.7665, 254.9229, 252.7404, 253.6735, 
    252.0789,
  275.5239, 274.8087, 273.8095, 272.0161, 266.0287, 258.2513, 256.7906, 
    254.2093, 252.5905, 253.4249, 254.2792, 257.0511, 255.8735, 254.4439, 
    253.9805,
  274.8053, 273.8088, 270.764, 260.3401, 254.8441, 254.9814, 254.3687, 
    257.1588, 254.0696, 251.356, 251.3942, 254.5425, 257.2469, 257.457, 
    256.0044,
  260.8344, 257.6029, 257.4727, 256.989, 252.5001, 249.8268, 249.5446, 
    251.1424, 251.8709, 249.826, 249.4869, 249.8641, 247.2825, 247.159, 
    246.6594,
  259.584, 257.1951, 259.2419, 258.5055, 254.995, 247.1465, 247.6621, 
    249.1485, 250.4962, 252.3519, 250.3378, 251.7066, 253.1434, 246.2754, 
    246.0483,
  267.9873, 258.7915, 256.3967, 258.5504, 258.7138, 246.9976, 247.9688, 
    249.2204, 250.0447, 250.4697, 251.5202, 251.9137, 252.4694, 253.841, 
    251.1201,
  272.7105, 271.1733, 266.0932, 257.7874, 260.1746, 256.6748, 245.4408, 
    249.0706, 251.0269, 253.6126, 253.6361, 252.9898, 252.7616, 254.2621, 
    252.8959,
  274.0734, 272.6405, 271.6358, 261.8291, 258.5529, 258.5706, 256.6526, 
    240.5637, 243.9038, 253.634, 253.5334, 252.3525, 252.373, 253.9891, 
    256.085,
  274.8615, 273.2952, 271.1035, 264.6456, 261.0267, 257.9079, 257.0345, 
    253.6899, 253.2227, 254.8023, 252.1051, 251.7582, 251.533, 253.9937, 
    255.5658,
  275.3037, 274.3824, 272.8051, 268.7818, 268.0089, 258.2939, 256.0163, 
    253.4427, 254.2536, 255.5894, 254.1889, 251.4771, 250.0098, 251.2697, 
    254.5042,
  275.5945, 274.6768, 273.3913, 271.9253, 269.9676, 258.4855, 255.3257, 
    253.7575, 253.785, 255.0414, 254.9641, 251.8834, 250.1987, 250.8887, 
    252.8329,
  275.4858, 274.7327, 273.7351, 270.9006, 261.1939, 254.0381, 253.8663, 
    253.9347, 253.9142, 255.2009, 254.9249, 253.143, 249.9451, 250.4862, 
    252.238,
  274.7397, 273.5959, 268.8953, 256.5496, 251.6212, 251.2423, 251.5301, 
    257.8227, 255.7282, 253.1616, 252.9024, 254.4777, 252.5429, 250.3473, 
    251.0837,
  257.9643, 256.359, 254.4302, 253.3769, 252.8536, 249.7096, 249.1526, 
    248.2792, 249.2503, 246.8241, 251.0113, 251.8082, 248.4862, 247.7899, 
    246.8901,
  257.239, 255.2402, 255.1535, 253.5363, 251.9892, 244.9232, 246.315, 
    247.3459, 248.2895, 250.9505, 251.7511, 253.5495, 253.918, 249.4822, 
    245.4434,
  265.3192, 255.3743, 255.4823, 255.8508, 255.3383, 243.9139, 246.1498, 
    246.4402, 246.9222, 249.1234, 251.9475, 252.8347, 252.7713, 252.3591, 
    248.9868,
  272.4302, 269.8875, 263.6051, 255.5347, 259.5165, 255.4169, 242.1294, 
    247.936, 249.2374, 250.8473, 252.5708, 253.6593, 253.6528, 253.7711, 
    251.9993,
  274.0398, 272.6067, 271.1606, 259.1046, 256.7083, 257.5324, 255.756, 
    239.0868, 242.7602, 253.8003, 254.8163, 253.5419, 252.9224, 253.3984, 
    254.386,
  274.8412, 273.2698, 270.6057, 263.1634, 259.7527, 256.633, 256.2057, 
    254.6437, 252.9848, 253.4457, 251.0191, 251.444, 251.7208, 252.4838, 
    253.2255,
  275.3129, 274.3712, 272.6871, 268.5099, 267.5318, 256.687, 253.9724, 
    252.9766, 252.977, 252.6774, 250.6256, 249.1362, 249.0186, 250.2803, 
    252.3838,
  275.6018, 274.6898, 273.3539, 271.8842, 269.1413, 256.8921, 253.1555, 
    252.2554, 251.2979, 250.6353, 249.5744, 248.8998, 248.2547, 250.378, 
    252.379,
  275.5175, 274.733, 273.7512, 270.5943, 261.1125, 254.7148, 252.7405, 
    252.4203, 251.4375, 250.5155, 248.8315, 249.1976, 248.7023, 251.0126, 
    252.3804,
  274.7895, 273.6048, 269.4061, 259.8495, 255.0423, 253.8687, 252.8767, 
    258.796, 254.8568, 248.3091, 245.4107, 248.0434, 248.8167, 251.0091, 
    252.069,
  255.8112, 253.9482, 252.1409, 252.0758, 249.7414, 245.9064, 246.9535, 
    247.6462, 248.3606, 245.8712, 248.4586, 251.3006, 249.8592, 250.5214, 
    251.0263,
  255.4733, 254.2256, 253.4666, 252.9279, 250.5595, 246.31, 248.1742, 
    248.6521, 249.7864, 249.805, 249.3891, 251.8441, 252.9238, 248.6076, 
    248.4859,
  264.5616, 256.9147, 255.8119, 257.0121, 256.6557, 248.4927, 249.3361, 
    249.1053, 249.2971, 249.907, 251.1833, 252.4292, 252.5819, 252.4088, 
    249.9982,
  272.3496, 269.9356, 265.4708, 259.5405, 261.3406, 258.4985, 251.289, 
    251.6786, 251.2949, 251.8883, 252.7626, 253.0576, 252.686, 252.4112, 
    250.581,
  274.0518, 272.6389, 271.9215, 263.5452, 262.331, 261.7618, 259.6518, 
    248.6517, 248.4271, 253.7717, 255.6631, 254.8245, 254.066, 254.0023, 
    253.7146,
  274.8823, 273.3126, 271.2852, 266.6805, 265.2756, 262.7704, 260.6389, 
    257.9575, 255.2596, 253.9191, 253.6432, 254.5516, 254.2392, 254.1185, 
    253.9785,
  275.3447, 274.4152, 272.8989, 269.8413, 269.5443, 263.157, 259.2749, 
    257.2768, 254.7863, 253.5305, 252.223, 252.4481, 253.3504, 253.3448, 
    253.819,
  275.6213, 274.7337, 273.3808, 271.9268, 270.3308, 262.5194, 258.1492, 
    255.7892, 253.6167, 252.1815, 251.3221, 250.5125, 250.6998, 252.0049, 
    252.8006,
  275.5439, 274.7465, 273.7694, 271.0026, 264.4467, 259.6198, 256.6027, 
    255.1492, 253.4284, 251.7658, 250.2079, 249.3562, 249.691, 250.9269, 
    251.3881,
  274.8233, 273.4397, 270.3768, 263.996, 260.3374, 257.3997, 254.6297, 
    257.4389, 254.9517, 250.0983, 248.5207, 248.7762, 248.2898, 249.5376, 
    250.1806,
  258.7963, 258.4424, 258.7744, 258.8214, 256.5471, 251.9182, 251.421, 
    250.0732, 249.6226, 245.7924, 246.9855, 248.3146, 246.1128, 247.1131, 
    245.2956,
  260.0986, 259.6239, 259.9375, 260.234, 257.425, 255.6631, 256.2794, 
    256.328, 254.1612, 253.4212, 253.2394, 253.5903, 252.6714, 248.5679, 
    247.1252,
  267.5082, 263.3466, 263.951, 265.5009, 262.9861, 261.469, 258.7087, 
    255.9414, 254.8333, 254.279, 253.7061, 254.9831, 253.8475, 252.7435, 
    251.1005,
  272.6729, 271.9062, 270.5418, 268.3108, 266.7047, 263.5661, 256.4066, 
    255.5265, 255.6537, 255.5367, 255.7432, 254.7532, 254.1599, 255.1386, 
    254.1912,
  274.0219, 272.6967, 272.7393, 268.8305, 266.0013, 263.7417, 261.2047, 
    250.926, 250.6951, 255.5913, 256.8593, 255.4624, 254.8844, 254.7421, 
    254.8843,
  274.8271, 273.368, 271.8315, 268.684, 266.3513, 262.5391, 261.0933, 
    257.6909, 253.7658, 250.1006, 252.2336, 253.2371, 253.4536, 253.9198, 
    254.3815,
  275.3047, 274.4081, 272.9798, 270.3276, 269.8531, 262.2134, 257.9666, 
    255.0224, 252.8186, 249.9873, 249.2574, 249.7389, 250.6322, 251.209, 
    252.2886,
  275.6078, 274.7161, 273.346, 271.9153, 269.8503, 258.5659, 252.9126, 
    250.5643, 249.9861, 249.1653, 249.0951, 249.2446, 249.6214, 249.6911, 
    250.6584,
  275.5302, 274.7365, 273.7358, 270.187, 260.7695, 254.5117, 251.1045, 
    250.9918, 251.4072, 251.9189, 250.0421, 248.9606, 248.8004, 249.1503, 
    249.1496,
  274.7581, 273.0882, 269.3007, 259.4597, 254.5565, 251.5212, 249.9803, 
    254.4348, 254.0123, 249.6079, 249.5217, 248.62, 246.4905, 247.0586, 
    247.9381,
  259.1216, 257.5306, 257.9857, 258.6227, 261.6372, 262.1972, 265.5913, 
    262.4041, 259.5857, 254.7055, 255.8359, 255.4968, 251.6699, 250.2198, 
    248.1423,
  259.2369, 258.7725, 259.0841, 260.6042, 261.8218, 260.8578, 265.2902, 
    260.3276, 259.739, 258.308, 258.2841, 259.5206, 258.728, 255.7382, 254.736,
  268.0066, 262.6867, 263.1107, 265.3153, 266.4744, 263.8415, 259.7612, 
    257.9323, 256.1799, 255.5114, 255.4023, 257.2383, 257.1549, 257.1472, 
    255.3228,
  272.8485, 272.6227, 271.6309, 268.4015, 266.5385, 262.1584, 252.2568, 
    253.8526, 253.9313, 253.5916, 254.6716, 254.7788, 255.1294, 255.913, 
    256.6478,
  274.0129, 272.7959, 272.887, 267.1522, 261.3809, 259.671, 257.4654, 
    247.555, 249.3093, 253.5344, 255.827, 254.7755, 254.2419, 254.7574, 
    256.081,
  274.8333, 273.3862, 271.7548, 266.4233, 262.4336, 255.339, 253.2961, 
    251.7136, 250.1312, 247.9436, 250.3282, 252.7641, 252.8152, 253.2641, 
    253.8721,
  275.3148, 274.4349, 272.9177, 269.6022, 268.7963, 255.0677, 250.8396, 
    249.7113, 248.8768, 248.1793, 248.1181, 248.8481, 249.2964, 249.2899, 
    249.5176,
  275.6248, 274.7191, 273.3468, 271.8697, 268.7473, 254.6362, 250.9795, 
    250.2059, 249.937, 249.2942, 248.6291, 248.7723, 248.4946, 248.2899, 
    248.8996,
  275.5365, 274.7294, 273.6751, 269.1196, 257.2006, 252.9794, 251.593, 
    251.9549, 252.4173, 252.4267, 248.9592, 247.4444, 248.5814, 249.4444, 
    248.7545,
  274.751, 272.6334, 267.6136, 256.0881, 252.6248, 252.1895, 251.7416, 
    255.1297, 255.1219, 249.2632, 248.8019, 247.1893, 247.9169, 249.5996, 
    247.7515,
  262.4104, 261.0229, 259.4676, 258.6266, 257.7945, 257.6598, 260.3863, 
    261.252, 260.2466, 255.7185, 253.0901, 250.92, 248.6836, 249.4995, 
    248.6963,
  262.7704, 261.5593, 260.292, 259.5471, 257.6307, 257.742, 259.9851, 
    258.453, 253.7752, 251.7405, 249.9082, 250.4205, 250.2093, 248.4793, 
    248.8636,
  268.8803, 263.7057, 261.9597, 261.5456, 261.7857, 259.2908, 258.2792, 
    255.4653, 251.8292, 251.3409, 250.9917, 250.7628, 250.8018, 250.2575, 
    249.7058,
  272.8828, 272.7766, 271.7002, 267.0188, 265.1195, 263.6876, 253.8304, 
    252.4568, 251.0893, 251.0664, 251.8647, 251.5507, 250.9413, 250.5944, 
    249.4793,
  274.0205, 272.83, 272.9242, 267.5908, 264.5459, 263.317, 258.731, 247.9903, 
    246.1197, 251.0813, 253.2518, 251.6353, 250.585, 250.6566, 250.7793,
  274.8338, 273.3404, 271.8057, 268.3794, 265.4282, 261.0051, 258.3695, 
    253.3687, 249.7478, 247.2105, 247.9314, 250.4727, 250.6619, 250.4483, 
    250.0412,
  275.332, 274.4733, 272.9844, 270.1606, 269.6948, 260.915, 254.3125, 
    250.6249, 249.9948, 249.3969, 250.8187, 250.851, 250.7431, 249.8194, 
    249.325,
  275.654, 274.7784, 273.4254, 271.9008, 269.721, 256.4568, 252.2749, 
    250.4474, 251.1293, 250.8879, 250.9124, 250.3441, 249.0898, 248.1821, 
    249.1798,
  275.6115, 274.7719, 273.6811, 269.9735, 260.0558, 254.3722, 252.1894, 
    252.1999, 253.4983, 252.9817, 248.9648, 247.446, 247.4494, 248.6012, 
    249.1032,
  274.854, 273.3583, 269.1545, 260.1382, 254.2358, 252.3631, 250.9503, 
    254.3257, 255.3372, 248.7723, 247.3183, 244.7065, 245.7459, 249.2017, 
    249.3094,
  264.5597, 263.5631, 262.5639, 261.7055, 259.9709, 259.2642, 259.4214, 
    258.5158, 258.2756, 257.705, 258.4965, 259.0467, 257.6158, 257.1524, 
    254.8467,
  264.6449, 263.3595, 262.5901, 260.7199, 259.1959, 259.0776, 259.6169, 
    258.6995, 258.3653, 258.6444, 257.848, 257.3604, 256.3411, 254.5927, 
    253.3005,
  268.8559, 264.3456, 262.4004, 261.5307, 260.9439, 256.7001, 259.071, 
    259.6631, 258.6336, 258.8668, 258.31, 257.5345, 256.5147, 255.3845, 
    254.4662,
  272.882, 272.451, 270.9302, 265.3814, 261.9087, 262.316, 256.0069, 
    258.9497, 259.6732, 259.425, 259.0225, 258.1902, 256.9239, 255.3506, 
    254.2507,
  274.0646, 272.8646, 272.9351, 267.9417, 262.6097, 262.8721, 261.7906, 
    256.1867, 256.4406, 258.8711, 260.2286, 258.7583, 256.8262, 255.4349, 
    254.2083,
  274.8525, 273.3274, 271.9633, 268.9623, 265.4322, 262.7557, 262.3697, 
    260.7576, 259.8803, 256.7237, 255.4726, 256.1982, 254.7438, 253.4625, 
    252.3048,
  275.3399, 274.4544, 273.0287, 270.3381, 269.6726, 264.4842, 262.6479, 
    261.0073, 258.5481, 255.8596, 254.5514, 253.4045, 253.0745, 250.8174, 
    249.5535,
  275.6346, 274.7586, 273.4129, 271.9176, 271.2283, 265.6425, 263.3476, 
    260.5003, 257.607, 254.7849, 253.6898, 252.2646, 249.8235, 248.7476, 
    248.9613,
  275.6441, 274.7978, 273.7301, 271.4501, 267.8158, 265.4121, 263.2662, 
    259.5625, 257.4221, 255.0138, 251.0081, 248.614, 247.6004, 246.9927, 
    247.4872,
  274.9017, 273.6321, 271.1395, 267.5251, 265.3915, 262.3197, 259.565, 
    258.0498, 256.4901, 248.8311, 244.1672, 244.3395, 244.589, 246.2788, 
    247.9898,
  265.2407, 264.655, 264.241, 263.4622, 262.3985, 261.3045, 261.1509, 
    261.8748, 260.889, 258.5152, 258.6937, 259.2385, 257.0804, 257.3098, 
    256.1159,
  265.8554, 265.4879, 265.1444, 263.7401, 262.3611, 261.5816, 260.8547, 
    260.6625, 260.6155, 260.0595, 259.5453, 259.9607, 258.8253, 256.1897, 
    255.6126,
  269.5488, 265.511, 264.7527, 264.9228, 264.1034, 260.4671, 261.1271, 
    260.4164, 260.6535, 259.6844, 259.1986, 258.8715, 258.311, 257.5377, 
    256.8464,
  272.8311, 272.342, 271.1923, 267.148, 265.0611, 264.0728, 257.884, 
    260.0178, 260.3773, 259.5041, 259.0091, 258.757, 258.3327, 257.3204, 
    257.3863,
  274.1109, 272.9225, 272.9753, 268.5276, 264.0911, 264.3839, 262.5997, 
    256.2508, 255.9038, 258.1102, 260.3705, 259.5936, 258.4316, 257.6749, 
    257.6768,
  274.9167, 273.416, 272.0124, 268.7128, 264.7787, 263.2885, 262.5927, 
    260.185, 257.8189, 255.7437, 256.5744, 257.8457, 257.4153, 257.6111, 
    257.5686,
  275.4204, 274.5158, 273.0392, 269.9416, 268.4223, 263.1436, 261.1203, 
    259.2512, 257.0551, 256.5127, 256.0602, 255.3411, 255.7601, 255.3629, 
    256.1335,
  275.6591, 274.794, 273.3772, 271.8714, 271.0383, 262.8331, 260.675, 
    259.137, 257.1339, 255.966, 255.4472, 256.2641, 255.6097, 254.0623, 
    253.8522,
  275.6313, 274.8133, 273.7004, 271.1104, 265.7036, 262.5968, 261.0765, 
    259.6352, 257.5172, 255.3708, 251.4986, 250.2571, 249.7628, 247.4077, 
    245.2555,
  274.8259, 273.4722, 269.4967, 262.8073, 260.3853, 258.5766, 256.8068, 
    257.1457, 253.0178, 246.4415, 243.1129, 243.0754, 242.4653, 242.8893, 
    243.6976,
  266.6662, 265.8494, 266.7137, 266.0796, 264.5416, 263.9706, 264.7679, 
    265.0001, 264.6272, 263.026, 262.164, 262.5446, 260.8984, 260.0053, 
    259.036,
  266.7181, 267.0807, 266.7684, 264.7794, 263.6586, 264.028, 263.735, 
    262.7918, 264.3935, 263.8695, 263.1497, 263.1228, 262.519, 258.9758, 
    257.2568,
  270.4225, 267.1086, 265.6111, 264.5765, 263.9777, 262.0739, 263.573, 
    263.3231, 262.46, 262.7432, 261.8461, 260.4107, 259.96, 259.2355, 258.4691,
  272.8213, 272.598, 271.3565, 266.1214, 264.1214, 264.1099, 259.5803, 
    262.3239, 261.2523, 260.6715, 259.6963, 259.7014, 259.2991, 259.8675, 
    258.9178,
  274.0953, 272.8992, 272.942, 266.2263, 262.4672, 263.5448, 263.4403, 
    255.926, 257.4993, 259.826, 260.855, 259.9257, 259.0993, 258.6923, 
    258.8838,
  274.845, 273.3827, 271.8083, 266.2119, 261.6289, 260.3186, 261.1981, 
    261.049, 260.3691, 259.7314, 259.4423, 259.9179, 259.6001, 259.3685, 
    258.5893,
  275.3443, 274.4104, 272.8641, 267.7722, 265.0426, 257.7712, 257.502, 
    258.1472, 258.5263, 258.4823, 258.2683, 258.1768, 258.2601, 257.8526, 
    258.1138,
  275.5777, 274.6741, 273.2542, 271.7759, 268.2446, 256.3762, 255.2922, 
    254.1641, 254.293, 253.7989, 253.6747, 254.0224, 253.9143, 254.1076, 
    254.2897,
  275.4993, 274.6783, 273.5836, 268.9317, 257.3884, 253.9603, 252.8754, 
    252.0845, 250.427, 248.5673, 246.4964, 247.2046, 247.4878, 247.3605, 
    246.3638,
  274.6461, 273.1447, 267.3923, 255.5079, 251.0011, 250.0111, 250.6884, 
    254.0674, 249.8515, 244.5471, 243.043, 244.005, 243.7451, 243.9005, 
    243.304,
  262.8457, 260.9058, 261.7915, 260.8709, 258.848, 258.6263, 259.3712, 
    258.6811, 259.2944, 259.7358, 260.9621, 262.2207, 262.0786, 261.9429, 
    261.5314,
  262.6438, 262.1123, 261.6675, 260.4267, 257.0616, 257.5588, 257.1198, 
    256.7075, 256.9452, 258.4185, 260.5415, 262.2247, 262.3345, 260.4638, 
    260.4189,
  270.2337, 264.4969, 261.838, 260.5218, 257.7277, 253.261, 256.0173, 
    255.6254, 256.387, 258.2184, 259.8706, 260.6726, 260.3238, 260.3566, 
    259.8286,
  272.8689, 272.7013, 271.3868, 264.7553, 259.555, 257.3508, 249.741, 
    253.5951, 256.5064, 256.6988, 257.8372, 258.1749, 258.6573, 258.9029, 
    258.966,
  274.1049, 272.873, 272.9084, 265.9138, 260.1693, 258.4537, 257.2456, 
    245.6997, 249.5348, 255.0329, 256.6074, 256.0188, 255.7166, 256.3931, 
    257.5929,
  274.8058, 273.3521, 271.8102, 266.684, 260.8587, 256.7111, 255.6729, 
    253.8008, 252.5063, 252.5381, 251.814, 253.4299, 253.7896, 254.9016, 
    256.0229,
  275.3073, 274.3656, 272.871, 268.6702, 264.5992, 255.3721, 252.5674, 
    252.248, 251.3647, 251.3456, 250.9316, 250.6158, 251.0038, 251.973, 
    253.6138,
  275.5743, 274.6795, 273.2563, 271.763, 266.9468, 253.4585, 250.9479, 
    249.9024, 249.8878, 249.6348, 249.0453, 249.4285, 247.9811, 249.3885, 
    250.7191,
  275.5232, 274.702, 273.6381, 269.6367, 257.5933, 252.2829, 250.9904, 
    250.8368, 250.3498, 249.1511, 247.5337, 247.7917, 245.999, 246.7149, 
    247.9374,
  274.6352, 273.3915, 269.7022, 259.8926, 252.4566, 250.6643, 251.2744, 
    253.3939, 251.1248, 246.9896, 245.6607, 245.7503, 244.1011, 244.8359, 
    245.2243,
  264.8893, 263.8517, 263.0027, 262.5679, 261.2498, 261.4761, 263.0127, 
    260.7621, 259.2281, 257.5973, 256.8898, 256.5677, 254.5369, 253.6516, 
    253.097,
  262.6357, 262.1246, 262.3506, 262.264, 261.3349, 262.11, 261.0873, 
    259.8036, 258.7809, 256.8547, 256.3398, 257.1352, 255.6349, 253.1065, 
    251.7918,
  270.0504, 266.0499, 262.3899, 262.046, 260.109, 257.2448, 258.6647, 
    258.042, 256.2415, 257.3542, 258.067, 257.4006, 256.2868, 254.3527, 
    252.4332,
  272.9554, 272.7169, 271.502, 266.3748, 261.0115, 260.4518, 257.5938, 
    258.5398, 259.4582, 258.135, 257.0754, 255.1962, 254.3393, 252.9578, 
    250.9723,
  274.1466, 272.8748, 272.9607, 268.1123, 263.7215, 265.0367, 264.6922, 
    254.2625, 248.722, 252.3008, 254.005, 252.3304, 251.8183, 250.9123, 
    250.7083,
  274.836, 273.3611, 271.926, 266.7899, 262.9958, 260.7258, 257.9347, 
    254.6561, 250.5364, 247.3195, 247.4725, 249.1021, 249.5267, 249.3947, 
    249.3484,
  275.2837, 274.3084, 272.5962, 264.6499, 260.5052, 254.9001, 252.6735, 
    249.9007, 247.6824, 246.9909, 247.0486, 247.4215, 247.4364, 247.0243, 
    247.8922,
  275.5087, 274.5955, 273.1731, 271.2973, 263.8176, 252.627, 249.8555, 
    247.5482, 247.3495, 247.307, 246.4454, 246.651, 245.1919, 245.7591, 
    247.0466,
  275.424, 274.5644, 273.5081, 267.9715, 254.8753, 250.7261, 249.0011, 
    248.3969, 248.1172, 246.7942, 245.1685, 245.1669, 244.6513, 244.8006, 
    245.7554,
  274.4088, 273.2493, 266.8887, 253.4785, 249.6702, 248.9576, 248.7456, 
    251.6105, 249.3391, 245.6894, 244.8634, 244.8186, 244.0981, 244.038, 
    244.3133,
  266.2425, 265.6275, 264.7428, 264.7109, 266.1557, 266.9893, 267.4908, 
    266.3989, 265.7478, 265.047, 264.7604, 264.7415, 263.2065, 262.3463, 
    260.6259,
  265.6638, 264.9796, 264.5334, 264.5434, 264.3059, 264.2355, 264.738, 
    264.7026, 264.6047, 264.7791, 263.7532, 264.342, 263.4007, 261.1355, 
    259.8646,
  270.2657, 266.1344, 264.4563, 263.7309, 263.0385, 259.9138, 261.4659, 
    261.7562, 262.0367, 263.4814, 263.9907, 263.1946, 262.6186, 262.2739, 
    260.6829,
  272.953, 272.617, 271.103, 265.7383, 262.2428, 262.1606, 259.6958, 
    260.6643, 260.884, 260.6547, 259.8384, 258.0534, 257.4886, 256.2997, 
    253.9946,
  274.1727, 272.8688, 272.9378, 266.7178, 261.8473, 263.3929, 264.1403, 
    255.8383, 253.0513, 253.9181, 255.2915, 253.5012, 252.4738, 251.6478, 
    250.4848,
  274.7953, 273.2926, 271.372, 262.5304, 259.0561, 257.3907, 258.2021, 
    257.3609, 252.4987, 249.0594, 248.3752, 249.5541, 249.0108, 248.4874, 
    247.555,
  275.2055, 274.1847, 271.6212, 261.0301, 258.1143, 253.8371, 252.5278, 
    251.1236, 248.4673, 248.1802, 247.3058, 247.0436, 247.4748, 247.5179, 
    247.4379,
  275.4654, 274.5112, 273.0882, 271.0057, 262.6296, 251.8745, 249.1712, 
    247.9184, 248.0765, 248.0498, 247.1755, 247.4229, 247.4781, 248.1214, 
    248.5841,
  275.4224, 274.5074, 273.5287, 269.2848, 258.017, 253.7244, 251.8431, 
    251.0189, 250.4655, 250.2706, 250.1235, 249.6905, 249.4557, 249.5574, 
    249.0586,
  274.3942, 273.3874, 269.2917, 259.7312, 256.0674, 254.53, 252.8325, 
    253.2884, 253.3216, 252.8206, 253.8773, 252.5094, 251.7712, 252.1113, 
    251.5562,
  264.6592, 262.6892, 262.9083, 264.006, 267.8942, 268.6088, 269.4053, 
    268.5178, 269.3113, 268.2831, 267.9532, 268.4333, 267.6087, 266.375, 
    266.124,
  263.661, 262.606, 262.8318, 264.1349, 265.5603, 267.5012, 268.0684, 
    268.4359, 269.0964, 268.7143, 268.0823, 268.1158, 267.3751, 265.0943, 
    264.5744,
  269.8364, 265.2261, 263.9928, 264.1202, 264.0514, 262.6792, 266.6181, 
    268.29, 268.9378, 268.807, 268.3284, 267.3642, 266.7735, 266.2789, 
    264.6499,
  272.9149, 272.666, 271.0306, 264.1982, 263.524, 264.8367, 263.2237, 
    265.8152, 267.323, 267.621, 267.662, 266.552, 266.1389, 264.868, 263.7723,
  274.1511, 272.8314, 272.5522, 263.2281, 261.5776, 263.2891, 265.4301, 
    261.1682, 260.0291, 265.1084, 266.2554, 265.1356, 264.5935, 263.6693, 
    262.8305,
  274.8324, 273.3003, 270.8427, 261.2659, 260.44, 260.5416, 261.9134, 
    263.3997, 262.4417, 263.0284, 263.2255, 263.0153, 262.7855, 261.8768, 
    260.538,
  275.2611, 274.2339, 271.7979, 263.3034, 261.1882, 258.8136, 258.7995, 
    259.5434, 260.7817, 261.2379, 260.5677, 260.4464, 260.1405, 259.6061, 
    257.9314,
  275.4991, 274.5634, 273.1455, 271.2862, 264.7582, 255.3759, 255.0181, 
    255.739, 256.2597, 257.7843, 258.203, 257.9756, 257.4809, 257.0959, 
    255.851,
  275.4832, 274.5391, 273.6133, 271.1758, 264.7645, 257.5627, 254.1616, 
    254.0769, 254.5583, 254.9308, 255.4182, 255.5841, 255.2631, 254.2342, 
    253.0265,
  274.3776, 273.4853, 272.048, 269.2463, 266.7564, 260.8561, 254.7614, 
    252.6691, 252.5695, 252.0809, 254.6939, 253.9027, 253.4246, 253.608, 
    252.6586,
  260.9147, 259.0072, 258.2674, 261.5195, 265.3336, 265.364, 264.3879, 
    262.19, 260.9261, 264.9815, 261.8655, 265.5195, 265.4269, 264.2748, 
    263.0304,
  262.608, 261.5587, 261.0428, 263.9178, 264.7466, 264.3844, 264.5199, 
    260.6625, 264.9725, 263.9795, 263.2829, 267.2099, 267.1518, 266.4273, 
    262.8465,
  270.6693, 266.3844, 264.3458, 264.8049, 263.502, 264.3238, 265.9572, 
    262.5645, 267.6724, 267.8365, 268.0863, 267.8283, 268.4877, 268.1825, 
    266.0997,
  272.916, 272.7374, 272.155, 266.0941, 263.937, 266.0278, 263.9316, 
    264.5284, 268.1406, 267.998, 267.9897, 267.0894, 267.2645, 266.7527, 
    264.6231,
  274.192, 272.8549, 272.7159, 264.2975, 263.218, 265.8365, 268.1992, 
    265.6404, 265.1392, 267.081, 267.7453, 265.94, 266.1771, 264.7171, 
    264.1661,
  274.8706, 273.3582, 271.4435, 264.257, 264.0308, 264.3765, 265.46, 
    266.4154, 266.3282, 266.34, 266.1547, 266.6581, 265.0673, 262.5366, 
    262.0996,
  275.3018, 274.2596, 272.4755, 267.8691, 265.4504, 263.3114, 265.2173, 
    264.6583, 265.9794, 266.7751, 265.8256, 266.195, 264.2882, 262.6982, 
    260.8703,
  275.4898, 274.5724, 273.1647, 271.6111, 267.0751, 262.0934, 261.7244, 
    262.1704, 264.6186, 265.5384, 265.4191, 265.9117, 264.0492, 261.9456, 
    259.4933,
  275.4741, 274.5065, 273.6378, 271.603, 268.2873, 265.4649, 259.8762, 
    262.4438, 263.0357, 263.7751, 265.3735, 265.549, 263.5808, 260.6349, 
    258.2123,
  274.0003, 272.3876, 269.2792, 266.2061, 268.4, 265.8689, 261.0811, 
    259.8312, 261.5498, 262.2865, 264.0797, 265.009, 262.8974, 260.0839, 
    258.7976,
  263.4403, 261.6751, 260.0878, 261.6962, 261.4827, 258.8357, 261.894, 
    262.5667, 262.6957, 264.527, 261.6078, 263.2551, 263.0839, 262.6795, 
    260.8434,
  264.6704, 263.7505, 263.0406, 261.813, 262.1452, 258.5176, 260.2926, 
    261.6534, 264.4206, 259.2783, 262.2247, 263.9424, 264.7364, 263.6223, 
    258.6528,
  271.02, 267.4683, 264.1356, 263.4605, 261.9326, 258.9397, 258.2966, 
    257.6553, 261.7146, 261.4873, 265.8653, 265.813, 265.442, 264.6101, 
    262.8092,
  273.0164, 272.78, 272.1509, 265.9778, 262.9641, 262.3266, 260.3213, 
    259.9283, 266.0942, 265.5008, 261.2643, 263.102, 264.8386, 265.8542, 
    265.2893,
  274.0905, 272.8073, 272.6193, 264.2244, 263.1494, 263.9582, 264.8078, 
    262.3922, 258.2354, 259.9085, 263.1689, 265.4453, 266.0268, 266.2816, 
    266.0745,
  274.7198, 273.2893, 271.2037, 264.496, 263.8439, 264.3376, 264.5679, 
    263.7266, 262.028, 264.2225, 260.9034, 265.0578, 266.0891, 265.9528, 
    263.8976,
  275.1939, 274.1296, 272.3307, 266.0507, 265.8204, 262.9761, 266.9414, 
    259.7493, 263.4819, 266.2628, 264.12, 264.6342, 265.3777, 263.8763, 
    258.5986,
  275.4001, 274.3998, 273.0263, 271.5958, 268.1662, 261.9098, 261.1832, 
    263.9034, 263.6337, 265.7884, 263.6854, 264.2231, 262.652, 257.8365, 
    253.0533,
  275.3804, 274.3777, 273.4512, 269.7448, 266.8981, 264.6774, 261.0375, 
    262.2039, 265.108, 264.5529, 263.3402, 262.7267, 257.9383, 253.8831, 
    252.1246,
  272.8926, 270.1717, 264.8889, 258.5331, 264.0257, 266.0149, 262.947, 
    264.6832, 263.5311, 263.3327, 262.3007, 259.1952, 255.4152, 253.3392, 
    252.8145,
  262.2574, 259.122, 256.9444, 257.7267, 261.6333, 262.2524, 260.897, 
    263.0356, 264.0122, 262.5397, 262.3483, 264.2555, 262.9067, 262.5276, 
    260.9782,
  263.5565, 260.048, 258.4686, 258.7066, 261.457, 260.8197, 262.2704, 
    263.1588, 263.1105, 262.9351, 261.9463, 264.5318, 264.5899, 260.4211, 
    258.8407,
  271.1882, 266.779, 261.6777, 259.7309, 259.1165, 260.2081, 259.7581, 
    260.6952, 257.143, 258.6623, 263.6471, 264.6555, 263.4528, 262.6112, 
    258.8833,
  273.0678, 272.8069, 272.2226, 263.5295, 260.5089, 261.616, 259.3052, 
    257.8394, 260.4238, 261.7011, 262.0603, 263.1744, 262.2415, 260.7239, 
    259.2201,
  274.028, 272.7515, 272.4825, 264.0121, 261.6508, 262.5047, 263.9442, 
    254.3123, 257.3996, 258.6238, 261.9427, 262.3348, 261.1125, 259.933, 
    258.4822,
  274.6693, 273.2456, 271.2025, 265.9889, 264.9541, 263.2461, 263.8572, 
    264.2258, 260.4338, 262.226, 260.0468, 261.4121, 259.8539, 257.9486, 
    256.0091,
  275.1227, 274.0446, 272.4166, 268.5388, 266.6567, 262.1749, 262.2153, 
    261.4163, 261.4292, 261.2323, 261.3437, 260.1652, 257.5839, 254.3658, 
    252.5477,
  275.3884, 274.3077, 272.8871, 271.6535, 268.9276, 262.2477, 260.0104, 
    260.9319, 259.5046, 260.7841, 259.0962, 256.1029, 253.243, 251.1884, 
    250.3297,
  275.3771, 274.3611, 273.172, 267.855, 264.8043, 263.4726, 259.5654, 
    259.4268, 261.6162, 258.1969, 254.9376, 252.7378, 250.7929, 250.3593, 
    250.3265,
  272.0804, 268.8717, 264.1064, 259.5811, 260.3958, 260.5273, 259.8206, 
    259.4169, 259.6479, 255.9136, 252.4089, 250.6224, 250.1293, 250.1175, 
    251.0812,
  264.1294, 260.8277, 259.5364, 262.2245, 261.4364, 259.1692, 257.8833, 
    260.0049, 260.7996, 259.5551, 259.3129, 260.856, 259.7747, 259.4532, 
    256.8244,
  265.6437, 262.2114, 261.7124, 262.1073, 260.7208, 256.0506, 256.8264, 
    258.7039, 258.1333, 259.2393, 258.1902, 260.7535, 261.595, 257.7089, 
    256.6306,
  271.6338, 268.193, 264.3646, 263.9204, 259.5689, 256.217, 254.5643, 
    257.3425, 256.7497, 257.5531, 257.9575, 259.2551, 260.5034, 261.0331, 
    258.9101,
  273.1191, 272.8336, 272.2304, 265.1183, 261.768, 259.9296, 251.6279, 
    254.5663, 255.7788, 255.7529, 255.4341, 256.1852, 257.6634, 258.6843, 
    259.6507,
  274.0688, 272.7872, 272.1478, 263.5208, 261.4596, 260.8348, 259.1836, 
    250.4274, 251.1048, 253.7672, 254.4035, 254.0018, 255.045, 255.8868, 
    257.5467,
  274.745, 273.2213, 271.0786, 266.4108, 264.2371, 260.4811, 259.4242, 
    259.1529, 255.4264, 256.0633, 252.7401, 253.1986, 252.7377, 253.1399, 
    254.5533,
  275.1872, 274.0844, 272.3992, 268.921, 265.1073, 259.4433, 255.5806, 
    254.3462, 254.3544, 253.4508, 252.0291, 251.7782, 251.6211, 251.211, 
    251.6167,
  275.5311, 274.4417, 272.8774, 271.5728, 268.263, 260.1887, 254.937, 
    252.6169, 251.1551, 250.8244, 249.9281, 250.0934, 249.9526, 250.1673, 
    249.9767,
  275.5401, 274.5079, 273.2482, 267.8585, 265.78, 263.5751, 255.8397, 
    252.7878, 250.5011, 248.9311, 248.2468, 248.8721, 248.5975, 249.2635, 
    249.8258,
  273.3187, 270.725, 266.4364, 262.8655, 262.6288, 262.1324, 256.9604, 
    254.386, 250.9953, 248.0397, 247.5218, 248.0659, 247.5214, 248.0967, 
    250.0058,
  270.4998, 266.5532, 263.4181, 263.7397, 261.9478, 258.9768, 257.3646, 
    256.4405, 256.1381, 255.6144, 255.2911, 257.6304, 255.6956, 255.7138, 
    255.4378,
  270.0447, 268.7886, 265.5664, 264.2931, 263.6129, 259.9294, 258.5184, 
    257.26, 256.704, 257.2002, 255.4273, 257.0789, 258.4174, 253.2897, 
    251.8337,
  272.0103, 270.798, 268.1245, 265.9231, 262.9731, 258.4762, 258.5525, 
    257.1342, 256.8359, 256.4509, 256.2523, 256.5207, 257.8075, 258.0726, 
    254.4865,
  273.1538, 272.8438, 272.414, 267.5108, 264.3133, 261.6074, 256.3464, 
    256.5428, 256.556, 256.0302, 255.6134, 255.1932, 255.974, 256.5534, 
    256.1791,
  274.173, 272.8095, 272.6024, 267.225, 264.6982, 262.4662, 260.6491, 
    252.6187, 251.3512, 255.4453, 255.5965, 254.8803, 254.5554, 254.8256, 
    256.4388,
  274.8683, 273.2365, 271.5502, 267.7016, 265.9932, 262.8187, 260.7298, 
    260.4902, 258.3291, 257.6855, 255.6397, 255.0722, 253.7192, 253.6135, 
    254.2335,
  275.3321, 274.1848, 272.6091, 269.4967, 265.7559, 261.8174, 260.0536, 
    259.2116, 258.5271, 257.9521, 255.7379, 255.0225, 253.4652, 252.3368, 
    253.1728,
  275.6438, 274.6377, 272.9908, 271.403, 266.9213, 260.855, 259.6012, 
    259.7151, 258.7914, 257.7456, 256.9133, 255.2727, 253.0551, 251.4269, 
    251.4857,
  275.6646, 274.6519, 273.3444, 266.9493, 261.9846, 259.3488, 259.1582, 
    260.1435, 259.5427, 258.3826, 257.1898, 255.8298, 253.0983, 251.403, 
    251.5346,
  273.7804, 271.249, 266.9095, 261.6762, 259.0417, 257.5297, 258.3316, 
    260.545, 260.6545, 258.5092, 257.6422, 255.6738, 252.5806, 251.4009, 
    251.3493,
  267.9629, 266.7784, 264.3719, 262.9966, 262.0818, 261.0293, 260.9873, 
    259.9811, 259.2471, 257.4353, 258.1735, 257.4659, 256.0557, 256.5949, 
    256.5068,
  268.0361, 266.8944, 264.1995, 262.3293, 261.3262, 259.0677, 259.5964, 
    259.0942, 257.8063, 257.9761, 255.2951, 256.5823, 257.6806, 255.394, 
    255.1049,
  271.9591, 269.9478, 266.6343, 262.2608, 259.4817, 257.3662, 258.901, 
    258.9432, 257.4883, 255.836, 255.8942, 256.818, 257.6245, 258.9578, 
    258.0712,
  273.1695, 272.856, 272.2545, 264.0477, 259.5402, 258.2601, 255.6287, 
    258.2789, 258.3665, 256.8822, 255.8669, 258.1512, 257.7426, 259.5071, 
    259.8441,
  274.1543, 272.7725, 271.9755, 262.4258, 260.2187, 259.2371, 258.493, 
    254.5225, 255.8629, 258.4485, 256.4085, 257.5789, 259.6024, 259.2866, 
    259.9688,
  274.8459, 273.2219, 270.6342, 262.4244, 261.7557, 260.6333, 259.5399, 
    259.7467, 259.7678, 259.26, 256.4224, 257.6994, 258.6422, 258.4415, 
    258.838,
  275.3422, 274.1572, 272.4617, 267.6754, 262.1852, 258.726, 259.4122, 
    259.3132, 258.9949, 258.1938, 256.8098, 256.8762, 256.9193, 256.6671, 
    255.9908,
  275.6406, 274.6266, 272.9155, 270.3514, 263.9144, 257.4711, 257.6954, 
    258.2103, 258.285, 258.2113, 255.1082, 256.3618, 255.4036, 254.3594, 
    254.0961,
  275.6718, 274.6534, 272.8435, 263.3535, 258.7525, 256.5816, 257.0243, 
    257.4457, 257.5882, 256.8704, 255.8356, 255.0105, 253.5452, 252.0606, 
    250.598,
  273.7513, 270.5625, 264.8357, 258.9409, 257.3997, 255.9411, 255.6714, 
    258.3981, 257.6754, 254.2409, 252.9433, 252.9975, 251.5294, 251.0046, 
    250.2126,
  266.2712, 264.5087, 262.0914, 260.7996, 261.0186, 258.2716, 257.2083, 
    256.969, 256.4764, 255.2878, 257.9663, 257.2467, 252.9974, 251.7706, 
    252.0722,
  267.0563, 266.4961, 264.3817, 262.6199, 262.3684, 259.2404, 259.2311, 
    258.4168, 257.8736, 257.2688, 254.677, 258.1101, 257.5477, 254.7076, 
    249.2683,
  271.9562, 270.4456, 268.5072, 265.0697, 262.3902, 258.9822, 260.8631, 
    259.9731, 259.1624, 257.391, 256.8906, 256.8954, 258.3883, 260.282, 
    254.7839,
  273.1615, 272.8456, 272.3747, 267.7554, 264.6897, 261.7737, 258.3517, 
    260.1555, 260.1322, 258.0615, 256.8111, 258.0725, 258.6368, 257.7196, 
    257.4978,
  274.161, 272.7655, 272.5156, 268.1001, 266.5025, 264.369, 261.3547, 
    255.7824, 256.3053, 259.0883, 256.8965, 255.9015, 256.803, 257.6907, 
    258.4803,
  274.8779, 273.3115, 271.7025, 269.4092, 268.885, 266.8217, 263.7952, 
    261.5648, 259.8686, 258.3352, 255.7048, 254.9542, 254.5043, 255.0961, 
    256.493,
  275.4174, 274.2625, 272.6596, 271.0648, 269.5866, 267.2784, 265.2447, 
    263.1816, 260.8658, 258.8808, 256.7211, 255.4382, 253.9815, 253.2546, 
    253.6265,
  275.7305, 274.7298, 273.0547, 271.6508, 270.7144, 268.4345, 266.1554, 
    264.5533, 262.3191, 260, 257.0186, 254.8783, 253.4573, 252.0645, 251.3608,
  275.7221, 274.7558, 273.4745, 271.9347, 270.9664, 269.3673, 267.4919, 
    265.9638, 264.044, 261.1582, 257.6751, 254.9928, 252.8305, 251.5773, 
    250.3658,
  274.2288, 273.1234, 272.3574, 271.9905, 271.1446, 269.8258, 268.1918, 
    267.1057, 265.4977, 261.1622, 257.4845, 254.8365, 251.8508, 250.0934, 
    251.0638,
  271.6324, 271.3039, 271.283, 271.4643, 271.2443, 270.4384, 269.6855, 
    267.9865, 265.4085, 261.6975, 261.7135, 261.02, 258.3385, 256.9769, 
    254.787,
  271.4671, 271.773, 271.8091, 272.0527, 272.0757, 271.2844, 270.5646, 
    269.6203, 267.9942, 264.9157, 262.7686, 262.1148, 261.2005, 258.4181, 
    255.39,
  272.2341, 271.8208, 271.7916, 272.1471, 272.3684, 271.0335, 270.909, 
    270.7761, 269.3991, 267.7673, 265.4146, 263.5037, 262.1815, 261.678, 
    260.1594,
  273.2578, 272.9193, 272.6422, 271.6818, 272.0329, 272.0127, 270.5396, 
    270.0525, 269.3518, 268.2069, 266.1874, 264.5212, 262.9262, 261.7917, 
    260.9164,
  274.1844, 272.8031, 272.8385, 271.0718, 271.3206, 271.4247, 271.302, 
    268.5738, 268.052, 269.701, 268.8488, 266.4608, 264.0062, 262.2094, 
    261.4095,
  274.8939, 273.3645, 271.9652, 270.4288, 270.712, 270.143, 270.1467, 
    270.1898, 270.049, 269.8733, 268.9166, 267.3048, 264.6393, 262.4395, 
    260.9646,
  275.393, 274.2977, 272.7029, 271.0853, 270.0209, 268.6955, 268.3815, 
    269.0722, 269.1212, 269.2562, 268.5125, 266.7482, 263.8146, 261.4726, 
    259.9552,
  275.7032, 274.7193, 273.0913, 271.127, 269.1124, 267.6096, 267.0103, 
    267.5292, 267.0915, 267.8106, 267.6212, 265.4853, 262.2576, 259.6841, 
    258.1754,
  275.6298, 274.7214, 273.2202, 268.1247, 265.7203, 265.6557, 265.1318, 
    265.2751, 265.5482, 265.6293, 264.6335, 262.1096, 259.0554, 257.3088, 
    255.5467,
  273.787, 271.9317, 269.1145, 266.3591, 263.8807, 263.2921, 262.4915, 
    263.4159, 263.1162, 261.0164, 259.9555, 257.1571, 255.3248, 253.6367, 
    251.6045,
  272.4596, 271.5997, 270.9995, 269.776, 267.6528, 266.0602, 265.7303, 
    265.1786, 268.8505, 268.7142, 268.9482, 268.1056, 264.3124, 261.489, 
    258.7935,
  272.2067, 271.8253, 271.1846, 269.6165, 266.5595, 264.0741, 264.0075, 
    262.7773, 263.5245, 266.0105, 267.0964, 268.2112, 266.6131, 262.1943, 
    259.7005,
  272.2659, 271.7318, 271.3937, 269.8713, 267.1731, 261.9691, 263.643, 
    261.8192, 262.6575, 265.6709, 266.9338, 267.9755, 267.8977, 266.0953, 
    262.4933,
  273.3202, 272.9538, 272.6368, 270.2154, 267.5792, 264.3812, 258.6301, 
    260.8528, 260.5041, 262.6954, 265.3351, 267.1226, 268.0351, 267.5221, 
    264.4298,
  274.1886, 272.8131, 272.8404, 269.968, 267.9786, 264.8994, 261.9405, 
    254.677, 257.067, 261.2842, 263.9611, 266.1966, 267.7681, 268.4279, 
    267.1399,
  274.9258, 273.354, 272.0211, 270.5083, 269.8557, 266.1922, 262.7203, 
    260.9218, 257.5494, 258.5655, 260.7787, 265.07, 266.8274, 267.8171, 
    265.782,
  275.4129, 274.338, 272.7156, 271.3125, 270.1924, 267.181, 263.8548, 
    261.2921, 258.5669, 256.954, 258.7262, 262.0004, 265.2544, 264.6584, 
    262.6757,
  275.7471, 274.7563, 273.1063, 271.623, 270.6003, 267.8008, 264.9394, 
    262.1764, 258.4287, 256.01, 257.9823, 257.2654, 258.8003, 259.2201, 
    258.6352,
  275.657, 274.7653, 273.4201, 271.7288, 270.0248, 267.9163, 265.176, 
    262.7052, 259.8239, 256.764, 255.5548, 256.9433, 255.102, 254.6893, 
    254.6283,
  274.1996, 273.3162, 272.48, 271.6348, 270.1624, 268.329, 265.9933, 
    264.0922, 261.7431, 257.3102, 254.461, 253.676, 252.7961, 252.2189, 
    252.1092,
  273.0796, 272.4509, 272.3637, 272.6858, 272.3289, 269.3365, 267.5626, 
    264.7215, 263.2098, 263.5432, 259.2875, 264.0744, 265.5887, 265.2071, 
    263.8026,
  272.6207, 272.2422, 272.0025, 272.2403, 272.3311, 270.3112, 268.0573, 
    264.6255, 261.4969, 260.8024, 261.6063, 264.4177, 265.6373, 264.1667, 
    262.3287,
  272.3326, 271.8331, 271.7316, 271.7566, 272.2755, 269.9303, 268.1984, 
    265.6429, 262.5739, 261.6035, 261.9782, 264.0118, 264.3506, 265.9223, 
    265.127,
  273.396, 273.011, 272.702, 271.4425, 271.7963, 271.8256, 268.1864, 
    265.8034, 263.8527, 262.7866, 262.6552, 261.3846, 262.4756, 264.565, 
    266.232,
  274.2325, 272.8451, 272.8869, 271.1067, 271.0972, 271.5826, 270.6469, 
    264.5916, 262.0725, 265.0544, 263.495, 262.0026, 262.9316, 264.6392, 
    266.1054,
  274.985, 273.3604, 272.0753, 270.8485, 270.8016, 270.7479, 270.7433, 
    269.5173, 267.0618, 264.2132, 262.5278, 262.2552, 261.844, 263.0703, 
    265.5786,
  275.4245, 274.3872, 272.7511, 271.2065, 270.4366, 269.6999, 269.9692, 
    269.6717, 268.2071, 265.648, 263.0215, 261.7811, 261.4033, 262.0831, 
    263.2088,
  275.7647, 274.7894, 273.1557, 271.0914, 269.3202, 268.0394, 268.4532, 
    268.969, 268.1479, 265.8555, 263.546, 261.9513, 260.7975, 259.9633, 
    261.4048,
  275.6445, 274.7802, 273.1397, 268.8, 266.2719, 266.2634, 266.7113, 
    267.0662, 266.5314, 265.0356, 263.0746, 261.7151, 260.8687, 259.4434, 
    258.4847,
  274.099, 272.6836, 270.9059, 267.8355, 264.8507, 264.4795, 264.5747, 
    264.7752, 264.782, 262.9632, 261.9831, 261.4899, 260.2283, 259.4645, 
    257.8573,
  273.004, 272.0264, 271.4937, 269.9207, 268.2594, 268.5684, 268.5517, 
    270.6173, 269.5021, 267.0661, 263.0072, 263.2569, 260.485, 264.2976, 
    265.6456,
  272.3794, 271.941, 270.9648, 269.2264, 265.8105, 264.9597, 266.7562, 
    268.7094, 269.4276, 267.7461, 265.8391, 264.8265, 262.6133, 260.46, 
    264.3622,
  272.4045, 271.8245, 271.3887, 268.797, 266.1307, 264.4929, 265.7836, 
    267.2866, 268.2964, 267.5254, 266.5516, 266.0961, 264.5383, 261.8435, 
    262.2845,
  273.4717, 273.0598, 272.6906, 268.5329, 265.3898, 264.968, 263.7174, 
    264.0534, 265.5497, 266.1781, 265.7224, 266.1321, 265.6078, 264.1588, 
    263.868,
  274.2237, 272.8575, 272.778, 267.7458, 264.7918, 263.4092, 263.9094, 
    261.0913, 261.3076, 264.644, 265.4136, 265.5833, 266.1309, 265.3413, 
    264.0559,
  274.9709, 273.3263, 271.9881, 268.3059, 266.6886, 261.2718, 261.7898, 
    262.03, 261.7839, 262.0044, 261.4289, 262.6393, 264.1204, 265.3431, 
    264.5633,
  275.3778, 274.369, 272.7284, 270.7158, 266.4495, 260.5146, 259.2389, 
    258.7979, 258.1723, 258.0004, 257.8876, 259.5547, 261.0368, 262.7711, 
    264.1546,
  275.7262, 274.7593, 273.1377, 269.5965, 264.082, 258.7634, 257.5067, 
    256.725, 256.0228, 255.2883, 255.1617, 256.3995, 258.4186, 260.4736, 
    262.8987,
  275.5856, 274.7518, 272.457, 263.994, 258.3517, 258.0456, 256.7824, 
    255.8443, 254.2678, 254.4369, 253.3744, 253.4497, 255.0105, 258.099, 
    260.7413,
  273.5169, 270.9178, 266.8714, 261.3337, 258.0386, 256.2104, 254.8168, 
    255.9016, 254.9674, 252.026, 250.8954, 251.6782, 252.3655, 255.1006, 
    258.3778,
  265.5678, 261.2939, 259.0284, 258.8555, 258.0294, 257.3604, 256.2166, 
    256.9847, 258.1767, 258.3463, 260.1208, 263.4817, 263.9135, 263.4058, 
    261.8929,
  269.1344, 264.3975, 259.8787, 258.3176, 257.5347, 254.3686, 254.5078, 
    255.2615, 255.8919, 256.2273, 256.8349, 261.2032, 262.8769, 261.4939, 
    260.8553,
  272.4056, 271.7608, 268.8876, 259.6206, 257.0319, 252.65, 254.8095, 
    253.3602, 253.1218, 253.5682, 254.4135, 257.3488, 260.5376, 262.9039, 
    263.3429,
  273.4739, 273.0233, 272.3392, 260.632, 257.5777, 255.3913, 250.6642, 
    253.1943, 253.4314, 252.9157, 252.6831, 254.4972, 257.6464, 260.8633, 
    263.1727,
  274.1773, 272.8236, 272.1996, 261.7539, 259.7793, 255.826, 254.1027, 
    247.5111, 249.5138, 254.4805, 253.283, 252.417, 254.0196, 257.6427, 
    262.4366,
  274.9459, 273.249, 271.6603, 265.4315, 264.3839, 256.2694, 254.138, 
    252.9567, 251.0756, 249.0057, 248.4575, 250.2777, 251.7903, 254.2785, 
    259.2756,
  275.338, 274.3228, 272.668, 269.5275, 264.2435, 256.6111, 254.4645, 
    253.3644, 252.4006, 250.3571, 249.0071, 249.1053, 250.7305, 251.8982, 
    256.057,
  275.6901, 274.7267, 273.105, 268.2637, 262.9548, 257.1605, 255.2429, 
    253.9747, 252.7978, 251.1538, 249.4908, 248.5315, 248.9864, 250.3547, 
    254.6932,
  275.5666, 274.7173, 271.7454, 262.2274, 258.405, 257.6218, 255.2342, 
    254.3321, 253.3785, 252.6337, 249.5316, 247.8519, 247.4977, 249.342, 
    253.6859,
  272.9431, 269.3895, 265.9796, 260.463, 258.0209, 257.1842, 254.9016, 
    255.5695, 255.3539, 250.9301, 248.4639, 247.0012, 246.2669, 248.0546, 
    251.9288,
  266.5688, 264.3759, 262.9661, 262.4084, 262.3802, 260.717, 257.763, 
    253.2284, 251.8416, 249.4835, 248.675, 251.1443, 255.7877, 260.1599, 
    263.098,
  269.8012, 267.2689, 264.6406, 263.2304, 262.6072, 260.2711, 256.7721, 
    253.4718, 252.4776, 251.7141, 248.7118, 250.6686, 253.1672, 254.3337, 
    258.8436,
  272.4227, 271.8224, 270.1371, 264.3048, 263.6396, 258.7159, 258.2115, 
    255.2329, 254.3358, 252.0855, 251.5608, 251.115, 252.4333, 255.3546, 
    258.371,
  273.5376, 273.0475, 272.445, 264.6822, 263.4133, 260.7733, 256.8062, 
    257.1905, 256.0132, 254.8274, 253.3506, 251.4114, 251.5405, 253.0319, 
    256.8259,
  274.1474, 272.8101, 272.3431, 263.5808, 263.2704, 262.51, 258.9848, 
    253.9577, 252.1067, 255.7744, 255.118, 251.841, 250.461, 251.4373, 
    254.4015,
  274.8999, 273.2306, 271.7749, 266.5141, 265.5345, 261.0495, 259.7552, 
    257.3482, 254.306, 251.4759, 251.4423, 251.5459, 249.832, 250.2114, 
    252.8791,
  275.2861, 274.2714, 272.6561, 269.2343, 264.7709, 258.4262, 258.0215, 
    256.5746, 255.2008, 252.4767, 252.5463, 251.7982, 250.4508, 249.2041, 
    251.5761,
  275.6322, 274.6635, 272.9759, 266.9547, 261.9042, 256.995, 255.8746, 
    255.7481, 254.5948, 253.241, 251.6864, 251.5872, 250.2834, 248.6053, 
    251.4656,
  275.4982, 274.4951, 269.9597, 260.5195, 257.5942, 255.7898, 255.4685, 
    255.7378, 254.6769, 252.7353, 250.8628, 250.8603, 249.19, 248.5074, 
    250.9494,
  271.8731, 266.8202, 263.2427, 258.5284, 256.5452, 255.6449, 254.8209, 
    256.4328, 255.4832, 252.1666, 250.186, 250.2325, 248.034, 247.4687, 249.57,
  265.4331, 262.2225, 260.3449, 259.5638, 259.9959, 262.0825, 263.1051, 
    261.2889, 258.8951, 256.7518, 254.8659, 251.6491, 252.6794, 257.5345, 
    261.9726,
  269.2459, 265.9123, 261.96, 259.7552, 261.0584, 262.9616, 261.8701, 
    259.2767, 257.7762, 256.0988, 252.763, 251.6375, 254.3012, 257.0725, 
    260.9395,
  272.4391, 271.8495, 269.9358, 261.2413, 262.1333, 259.6032, 260.5458, 
    257.8774, 255.8885, 253.9258, 252.7342, 251.9541, 255.0867, 259.2569, 
    262.304,
  273.561, 273.0447, 272.3597, 261.894, 261.3588, 260.7733, 255.6193, 
    256.1195, 254.6065, 253.5188, 252.4182, 251.945, 255.7908, 258.97, 
    261.6917,
  274.04, 272.7445, 272.024, 259.9817, 260.4264, 260.3793, 259.1977, 
    252.1492, 249.112, 253.1942, 253.0557, 252.1623, 254.8533, 257.9612, 
    260.5667,
  274.7899, 273.1429, 271.6326, 264.264, 262.6223, 258.1986, 259.5781, 
    258.7417, 254.7974, 252.9281, 251.0202, 252.3539, 253.6606, 257.0692, 
    259.6796,
  275.1676, 274.1366, 272.5185, 267.1819, 262.7788, 257.8483, 259.2163, 
    257.8886, 255.6894, 253.7244, 253.731, 253.291, 254.1976, 257.1319, 
    260.0213,
  275.5217, 274.507, 272.2615, 265.5664, 261.6176, 258.9225, 258.0486, 
    256.3205, 254.0208, 253.9545, 253.2143, 253.5253, 254.7215, 256.8365, 
    259.9364,
  275.4052, 274.057, 267.4467, 259.9704, 259.0703, 257.8808, 257.229, 
    254.8125, 252.9152, 252.3891, 251.9412, 252.6357, 253.7778, 256.4659, 
    258.9464,
  270.7278, 265.0205, 261.0887, 258.1487, 256.9404, 256.5794, 255.1591, 
    255.5409, 253.0135, 250.8527, 250.8045, 251.7281, 252.5118, 255.6784, 
    259.4039,
  262.9224, 259.2565, 257.5345, 256.2971, 257.3144, 257.0507, 256.0577, 
    254.9044, 258.5677, 262.8305, 263.6501, 262.225, 259.9098, 258.6584, 
    255.4809,
  268.8197, 264.9309, 259.774, 256.9202, 258.1595, 257.9413, 258.8973, 
    257.1017, 259.9859, 263.1914, 262.7778, 261.2563, 260.1078, 255.8154, 
    254.6879,
  272.4308, 271.7027, 268.7384, 258.4503, 258.3854, 256.1313, 258.8834, 
    258.569, 260.3019, 262.1667, 261.3251, 260.3324, 259.2499, 257.546, 
    256.4169,
  273.5548, 273.0569, 272.0215, 260.1152, 258.7231, 259.0836, 255.3081, 
    257.9124, 259.3454, 260.264, 258.5654, 258.2762, 259.1197, 257.7669, 
    257.819,
  273.983, 272.7293, 271.5421, 259.5219, 258.7583, 258.8642, 260.0253, 
    251.9449, 251.1087, 257.928, 257.6068, 254.3563, 256.7789, 258.9779, 
    258.8822,
  274.7801, 273.1134, 271.3786, 263.9816, 260.8477, 256.9506, 256.8019, 
    257.5837, 253.2749, 252.6988, 251.5481, 253.5641, 259.2676, 260.3279, 
    259.9906,
  275.1242, 274.08, 272.2512, 266.3872, 261.0217, 255.6577, 254.4093, 
    253.9016, 253.0359, 251.0117, 251.8646, 256.6381, 261.9817, 263.1532, 
    262.6781,
  275.5082, 274.4698, 271.3953, 265.2824, 260.1777, 256.0002, 253.8365, 
    252.6324, 251.338, 252.3239, 255.6312, 260.7573, 262.9539, 263.4315, 
    264.1967,
  275.4556, 274.1914, 266.7271, 260.7746, 257.6503, 256.1703, 254.9207, 
    254.059, 253.645, 255.0576, 258.7574, 262.4013, 262.8734, 262.5997, 
    263.3366,
  271.1384, 265.5701, 261.3153, 258.764, 256.5055, 255.8689, 255.4621, 
    257.0471, 257.2872, 257.2576, 258.8794, 261.2069, 261.496, 262.8839, 
    264.1061,
  264.8289, 258.7737, 256.663, 256.4896, 258.6392, 259.7493, 261.3888, 
    261.796, 262.3678, 261.7625, 261.8768, 262.93, 263.2613, 263.4202, 
    262.5866,
  269.2398, 263.1942, 259.3157, 257.7899, 258.9247, 259.3901, 261.9821, 
    262.1827, 263.1653, 264.191, 264.6466, 265.6638, 265.7126, 263.0924, 
    262.8982,
  272.5125, 271.553, 267.7844, 258.9467, 258.4926, 257.4811, 261.0891, 
    261.5987, 261.773, 262.217, 262.5659, 263.3565, 263.9716, 264.6484, 
    263.773,
  273.5276, 273.0583, 271.5497, 259.9957, 259.1816, 260.1873, 259.254, 
    260.9856, 260.3329, 260.3678, 260.2019, 260.6254, 261.6362, 262.3808, 
    262.6377,
  274.0425, 272.7548, 271.0006, 259.771, 259.5549, 259.8556, 261.6273, 
    256.5574, 255.9823, 259.9211, 259.3234, 258.0045, 258.6094, 259.8763, 
    261.0697,
  274.8515, 273.0818, 271.0179, 263.7743, 261.7552, 258.8523, 259.2209, 
    259.717, 256.3279, 257.2573, 256.9336, 257.7666, 257.8685, 257.6317, 
    258.702,
  275.1523, 274.0702, 271.9162, 266.1227, 261.6807, 259.2796, 258.1819, 
    258.0301, 257.2612, 255.4872, 256.2351, 257.617, 258.4142, 256.8228, 
    259.0505,
  275.5241, 274.5176, 270.9398, 264.5112, 260.7328, 259.2429, 258.062, 
    259.88, 259.3404, 257.8473, 258.0567, 256.772, 256.4615, 259.9711, 
    261.5803,
  275.5351, 274.3012, 265.7678, 260.3455, 258.4181, 257.7898, 259.1076, 
    258.8696, 261.0014, 260.3498, 260.6391, 260.5095, 260.7881, 259.6796, 
    263.0858,
  271.3733, 265.7154, 260.5654, 258.2099, 258.1538, 258.4989, 259.959, 
    263.3842, 262.5783, 262.9738, 263.718, 264.0334, 263.4646, 263.1224, 
    263.3861,
  263.1146, 260.264, 259.1088, 259.3197, 260.9997, 258.463, 257.3599, 
    257.3499, 259.2878, 261.4538, 262.6483, 260.2083, 254.2193, 256.3394, 
    255.2554,
  268.3987, 263.8734, 261.3997, 260.3949, 261.0691, 258.036, 257.6557, 
    257.2346, 258.1402, 261.1021, 261.6917, 263.6595, 260.9525, 253.9549, 
    254.3364,
  272.4818, 271.5287, 268.5902, 261.3509, 258.9988, 256.499, 258.0798, 
    257.6437, 258.0279, 258.7343, 260.1754, 263.3601, 262.302, 259.3235, 
    256.9428,
  273.4603, 273.0267, 271.6052, 262.3531, 260.0797, 259.1687, 256.3397, 
    257.0371, 258.1252, 258.2524, 258.58, 261.5667, 264.6292, 262.7887, 
    258.6578,
  274.0781, 272.7362, 271.2475, 262.2071, 261.6562, 260.8194, 260.4108, 
    256.3673, 256.6302, 259.6693, 259.0844, 259.6458, 262.8114, 263.9437, 
    261.7684,
  274.8983, 273.0894, 271.1735, 266.2833, 263.5358, 260.8676, 260.4786, 
    261.793, 261.3839, 260.4308, 258.7155, 258.9676, 260.9755, 263.0161, 
    263.808,
  275.2755, 274.1144, 272.0805, 267.5629, 262.8002, 260.7024, 260.1451, 
    261.7377, 262.7223, 261.6907, 259.5614, 259.2019, 260.6072, 263.1434, 
    264.4569,
  275.6122, 274.629, 271.5901, 266.0526, 262.408, 259.6975, 259.4246, 
    262.0988, 263.8627, 263.6167, 261.1852, 260.1938, 260.6135, 262.6165, 
    264.0642,
  275.6644, 274.4819, 269.3436, 264.3114, 261.0353, 258.5242, 258.8655, 
    261.617, 264.0198, 264.4742, 263.1576, 262.0676, 261.8641, 262.5905, 
    262.0606,
  273.0327, 269.8184, 266.2553, 263.1768, 260.8419, 257.6458, 258.1565, 
    262.2934, 264.163, 264.4337, 264.2425, 263.4423, 263.4478, 263.7328, 
    263.4362,
  266.2335, 265.3088, 265.3501, 264.1474, 263.0832, 263.0704, 262.2311, 
    260.1571, 258.354, 259.5608, 260.2862, 258.4133, 257.9007, 258.2858, 
    258.7175,
  269.8418, 268.3527, 266.4094, 265.5476, 265.528, 264.3502, 263.5409, 
    260.5603, 257.338, 260.6025, 260.9934, 259.6624, 259.9886, 256.428, 
    257.218,
  272.5475, 271.7992, 270.4461, 266.9377, 265.3478, 264.4486, 264.7978, 
    261.8543, 257.7495, 261.8857, 261.5217, 261.653, 258.9273, 259.5449, 
    258.0392,
  273.5401, 273.0859, 272.3465, 268.7768, 267.8928, 267.1648, 263.6712, 
    259.1834, 256.8013, 260.9504, 262.3183, 262.5904, 261.6672, 259.7401, 
    257.1674,
  274.1934, 272.832, 272.3981, 269.6283, 268.85, 266.3746, 264.5766, 253.167, 
    253.9677, 260.4031, 262.7324, 263.0007, 264.3415, 260.8756, 259.7398,
  275.0196, 273.2922, 271.8673, 270.3536, 268.7023, 264.881, 259.7509, 
    257.7041, 256.2721, 260.8896, 262.0851, 262.6838, 264.4594, 262.9882, 
    262.5041,
  275.4374, 274.2528, 272.5655, 269.9424, 266.7156, 261.9562, 258.7858, 
    259.6694, 260.5366, 263.2982, 262.8729, 262.7226, 263.8015, 265.321, 
    264.6647,
  275.7069, 274.7485, 272.5807, 268.1159, 264.2169, 259.0583, 259.1005, 
    260.5234, 261.9431, 263.8412, 263.1612, 262.3615, 263.244, 264.4362, 
    265.2776,
  275.741, 274.5941, 270.9568, 265.1685, 261.201, 257.5909, 259.0809, 
    260.4842, 263.6831, 264.9462, 263.7114, 262.5851, 262.6853, 263.3829, 
    263.8184,
  273.5663, 271.5825, 269.5353, 264.439, 262.3588, 256.4705, 258.7192, 
    262.7761, 264.5321, 264.1199, 263.4034, 262.9695, 263.7485, 263.8239, 
    264.114,
  268.8901, 268.4638, 269.2775, 268.1565, 267.933, 268.5788, 268.7025, 
    268.937, 267.0258, 261.5115, 257.4364, 261.0507, 260.4634, 259.5105, 
    259.1546,
  270.96, 270.4647, 268.8625, 267.3304, 265.8146, 266.4774, 268.0849, 
    267.4554, 264.7491, 258.9729, 257.3407, 262.418, 261.2827, 258.9667, 
    258.7477,
  272.6295, 271.9315, 270.4437, 265.3108, 264.0425, 262.2029, 264.232, 
    263.6559, 258.7183, 257.341, 260.6284, 262.3046, 262.2148, 262.7856, 
    261.6454,
  273.6205, 273.1252, 272.3066, 264.4813, 262.6042, 261.9077, 258.6115, 
    259.5579, 256.6727, 257.9183, 258.9472, 262.2851, 263.0403, 263.2287, 
    261.6672,
  274.3681, 272.9029, 272.241, 263.7742, 262.5876, 259.8319, 260.2379, 
    254.1767, 252.4258, 258.5881, 262.5816, 262.5267, 263.3041, 262.7521, 
    263.7011,
  275.2757, 273.4576, 271.7143, 266.4415, 264.3562, 260.433, 259.8563, 
    260.2646, 259.4381, 258.9598, 262.4027, 261.0113, 263.0511, 263.1483, 
    263.0412,
  275.6413, 274.4007, 272.5144, 268.2284, 264.8783, 260.554, 259.6168, 
    260.9137, 261.7873, 262.9791, 263.2071, 261.7805, 263.9822, 263.4146, 
    262.4637,
  275.89, 274.8363, 272.5361, 268.4245, 265.6317, 260.1191, 259.4145, 
    261.4793, 263.3357, 264.0297, 264.0866, 262.8179, 264.4952, 263.6563, 
    262.8438,
  275.9028, 274.642, 271.3777, 268.4379, 266.3928, 261.5309, 259.271, 
    261.9998, 263.668, 265.0199, 264.5289, 263.9141, 265.0889, 265.1643, 
    265.1969,
  273.8026, 271.9905, 270.1974, 269.3488, 266.8406, 260.7952, 258.889, 
    264.0885, 265.0849, 264.559, 265.0276, 265.5339, 265.8744, 265.5094, 
    263.1521,
  268.0151, 263.5781, 263.569, 262.0294, 260.3197, 260.8073, 258.8292, 
    261.6501, 262.1783, 262.2623, 261.9235, 263.1261, 262.4112, 261.5862, 
    260.7566,
  270.8189, 267.2523, 266.0076, 264.2726, 262.6527, 260.2202, 259.0439, 
    257.0197, 259.5187, 261.325, 261.5841, 262.7516, 261.9612, 259.2154, 
    259.5318,
  272.7271, 271.9615, 270.6349, 266.249, 264.5664, 261.0312, 258.6096, 
    258.8748, 260.6553, 260.3941, 261.1312, 263.3781, 263.0649, 262.7276, 
    261.9609,
  273.6041, 273.1164, 272.4977, 267.8557, 267.787, 265.3095, 259.1901, 
    257.1638, 260.7358, 262.2207, 263.0271, 263.9658, 264.0046, 264.5041, 
    264.2512,
  274.5017, 272.9302, 272.635, 269.0119, 268.9951, 266.7992, 261.428, 
    257.4167, 259.2246, 264.0095, 264.5773, 263.9256, 264.1704, 264.1535, 
    264.5631,
  275.4318, 273.5728, 271.9635, 270.7944, 269.0336, 266.0402, 262.4764, 
    262.8418, 263.0513, 263.9798, 263.7081, 262.9694, 264.097, 263.592, 
    263.8536,
  275.8579, 274.5467, 272.6559, 270.9945, 267.3816, 263.7236, 261.4832, 
    263.1921, 264.3811, 264.0122, 263.364, 263.1368, 263.8627, 263.9275, 
    264.3161,
  276.1682, 274.9383, 272.5764, 270.1592, 265.2383, 262.4072, 261.6497, 
    264.2484, 263.8245, 263.6548, 262.8225, 263.6528, 264.1755, 264.837, 
    264.7079,
  276.1449, 274.7163, 270.5421, 268.2893, 262.3456, 260.0002, 261.901, 
    264.7497, 264.177, 263.0822, 262.8664, 263.4496, 263.7949, 264.9561, 
    265.7466,
  273.9952, 271.7804, 268.3294, 266.9213, 260.0687, 260.1709, 262.1488, 
    266.2551, 264.9153, 262.4313, 261.955, 262.4365, 263.252, 263.8178, 
    265.1867,
  268.8049, 269.2992, 270.374, 268.1164, 264.8791, 264.3607, 260.6353, 
    261.0582, 261.9038, 262.6039, 261.9936, 262.2327, 262.7127, 260.7356, 
    259.1028,
  270.752, 271.3704, 270.3431, 266.8257, 265.1938, 261.4177, 261.522, 
    258.997, 259.1765, 259.7603, 261.535, 262.8053, 263.2652, 262.0092, 
    260.7644,
  273.0499, 272.1148, 271.119, 267.2068, 263.9258, 262.2752, 260.2226, 
    260.8321, 260.3318, 261.9243, 262.153, 262.8177, 262.8541, 261.9548, 
    261.2101,
  273.7527, 273.2203, 272.5393, 268.0625, 263.5852, 261.7308, 257.4505, 
    260.4218, 261.6065, 262.0932, 262.0652, 262.4898, 262.5879, 262.4839, 
    262.8531,
  274.6702, 273.0783, 272.5764, 267.2412, 263.0924, 261.6039, 261.2313, 
    256.3255, 258.2193, 262.6198, 262.8761, 262.0706, 262.7409, 263.0235, 
    262.511,
  275.5861, 273.7318, 271.8719, 268.6719, 265.5439, 261.0524, 260.256, 
    260.3522, 258.363, 259.4599, 260.913, 262.7525, 263.8529, 263.517, 
    263.7181,
  276.0208, 274.7154, 272.647, 268.8574, 264.7274, 261.5854, 260.1239, 
    259.8841, 259.3007, 259.8466, 260.541, 262.399, 263.7126, 264.4538, 
    264.2459,
  276.336, 275.0804, 271.8783, 267.771, 263.5989, 263.6424, 259.9038, 
    259.3161, 259.8558, 260.2026, 260.5179, 262.1296, 263.3557, 264.8025, 
    264.7692,
  276.2958, 274.7961, 268.6644, 263.7905, 264.1859, 261.843, 259.4965, 
    260.1853, 260.7975, 261.3574, 260.6244, 261.1093, 262.7014, 264.2739, 
    266.1928,
  274.2028, 271.8036, 268.1715, 264.7654, 263.8296, 263.9572, 259.9808, 
    263.6527, 262.8519, 259.7837, 258.7492, 260.4033, 262.0036, 263.7052, 
    266.084,
  266.4561, 263.6903, 263.5316, 259.1304, 256.8217, 256.1964, 255.6992, 
    256.5832, 257.1176, 258.2731, 258.3896, 257.4938, 261.1264, 261.6558, 
    260.4976,
  269.8577, 266.5051, 264.8519, 260.5692, 258.7721, 256.8833, 256.5014, 
    257.4395, 258.1725, 258.0072, 256.8766, 258.3768, 259.3255, 259.9591, 
    258.6166,
  273.0758, 272.1792, 270.2165, 262.9545, 259.9817, 257.1015, 258.326, 
    258.1076, 258.2448, 259.0738, 258.4446, 258.7269, 261.1876, 261.5503, 
    261.1173,
  273.7996, 273.2103, 272.548, 267.6256, 262.8508, 260.7581, 257.8915, 
    259.22, 259.6093, 259.8973, 259.587, 259.7084, 261.2458, 261.7147, 
    260.6337,
  274.847, 273.1186, 272.7277, 269.1567, 265.3321, 263.032, 262.6948, 
    257.2541, 256.9512, 261.9893, 261.5236, 260.5399, 261.039, 260.5942, 
    261.1083,
  275.6441, 273.8902, 272.0184, 270.1394, 268.4817, 265.5133, 263.4565, 
    261.7495, 260.5858, 260.5135, 260.6574, 260.7994, 261.6146, 260.2866, 
    261.212,
  276.0604, 274.8609, 272.828, 270.3348, 268.5364, 266.4335, 264.3955, 
    263.4956, 262.7094, 261.9785, 261.8114, 261.1382, 260.5323, 260.9964, 
    262.234,
  276.4178, 275.2261, 272.8334, 270.637, 269.1281, 267.8113, 266.6405, 
    265.2837, 264.4927, 263.9774, 263.0631, 261.0887, 260.0408, 261.775, 
    263.2029,
  276.3911, 274.9021, 271.9648, 270.3473, 269.2841, 268.691, 267.6947, 
    266.8912, 266.1795, 265.4388, 263.798, 261.5365, 260.8476, 261.1989, 
    264.4763,
  274.4162, 272.4772, 272.1696, 271.7711, 270.4003, 269.868, 268.7457, 
    268.9641, 268.173, 265.9432, 262.7835, 260.7303, 259.0099, 260.7282, 
    263.3207,
  269.8727, 268.5649, 267.9281, 266.5438, 265.9112, 263.684, 261.8983, 
    260.1941, 260.9402, 260.4754, 260.8047, 258.1201, 257.7158, 257.2498, 
    254.6543,
  271.5341, 270.4908, 268.8662, 267.0675, 264.8542, 265.1109, 262.4364, 
    262.8596, 263.0436, 261.3319, 261.9402, 260.2869, 259.5766, 258.5959, 
    256.9376,
  273.0973, 272.2392, 271.1962, 267.8636, 268.0918, 265.8503, 266.7121, 
    265.8436, 265.2841, 264.7328, 264.3252, 263.1898, 262.7854, 261.9732, 
    260.7137,
  274.0305, 273.5017, 272.8547, 270.4381, 270.4108, 267.718, 266.2221, 
    267.6121, 266.6548, 266.541, 265.6187, 264.518, 264.3247, 263.9092, 
    262.4887,
  275.272, 273.4773, 273.1245, 271.8449, 271.6366, 271.2803, 270.324, 
    267.0752, 266.6609, 269.0688, 269.3027, 268.5516, 267.5426, 266.2367, 
    264.6087,
  276.007, 274.3227, 272.2825, 271.7551, 272.0305, 272.2816, 272.0238, 
    271.661, 271.3405, 270.9919, 270.1831, 269.2503, 268.7173, 267.8275, 
    266.8737,
  276.1671, 275.018, 273.0276, 271.9352, 272.228, 272.4637, 272.3287, 
    271.7841, 270.5282, 269.1877, 267.9594, 267.6552, 267.9081, 267.6689, 
    267.5416,
  276.5387, 275.3982, 273.2429, 272.2297, 272.5628, 272.3734, 271.3137, 
    269.4334, 267.4341, 266.5861, 266.2515, 266.7782, 266.4589, 266.6982, 
    266.8648,
  276.5015, 275.0326, 272.257, 272.3339, 271.7246, 270.1196, 268.0467, 
    266.3218, 265.832, 266.0918, 263.9911, 264.5287, 264.8301, 265.1568, 
    266.0056,
  274.6008, 272.4524, 272.0253, 271.4086, 269.77, 266.7341, 264.2835, 
    264.8855, 265.8923, 263.5471, 262.5258, 262.7922, 263.244, 263.9996, 
    264.9387,
  270.9253, 270.5065, 271.9164, 270.9489, 270.9445, 270.7528, 270.0503, 
    267.5896, 266.4431, 265.5953, 266.3155, 266.9157, 266.0329, 266.1896, 
    264.7422,
  271.9331, 271.7192, 271.4276, 271.584, 271.895, 271.7949, 270.2732, 
    268.9719, 267.7522, 267.1535, 267.4799, 267.919, 267.8406, 265.9691, 
    264.7925,
  273.3456, 272.5092, 272.0634, 271.3611, 271.9271, 269.7272, 270.098, 
    269.068, 267.6406, 268.0923, 268.488, 269.3552, 269.6833, 269.3674, 
    267.2403,
  274.4014, 273.7803, 273.0589, 270.963, 270.5981, 269.0258, 267.3157, 
    266.2904, 266.5419, 267.5785, 267.48, 268.4877, 268.8654, 268.9314, 
    268.0008,
  275.5062, 273.6254, 273.1808, 269.738, 268.4117, 267.9043, 267.1362, 
    263.4624, 264.3498, 265.1588, 264.4232, 264.0804, 263.9866, 264.1329, 
    265.3847,
  276.13, 274.4628, 272.3086, 269.4733, 267.0543, 265.0099, 265.2602, 
    265.724, 264.9664, 261.5561, 259.5618, 258.9318, 258.7169, 258.2762, 
    260.5711,
  276.2597, 275.0915, 273.061, 269.2642, 264.6833, 262.2605, 261.1669, 
    262.1145, 261.7284, 260.8074, 259.3954, 258.0195, 259.495, 258.6454, 
    258.9049,
  276.5587, 275.423, 272.515, 266.7552, 263.1996, 260.401, 259.2958, 
    259.8438, 260.9807, 261.5216, 261.1758, 261.3332, 261.6049, 262.3866, 
    262.625,
  276.4572, 275.0598, 268.8943, 262.6138, 262.08, 259.617, 259.3647, 
    261.0354, 261.8871, 263.1044, 262.0089, 261.2786, 262.0398, 262.5584, 
    263.3888,
  274.6488, 271.3924, 265.7441, 261.7276, 259.9581, 259.1736, 259.877, 
    261.9281, 264.581, 263.0174, 262.06, 261.285, 261.347, 262.1295, 262.6349,
  269.6098, 267.2549, 265.8859, 265.0887, 264.9182, 265.0069, 262.3267, 
    261.8599, 261.8057, 262.8011, 263.3201, 263.92, 265.0497, 266.9301, 
    268.1846,
  271.03, 269.0084, 264.7434, 263.6618, 264.202, 261.428, 260.1796, 260.2935, 
    260.4298, 260.743, 262.0165, 263.2536, 264.1035, 264.7493, 266.9508,
  273.2937, 272.4319, 269.6185, 261.9285, 260.8518, 258.1308, 259.2657, 
    259.8246, 260.7263, 259.6605, 259.5195, 260.9547, 261.7948, 262.9034, 
    266.1181,
  274.2296, 273.4535, 272.441, 264.5188, 261.4399, 258.9763, 256.6291, 
    257.8973, 259.5027, 260.6846, 259.437, 259.269, 258.9733, 260.9862, 
    263.0801,
  275.3383, 273.3536, 272.8976, 266.0101, 262.5095, 261.9274, 259.5865, 
    255.2617, 258.1665, 261.2965, 260.3644, 259.1129, 258.5021, 257.923, 
    258.5507,
  275.9845, 274.2517, 272.2033, 268.0975, 264.4207, 260.3002, 261.2596, 
    261.8785, 262.0281, 259.9901, 258.5669, 258.8119, 260.0464, 257.9776, 
    257.1875,
  276.2264, 275.0598, 273.0247, 269.275, 264.2771, 259.5628, 260.2867, 
    261.6735, 261.5176, 261.2639, 260.2981, 259.6159, 261.4287, 261.0594, 
    260.0461,
  276.4981, 275.3796, 272.7624, 268.0583, 265.1882, 260.8246, 259.7333, 
    261.6094, 262.0145, 261.6018, 261.4417, 260.8649, 261.578, 263.0412, 
    263.2825,
  276.3736, 275.0536, 270.7118, 265.2556, 265.6958, 261.4448, 260.7157, 
    262.5144, 262.9457, 264.2457, 262.0702, 261.8386, 260.543, 261.3727, 
    263.111,
  274.6648, 272.2844, 269.9437, 266.8659, 266.3659, 263.3453, 260.8845, 
    263.1591, 265.3369, 263.2495, 261.6785, 261.306, 259.6376, 260.9609, 
    262.2558,
  270.1974, 267.5602, 265.9548, 264.2289, 263.745, 264.0562, 261.4032, 259.6, 
    259.1188, 259.5853, 260.499, 256.9057, 258.0073, 260.8028, 262.3888,
  271.4098, 270.1723, 268.3004, 266.4016, 265.7592, 264.2221, 262.9418, 
    261.6569, 260.4185, 259.2197, 258.3453, 255.9025, 256.3632, 260.3447, 
    259.1605,
  273.2987, 272.4475, 271.3328, 268.3561, 266.7898, 264.7089, 263.9614, 
    263.2425, 262.4029, 260.7947, 259.4619, 257.6064, 257.0912, 260.5232, 
    259.3202,
  274.2433, 273.4408, 272.7499, 270.6495, 269.2776, 266.9896, 263.4305, 
    262.8374, 262.508, 261.3975, 260.7985, 258.0229, 257.4337, 260.9445, 
    258.9424,
  275.3916, 273.3957, 273.0349, 271.5221, 270.6405, 269.4526, 267.3129, 
    261.6013, 260.1178, 262.77, 260.8045, 258.2594, 257.9397, 260.932, 
    260.7392,
  276.0151, 274.3625, 272.2856, 271.6753, 271.6738, 270.3537, 268.6582, 
    266.1435, 263.7418, 262.4059, 260.666, 257.9389, 257.8023, 258.1259, 
    262.0804,
  276.2876, 275.1555, 273.139, 271.8995, 272.0364, 270.5778, 269.1029, 
    266.7183, 263.5498, 261.2238, 260.5076, 259.2125, 257.8161, 259.3421, 
    261.4219,
  276.5567, 275.4414, 273.2881, 272.3442, 272.1614, 270.7754, 268.5409, 
    266.2709, 263.3936, 262.0982, 261.218, 259.1313, 258.3589, 260.9554, 
    261.4475,
  276.4352, 275.1185, 272.3918, 272.6656, 271.8818, 269.8889, 268.8719, 
    266.3733, 264.2707, 263.727, 259.3694, 258.2647, 257.6277, 258.9957, 
    263.0751,
  274.7655, 272.6353, 272.3732, 272.2305, 271.1396, 269.5807, 268.5169, 
    266.6411, 265.485, 261.1137, 257.6363, 257.741, 257.0908, 258.0859, 
    262.6339,
  272.1523, 271.6287, 271.4777, 270.5608, 270.1147, 269.9312, 269.7804, 
    269.999, 269.0876, 267.1027, 266.3655, 264.1939, 262.4728, 260.4831, 
    256.4771,
  272.4018, 272.0091, 271.921, 271.6706, 271.1989, 270.6863, 269.9544, 
    269.9766, 269.5648, 268.0387, 266.6731, 264.7352, 262.074, 260.3093, 
    256.8995,
  273.3425, 272.5175, 272.0703, 271.5187, 271.0445, 270.3918, 270.5931, 
    269.291, 268.2653, 266.4808, 265.3161, 264.3144, 261.6154, 261.4086, 
    260.5372,
  274.3496, 273.5178, 272.874, 271.0964, 270.4589, 270.3824, 268.0799, 
    266.8364, 266.1535, 266.2273, 265.0447, 262.7448, 260.8574, 261.0807, 
    260.8249,
  275.5326, 273.5194, 273.133, 270.4698, 269.4457, 269.0678, 267.2264, 
    263.0932, 262.9693, 265.0221, 263.0884, 261.5777, 261.0462, 260.3647, 
    261.7446,
  276.1602, 274.5607, 272.3818, 270.4669, 269.0772, 267.5316, 266.4312, 
    265.3909, 264.1025, 263.313, 261.9937, 260.7484, 260.4492, 259.9546, 
    259.3484,
  276.4449, 275.2501, 273.1839, 270.3569, 268.1302, 266.3639, 264.4115, 
    263.4532, 262.6596, 258.9906, 259.295, 260.3698, 260.2442, 260.1409, 
    259.5583,
  276.6981, 275.5049, 272.863, 268.9397, 266.5988, 265.0292, 264.3437, 
    263.2432, 261.7765, 259.6185, 258.3843, 259.0811, 260.7023, 260.7834, 
    261.3021,
  276.508, 275.1635, 270.4813, 266.744, 264.8945, 264.1686, 263.997, 
    263.5369, 262.4691, 261.3225, 258.2686, 257.8777, 257.7486, 258.7682, 
    261.6939,
  274.8829, 271.9314, 268.5009, 264.9784, 262.7971, 261.3602, 261.2598, 
    262.9247, 262.8396, 258.878, 255.5392, 256.0227, 256.1838, 257.4395, 
    260.1292,
  269.5051, 268.1059, 267.3565, 266.9397, 266.0316, 262.4323, 260.3944, 
    261.361, 262.9755, 264.4471, 265.9392, 266.8486, 267.0934, 267.0272, 
    265.1378,
  271.0931, 269.091, 266.1112, 265.8511, 264.2396, 260.3205, 259.3066, 
    259.9741, 261.0396, 263.3625, 265.22, 268.6173, 268.0582, 265.935, 
    264.3163,
  273.3271, 272.5207, 269.9554, 264.3074, 262.0367, 259.3747, 259.3127, 
    259.5242, 260.5631, 262.426, 264.6282, 267.562, 268.5357, 266.4742, 
    264.3423,
  274.331, 273.4635, 272.529, 264.8364, 261.1385, 260.1491, 256.8887, 
    258.4472, 259.3379, 260.9735, 263.0661, 265.2903, 265.826, 264.7052, 
    264.0735,
  275.5419, 273.4728, 272.9754, 265.6255, 263.0822, 262.393, 261.9702, 
    256.6145, 257.4059, 260.7223, 261.9488, 263.3376, 264.0967, 264.3766, 
    265.1255,
  276.1256, 274.506, 272.316, 268.0687, 264.0393, 262.0141, 262.0501, 
    261.7455, 259.8527, 259.4023, 260.0432, 261.6573, 262.9441, 263.1103, 
    262.6212,
  276.382, 275.1766, 273.0737, 267.7167, 262.8705, 262.1982, 261.6562, 
    261.7761, 261.5649, 258.8212, 259.3755, 260.8793, 260.8922, 261.2673, 
    261.0488,
  276.6285, 275.3931, 272.0586, 265.0505, 262.2982, 261.845, 261.5594, 
    261.4554, 261.6329, 259.2107, 258.3681, 260.1113, 261.2592, 260.9469, 
    261.9716,
  276.3788, 275.0165, 268.712, 263.6773, 262.1866, 261.4532, 261.6602, 
    262.359, 262.4405, 261.6199, 259.4873, 258.7909, 259.308, 260.2032, 
    260.4716,
  274.7679, 271.4593, 267.4296, 264.2202, 262.3181, 260.9695, 261.2511, 
    263.0027, 263.1078, 259.8488, 257.0806, 255.7541, 259.1035, 259.3323, 
    259.5542,
  268.028, 266.6659, 265.758, 264.8412, 263.8542, 259.8628, 257.9849, 
    256.1796, 256.2798, 258.8544, 260.565, 262.6745, 264.0864, 265.7603, 
    265.6105,
  270.771, 269.2477, 266.6789, 265.6491, 262.7686, 259.183, 258.5045, 
    257.408, 256.9409, 257.1967, 260.4981, 263.8016, 265.8886, 265.512, 
    264.5629,
  273.2285, 272.4962, 270.3327, 265.4567, 261.7835, 259.7703, 258.7298, 
    259.3191, 258.1253, 259.0081, 260.9038, 264.7625, 267.8219, 266.5963, 
    266.5073,
  274.2089, 273.417, 272.5163, 266.4609, 262.3689, 259.4349, 255.9573, 
    258.6032, 259.658, 260.5763, 261.1157, 264.2661, 267.4395, 267.7329, 
    267.2565,
  275.3551, 273.3427, 272.9527, 267.1544, 263.5914, 260.4765, 259.116, 
    254.9106, 256.8423, 261.0681, 260.9647, 262.7475, 265.1513, 267.1701, 
    267.3148,
  275.8906, 274.3433, 272.2598, 268.5656, 264.0144, 262.2791, 259.8135, 
    258.9074, 258.532, 259.7544, 260.0228, 261.062, 262.6543, 264.206, 265.478,
  276.1552, 275.0192, 272.9073, 267.7273, 263.9389, 262.7235, 259.9364, 
    260.034, 259.019, 258.9343, 259.8365, 260.6182, 261.588, 262.4317, 
    263.0743,
  276.4403, 275.2474, 271.7517, 266.1157, 263.8492, 262.6984, 260.9828, 
    260.8095, 260.2646, 259.83, 259.091, 259.7057, 261.3448, 262.2174, 
    263.4175,
  276.2156, 274.8855, 269.0988, 265.1841, 263.1546, 261.7012, 261.8171, 
    262.5351, 262.0041, 261.0075, 261.1092, 260.3994, 260.5001, 261.9657, 
    263.2637,
  274.6413, 271.6412, 267.2182, 264.8372, 262.9915, 261.8633, 261.4153, 
    263.7704, 263.7079, 260.7894, 259.5749, 260.4605, 261.0264, 261.5694, 
    262.9966,
  271.4783, 268.1287, 262.7965, 263.9868, 263.1554, 261.5782, 256.8496, 
    257.5137, 257.0859, 259.9352, 260.3451, 260.3897, 262.5233, 265.0368, 
    267.4225,
  271.9494, 269.4334, 264.1994, 263.2518, 262.9188, 259.7314, 257.5251, 
    258.1071, 258.1442, 257.3359, 259.2657, 262.6576, 263.8713, 264.3252, 
    265.4596,
  273.21, 272.563, 269.8335, 262.9477, 261.0205, 259.5255, 258.2751, 
    259.7805, 260.4313, 259.3082, 258.8208, 263.4076, 264.5181, 265.2086, 
    265.4718,
  274.1873, 273.4948, 272.5374, 265.2333, 261.6894, 258.0001, 257.0509, 
    259.9503, 261.0231, 261.6496, 260.722, 262.0511, 263.3761, 264.1001, 
    263.658,
  275.2324, 273.3194, 272.9534, 266.2266, 262.8588, 261.177, 258.2224, 
    256.4277, 257.54, 262.2218, 262.4999, 262.5162, 263.043, 265.1509, 
    267.3752,
  275.7518, 274.2651, 272.2456, 267.7186, 264.1224, 263.0877, 260.8698, 
    260.6413, 260.9499, 261.3937, 262.0377, 263.4374, 263.3935, 262.4393, 
    266.8405,
  276.0443, 274.9311, 272.6459, 266.3681, 263.5759, 263.3376, 262.4766, 
    262.3139, 261.7428, 261.5142, 262.3717, 263.7599, 265.1243, 264.007, 
    264.5121,
  276.3566, 275.1519, 270.9434, 264.294, 263.1133, 263.0827, 263.0107, 
    263.0621, 262.6502, 261.8529, 262.3731, 263.9811, 265.6158, 266.6118, 
    265.552,
  276.1412, 274.8317, 267.9231, 263.543, 262.6761, 262.9754, 263.518, 
    264.1303, 263.3796, 262.9366, 262.8099, 263.8694, 265.762, 267.2462, 
    267.437,
  274.6133, 271.3893, 264.8996, 264.4876, 263.2014, 263.2248, 263.8013, 
    265.7306, 265.0331, 262.9732, 262.5448, 263.5616, 265.3101, 267.3247, 
    268.6712,
  271.4696, 266.7993, 263.4125, 260.4735, 258.193, 257.77, 259.8994, 
    261.0974, 260.9506, 261.9272, 262.2903, 261.4519, 261.8548, 264.9428, 
    268.4324,
  270.7713, 267.0736, 262.5889, 259.7926, 259.369, 258.2012, 261.4723, 
    261.3105, 261.1668, 258.4611, 261.4572, 263.8253, 261.9623, 263.496, 
    266.8607,
  273.0701, 272.401, 268.3355, 262.941, 260.1972, 257.9664, 261.7821, 
    263.3157, 263.6435, 262.4954, 260.4164, 264.5666, 263.2967, 264.1236, 
    267.3006,
  274.0765, 273.3964, 272.3536, 265.328, 262.983, 260.178, 260.3229, 
    263.3932, 264.112, 264.4972, 262.932, 265.5431, 264.863, 261.3011, 
    266.6824,
  275.144, 273.2745, 272.8625, 266.3102, 263.7951, 263.0723, 262.6951, 
    259.3091, 260.7466, 265.1404, 265.2663, 266.8264, 265.9714, 261.1193, 
    265.9534,
  275.6791, 274.2105, 272.2214, 267.4861, 264.401, 263.1364, 262.983, 
    262.7726, 262.8983, 264.2027, 265.6567, 268.042, 267.3279, 264.8899, 
    265.1295,
  275.9918, 274.9279, 272.5992, 266.2591, 264.1157, 263.0954, 262.6894, 
    262.6668, 262.9219, 264.2067, 265.8171, 268.1017, 268.4717, 265.9439, 
    262.8603,
  276.3154, 275.179, 270.7427, 264.88, 264.0987, 263.6399, 262.7816, 
    261.8838, 262.1713, 263.7204, 265.5941, 266.695, 268.7001, 266.3709, 
    265.6323,
  276.1299, 274.7948, 266.9728, 263.9668, 264.2198, 262.5651, 262.2561, 
    262.9548, 262.8721, 264.166, 264.9226, 266.3335, 267.5389, 267.4844, 
    266.2669,
  274.6561, 271.4349, 263.985, 264.8459, 264.2575, 261.1354, 261.8661, 
    265.0412, 264.5537, 262.9551, 263.7319, 264.9743, 266.9847, 269.4731, 
    266.2866,
  267.6889, 265.4979, 262.8187, 259.5331, 258.9016, 257.5718, 259.0409, 
    260.6849, 262.8654, 264.3479, 265.8406, 265.977, 265.0783, 265.3708, 
    265.0965,
  268.4966, 265.2973, 262.4754, 260.9275, 260.5718, 259.5097, 261.2776, 
    263.5266, 264.1745, 261.8396, 266.3795, 267.0039, 266.5627, 264.4444, 
    264.9511,
  272.9338, 272.1741, 267.8148, 263.1199, 261.4907, 259.0813, 262.5807, 
    264.0272, 264.855, 265.7033, 266.2684, 267.4274, 267.0509, 265.5106, 
    266.4871,
  273.9908, 273.3442, 272.0104, 264.2664, 261.968, 261.2291, 260.1473, 
    263.3598, 265.2732, 266.5471, 266.7809, 267.0042, 266.6406, 265.1432, 
    268.125,
  275.0867, 273.2537, 272.6678, 265.6078, 263.3241, 262.3207, 261.1555, 
    260.7399, 262.8376, 267.203, 267.012, 266.7259, 266.3916, 265.8622, 
    268.9469,
  275.6424, 274.2311, 272.1625, 267.077, 263.6447, 262.0585, 261.4558, 
    262.4967, 264.5939, 265.9796, 266.9209, 267.2187, 266.5299, 266.2938, 
    268.6138,
  276.0287, 275.0382, 272.552, 265.907, 263.8153, 262.1466, 262.361, 262.753, 
    264.2497, 265.7147, 266.5656, 267.9231, 266.9526, 266.5347, 267.9124,
  276.3563, 275.3497, 270.0749, 262.7552, 263.6837, 262.4562, 262.7281, 
    262.7386, 263.1528, 264.7963, 265.8856, 267.5252, 267.9726, 267.0819, 
    267.5954,
  276.1853, 274.8603, 267.0324, 262.0805, 261.628, 262.1007, 262.7054, 
    264.8644, 264.9212, 265.7844, 265.0223, 267.0526, 268.3684, 267.8946, 
    266.9802,
  274.7419, 271.9193, 264.4446, 263.538, 261.4478, 261.5509, 261.9868, 
    266.5074, 266.5958, 264.9047, 262.9894, 265.008, 268.2803, 268.889, 
    267.1617,
  265.9352, 264.885, 260.8197, 261.8116, 259.8789, 259.5086, 260.9569, 
    264.8745, 266.2406, 266.0179, 267.5265, 267.473, 266.9507, 266.886, 
    266.3991,
  267.3902, 264.1004, 263.5823, 263.4414, 263.1088, 259.8885, 260.0909, 
    265.1693, 265.8154, 266.6323, 267.7541, 267.7484, 267.3734, 265.8266, 
    265.5318,
  273.0801, 272.26, 268.1657, 264.5055, 262.5232, 260.7003, 260.5763, 
    262.6329, 265.7709, 267.067, 267.8818, 267.9761, 267.5054, 267.2245, 
    266.5968,
  274.1683, 273.3963, 271.9833, 265.0835, 262.8214, 259.7456, 260.418, 
    261.8947, 265.1702, 266.7219, 267.5093, 268.5039, 268.2288, 268.123, 
    268.2792,
  275.2217, 273.4887, 272.6898, 266.5461, 263.7119, 263.1427, 264.1329, 
    261.4425, 262.8503, 267.044, 267.3408, 268.688, 268.4353, 268.5865, 
    269.0891,
  275.6927, 274.5, 272.3213, 267.2824, 264.2249, 263.445, 264.3786, 264.8481, 
    265.1762, 265.8015, 266.8319, 268.588, 268.8216, 268.6556, 269.4568,
  276.0323, 275.2397, 272.7559, 264.4365, 264.4673, 263.6328, 264.3119, 
    264.8475, 265.1744, 265.5746, 266.3743, 268.3701, 268.9461, 268.8948, 
    269.393,
  276.3364, 275.5027, 269.9498, 261.4952, 264.7697, 263.3679, 264.3939, 
    264.9358, 264.9394, 264.9695, 265.6225, 267.8546, 268.8905, 269.099, 
    269.2867,
  276.1885, 274.9609, 267.8936, 261.5996, 262.7845, 263.5123, 264.2685, 
    265.5844, 265.7014, 265.6377, 264.9127, 266.9787, 268.8245, 269.0482, 
    269.3448,
  274.7858, 272.1466, 266.3962, 261.9667, 264.0264, 263.4332, 262.739, 
    267.0561, 266.8182, 264.6313, 263.8057, 265.6083, 268.4757, 269.0343, 
    268.9771,
  265.9851, 266.472, 264.5549, 264.0268, 263.3854, 263.3695, 264.4742, 
    264.9229, 265.1423, 266.1425, 266.4668, 267.7731, 268.5002, 268.4709, 
    268.5283,
  268.7484, 267.5735, 266.2137, 264.6276, 263.6782, 263.8359, 263.5358, 
    261.5053, 261.2948, 265.382, 266.0616, 267.0094, 268.5481, 268.2126, 
    268.6777,
  273.1102, 272.4328, 268.7001, 265.3652, 263.8457, 262.2669, 261.3794, 
    260.6583, 263.1209, 265.5205, 265.4854, 266.8509, 268.2921, 269.1848, 
    269.4328,
  274.0768, 273.5421, 272.102, 266.1142, 264.5405, 263.5346, 261.8224, 
    260.0342, 261.5923, 264.6129, 264.9137, 266.1507, 268.2419, 268.4521, 
    269.0042,
  275.2074, 273.7119, 272.752, 267.0502, 264.5534, 264.4906, 264.6395, 
    260.3174, 261.2818, 264.5934, 264.6399, 266.0887, 268.1861, 268.0993, 
    268.9227,
  275.7106, 274.7584, 272.5411, 267.3983, 264.1589, 264.0444, 264.7148, 
    264.498, 263.2153, 263.3588, 264.093, 266.0651, 268.1575, 268.6272, 
    269.4679,
  276.0203, 275.3816, 272.9072, 265.4131, 264.3009, 263.903, 264.7569, 
    264.3997, 263.7044, 263.3703, 264.1387, 266.0562, 268.3097, 269.0006, 
    268.2497,
  276.3282, 275.6121, 270.9212, 264.4743, 263.9803, 263.6474, 264.6256, 
    264.6408, 263.846, 263.3562, 263.7624, 266.267, 268.1666, 267.6378, 
    268.6803,
  276.2494, 275.0401, 268.5915, 266.6253, 265.0323, 263.3053, 263.878, 
    265.3197, 265.0379, 264.5654, 264.0628, 266.3172, 267.9745, 265.8385, 
    266.6004,
  274.943, 272.4952, 270.0247, 268.133, 266.9393, 262.9637, 262.8952, 
    267.1182, 266.2815, 263.726, 263.4766, 266.1468, 267.0918, 265.3766, 
    266.3591,
  266.0878, 266.9652, 265.8599, 265.2761, 264.8363, 263.5026, 264.703, 
    264.1629, 261.037, 263.7296, 263.8911, 263.9071, 264.3846, 266.1194, 
    265.9503,
  268.1299, 268.6582, 267.5973, 266.2438, 265.3646, 264.3645, 264.1171, 
    259.65, 259.1276, 261.1484, 262.5344, 263.4656, 262.7519, 265.0578, 
    265.3004,
  273.294, 272.4554, 270.1468, 267.8695, 265.0755, 263.8847, 262.4608, 
    262.5647, 260.7649, 264.0856, 261.5309, 263.9857, 264.6962, 266.0276, 
    266.0379,
  274.2226, 273.4975, 272.2813, 268.877, 267.257, 266.0681, 262.9014, 
    261.8741, 261.6951, 262.2955, 263.3483, 263.5416, 264.7176, 266.2274, 
    266.9352,
  275.2611, 273.6862, 272.8485, 269.8291, 267.7642, 266.9699, 265.4835, 
    261.4258, 260.9226, 263.4912, 263.543, 262.9526, 264.8799, 265.4148, 
    265.0898,
  275.7232, 274.7236, 272.5422, 270.1376, 267.7785, 266.7209, 266.7497, 
    265.5487, 264.1141, 263.3677, 263.344, 263.3253, 264.7383, 264.2668, 
    264.9719,
  276.0005, 275.3205, 273.1002, 269.6455, 267.5745, 266.1884, 266.723, 
    266.6931, 265.6562, 263.81, 262.7174, 262.742, 265.4444, 265.0497, 
    265.3271,
  276.2945, 275.5107, 272.0744, 268.8888, 266.8612, 265.9693, 266.3073, 
    267.6841, 266.6554, 264.458, 262.8877, 263.6742, 265.8317, 266.4676, 
    267.4597,
  276.19, 274.8499, 270.2898, 268.2415, 267.6444, 266.6683, 266.2923, 
    267.538, 266.4385, 264.5871, 262.1739, 263.8049, 266.0192, 266.8087, 
    267.8838,
  274.8445, 272.4244, 269.4471, 268.4465, 267.0297, 265.5144, 265.3472, 
    267.6974, 266.0848, 264.6312, 263.0553, 265.7377, 266.0639, 267.7549, 
    268.5748,
  269.027, 267.1266, 267.0247, 266.4413, 266.5377, 266.5615, 264.8747, 
    264.4294, 265.1523, 265.1786, 265.5197, 264.6809, 263.9294, 264.6996, 
    265.7882,
  269.9394, 268.113, 269.1479, 268.6023, 268.3999, 268.3617, 266.5638, 
    265.7433, 264.6785, 264.1452, 263.4711, 263.2673, 261.3029, 263.3143, 
    264.2969,
  273.2441, 272.5256, 270.8027, 269.1957, 269.4117, 267.9137, 269.2457, 
    268.433, 267.2784, 265.885, 264.2276, 263.3907, 261.7024, 263.9764, 
    264.8506,
  274.1443, 273.4016, 272.5301, 269.4092, 267.7433, 268.3305, 266.6024, 
    268.053, 267.4202, 267.5742, 266.8989, 264.916, 262.4088, 263.9249, 
    264.192,
  275.2104, 273.4814, 272.9681, 269.0366, 266.5403, 266.4694, 266.4815, 
    263.498, 261.876, 266.3236, 266.9393, 265.8241, 263.2234, 263.0157, 
    262.3776,
  275.6427, 274.5303, 272.445, 267.6086, 265.4618, 265.171, 265.162, 
    265.3666, 263.8805, 264.0894, 265.8147, 266.2559, 264.3705, 262.1598, 
    262.8284,
  275.9202, 275.1571, 272.4092, 265.5617, 264.8799, 264.6089, 264.4187, 
    265.0418, 265.0556, 264.1787, 266.9161, 266.1798, 264.1657, 262.4758, 
    263.953,
  276.2014, 275.3347, 270.1581, 265.2217, 264.9811, 265.7005, 265.3211, 
    266.3278, 267.5693, 266.1593, 266.7514, 265.4686, 264.2019, 264.3636, 
    265.6627,
  276.0427, 274.6601, 268.2453, 265.4019, 265.7719, 266.5732, 267.0214, 
    267.2705, 266.8523, 265.3125, 266.3134, 264.7878, 263.9326, 265.1577, 
    265.7994,
  274.6943, 272.0785, 267.5938, 266.2057, 266.0983, 266.7067, 267.2534, 
    268.8813, 267.6928, 267.0648, 265.5466, 265.4875, 264.5957, 265.3199, 
    266.2518,
  269.4489, 265.2569, 268.1471, 264.4727, 263.4208, 262.7209, 264.0256, 
    265.8222, 264.745, 263.7023, 264.7202, 265.0408, 263.6896, 264.0993, 
    265.2648,
  270.8424, 268.0491, 268.4863, 267.3737, 267.5227, 267.8258, 267.6867, 
    267.3871, 266.4941, 264.6984, 264.6364, 265.4154, 264.3742, 262.94, 
    264.5643,
  273.3492, 272.6498, 270.6476, 267.5085, 267.1341, 266.5075, 266.4227, 
    265.7945, 267.8838, 267.2892, 265.175, 265.7868, 264.1986, 264.6605, 
    264.9041,
  274.2081, 273.4681, 272.6268, 269.3467, 267.6891, 267.6427, 264.7621, 
    265.0414, 262.5645, 267.5735, 266.0037, 266.5376, 265.7781, 265.1966, 
    264.6599,
  275.24, 273.5273, 273.0512, 270.2582, 267.5251, 267.1124, 266.1407, 
    262.2803, 261.1843, 263.3401, 268.1315, 267.2535, 266.0527, 266.0523, 
    260.7703,
  275.6469, 274.5444, 272.5388, 269.4497, 266.9262, 265.2602, 266.2268, 
    265.2986, 263.2422, 261.655, 267.6552, 268.3003, 266.7401, 263.2075, 
    262.6539,
  275.9051, 275.131, 272.3499, 267.9796, 265.6071, 265.7041, 266.5403, 
    267.4463, 265.8405, 262.1049, 265.3679, 268.5029, 266.8488, 263.2363, 
    265.3297,
  276.1891, 275.2916, 270.3396, 267.0365, 268.055, 267.4232, 267.5024, 
    268.4432, 265.8495, 265.757, 265.1773, 267.6952, 266.2593, 263.6686, 
    266.2512,
  276.0058, 274.5733, 268.7167, 266.8898, 266.7612, 266.2412, 269.4051, 
    269.2053, 266.868, 266.0885, 264.6752, 267.4344, 265.1618, 264.2442, 
    266.2081,
  274.5829, 271.8715, 267.8812, 267.59, 267.5442, 268.6977, 269.1682, 
    268.9185, 266.7501, 265.9442, 265.9725, 267.1462, 263.8532, 264.2299, 
    265.4101,
  270.6638, 268.5655, 269.8188, 269.8256, 268.2213, 265.4424, 266.2448, 
    266.7244, 266.5526, 268.011, 266.7093, 263.7506, 263.6189, 263.2601, 
    265.926,
  270.6129, 269.2926, 268.7251, 269.8061, 270.1979, 269.3672, 267.0266, 
    266.9186, 266.3718, 268.5387, 267.3775, 265.4645, 262.8099, 260.7007, 
    263.5393,
  273.6299, 272.9586, 271.4042, 271.2552, 271.2815, 269.6047, 268.6595, 
    267.973, 266.6434, 268.3918, 266.8051, 265.8178, 264.8555, 262.0302, 
    263.6427,
  274.4342, 273.6646, 272.8761, 269.6446, 269.339, 271.4948, 268.8481, 
    268.6308, 265.7898, 266.9693, 266.6771, 265.3239, 265.6053, 262.0525, 
    262.8098,
  275.3828, 273.7416, 273.2492, 270.0667, 266.9813, 267.6239, 266.0987, 
    265.7102, 263.581, 265.0302, 267.3139, 265.4375, 264.4674, 263.1295, 
    261.7831,
  275.7224, 274.704, 272.9172, 270.4276, 267.5866, 262.584, 267.1401, 
    266.7884, 265.321, 264.8338, 266.9456, 266.1032, 265.9863, 262.3311, 
    263.3857,
  275.9686, 275.2713, 272.4344, 268.7932, 267.8793, 262.6231, 266.651, 
    266.0469, 265.6782, 264.9936, 266.6337, 265.9061, 265.5525, 262.7793, 
    266.8637,
  276.2415, 275.3788, 270.8451, 268.1075, 268.7581, 265.649, 264.5673, 
    266.8313, 265.0021, 265.5121, 266.4567, 266.078, 264.305, 264.7341, 
    268.2462,
  276.0445, 274.5604, 268.4894, 269.0024, 268.5667, 266.5256, 267.3226, 
    267.4321, 266.2485, 265.6863, 265.1386, 265.6165, 263.4591, 267.1392, 
    268.5049,
  274.5568, 271.6647, 267.008, 268.5209, 267.4164, 267.278, 267.4061, 
    268.0737, 266.124, 265.7252, 265.5764, 266.3123, 263.4999, 267.0368, 
    268.5699,
  272.9221, 267.877, 267.4823, 267.8111, 268.8097, 267.8058, 266.3609, 
    268.1106, 267.7713, 269.5461, 267.4031, 263.5233, 265.7729, 267.0743, 
    269.4999,
  271.4517, 269.4409, 267.9539, 270.0539, 270.6339, 268.5485, 268.1581, 
    268.0783, 265.8504, 265.5888, 269.1061, 264.1056, 265.5918, 266.3349, 
    268.9795,
  273.9622, 273.1935, 271.4157, 269.2137, 269.089, 268.3493, 268.7021, 
    268.1528, 265.6997, 266.6655, 267.4261, 264.4278, 266.2431, 266.182, 
    268.3719,
  274.6399, 273.8395, 273.0579, 269.4849, 267.787, 269.0446, 268.4252, 
    269.3797, 265.915, 267.4804, 266.1617, 264.3623, 264.9435, 265.4589, 
    267.2664,
  275.5047, 273.9148, 273.469, 270.0468, 269.2166, 268.9691, 270.0488, 
    266.7235, 265.9366, 266.6954, 265.7986, 266.4614, 265.2254, 265.1115, 
    266.3893,
  275.8059, 274.8563, 273.2699, 269.7749, 267.4436, 264.8679, 269.1909, 
    270.1249, 267.5419, 266.6576, 267.6915, 266.5751, 265.9706, 264.5457, 
    266.463,
  276.0212, 275.431, 272.4353, 270.1275, 267.0606, 265.2237, 268.6883, 
    269.5787, 268.0154, 266.2921, 267.5727, 266.562, 266.5725, 266.1383, 
    267.8199,
  276.2792, 275.5171, 271.314, 266.5129, 267.9331, 265.2817, 265.0943, 
    268.3397, 267.279, 265.3813, 266.2953, 266.2701, 265.2068, 266.5693, 
    268.5743,
  276.0838, 274.5556, 267.3016, 266.3599, 266.3057, 265.4512, 267.4411, 
    268.4511, 267.7339, 265.1056, 266.3445, 265.9539, 264.5012, 267.0351, 
    268.3853,
  274.5694, 271.7184, 267.374, 267.4566, 266.7913, 267.4092, 268.0235, 
    268.5784, 267.0208, 265.5111, 266.1913, 266.0124, 264.4534, 267.299, 
    268.0939,
  273.4731, 268.1487, 267.3972, 269.6488, 268.9683, 269.1721, 270.0068, 
    270.6644, 270.7656, 270.3799, 269.3828, 267.6674, 267.2619, 267.0279, 
    268.6591,
  271.1006, 269.3916, 268.3063, 268.7599, 271.8575, 271.6331, 270.9995, 
    270.6165, 269.5974, 268.1322, 269.8849, 267.426, 266.7699, 267.4848, 
    269.892,
  274.5657, 273.5961, 271.8085, 268.179, 271.4786, 268.6595, 268.6287, 
    267.3809, 269.6393, 267.8876, 269.1332, 266.9082, 266.4498, 268.1242, 
    271.3295,
  274.8933, 273.9949, 273.2122, 270.3311, 266.9455, 268.5154, 270.116, 
    266.3372, 268.0435, 265.1484, 263.1735, 263.7421, 267.5229, 269.8027, 
    271.4174,
  275.5854, 274.0267, 273.6472, 270.6031, 269.7424, 270.6123, 270.4946, 
    264.9835, 262.8425, 267.4494, 265.0206, 266.5862, 269.4066, 270.4836, 
    270.5422,
  275.869, 275.0226, 273.7133, 269.1425, 270.4141, 269.3468, 268.459, 
    266.2868, 266.432, 266.3555, 267.4465, 268.4417, 270.0555, 270.4699, 
    270.5209,
  276.1021, 275.6511, 272.6648, 268.246, 268.8544, 269.3573, 270.4591, 
    266.8658, 266.5529, 266.776, 268.4394, 269.4614, 269.8225, 270.1223, 
    269.9571,
  276.39, 275.7343, 271.1808, 264.5091, 268.9099, 267.808, 269.2736, 
    268.4235, 266.5366, 267.2351, 268.8649, 269.4948, 269.5745, 269.4264, 
    269.2157,
  276.2007, 274.6503, 268.3327, 268.2819, 268.7418, 267.8437, 269.1478, 
    268.2152, 267.0836, 266.8839, 268.2402, 268.9331, 268.8831, 268.9276, 
    268.5653,
  274.6642, 271.7563, 267.0447, 267.9838, 268.4926, 268.5821, 268.6456, 
    268.2563, 267.1022, 267.3036, 267.8028, 268.1047, 268.3476, 268.1669, 
    268.1615,
  272.6473, 270.232, 268.8002, 271.177, 270.1617, 270.7248, 271.2828, 
    271.3394, 270.637, 270.5875, 270.2822, 270.7537, 270.4771, 270.0037, 
    269.3128,
  272.1346, 269.3157, 268.706, 270.6793, 271.1613, 271.6906, 271.4935, 
    270.8832, 269.9333, 270.4035, 269.4164, 270.9996, 270.7712, 269.6713, 
    269.2214,
  274.4532, 273.9581, 272.2756, 270.0095, 270.4467, 267.6527, 267.1029, 
    267.9774, 268.5237, 268.0404, 268.6517, 270.5034, 269.1752, 267.6377, 
    267.2145,
  275.3692, 274.4745, 273.4796, 270.0052, 265.3225, 266.9691, 266.6849, 
    265.3246, 268.1259, 269.8515, 269.0458, 268.454, 266.619, 266.7353, 
    267.7269,
  275.9023, 274.2761, 273.9803, 270.5222, 264.6571, 269.2817, 268.8394, 
    266.218, 264.4141, 265.632, 266.9968, 266.2204, 266.0435, 266.264, 
    269.9039,
  276.0576, 275.3156, 274.233, 269.1822, 266.718, 267.6759, 267.8882, 
    265.7199, 267.0527, 264.1212, 264.3336, 265.9418, 267.1639, 269.6585, 
    270.2956,
  276.313, 276.0401, 273.0672, 267.9919, 267.0029, 267.2992, 267.8776, 
    264.8752, 267.8618, 268.6632, 269.1774, 269.9811, 270.1019, 270.3398, 
    269.8647,
  276.6882, 275.9587, 270.7992, 266.5908, 267.6351, 267.7262, 267.2949, 
    266.33, 266.2534, 269.4848, 269.9368, 270.0414, 270.1089, 269.3933, 
    268.9639,
  276.4058, 274.653, 268.286, 268.9464, 268.965, 268.6227, 268.1424, 
    267.7723, 268.3616, 270.1459, 270.0925, 269.0177, 268.9739, 268.7476, 
    269.1761,
  274.7991, 271.9609, 268.3804, 268.6206, 268.3787, 268.4066, 268.3177, 
    268.5802, 269.8524, 269.7111, 269.3554, 268.6, 268.6688, 269.0477, 
    269.7583,
  274.4339, 272.1394, 271.68, 271.4691, 270.962, 269.8457, 268.9516, 
    268.5057, 267.5307, 268.4105, 270.6135, 268.33, 268.2534, 269.0453, 
    270.0334,
  272.3277, 270.8148, 270.5168, 271.3683, 270.8246, 271.4018, 269.3964, 
    268.3405, 267.1782, 267.6859, 269.5643, 268.7959, 267.2201, 269.5142, 
    267.9661,
  274.1299, 273.8724, 272.6491, 270.8758, 270.5477, 267.4453, 266.7316, 
    266.3992, 265.9341, 266.5083, 266.9558, 268.6107, 267.5745, 266.3505, 
    268.082,
  275.1544, 274.4158, 273.6088, 271.5437, 268.464, 268.0702, 264.379, 
    263.8116, 263.5464, 267.3777, 269.3415, 268.8735, 268.9823, 268.2769, 
    268.3715,
  275.8847, 274.4927, 274.2518, 271.4622, 266.0967, 266.4146, 265.4852, 
    264.7472, 262.2778, 266.4828, 269.0989, 269.2877, 270.0872, 267.3518, 
    267.1282,
  276.2243, 275.5777, 274.3176, 269.501, 265.572, 266.4094, 266.9859, 
    265.9974, 265.2463, 264.7664, 265.3293, 266.1313, 267.6996, 268.466, 
    269.6288,
  276.5531, 276.1909, 272.507, 267.0213, 265.9757, 267.1717, 267.1117, 
    266.529, 268.387, 266.7154, 269.547, 269.5259, 269.4589, 268.9221, 
    269.8483,
  276.899, 276.0442, 269.5274, 265.8671, 266.9332, 267.1381, 265.7169, 
    266.7844, 263.9851, 265.104, 267.1664, 268.8856, 269.659, 269.6458, 
    269.763,
  276.5717, 274.6494, 267.8175, 267.1764, 268.472, 265.8087, 264.6033, 
    264.6275, 268.362, 268.1854, 265.2947, 267.8985, 269.4174, 269.6028, 
    269.718,
  274.8551, 271.8864, 267.9578, 268.6208, 267.187, 268.8713, 267.3215, 
    268.1926, 269.4051, 269.1695, 266.7812, 269.5479, 269.6132, 269.5696, 
    269.9175,
  277.8656, 272.8303, 272.89, 272.9839, 273.0418, 272.691, 272.1966, 
    271.6826, 271.0173, 270.8149, 271.1079, 270.4245, 270.6152, 270.0578, 
    270.3928,
  272.7811, 272.8274, 272.9152, 273.0723, 272.9742, 272.4456, 271.8974, 
    271.5485, 270.9491, 269.8548, 270.2163, 269.4138, 268.5699, 269.7602, 
    268.8499,
  273.8852, 273.439, 272.8838, 272.8058, 272.4842, 271.6419, 270.5131, 
    269.894, 269.597, 268.5269, 268.139, 267.9932, 267.9578, 266.5793, 268.464,
  274.8787, 274.111, 273.3336, 272.5545, 271.8828, 271.0042, 267.3845, 
    267.8862, 267.815, 267.3771, 267.4724, 266.5267, 269.7398, 270.368, 
    267.4349,
  275.6814, 274.0036, 273.5945, 271.8785, 269.9375, 268.6939, 267.8434, 
    265.9618, 264.8687, 267.2596, 266.4984, 267.5964, 268.9157, 269.8187, 
    270.1369,
  275.6996, 274.7312, 273.173, 270.3527, 268.5087, 267.3436, 266.3906, 
    266.4072, 266.6837, 265.4058, 265.3401, 264.5211, 269.4492, 269.7728, 
    269.3949,
  276.0081, 275.4105, 272.4195, 268.0346, 266.8408, 266.3272, 265.6366, 
    265.6507, 267.7355, 268.439, 269.1674, 267.6862, 268.6392, 269.1161, 
    269.1693,
  276.416, 275.7113, 270.3046, 266.782, 266.2291, 268.4746, 266.3022, 
    267.6482, 267.0696, 268.3069, 267.3934, 267.0586, 268.062, 269.732, 
    270.1526,
  276.3662, 274.6511, 268.6423, 267.607, 269.2767, 267.0476, 266.7238, 
    267.7598, 268.4757, 268.7751, 267.2112, 269.2377, 269.651, 269.9272, 
    270.2083,
  274.8631, 272.1831, 269.2994, 269.4275, 268.2194, 268.696, 268.5045, 
    268.6829, 268.7461, 269.1656, 267.4014, 269.0327, 269.3639, 269.3569, 
    269.9317,
  275.5893, 271.8321, 271.5572, 272.0122, 272.2462, 272.3168, 272.3054, 
    272.4585, 272.6675, 272.837, 272.9664, 272.9773, 273.0798, 272.785, 
    272.4225,
  272.4711, 272.121, 272.0113, 272.1887, 272.4698, 272.5488, 272.5502, 
    272.6473, 272.7574, 272.8967, 272.9857, 272.9984, 272.7923, 272.3509, 
    271.8189,
  273.7861, 273.3622, 272.6157, 272.1126, 272.4621, 272.4096, 272.3235, 
    271.449, 271.6229, 272.0627, 272.3517, 272.4957, 272.1996, 271.7953, 
    271.375,
  274.821, 274.0681, 273.3397, 272.1519, 271.502, 271.4738, 268.9185, 
    269.0903, 269.5712, 270.4318, 270.8996, 271.2606, 271.2558, 270.7787, 
    270.4042,
  275.5162, 273.8838, 273.4938, 270.406, 269.1204, 268.9252, 269.0441, 
    266.5298, 265.4501, 269.413, 269.6456, 269.7326, 269.9092, 269.9792, 
    270.0497,
  275.5381, 274.3419, 272.5472, 268.5449, 267.1972, 266.8246, 266.8403, 
    268.0059, 268.5621, 268.7495, 268.9378, 268.8768, 269.056, 269.2071, 
    269.2274,
  275.8123, 274.9837, 271.3886, 266.9377, 266.2051, 265.7568, 265.4357, 
    265.6228, 266.502, 268.1898, 268.5648, 268.4823, 268.5316, 268.5434, 
    268.5766,
  276.2377, 275.4029, 269.8911, 267.5688, 266.5166, 266.4653, 265.7935, 
    265.6398, 265.5619, 266.3442, 267.4659, 267.7416, 268.0506, 268.3695, 
    268.3607,
  276.2261, 274.5503, 269.0369, 268.3045, 267.9481, 267.834, 266.5588, 
    266.8072, 266.6967, 266.4478, 266.7031, 267.2795, 267.5851, 267.6299, 
    269.5934,
  274.8497, 272.47, 269.4732, 268.7723, 267.9708, 267.9772, 268.1444, 266.61, 
    266.632, 266.7685, 267.1041, 267.8816, 268.0633, 268.8677, 269.8582,
  275.1505, 272.2234, 271.5662, 270.4087, 271.3055, 270.941, 270.7544, 
    266.7937, 266.4386, 267.3123, 269.3043, 270.0685, 270.8922, 271.4802, 
    272.1526,
  272.4484, 271.9355, 271.299, 270.0883, 270.4642, 271.2475, 270.3102, 
    265.8422, 265.6718, 266.347, 268.4371, 270.1438, 270.4912, 271.2237, 
    272.1786,
  273.6659, 273.2979, 272.5398, 269.9136, 269.1084, 269.7325, 269.9647, 
    265.0145, 264.998, 265.816, 267.2059, 269.2965, 270.8048, 271.7087, 
    272.4626,
  274.7532, 274.0355, 273.3506, 270.8522, 267.6688, 269.0504, 266.6783, 
    264.8118, 265.028, 266.0605, 266.7236, 268.5218, 270.7477, 271.9237, 
    272.4912,
  275.4332, 273.8318, 273.4971, 269.2151, 266.4536, 265.1775, 269.7617, 
    265.645, 265.183, 266.9105, 266.9958, 268.0268, 270.4883, 271.9358, 
    272.6301,
  275.5296, 274.2998, 272.5528, 267.5771, 265.3777, 264.6291, 269.5013, 
    269.4568, 268.9615, 267.6675, 266.3625, 268.4978, 269.8728, 270.9886, 
    271.9796,
  275.8187, 274.9866, 271.8236, 268.4653, 265.439, 265.6949, 264.4511, 
    268.1559, 267.753, 266.4417, 265.5403, 268.4888, 269.5587, 270.1146, 
    270.7583,
  276.2529, 275.4455, 270.8577, 269.1948, 268.0547, 267.4534, 264.4361, 
    264.5682, 267.0166, 264.6558, 266.1269, 268.6241, 269.6069, 269.927, 
    270.1992,
  276.3358, 274.6036, 269.8661, 269.0381, 268.4709, 268.2362, 265.4065, 
    264.857, 264.5726, 264.5085, 265.7734, 268.88, 269.7539, 270.1382, 
    270.4075,
  274.9014, 272.6025, 269.9039, 269.2976, 268.9356, 266.2763, 266.692, 
    265.355, 264.4954, 264.9313, 266.8832, 269.2698, 270.1127, 270.3943, 
    270.6928,
  273.762, 271.5305, 271.2699, 271.8176, 271.9525, 271.8871, 271.8578, 
    271.0617, 269.9031, 269.9068, 269.8172, 268.6317, 267.7192, 266.0183, 
    265.0982,
  272.1912, 271.7954, 271.6451, 271.6977, 272.0429, 271.9491, 271.5884, 
    269.903, 268.7236, 268.4675, 269.0451, 267.8057, 265.0626, 264.2186, 
    264.7812,
  273.5456, 273.1957, 272.5397, 271.3954, 271.4949, 270.4321, 270.1658, 
    268.6023, 267.9025, 267.3172, 267.2219, 266.7988, 264.6609, 264.6769, 
    267.7532,
  274.6894, 273.9798, 273.2523, 271.397, 270.2062, 269.9834, 266.9648, 
    267.9521, 267.5594, 266.9604, 266.0739, 264.5042, 264.7688, 268.1364, 
    270.2362,
  275.2002, 273.6436, 273.2956, 269.5797, 268.7982, 268.5663, 269.2522, 
    265.463, 265.2094, 266.8381, 264.9402, 263.8223, 267.028, 270.4048, 
    272.167,
  275.4449, 274.1661, 272.2422, 268.2664, 267.5356, 267.6837, 268.4409, 
    268.881, 268.1951, 268.6669, 267.5353, 266.74, 269.728, 271.5522, 272.7938,
  275.8504, 274.9544, 271.1903, 267.3621, 267.4731, 267.811, 267.4293, 
    267.6843, 268.3787, 268.5569, 264.9007, 269.3815, 270.8946, 271.9558, 
    272.7876,
  276.3896, 275.4053, 269.8579, 268.3763, 268.2954, 268.1841, 266.6398, 
    264.7443, 268.5661, 264.4819, 266.9087, 270.7022, 271.176, 271.2412, 
    271.6643,
  276.5786, 274.5882, 269.5614, 269.4304, 269.6003, 269.5045, 269.0498, 
    263.9268, 263.9753, 266.0303, 269.5542, 271.2842, 270.844, 270.8749, 
    271.0834,
  275.0961, 272.7882, 270.6124, 269.3846, 270.112, 263.8595, 264.0766, 
    264.7361, 264.4154, 268.0384, 270.1413, 271.1196, 270.2555, 270.389, 
    270.5244,
  276.5512, 272.1715, 271.5729, 269.5234, 267.5974, 267.2228, 267.8537, 
    269.2151, 270.6751, 271.5167, 271.9098, 270.8034, 269.8889, 269.2818, 
    269.8195,
  272.4972, 272.0956, 271.4135, 268.9095, 266.8508, 267.0207, 267.4083, 
    268.2339, 269.6221, 270.1749, 270.0099, 269.331, 268.8456, 268.0186, 
    268.1021,
  273.5631, 273.3004, 272.5722, 268.2912, 266.104, 266.7851, 266.9005, 
    267.3434, 267.9495, 268.4698, 268.088, 267.8439, 267.1292, 266.8252, 
    268.0637,
  274.6907, 274.0492, 273.3475, 269.4129, 266.307, 268.2648, 266.7614, 
    267.0693, 267.1999, 267.9817, 268.4915, 268.0585, 267.4772, 267.8209, 
    270.853,
  275.3121, 273.6663, 273.4922, 268.0374, 266.608, 268.4642, 269.1729, 
    264.9891, 264.5889, 268.6315, 269.097, 269.7816, 270.9787, 271.9656, 
    272.3401,
  275.8661, 274.2515, 272.5975, 269.8765, 268.7792, 268.21, 267.8275, 
    268.5118, 268.4276, 269.6013, 270.1952, 271.0052, 272.24, 272.4796, 
    272.4789,
  276.4026, 275.0954, 272.5062, 270.3637, 269.7987, 269.1871, 268.4157, 
    268.2054, 268.5651, 269.7479, 270.6083, 271.7834, 272.5621, 272.6642, 
    272.7155,
  276.6949, 275.544, 272.1703, 271.0489, 270.5502, 270.0022, 269.1448, 
    268.6662, 268.5625, 268.9802, 270.9115, 271.873, 272.5521, 272.7444, 
    272.6251,
  276.6805, 274.7268, 270.7006, 270.4897, 270.9471, 270.4856, 269.8089, 
    265.8671, 267.6941, 269.9864, 270.8708, 271.3343, 271.663, 271.6545, 
    271.6708,
  275.1983, 272.909, 270.5266, 269.2862, 270.0642, 269.666, 267.9685, 
    265.9159, 269.2648, 270.5777, 270.5334, 270.5213, 270.5316, 270.899, 
    271.1752,
  278.927, 272.8116, 272.7104, 271.0758, 268.1495, 265.0035, 262.3561, 
    264.3937, 269.1754, 270.9044, 271.8872, 272.0394, 271.8209, 271.6017, 
    271.8227,
  273.0515, 272.7296, 272.139, 270.2454, 268.1453, 264.9627, 262.3462, 
    264.4752, 267.3019, 270.968, 272.0481, 272.0872, 271.4164, 271.2793, 
    271.9814,
  274.109, 273.7713, 272.7294, 269.4062, 266.581, 264.9511, 263.3729, 
    264.2441, 266.9268, 270.6189, 271.8304, 272.3534, 272.1276, 271.9911, 
    272.1153,
  275.1367, 274.5688, 273.3708, 270.821, 264.8977, 267.031, 265.8045, 
    264.7083, 266.6883, 269.6341, 271.4214, 272.326, 272.3564, 272.2473, 
    272.0433,
  275.7537, 274.2461, 273.5739, 269.8896, 266.9943, 269.1828, 269.773, 
    265.5474, 265.1526, 269.3229, 271.148, 272.091, 272.2128, 271.9621, 
    271.8864,
  276.3818, 274.7505, 273.0456, 271.0264, 269.7906, 269.3942, 269.5671, 
    269.5847, 267.846, 269.7581, 271.1459, 272.0304, 271.8391, 271.3733, 
    271.5179,
  276.8919, 275.3756, 273.0018, 271.8182, 270.8156, 270.4456, 270.3979, 
    270.0469, 267.2477, 269.6995, 270.7205, 271.567, 271.4698, 271.2706, 
    271.3098,
  277.1143, 275.8942, 271.5266, 271.1609, 270.2186, 271.885, 271.3875, 
    270.1624, 269.2777, 269.4495, 270.4487, 271.1289, 271.1994, 270.9227, 
    271.0659,
  276.867, 274.8521, 269.9768, 269.805, 271.6829, 271.7041, 270.7324, 
    267.4147, 269.2628, 269.4674, 270.3926, 270.8857, 270.9721, 270.8238, 
    271.2493,
  275.3699, 273.0612, 270.2385, 269.7219, 269.6066, 270.5213, 269.5112, 
    267.3339, 269.6216, 269.9421, 270.5972, 270.7669, 270.9951, 271.0727, 
    271.3567,
  275.3833, 272.3206, 271.3403, 269.0782, 266.6301, 264.7541, 262.8832, 
    263.1219, 266.1242, 270.0351, 271.4331, 271.7574, 271.7838, 271.7358, 
    271.5295,
  272.8431, 272.453, 271.487, 268.7591, 267.4744, 265.1384, 263.2982, 
    264.0806, 264.1912, 269.7346, 270.8028, 271.4578, 271.8766, 270.9266, 
    270.7777,
  273.8986, 273.5408, 272.7378, 269.2107, 267.7163, 265.9895, 265.7228, 
    268.2157, 265.0523, 269.5168, 270.5897, 271.4443, 271.8142, 271.2961, 
    271.3374,
  274.9657, 274.3672, 273.4338, 270.5984, 266.1196, 268.2334, 267.8021, 
    266.859, 266.3434, 269.408, 270.6033, 271.2486, 271.7665, 271.6777, 
    271.6759,
  275.5002, 274.0798, 273.6761, 271.041, 267.4668, 270.0043, 270.6091, 
    266.9914, 265.7662, 269.3344, 270.4952, 271.171, 271.9427, 271.9797, 
    272.1283,
  275.9968, 274.6931, 273.1505, 271.6095, 271.4576, 270.8253, 269.1385, 
    269.8135, 268.9324, 269.9105, 270.9362, 271.4192, 272.128, 272.1892, 
    272.3571,
  276.4839, 275.3339, 272.4948, 269.6249, 269.5814, 270.4591, 270.5129, 
    269.956, 268.6684, 270.068, 270.2363, 271.0722, 272.1338, 272.2655, 
    272.3932,
  276.9158, 275.8029, 271.2945, 269.9065, 269.9247, 269.6691, 269.4481, 
    269.1246, 270.1285, 269.9684, 270.9434, 271.5443, 272.2038, 272.3597, 
    272.4257,
  276.7469, 274.7768, 270.7913, 270.05, 269.7533, 269.3943, 268.637, 
    269.2438, 270.3038, 270.4142, 271.0215, 271.6631, 272.306, 272.4198, 
    272.1785,
  275.3684, 273.2361, 270.939, 269.9786, 269.3785, 268.3658, 268.6353, 
    269.7092, 270.275, 270.6971, 271.2189, 271.9981, 272.4346, 272.5326, 
    272.2263,
  273.7144, 271.0298, 269.6036, 267.8382, 268.5753, 267.4148, 266.7014, 
    267.0469, 268.8743, 270.241, 271.2254, 272.0122, 272.2278, 272.1431, 
    272.2593,
  272.2625, 271.8749, 271.1211, 269.5236, 269.8896, 269.6927, 268.3398, 
    268.9199, 268.2212, 270.2498, 271.2013, 271.95, 271.9478, 271.7224, 
    271.9041,
  273.7815, 273.4599, 272.7976, 270.1497, 269.1106, 268.2764, 269.7012, 
    269.8997, 269.7715, 270.315, 271.0903, 271.7264, 271.9709, 271.6924, 
    271.8185,
  274.8811, 274.3274, 273.4699, 271.3036, 269.2344, 269.8163, 267.8147, 
    268.2304, 269.3271, 270.2125, 270.4994, 271.5726, 271.4542, 271.6265, 
    271.9681,
  275.4123, 274.0129, 273.7428, 270.2868, 269.131, 269.3332, 270.0277, 
    266.6031, 266.3297, 270.3292, 270.7358, 271.2619, 271.616, 272.0668, 
    272.1635,
  275.7862, 274.5873, 273.1523, 269.7998, 269.3148, 269.4463, 269.5557, 
    269.4028, 269.731, 270.4582, 271.4642, 271.2358, 271.8497, 272.2334, 
    272.4591,
  276.1872, 275.2466, 272.17, 269.3525, 269.3346, 269.4789, 269.4449, 
    269.5028, 269.8919, 270.6342, 271.0081, 271.7663, 272.2661, 272.4982, 
    272.5532,
  276.6614, 275.6668, 271.0373, 269.6252, 269.5198, 269.3463, 269.3189, 
    269.4396, 270.1044, 270.4665, 271.0621, 271.9464, 272.366, 272.4883, 
    272.4187,
  276.575, 274.7312, 270.1038, 269.7024, 269.5532, 269.2429, 268.8631, 
    269.3409, 270.1456, 270.6302, 270.8801, 271.9844, 272.4412, 272.3327, 
    272.1308,
  275.3669, 273.2621, 270.9169, 269.9096, 269.4939, 268.9758, 268.9175, 
    269.5233, 270.215, 270.4886, 271.0621, 271.8967, 272.2929, 272.4593, 
    272.2092,
  273.3308, 271.487, 270.5279, 269.6464, 270.2054, 270.045, 269.3924, 
    269.4818, 269.9434, 270.2455, 270.771, 270.8609, 271.4082, 271.985, 
    272.0325,
  272.1537, 271.9752, 271.4077, 270.2057, 270.3762, 270.2957, 269.5151, 
    269.5545, 270.2301, 270.4509, 270.6439, 271.0532, 271.4648, 271.3586, 
    272.0831,
  273.819, 273.5212, 272.8695, 270.6857, 269.727, 267.977, 269.3131, 
    269.8872, 269.9229, 270.1701, 270.5473, 271.2096, 271.7362, 272.0247, 
    272.4285,
  274.912, 274.4008, 273.513, 271.2032, 269.1872, 269.6835, 267.5082, 
    269.0685, 269.4438, 270.211, 270.3931, 271.7437, 272.2156, 272.2602, 
    272.6761,
  275.5275, 274.1454, 273.7714, 270.155, 269.366, 268.9596, 269.5091, 
    265.8454, 266.2209, 270.2259, 270.9342, 272.1339, 272.3896, 272.3279, 
    272.4705,
  275.8692, 274.6662, 273.1161, 269.6966, 269.4583, 269.0003, 268.7694, 
    268.9815, 269.4395, 270.1195, 271.8403, 272.6375, 272.6569, 272.3318, 
    272.2664,
  276.2604, 275.3228, 272.2017, 269.4066, 269.541, 269.0797, 268.5882, 
    269.1415, 269.9712, 270.7151, 272.175, 272.7792, 272.4824, 272.3796, 
    272.3005,
  276.7117, 275.6948, 271.1494, 269.8669, 269.563, 269.0505, 268.9032, 
    269.5211, 270.4821, 271.2383, 272.3691, 272.7385, 272.5884, 272.3536, 
    271.9713,
  276.6557, 274.6809, 270.915, 270.136, 269.4811, 269.1004, 269.3184, 
    270.0352, 270.6825, 271.5418, 272.3676, 272.7133, 272.6323, 272.3444, 
    271.9878,
  275.4164, 273.3827, 271.4815, 270.4404, 269.5462, 269.1598, 269.5481, 
    270.5272, 271.1843, 272.1785, 272.6064, 272.7635, 272.6631, 272.5354, 
    272.022,
  273.5918, 271.7981, 271.2368, 270.2858, 269.3383, 270.2611, 269.4415, 
    269.9101, 270.4402, 270.8337, 271.4204, 271.8644, 272.3478, 272.5089, 
    272.7188,
  272.2839, 272.1509, 271.8029, 270.6485, 270.6492, 270.4213, 269.6626, 
    269.1962, 269.3944, 270.6344, 271.1501, 271.7079, 271.9324, 272.0403, 
    272.5643,
  274.1119, 273.7001, 272.9109, 271.0956, 270.3653, 268.5046, 269.8594, 
    269.7796, 269.8728, 270.3611, 270.9614, 271.3737, 271.7244, 272.0738, 
    272.5176,
  275.1376, 274.5998, 273.5279, 271.7332, 270.2946, 270.1516, 268.2752, 
    270.3208, 270.3233, 270.2581, 270.5764, 271.0091, 271.644, 272.0106, 
    272.2392,
  275.7815, 274.2678, 273.7472, 271.2972, 270.4469, 270.4388, 270.5818, 
    267.3527, 267.5096, 270.961, 270.7129, 270.6855, 271.507, 271.8939, 
    272.3008,
  276.1597, 274.7252, 273.0523, 271.3425, 270.7645, 270.7014, 270.9983, 
    270.9943, 270.9917, 270.9275, 271.0586, 271.0316, 271.4124, 271.8627, 
    272.164,
  276.4036, 275.334, 272.6505, 271.254, 271.1017, 271.4003, 271.4066, 
    271.4681, 271.3019, 271.4446, 271.5077, 271.4564, 271.7267, 271.9247, 
    272.0721,
  276.7382, 275.6374, 272.0694, 271.2808, 271.2799, 271.7096, 271.6335, 
    271.6497, 271.4974, 271.6255, 271.7952, 272.0478, 271.8627, 271.8974, 
    272.0743,
  276.6384, 274.5873, 271.7231, 271.7765, 271.5466, 271.9051, 271.7246, 
    271.7398, 271.6376, 271.7249, 272.4535, 272.6836, 271.0881, 271.3143, 
    272.1602,
  275.3812, 273.3088, 271.9477, 271.8173, 271.369, 271.9941, 271.8873, 
    271.8426, 271.9343, 272.2762, 272.7239, 272.8661, 272.6469, 272.2613, 
    272.282,
  274.7122, 271.7315, 271.6263, 271.4357, 271.3569, 271.4718, 271.3738, 
    271.5663, 271.5238, 271.9127, 272.25, 271.4272, 272.0383, 272.1853, 
    272.391,
  272.297, 272.4356, 272.0596, 271.5904, 271.8047, 271.7503, 271.6432, 
    271.7302, 271.8127, 272.0122, 272.4442, 272.0048, 271.5378, 271.4138, 
    272.3882,
  274.3512, 273.8821, 272.9392, 271.8701, 271.8521, 270.253, 271.7299, 
    271.6983, 272.1945, 271.9517, 272.0514, 272.1605, 271.7773, 271.4384, 
    272.2021,
  275.4589, 274.6691, 273.537, 272.2429, 271.8202, 272.2137, 270.5879, 
    271.2826, 272.1501, 272.1926, 272.1532, 272.2932, 271.9014, 271.3117, 
    271.7074,
  275.9272, 274.3089, 273.7394, 271.9931, 271.9054, 272.2025, 272.084, 
    269.7947, 269.5282, 272.2159, 272.3795, 272.2236, 271.9036, 271.2705, 
    271.356,
  276.3037, 274.7787, 273.0155, 271.821, 272.0901, 272.5052, 272.5758, 
    272.6023, 272.7373, 272.6843, 272.8665, 272.1999, 272.0653, 271.4436, 
    271.4514,
  276.46, 275.3594, 272.5444, 272.0232, 272.3142, 272.5957, 272.6, 272.5552, 
    272.6457, 272.6266, 272.9109, 272.2036, 272.1649, 271.3109, 271.2212,
  276.7669, 275.586, 272.164, 272.1334, 272.3317, 272.4658, 272.4929, 
    272.5411, 272.6205, 272.7834, 272.8757, 272.8203, 272.1086, 271.266, 
    271.2532,
  276.6749, 274.5862, 272.0718, 272.2994, 272.4413, 272.5751, 272.4338, 
    272.2388, 272.2019, 272.2777, 272.4577, 272.7386, 272.0263, 271.2483, 
    271.5434,
  275.4984, 273.4508, 272.27, 272.3134, 272.4707, 272.5727, 272.5603, 
    272.1315, 272.187, 272.6108, 272.7775, 272.7505, 272.1582, 271.1736, 
    271.5721,
  274.4668, 271.9319, 271.9815, 271.8844, 271.8225, 272.0663, 271.8944, 
    271.9319, 271.7784, 272.1227, 272.7431, 272.0119, 272.2377, 270.0109, 
    271.0262,
  272.2483, 272.5574, 272.3236, 271.4666, 272.2567, 272.3631, 272.1391, 
    271.8692, 271.9373, 272.1653, 271.6108, 271.0013, 272.0526, 272.013, 
    271.4776,
  274.3677, 273.9583, 272.9971, 272.0935, 272.4992, 270.9192, 271.9911, 
    271.7021, 271.5429, 272.2046, 271.2195, 272.3347, 272.1592, 272.2355, 
    272.2296,
  275.4656, 274.697, 273.5617, 272.4029, 272.3747, 272.6295, 271.0738, 
    271.8503, 271.1947, 271.9982, 271.9283, 272.4565, 271.8269, 271.2751, 
    270.7661,
  276.0187, 274.3875, 273.7568, 272.1609, 272.5348, 272.8335, 272.8633, 
    270.0983, 269.8134, 271.7498, 272.6111, 272.4376, 271.8571, 270.8661, 
    269.6723,
  276.3781, 274.843, 273.0133, 272.175, 272.6387, 272.8927, 272.9708, 
    272.3428, 271.6495, 272.5558, 272.8165, 272.1946, 271.6625, 271.2523, 
    270.5023,
  276.503, 275.3891, 272.803, 272.3716, 272.6475, 272.8564, 272.6691, 
    271.7435, 272.0041, 272.7715, 272.505, 272.1409, 271.9148, 271.848, 
    270.8079,
  276.8059, 275.5299, 272.4691, 272.4482, 272.5594, 272.6574, 272.6797, 
    272.6554, 272.7177, 272.8002, 272.6048, 272.1607, 271.7863, 271.8178, 
    271.3204,
  276.6926, 274.5329, 272.212, 272.5407, 272.5888, 272.4499, 272.4806, 
    272.3743, 272.3908, 272.5013, 272.5489, 272.0662, 271.8489, 271.6957, 
    271.8071,
  275.5024, 273.6176, 272.3721, 272.5637, 272.6921, 272.6518, 272.5955, 
    272.1217, 272.3035, 272.7761, 272.6603, 272.178, 271.7561, 271.7014, 
    271.9761,
  274.4258, 272.4156, 272.4321, 272.1924, 271.5922, 271.0398, 272.0684, 
    272.3885, 271.3759, 271.8194, 272.5172, 272.2759, 272.3842, 270.1573, 
    272.5066,
  272.5284, 272.7429, 272.5063, 271.9134, 272.3523, 272.332, 272.2586, 
    272.458, 272.2133, 271.9763, 271.8495, 271.9925, 269.0498, 272.1218, 
    272.6149,
  274.5649, 274.1163, 273.1067, 272.1454, 271.4941, 272.2979, 272.3047, 
    272.614, 272.2346, 272.0578, 271.4378, 271.8378, 268.5228, 270.5839, 
    272.7371,
  275.5524, 274.8285, 273.6525, 272.5849, 272.1844, 272.3978, 272.1593, 
    272.5404, 272.0917, 272.1859, 271.6606, 272.0126, 272.3323, 272.2101, 
    272.6306,
  276.1417, 274.5678, 273.8545, 272.4723, 272.7508, 271.8766, 272.5734, 
    270.1094, 268.8986, 272.2484, 271.7609, 272.2213, 271.0667, 271.9666, 
    272.4401,
  276.43, 274.9373, 273.093, 272.3871, 272.5573, 272.4391, 272.3475, 
    271.0193, 271.1815, 272.0706, 272.1811, 272.2702, 272.5017, 272.0201, 
    272.4929,
  276.519, 275.4382, 272.8747, 272.3998, 272.3613, 272.2902, 271.0108, 
    270.7042, 271.915, 272.2903, 272.4738, 272.6267, 272.6174, 272.3167, 
    272.5417,
  276.7738, 275.5287, 272.5016, 271.7754, 272.1198, 272.2076, 272.3785, 
    272.2482, 272.157, 272.3491, 272.3336, 272.3991, 272.4627, 272.1455, 
    272.4018,
  276.6234, 274.5508, 272.0637, 271.9744, 272.1431, 272.2776, 272.0598, 
    272.1049, 272.2612, 272.2665, 272.3094, 272.3144, 272.3914, 272.442, 
    272.363,
  275.5194, 273.7306, 272.3019, 272.3651, 272.5296, 272.5525, 272.4778, 
    272.0336, 272.1721, 272.4855, 272.5762, 272.338, 272.3203, 272.3188, 
    272.2831,
  277.0735, 272.727, 273.1712, 272.1984, 271.7218, 271.8544, 271.9337, 
    271.9602, 271.9896, 269.5778, 273.252, 271.8145, 271.972, 270.0745, 
    272.4409,
  272.5638, 272.8018, 272.7068, 271.9363, 272.2245, 272.047, 271.7841, 
    272.1074, 271.5534, 271.9695, 272.3726, 272.2826, 267.2344, 271.7552, 
    272.1725,
  274.3676, 274.1567, 273.2983, 272.0465, 272.0185, 272.1003, 271.9296, 
    271.9276, 272.0277, 272.3734, 272.3822, 272.061, 267.1994, 268.6813, 
    272.3692,
  275.2785, 274.8431, 273.8421, 272.6578, 272.1516, 272.5518, 270.0955, 
    272.7745, 272.2686, 271.4318, 272.2987, 271.9897, 268.6005, 270.1673, 
    272.7712,
  276.0078, 274.7242, 274.1344, 272.4105, 272.3761, 272.3108, 272.1942, 
    271.0721, 270.0917, 270.1694, 272.1742, 270.0349, 269.3889, 271.7406, 
    272.945,
  276.296, 275.0078, 273.2466, 272.1957, 271.2124, 271.672, 271.7, 270.2493, 
    270.0671, 269.3256, 269.531, 268.841, 271.114, 272.8136, 272.9349,
  276.4341, 275.4872, 272.696, 272.0736, 272.1591, 272.026, 271.5656, 
    271.9542, 269.5306, 268.9164, 271.92, 272.287, 272.7072, 272.9321, 
    272.9347,
  276.7214, 275.6316, 272.0933, 270.1238, 271.5458, 271.7886, 272.0316, 
    272.0155, 271.6487, 272.4747, 272.1664, 272.7379, 272.8345, 272.8238, 
    272.7758,
  276.6109, 274.6237, 271.9164, 271.8097, 271.8565, 272.0219, 272.2375, 
    272.2772, 272.3954, 272.442, 272.8232, 272.8621, 272.795, 272.6775, 
    272.4989,
  275.6119, 273.9186, 272.1729, 271.618, 272.1661, 272.3418, 271.6628, 
    272.0129, 272.4145, 272.7879, 272.9887, 272.8972, 272.7003, 272.6081, 
    272.3857,
  279.2921, 273.0654, 275.1376, 272.3711, 271.9095, 271.4294, 270.481, 
    270.2238, 270.607, 272.1327, 272.8759, 272.4117, 268.6522, 272.3218, 
    272.455,
  272.7846, 272.8493, 272.7125, 271.9518, 272.0634, 271.6748, 271.5138, 
    271.3443, 271.5718, 270.0969, 269.4746, 268.2523, 268.1786, 271.8232, 
    271.9871,
  274.2144, 273.9681, 273.2253, 272.0292, 271.9846, 270.5249, 271.2299, 
    271.3232, 271.5114, 272.1094, 272.1601, 269.0616, 270.9968, 270.6539, 
    272.5541,
  275.0371, 274.5853, 273.7112, 272.655, 272.0382, 272.0502, 269.7779, 
    271.5265, 271.8387, 271.9564, 269.2071, 270.3598, 271.1068, 271.7093, 
    272.9404,
  275.7684, 274.587, 274.0681, 272.3478, 272.0056, 272.1623, 271.5018, 
    269.8302, 268.4066, 269.4719, 272.2094, 271.5437, 271.2026, 272.5851, 
    273.0232,
  276.1263, 274.9661, 273.3407, 271.903, 271.3043, 272.0956, 272.0589, 
    269.8793, 268.6453, 268.1036, 271.9527, 271.3412, 271.8897, 272.9001, 
    272.9307,
  276.3665, 275.5082, 272.6547, 271.5701, 271.8422, 271.8012, 271.6276, 
    269.5694, 268.2587, 270.4555, 271.8867, 271.8722, 272.7583, 272.8805, 
    272.8986,
  276.7386, 275.7705, 271.7685, 270.9903, 271.657, 271.9482, 272.3183, 
    270.3429, 272.0212, 272.2048, 271.9132, 272.6908, 272.7892, 272.8007, 
    272.797,
  276.9352, 275.022, 272.1631, 271.8477, 272.0211, 271.4298, 271.7767, 
    271.1498, 272.2219, 272.2357, 272.6898, 272.8379, 272.7682, 272.6977, 
    272.5469,
  275.9021, 274.0768, 272.3626, 272.2512, 272.0376, 271.6791, 271.6883, 
    271.3885, 271.2455, 272.1794, 272.9336, 272.8743, 272.7, 272.6037, 
    272.4067,
  281.0798, 273.3346, 276.3502, 272.9138, 272.801, 272.5612, 272.2028, 
    271.9379, 271.4286, 272.0497, 273.3256, 272.4377, 271.928, 272.2927, 
    272.3906,
  273.1426, 272.8526, 272.7195, 272.4477, 272.6991, 272.9136, 272.6664, 
    271.6313, 271.0453, 271.308, 271.2848, 270.766, 271.8136, 271.9052, 
    272.0809,
  274.4266, 274.0204, 273.2068, 272.2733, 272.2191, 271.8762, 272.2286, 
    272.0732, 271.5824, 271.2978, 271.6193, 271.6276, 272.0638, 271.502, 
    272.4303,
  275.0935, 274.4594, 273.5877, 272.9034, 272.1747, 271.8902, 270.1898, 
    271.1822, 271.1901, 271.791, 267.9552, 271.9294, 271.7853, 272.3953, 
    273.0195,
  275.6687, 274.3661, 273.8726, 272.6602, 272.4024, 271.5466, 270.7581, 
    268.4214, 268.3351, 268.1869, 269.4278, 272.371, 272.7121, 272.9846, 
    273.0477,
  275.9384, 274.7592, 273.2486, 272.0719, 272.0392, 271.0492, 270.5219, 
    269.9257, 269.1542, 268.6175, 272.2696, 272.4257, 272.9116, 272.9321, 
    272.9241,
  276.2048, 275.381, 272.8139, 271.8035, 271.5701, 271.2513, 270.9123, 
    270.1803, 269.6833, 270.993, 272.2652, 272.8535, 272.8545, 272.8249, 
    272.8588,
  276.6299, 275.6384, 272.1959, 271.42, 271.2153, 271.0409, 270.7611, 
    269.232, 269.5349, 270.5751, 272.7263, 272.8418, 272.7319, 272.7746, 
    272.772,
  276.7951, 274.8651, 271.994, 271.2895, 271.1425, 270.9088, 270.782, 
    268.4269, 269.6533, 270.3046, 272.7629, 272.7985, 272.7376, 272.7011, 
    272.5926,
  275.9264, 274.1504, 272.3235, 271.3852, 271.145, 271.0929, 271.2024, 
    270.5662, 270.1899, 272.0131, 272.8849, 272.8237, 272.6739, 272.5832, 
    272.3945,
  277.8991, 273.1069, 275.5708, 272.9222, 273.029, 273.0853, 273.0492, 
    272.9716, 272.5315, 272.8619, 273.9372, 272.5132, 271.6312, 271.8383, 
    269.768,
  273.3475, 272.8076, 272.691, 272.666, 272.9539, 273.1514, 273.1287, 
    273.028, 272.705, 272.6463, 272.512, 271.9106, 270.3636, 271.4787, 
    271.9661,
  274.6679, 274.1666, 273.3174, 272.4746, 272.5083, 273.0948, 273.0476, 
    272.9848, 272.6778, 272.1324, 271.8062, 270.8068, 269.6624, 269.6518, 
    272.5835,
  275.2489, 274.5229, 273.6543, 273.1573, 272.5576, 272.524, 271.763, 
    271.9835, 271.9382, 272.0021, 269.8152, 270.0072, 271.525, 272.1935, 
    272.5663,
  275.7661, 274.3861, 273.8619, 273.0683, 272.89, 272.5235, 272.0963, 270.51, 
    268.7574, 270.3612, 271.6615, 271.7431, 271.9834, 272.4135, 272.808,
  275.9515, 274.7054, 273.2581, 272.7395, 272.6709, 272.4151, 271.7825, 
    271.485, 270.5977, 270.3099, 270.5246, 271.7699, 272.6423, 272.8604, 
    272.9357,
  276.1542, 275.2837, 273.1174, 272.3448, 271.6505, 270.4502, 270.3256, 
    270.2154, 270.9191, 271.2927, 272.4911, 272.8016, 272.8086, 272.7843, 
    272.8018,
  276.5249, 275.5829, 272.7491, 271.3941, 270.417, 270.0576, 270.6729, 
    271.176, 271.5983, 272.734, 272.8913, 272.8276, 272.7061, 272.7234, 
    272.7321,
  276.4942, 274.7875, 271.868, 270.6833, 270.6877, 270.7954, 270.8096, 
    271.2916, 272.2262, 272.8326, 272.8411, 272.7813, 272.716, 272.6816, 
    272.6596,
  275.6644, 274.1575, 272.4275, 270.6809, 270.7332, 270.8526, 270.7393, 
    271.8517, 272.593, 272.8926, 272.9146, 272.8212, 272.6488, 272.5425, 
    272.4556,
  277.7828, 273.1527, 275.4878, 272.846, 272.9696, 272.9088, 272.8842, 
    272.9868, 272.811, 272.9741, 274.0854, 273.4173, 272.5867, 273.0333, 
    273.158,
  273.2221, 272.8796, 272.6443, 272.6255, 273.0276, 272.1937, 272.7875, 
    273.002, 272.9466, 272.8177, 273.1302, 272.9083, 272.5749, 272.4183, 
    273.1138,
  274.6933, 274.2636, 273.4304, 272.4031, 272.4019, 271.9291, 271.4, 
    272.5993, 273.0682, 273.0158, 273.0226, 272.9933, 272.4303, 271.9814, 
    272.6761,
  275.3332, 274.6135, 273.7448, 273.1471, 272.4315, 271.8675, 273.1117, 
    273.097, 273.0981, 273.0709, 272.9648, 272.7351, 273.0039, 272.8641, 
    272.1894,
  275.8112, 274.4711, 273.9347, 273.1057, 272.8338, 271.3833, 271.6093, 
    272.9498, 272.4329, 273.0237, 272.906, 272.7675, 272.4881, 272.465, 
    272.4711,
  275.8856, 274.6912, 273.3439, 272.8376, 272.9033, 272.9221, 272.766, 
    272.4359, 272.3342, 272.4524, 272.4857, 272.4353, 272.6545, 272.5673, 
    272.4832,
  276.1193, 275.2519, 273.1787, 272.7205, 272.7289, 272.6387, 272.5887, 
    272.2421, 271.7978, 271.995, 272.4953, 272.6031, 272.4797, 272.3462, 
    272.6329,
  276.4918, 275.5627, 272.73, 272.0061, 272.2573, 272.3907, 272.049, 
    272.0118, 272.2792, 272.3817, 272.5047, 272.2974, 272.5074, 272.5747, 
    272.6729,
  276.4348, 274.8174, 272.3163, 272.1685, 272.4272, 272.5089, 272.2614, 
    272.2186, 272.6398, 272.6988, 272.4167, 272.5615, 272.6916, 272.6754, 
    272.8126,
  275.5827, 274.2703, 272.7865, 272.2589, 272.5127, 272.7721, 272.7359, 
    272.6017, 272.8416, 272.9023, 272.9414, 272.8103, 272.6104, 272.5066, 
    272.6718,
  277.4021, 273.0647, 275.8088, 272.823, 272.7101, 273.3692, 272.6576, 
    272.2553, 271.941, 272.5287, 274.1871, 273.7255, 273.0603, 273.2315, 
    273.0784,
  273.445, 272.9901, 272.9433, 272.4861, 272.9212, 272.9924, 273.0627, 
    272.4652, 271.9956, 272.1986, 273.2295, 273.256, 272.7017, 273.1024, 
    273.1595,
  274.7505, 274.4369, 273.5911, 272.316, 272.7459, 273.1086, 272.9753, 
    272.6111, 272.5028, 272.2973, 272.9789, 272.9726, 272.4888, 272.9411, 
    272.8829,
  275.4625, 274.8104, 273.9588, 273.1245, 272.4501, 272.761, 273.1321, 
    272.915, 272.8983, 273.0021, 273.0584, 272.9344, 272.3086, 273.081, 
    273.0071,
  275.9711, 274.7036, 274.1456, 273.0805, 272.7794, 272.6691, 272.5842, 
    273.0706, 273.1285, 273.1061, 273.0892, 272.7496, 273.0761, 273.0612, 
    272.9442,
  276.0323, 274.873, 273.6024, 272.7302, 272.8456, 272.8945, 272.8206, 
    272.5979, 272.6898, 272.7289, 272.9308, 273.0039, 273.0339, 272.9994, 
    272.9381,
  276.2404, 275.3758, 273.3112, 272.6609, 272.7873, 272.8338, 272.8238, 
    272.8143, 272.7414, 272.725, 272.8071, 272.9216, 272.8449, 272.5976, 
    272.6013,
  276.5096, 275.5707, 273.0471, 272.5883, 272.7658, 272.8007, 272.751, 
    272.7764, 272.8171, 272.8481, 272.822, 272.7342, 272.474, 272.3075, 
    272.4168,
  276.4127, 274.8355, 272.6691, 272.5972, 272.7044, 272.7174, 272.7737, 
    272.7426, 272.8037, 272.8919, 272.7285, 272.6547, 272.4804, 272.5145, 
    272.823,
  275.5783, 274.386, 273.0343, 272.7216, 272.7153, 272.6933, 272.5856, 
    272.5482, 272.8649, 272.9501, 272.9656, 272.6807, 272.4924, 272.4302, 
    273.0064,
  277.2542, 273.2037, 275.2691, 272.7369, 273.0398, 274.2664, 272.9626, 
    272.8249, 272.8492, 272.6248, 273.5771, 273.8486, 273.1631, 273.4089, 
    273.1104,
  273.6978, 273.0707, 273.1883, 272.5714, 273.0929, 273.0623, 272.9841, 
    272.9325, 272.6129, 271.9143, 272.8668, 273.3677, 273.1268, 273.1564, 
    273.1217,
  274.8447, 274.5327, 273.6365, 272.353, 272.7766, 273.1314, 272.8767, 
    272.9215, 272.9863, 271.7072, 272.6241, 273.1066, 273.0761, 273.041, 
    273.0093,
  275.5036, 274.8442, 273.93, 273.0784, 272.4908, 272.7628, 273.1284, 
    272.7821, 272.963, 271.8375, 272.9416, 273.0641, 273.0405, 273.0267, 
    272.937,
  275.9319, 274.6711, 274.09, 272.9492, 272.7429, 272.5886, 272.5948, 
    273.0682, 273.0952, 272.2314, 272.9502, 273.0001, 273.0296, 272.9889, 
    272.9217,
  275.9513, 274.7829, 273.5116, 272.496, 272.7339, 272.8282, 272.7489, 
    272.5316, 272.7245, 272.6127, 272.8316, 272.9506, 272.9952, 272.9198, 
    272.8761,
  276.1307, 275.2816, 273.1681, 272.4247, 272.6209, 272.8189, 272.8529, 
    272.8196, 272.6949, 272.2738, 272.5677, 272.4549, 272.8898, 272.879, 
    272.8387,
  276.4535, 275.4979, 272.8231, 272.5292, 272.6913, 272.8146, 272.7635, 
    272.7711, 272.7271, 272.2181, 272.3928, 272.4781, 272.7491, 272.6274, 
    272.5867,
  276.3761, 274.7826, 272.4377, 272.5608, 272.799, 272.8341, 272.837, 
    272.4727, 272.1699, 272.2858, 272.9111, 272.6713, 272.7205, 272.7143, 
    272.8349,
  275.5514, 274.3994, 272.6319, 272.312, 272.6501, 272.7461, 272.5612, 
    272.3851, 272.3369, 272.5802, 272.4791, 272.8258, 272.6639, 272.5967, 
    272.907,
  277.4802, 273.3079, 274.6265, 272.4947, 273.1168, 273.7265, 272.8964, 
    272.8244, 272.9382, 273.0951, 274.3402, 273.9676, 273.1925, 273.5111, 
    273.1595,
  273.915, 273.1826, 273.1902, 272.4579, 273.1128, 272.938, 272.817, 
    272.8632, 272.7965, 272.9353, 273.5921, 273.2923, 273.1387, 273.157, 
    273.1595,
  274.8413, 274.5139, 273.6596, 272.3453, 272.7713, 273.0143, 272.9969, 
    272.9724, 272.9601, 272.785, 272.7415, 272.6659, 273.0553, 273.0226, 
    273.0585,
  275.4706, 274.8197, 273.9208, 273.1015, 272.5033, 272.7753, 272.9747, 
    272.6016, 272.9257, 272.4629, 272.6159, 272.9087, 273.0262, 272.9855, 
    272.9185,
  275.8342, 274.5969, 274.0807, 272.898, 272.7464, 272.553, 272.5983, 
    272.7128, 273.0953, 272.3319, 272.5447, 272.933, 272.9819, 272.9765, 
    272.9128,
  275.8658, 274.7346, 273.5164, 272.4359, 272.7037, 272.8217, 272.7531, 
    272.541, 272.3674, 272.1202, 272.9011, 272.937, 272.955, 272.9754, 
    272.9793,
  276.0348, 275.2382, 273.103, 272.1606, 272.5728, 272.7998, 272.8558, 
    272.7643, 271.9809, 272.1727, 272.7115, 272.8909, 272.8838, 272.7773, 
    272.6944,
  276.392, 275.4448, 272.6805, 272.3296, 272.6084, 272.7957, 272.7573, 
    272.5606, 272.3255, 272.5717, 272.8432, 272.8212, 272.7564, 272.5768, 
    272.557,
  276.336, 274.7246, 272.5617, 272.7061, 272.795, 272.8309, 272.8216, 
    272.5915, 272.6632, 272.6546, 272.9295, 272.8112, 272.7093, 272.6767, 
    272.8014,
  275.5083, 274.3917, 273.0925, 272.9531, 272.8946, 272.8318, 272.5859, 
    272.4994, 272.6011, 272.9684, 272.9345, 272.8433, 272.6612, 272.6067, 
    272.8925,
  280.3813, 273.7885, 276.4903, 272.5037, 273.3355, 274.5049, 272.9293, 
    272.9308, 273.0469, 273.1404, 274.4956, 274.1579, 273.2041, 273.4029, 
    272.824,
  274.576, 273.6268, 273.5016, 272.4511, 273.3767, 273.5597, 272.8662, 
    272.9422, 272.9235, 273.0238, 273.8923, 273.4922, 273.122, 273.1362, 
    273.1595,
  275.4418, 274.8763, 273.8126, 272.4193, 272.7764, 273.0738, 272.653, 
    272.9181, 272.915, 272.6344, 272.6562, 273.0386, 273.0414, 273.0492, 
    273.0617,
  275.731, 274.9634, 273.9892, 273.2466, 272.4023, 272.819, 273.0736, 
    272.9562, 272.5934, 272.6713, 272.756, 272.8794, 272.8958, 272.7773, 
    272.7809,
  275.872, 274.6136, 274.0875, 272.7894, 272.6944, 272.5857, 272.6722, 
    272.275, 272.5851, 272.8806, 272.5735, 272.8578, 272.9271, 272.7789, 
    272.8436,
  275.8758, 274.7018, 273.519, 272.2215, 272.5929, 272.7717, 272.738, 
    272.6267, 272.8607, 272.7037, 272.845, 272.8747, 272.8314, 272.864, 
    272.8925,
  276.0302, 275.2448, 273.0443, 271.7744, 272.241, 272.6579, 272.7971, 
    272.813, 272.7108, 272.5293, 272.718, 272.8138, 272.805, 272.6768, 
    272.6924,
  276.3979, 275.4312, 272.5934, 271.9436, 272.4569, 272.6853, 272.7233, 
    272.7248, 272.7477, 272.8389, 272.7622, 272.8004, 272.75, 272.5945, 
    272.5528,
  276.3563, 274.6372, 272.5097, 272.6238, 272.7221, 272.809, 272.7938, 
    272.8388, 272.899, 272.9583, 272.9235, 272.8179, 272.7026, 272.6507, 
    272.7908,
  275.5302, 274.3795, 273.0237, 272.9474, 272.9131, 272.8484, 272.6184, 
    272.5673, 272.8413, 272.9647, 272.9297, 272.8608, 272.6626, 272.6367, 
    272.8543,
  280.078, 274.1122, 277.5517, 272.5692, 273.4569, 275.3118, 272.9023, 
    272.9136, 273.1768, 276.2174, 277.0322, 275.7378, 272.7825, 274.5161, 
    273.7459,
  274.7283, 273.9249, 273.8417, 272.6297, 274.7914, 275.6909, 272.8419, 
    272.9003, 272.924, 273.6738, 274.3851, 272.9101, 272.6662, 272.8321, 
    272.9258,
  275.489, 275.0865, 274.0002, 272.6064, 272.8672, 273.1119, 272.5892, 
    272.6012, 272.3997, 272.0231, 271.6277, 271.8057, 272.8223, 273.0052, 
    273.0929,
  275.9742, 275.3848, 274.372, 273.683, 272.3734, 272.9255, 273.1015, 
    272.2021, 271.6153, 271.2524, 271.37, 271.5874, 272.7317, 272.9219, 
    272.8236,
  276.3105, 275.0096, 274.3311, 272.8315, 272.558, 272.313, 272.6356, 
    273.0327, 272.8911, 271.2309, 271.3636, 271.4492, 272.6209, 272.9058, 
    272.2903,
  276.0833, 274.9633, 273.6479, 272.1928, 272.412, 272.6398, 272.435, 
    272.6408, 272.6153, 272.0232, 271.6056, 272.6942, 272.5508, 272.7904, 
    272.5298,
  276.2142, 275.379, 273.0298, 271.8017, 271.9811, 272.6111, 272.7655, 
    272.8099, 272.6896, 271.9633, 272.7072, 272.8153, 272.8314, 272.7111, 
    272.453,
  276.5185, 275.5131, 272.6931, 272.1204, 272.3964, 272.6396, 272.711, 
    272.6646, 272.7788, 272.6955, 272.8071, 272.7976, 272.7253, 272.4609, 
    272.2885,
  276.4568, 274.5331, 272.5327, 272.6771, 272.7172, 272.7653, 272.757, 
    272.8034, 272.9181, 272.9831, 272.9245, 272.737, 272.6461, 272.4698, 
    272.4923,
  275.6086, 274.3764, 272.9533, 272.942, 272.9215, 272.8577, 272.6456, 
    272.6225, 272.9206, 272.9917, 272.881, 272.8165, 272.6483, 272.4889, 
    272.7927,
  277.4829, 274.2249, 277.2755, 272.5737, 273.4837, 275.2364, 272.8642, 
    272.8835, 273.1975, 278.3717, 278.6306, 277.0446, 275.0968, 275.3087, 
    275.1062,
  274.4363, 274.1322, 274.0418, 272.7277, 275.695, 275.7222, 272.8767, 
    272.9234, 272.9286, 274.0445, 276.7812, 273.6413, 272.9386, 273.0575, 
    273.1595,
  275.2946, 275.1934, 274.1448, 272.7014, 273.1462, 273.1445, 272.9479, 
    272.9193, 272.9348, 272.7709, 272.5849, 272.3712, 272.5362, 273.0432, 
    273.1065,
  275.8025, 275.3954, 274.3638, 273.7, 272.2982, 273.0214, 273.1211, 
    272.9458, 272.7035, 272.1809, 272.0075, 272.178, 272.5666, 272.9752, 
    272.9933,
  275.9692, 274.8612, 274.3534, 272.9249, 272.5624, 272.5762, 272.8052, 
    273.1239, 272.6092, 271.9975, 271.8853, 272.1943, 272.646, 272.8148, 
    272.8149,
  276.0424, 274.865, 273.6835, 272.2896, 272.3535, 272.685, 272.6832, 
    272.6293, 272.9033, 272.3338, 272.1591, 272.2976, 272.6448, 272.6128, 
    272.5585,
  276.4406, 275.4367, 273.0027, 271.8257, 271.7776, 272.5694, 272.7685, 
    272.8046, 272.4621, 272.1461, 272.2277, 272.4528, 272.4236, 272.1998, 
    272.0982,
  277.0899, 275.7034, 272.7076, 271.9608, 272.1703, 272.6476, 272.7015, 
    272.6422, 272.2882, 272.5457, 272.2952, 272.2819, 272.2343, 271.9282, 
    271.9103,
  276.8578, 274.6836, 272.54, 272.7134, 272.7159, 272.752, 272.7597, 
    272.7967, 272.8453, 272.8974, 272.5079, 272.3206, 272.1169, 271.9037, 
    272.0006,
  275.7964, 274.4902, 272.9314, 272.9239, 272.9103, 272.877, 272.7079, 
    272.7043, 272.9775, 273.0024, 272.6445, 272.3292, 272.1283, 271.8421, 
    272.5422,
  277.6225, 273.2487, 275.3552, 272.4922, 273.2926, 274.7328, 272.8897, 
    272.8784, 273.0069, 276.1583, 278.1846, 276.8491, 275.6223, 276.1849, 
    277.0156,
  273.8687, 273.6449, 273.9374, 272.7805, 275.0074, 274.9987, 273.0139, 
    272.9732, 272.8813, 273.4633, 276.8913, 274.2543, 273.6129, 273.1988, 
    273.6466,
  274.9979, 274.8626, 274.2088, 272.9085, 273.8365, 273.1766, 273.126, 
    273.0428, 272.9455, 272.8857, 273.2931, 273.0485, 273.0428, 273.2133, 
    273.0964,
  275.8553, 275.3617, 274.499, 273.9244, 272.3151, 273.1908, 272.8431, 
    272.9223, 272.5084, 272.637, 272.7693, 272.8947, 273.0255, 272.9823, 
    272.9578,
  276.0724, 274.8618, 274.5494, 273.2002, 272.5343, 272.4566, 272.8764, 
    272.2452, 270.5597, 272.6326, 272.5893, 272.8023, 272.7462, 272.4646, 
    272.383,
  276.23, 274.8969, 273.938, 272.5838, 272.4249, 272.5988, 272.4619, 
    272.3643, 272.7469, 272.4098, 272.3925, 272.4383, 272.2586, 272.1039, 
    271.8972,
  276.6676, 275.4913, 273.1216, 272.0234, 271.8857, 272.414, 272.5987, 
    272.5974, 272.0535, 271.8073, 272.0949, 272.0159, 271.7938, 270.874, 
    271.6342,
  277.2235, 275.7562, 272.6837, 271.8909, 271.8941, 272.5064, 272.5409, 
    272.3269, 271.9035, 271.9803, 271.6664, 271.6754, 271.5423, 271.6524, 
    271.696,
  277.3566, 274.7302, 272.2124, 272.5416, 272.4949, 272.6788, 272.5762, 
    272.2686, 272.2577, 272.005, 271.8077, 271.7408, 271.6421, 271.6953, 
    271.9101,
  276.3673, 274.6925, 272.8662, 272.9006, 272.9063, 272.8678, 272.418, 
    272.2749, 271.8727, 272.3254, 271.9345, 271.6787, 271.6968, 271.4205, 
    272.4687,
  280.7637, 273.4165, 275.6207, 272.54, 273.3736, 274.9236, 273.0414, 
    272.9306, 273.0971, 278.2652, 279.7242, 277.5707, 277.3481, 277.36, 
    277.0659,
  274.0148, 273.6371, 273.896, 272.9069, 275.7463, 275.1926, 273.0829, 
    273.031, 272.6332, 274.0144, 277.5831, 274.6515, 274.0124, 273.1117, 
    275.2844,
  275.0795, 274.8509, 274.2433, 273.0965, 275.0074, 273.1911, 273.3742, 
    273.081, 272.987, 272.8598, 273.9595, 272.863, 272.4184, 272.413, 272.808,
  275.9083, 275.4234, 274.5255, 274.0474, 272.4626, 273.3979, 273.101, 
    273.0981, 273.0374, 273.0129, 272.984, 272.8787, 272.3008, 272.3242, 
    272.6487,
  276.032, 274.9218, 274.5508, 273.2862, 272.454, 272.405, 273.1075, 
    272.3364, 271.7934, 273.0686, 272.9068, 272.5228, 272.3539, 272.0461, 
    272.4096,
  276.1551, 274.9294, 273.9627, 272.5667, 272.3421, 272.611, 272.5718, 
    272.6204, 272.887, 272.8424, 272.6635, 272.0137, 271.9534, 271.9763, 
    272.3952,
  276.5726, 275.5217, 273.1495, 272.1114, 271.98, 272.2558, 272.6806, 
    272.7221, 272.534, 272.1815, 272.0322, 271.5816, 271.6272, 271.8105, 
    272.3032,
  277.0966, 275.7927, 272.7841, 271.9696, 271.8982, 272.2888, 272.6042, 
    272.4533, 272.2378, 272.0264, 271.7528, 271.3823, 271.8668, 272.2121, 
    272.4376,
  277.2799, 274.7107, 272.3165, 272.2597, 272.3104, 272.5409, 272.4735, 
    272.3768, 272.2022, 271.6862, 271.1803, 271.7073, 272.0432, 272.4477, 
    272.263,
  276.4577, 274.6862, 272.7604, 272.8313, 272.8292, 272.6681, 272.1931, 
    271.9617, 271.6678, 271.5256, 271.6664, 271.7298, 272.2387, 272.5181, 
    272.947,
  277.2579, 273.5791, 275.6911, 272.5902, 273.2861, 274.866, 273.026, 
    272.9546, 273.1756, 279.3677, 280.3901, 277.7664, 277.4262, 277.1878, 
    277.244,
  274.1517, 273.8064, 273.9797, 273.0117, 275.3692, 275.2224, 272.7182, 
    272.9992, 272.9095, 274.2241, 278.43, 275.0877, 274.4089, 273.4264, 
    274.9189,
  275.2119, 275.0014, 274.3602, 273.2314, 274.64, 272.626, 273.2536, 
    272.9676, 272.9767, 272.8985, 274.4887, 273.4854, 273.0199, 273.1108, 
    273.1515,
  276.0671, 275.6948, 274.5885, 274.1452, 272.6302, 273.729, 272.6751, 
    272.9436, 272.5643, 272.99, 272.9874, 273.0251, 273.0041, 272.6747, 
    272.8498,
  276.2652, 275.0289, 274.5155, 273.3224, 272.2988, 272.341, 273.0606, 
    272.3601, 271.9756, 272.9119, 273.0015, 272.9062, 272.7691, 272.4696, 
    272.6606,
  276.2168, 274.9603, 273.8706, 272.5396, 272.1357, 272.5638, 272.5779, 
    272.6417, 272.9628, 272.8474, 272.8703, 272.707, 272.3365, 272.269, 
    272.6104,
  276.5042, 275.4936, 273.0984, 271.9978, 271.9551, 272.0184, 272.7244, 
    272.7377, 272.5179, 272.3599, 272.311, 272.1125, 271.7965, 272.2295, 
    272.473,
  276.886, 275.6464, 272.8051, 271.8991, 271.9523, 272.1191, 272.6383, 
    272.5094, 272.5222, 272.6055, 272.3598, 271.6498, 271.8857, 272.1853, 
    272.3587,
  276.8615, 274.6103, 272.424, 272.2945, 272.111, 272.2624, 272.5952, 
    272.719, 272.8725, 272.6011, 271.7117, 271.433, 271.999, 272.2047, 
    272.6362,
  275.9643, 274.5164, 272.8759, 272.6106, 272.6925, 272.6432, 272.4842, 
    272.516, 272.4908, 271.9386, 271.4854, 271.4188, 272.1585, 272.4953, 
    273.1761,
  280.1588, 274.176, 278.0297, 272.66, 273.0822, 274.1313, 273.0038, 
    272.9218, 273.1395, 277.5391, 280.1473, 278.3629, 279.101, 278.3588, 
    278.2272,
  274.2304, 273.8118, 274.0242, 273.0631, 274.1201, 273.6858, 273.0042, 
    272.9723, 272.8795, 273.926, 278.0524, 275.2498, 274.7857, 275.3572, 
    276.855,
  275.1786, 274.9709, 274.3713, 273.334, 274.729, 272.4655, 272.9485, 
    272.8742, 272.3843, 272.6693, 274.4673, 273.7037, 273.0596, 273.2854, 
    274.4349,
  276.0043, 275.6909, 274.6537, 274.2845, 273.0186, 274.5073, 272.2803, 
    272.6971, 271.9184, 272.7818, 272.8374, 272.9649, 273.0048, 272.9278, 
    272.9681,
  276.3297, 275.2707, 274.7897, 273.634, 272.4017, 272.4799, 273.2065, 
    271.8477, 271.9982, 273.3914, 272.8074, 272.7874, 272.9247, 272.8288, 
    272.8052,
  276.5244, 275.2671, 274.1126, 272.759, 272.0259, 272.3738, 272.5985, 
    272.6744, 273.0042, 272.8654, 272.7668, 272.7313, 272.8709, 272.7706, 
    272.7727,
  276.7728, 275.6684, 273.2332, 272.1085, 272.0391, 271.8868, 272.5393, 
    272.71, 272.5751, 272.3438, 272.4221, 272.694, 272.8102, 272.7458, 
    272.6889,
  277.0497, 275.6906, 272.9044, 272.0113, 272.0739, 271.9632, 272.4449, 
    272.5046, 272.496, 272.7203, 272.7556, 272.6693, 272.7707, 272.4893, 
    272.3226,
  276.938, 274.7628, 272.5117, 272.3428, 272.2399, 272.0495, 272.4564, 
    272.7675, 272.9336, 272.9336, 272.9155, 272.8222, 272.677, 272.1509, 
    272.3725,
  275.9918, 274.5935, 272.9892, 272.688, 272.6925, 272.6831, 272.5568, 
    272.8741, 273.0212, 273.0042, 272.8856, 272.6606, 272.4107, 272.0657, 
    273.0229,
  277.2008, 273.6194, 275.5648, 272.5146, 273.2099, 274.6242, 272.9715, 
    272.8744, 273.0703, 277.9944, 280.4358, 279.2127, 280.8711, 280.2487, 
    279.0269,
  274.2906, 273.8185, 273.9114, 272.9977, 275.0448, 274.8438, 272.986, 
    272.9479, 272.8454, 273.8584, 278.0948, 275.3691, 275.3576, 277.8404, 
    278.0978,
  275.0034, 274.8765, 274.2767, 273.2495, 274.5592, 272.7921, 273.2799, 
    272.9625, 272.9351, 272.8881, 274.5621, 273.8968, 273.0582, 273.4239, 
    275.1157,
  275.8433, 275.4332, 274.3457, 274.0514, 272.8384, 274.2225, 272.52, 
    272.8057, 272.6066, 272.8732, 272.9754, 273.0038, 272.9763, 272.8935, 
    272.9742,
  276.1061, 275.0228, 274.5451, 273.4215, 272.1509, 272.3193, 273.3135, 
    272.2834, 271.6009, 272.9759, 272.8522, 272.9238, 272.9212, 272.8288, 
    272.7289,
  276.4105, 275.1063, 274.0463, 272.7698, 272.0009, 272.1797, 272.4621, 
    272.7685, 273.2967, 272.6258, 272.6081, 272.7214, 272.8164, 272.8163, 
    272.735,
  276.7874, 275.6483, 273.2714, 272.2284, 272.1737, 272.0038, 272.3352, 
    272.5113, 272.3572, 272.1033, 272.2296, 272.3141, 272.4324, 272.658, 
    272.7393,
  277.1458, 275.7407, 273.032, 272.1569, 272.2008, 272.0883, 272.3379, 
    272.493, 272.464, 272.4005, 272.532, 272.7513, 272.7972, 272.7285, 
    272.6832,
  277.0294, 274.8671, 272.6943, 272.2971, 272.33, 272.134, 272.4897, 
    272.7726, 272.8688, 272.9026, 272.8937, 272.8665, 272.7997, 272.668, 
    272.58,
  276.0444, 274.64, 272.9167, 272.6556, 272.6721, 272.6385, 272.5249, 
    272.7017, 272.9188, 272.9828, 272.9156, 272.8096, 272.7026, 272.3766, 
    272.9654,
  275.5519, 273.5087, 274.8569, 272.5398, 273.0481, 274.2663, 272.2022, 
    271.9519, 272.1597, 274.7657, 276.8483, 275.9606, 275.9751, 277.4948, 
    278.8025,
  274.3099, 273.8723, 273.8364, 272.9428, 274.4138, 274.5631, 271.9526, 
    272.0846, 272.086, 272.9352, 275.6558, 275.0893, 274.0619, 274.7299, 
    276.6468,
  275.1906, 275.0038, 274.3994, 273.2411, 274.1623, 272.0884, 272.9337, 
    272.0728, 272.1328, 272.048, 272.9982, 273.5262, 273.0062, 273.2358, 
    274.3709,
  276.2, 275.6939, 274.4896, 274.0186, 272.8241, 274.0147, 271.9152, 
    272.0824, 272.3615, 272.1242, 272.8343, 272.8994, 272.8726, 272.8676, 
    273.1008,
  276.4092, 275.3236, 274.6637, 273.3875, 272.1766, 272.447, 273.3474, 
    271.0501, 270.5595, 273.0949, 272.9267, 272.9099, 272.8578, 272.779, 
    272.6591,
  276.6902, 275.3759, 274.2026, 272.8372, 272.0442, 272.1475, 272.5086, 
    272.826, 273.0505, 272.9058, 272.9455, 272.9361, 272.8938, 272.8056, 
    272.6978,
  276.9845, 275.888, 273.4469, 272.321, 272.2641, 272.1404, 272.1902, 
    272.6076, 272.5228, 272.4341, 272.6521, 272.9124, 272.8381, 272.7802, 
    272.7375,
  277.4921, 276.0341, 273.2512, 272.2963, 272.314, 272.2553, 272.2797, 
    272.5009, 272.6027, 272.8034, 272.914, 272.907, 272.7994, 272.7217, 
    272.7076,
  277.2783, 275.0465, 272.8667, 272.37, 272.3438, 272.0696, 272.5262, 
    272.7784, 272.8352, 272.9438, 272.9833, 272.9164, 272.8221, 272.6936, 
    272.7287,
  276.0869, 274.6623, 272.8804, 272.7026, 272.6719, 272.6699, 272.4599, 
    272.6686, 272.9073, 272.9883, 273.0289, 272.8914, 272.7362, 272.6908, 
    273.0596,
  279.2404, 274.0419, 278.0646, 272.6987, 273.5706, 276.0883, 272.9312, 
    272.874, 273.0444, 277.1561, 279.2295, 276.886, 276.1609, 276.8831, 
    276.5498,
  274.0646, 273.7154, 273.7238, 272.9438, 275.7325, 275.2671, 272.8848, 
    272.7101, 272.7545, 273.7474, 277.3479, 275.5177, 273.8887, 274.8721, 
    275.382,
  274.9185, 274.781, 274.2178, 273.1653, 274.2356, 272.548, 272.9383, 
    272.7499, 272.7897, 272.7618, 273.4618, 273.2718, 272.9733, 273.3051, 
    274.4591,
  275.9454, 275.4562, 274.309, 273.9332, 272.8382, 273.8748, 272.3533, 
    272.4243, 272.825, 272.7999, 272.9508, 272.8489, 272.7742, 272.8948, 
    273.715,
  276.3643, 275.2339, 274.6266, 273.4445, 272.2048, 272.4396, 273.4819, 
    271.9206, 271.487, 273.6219, 272.8186, 272.8787, 272.7879, 272.665, 
    272.5956,
  276.8567, 275.4499, 274.3016, 273.0205, 272.2043, 272.1923, 272.4937, 
    272.9746, 273.6288, 272.9687, 272.7876, 272.8961, 272.8404, 272.2642, 
    272.3685,
  277.2607, 276.0008, 273.5645, 272.5103, 272.4562, 272.3557, 272.1783, 
    272.6097, 272.5198, 272.4233, 272.6297, 272.2721, 271.8097, 271.9138, 
    272.684,
  277.7109, 276.1736, 273.5394, 272.5514, 272.5417, 272.5219, 272.1311, 
    272.4434, 272.6661, 272.7968, 272.4902, 272.3257, 271.6138, 272.6195, 
    272.7007,
  277.4166, 275.1023, 273.1573, 272.4358, 272.3214, 272.1212, 272.4252, 
    272.7014, 272.7926, 272.8782, 272.8218, 272.7372, 272.7314, 272.6955, 
    272.7379,
  276.1703, 274.6893, 272.9687, 272.5559, 272.6228, 272.5614, 272.3929, 
    272.5765, 272.4561, 272.9669, 272.9551, 272.8679, 272.723, 272.697, 
    273.0753,
  276.713, 274.2551, 276.8753, 273.3724, 273.7264, 277.6549, 272.9287, 
    272.903, 273.4205, 284.4755, 285.1221, 280.0549, 280.0976, 278.7163, 
    278.9743,
  274.0962, 273.7991, 273.9782, 273.3164, 277.9975, 279.6996, 272.9338, 
    272.9265, 272.8857, 275.4826, 282.4899, 276.4921, 274.5232, 276.9482, 
    277.8785,
  274.8137, 274.7716, 274.3521, 273.3762, 276.2747, 273.1876, 274.1651, 
    272.9625, 272.9232, 272.8518, 274.0307, 273.8061, 273.0268, 273.3972, 
    275.3516,
  275.8213, 275.3491, 274.2747, 274.0871, 273.0098, 276.102, 273.2011, 
    273.3167, 272.9712, 272.9666, 272.9488, 272.8777, 272.8269, 272.9822, 
    274.1599,
  276.1573, 275.0194, 274.5098, 273.491, 272.4723, 272.5841, 273.5896, 
    273.2717, 273.0194, 274.5382, 272.9557, 272.9127, 272.8313, 272.6992, 
    272.6822,
  276.5231, 275.1678, 274.113, 272.935, 272.2144, 272.3583, 272.5122, 
    272.9865, 274.4525, 273.0147, 273.0248, 272.8941, 272.8812, 272.7246, 
    272.6216,
  277.0439, 275.7812, 273.3415, 272.4027, 272.4099, 272.3149, 272.2412, 
    272.6774, 272.5215, 272.3784, 272.6829, 272.8352, 272.7612, 272.6753, 
    272.6559,
  277.5981, 276.0219, 273.3214, 272.4237, 272.4092, 272.3829, 272.0461, 
    272.4977, 272.5637, 272.7036, 272.7951, 272.7589, 272.5011, 272.5865, 
    272.6597,
  277.4576, 275.0083, 272.9706, 272.0711, 271.9678, 271.909, 272.3496, 
    272.7827, 272.7975, 272.849, 272.7616, 272.7053, 272.6742, 272.6002, 
    272.8133,
  276.2198, 274.5854, 272.6932, 272.1703, 272.244, 272.1089, 272.2468, 
    272.5148, 272.7076, 272.762, 272.7728, 272.7143, 272.5624, 272.5721, 
    273.1899,
  275.4336, 274.0086, 275.9201, 273.4407, 273.7078, 277.4742, 272.9205, 
    272.886, 273.485, 286.714, 288.477, 283.3762, 285.9019, 283.8677, 283.9285,
  274.1101, 273.7782, 273.9411, 273.4574, 277.122, 277.8047, 272.9232, 
    272.9029, 272.9046, 275.9063, 286.0387, 278.509, 276.0206, 283.7354, 
    282.7821,
  274.8278, 274.7649, 274.3235, 273.4651, 275.2802, 273.1886, 273.7702, 
    272.9283, 272.9143, 272.896, 274.7279, 274.8071, 273.0949, 273.8529, 
    277.8012,
  275.8635, 275.3487, 274.2906, 274.0842, 273.1297, 275.2067, 273.2307, 
    273.863, 272.9311, 272.9163, 272.9113, 272.8837, 272.8893, 273.3019, 
    275.2271,
  276.2364, 275.0278, 274.5235, 273.5851, 272.4673, 272.6155, 273.944, 
    273.3405, 273.0652, 275.8068, 273.0161, 272.8571, 272.8399, 272.767, 
    272.686,
  276.5691, 275.168, 274.1138, 273.0028, 272.3221, 272.299, 272.4404, 
    273.0557, 274.6088, 273.1491, 274.4776, 272.8594, 272.8739, 272.759, 
    272.6557,
  277.0863, 275.7628, 273.3215, 272.4481, 272.4893, 272.423, 272.2064, 
    272.5344, 272.4557, 272.3837, 272.6209, 272.8509, 272.8457, 272.7838, 
    272.7194,
  277.6838, 275.9642, 273.2478, 272.4821, 272.4613, 272.4755, 272.071, 
    272.4158, 272.5591, 272.7409, 272.8023, 272.857, 272.8217, 272.749, 
    272.7677,
  277.6046, 275.0263, 272.9072, 272.4016, 272.2497, 271.9834, 272.3502, 
    272.6757, 272.8276, 272.9626, 272.9636, 272.8976, 272.8353, 272.7233, 
    272.8134,
  276.3275, 274.6617, 272.9213, 272.6278, 272.634, 272.2666, 272.3486, 
    272.5835, 272.8025, 272.982, 273.0547, 272.8732, 272.7328, 272.6702, 
    273.1586,
  274.4872, 273.7008, 276.5768, 273.5479, 274.0886, 277.2379, 272.9171, 
    272.8792, 273.5482, 287.1035, 289.3036, 284.4927, 288.3771, 287.4292, 
    289.3368,
  273.9216, 273.5502, 273.7532, 273.4533, 279.35, 278.4798, 272.9619, 
    272.8958, 272.8965, 276.3719, 287.339, 279.4685, 277.2531, 288.0512, 
    288.3449,
  274.7598, 274.6783, 274.2009, 273.4413, 276.0672, 273.1891, 273.7706, 
    272.9713, 272.9027, 272.8897, 275.5143, 275.9037, 273.1689, 274.0156, 
    280.7956,
  275.8483, 275.3091, 274.2424, 273.9987, 273.0961, 275.8153, 273.2364, 
    273.9287, 272.9728, 272.887, 272.8834, 272.8724, 272.8864, 273.341, 
    276.5064,
  276.3148, 275.077, 274.5182, 273.5983, 272.4299, 272.5747, 274.3952, 
    273.3811, 273.0739, 274.2151, 272.9402, 272.8436, 272.8246, 272.7687, 
    272.7121,
  276.8001, 275.2876, 274.1645, 273.0504, 272.332, 272.1989, 272.3242, 
    273.1702, 274.1125, 273.738, 274.1162, 272.8431, 272.8441, 272.7446, 
    272.6759,
  277.4709, 276.1354, 273.5971, 272.5922, 272.5344, 272.4718, 272.1312, 
    272.4144, 272.4233, 272.4701, 272.6684, 272.8439, 272.7732, 272.7545, 
    272.6941,
  277.9716, 276.3522, 273.7386, 272.8255, 272.5804, 272.5979, 272.0271, 
    272.3206, 272.4377, 272.6518, 272.8136, 272.8629, 272.7189, 272.6264, 
    272.7491,
  277.7479, 275.3229, 273.2059, 272.4334, 272.2861, 272.2143, 272.0943, 
    272.437, 272.6074, 272.6844, 272.7503, 272.5656, 272.6796, 272.6611, 
    272.6984,
  276.4928, 274.7937, 273.0494, 272.7394, 272.7116, 272.1305, 272.2337, 
    272.3926, 272.5624, 272.682, 272.784, 272.6776, 272.574, 272.4937, 
    273.0894,
  274.9123, 273.8353, 276.6247, 273.9548, 274.7001, 276.8957, 272.8669, 
    272.8712, 273.5131, 286.9084, 289.1698, 284.4406, 288.1957, 287.6051, 
    290.554,
  273.5962, 273.4921, 273.8503, 273.8041, 281.0034, 279.2492, 272.9693, 
    272.9469, 272.9153, 276.3768, 287.6616, 280.4707, 279.068, 288.4808, 
    290.2241,
  274.4449, 274.5237, 274.3229, 273.8281, 278.7845, 273.2062, 273.9697, 
    273.0061, 272.9619, 272.9712, 276.6014, 277.6299, 273.625, 274.096, 
    281.9715,
  275.6748, 275.1413, 274.2346, 274.39, 273.6494, 277.5532, 273.2656, 
    274.7911, 272.9958, 272.9309, 272.8997, 272.9347, 272.9439, 273.4577, 
    277.1407,
  276.1445, 274.9131, 274.3941, 273.662, 272.8549, 272.8338, 275.2036, 
    273.4712, 273.0829, 275.8973, 273.1108, 272.8493, 272.8509, 272.8152, 
    272.7469,
  276.56, 275.1211, 274.0614, 272.8746, 272.4323, 272.4987, 272.4169, 
    273.5133, 276.3528, 275.2004, 275.3004, 272.8325, 272.8399, 272.7469, 
    272.6756,
  277.3025, 275.8415, 273.358, 272.4226, 272.4703, 272.5673, 272.3743, 
    272.6333, 272.5634, 272.5389, 272.6918, 272.8391, 272.8391, 272.7629, 
    272.6832,
  277.9917, 276.2326, 273.5077, 272.5996, 272.4897, 272.5493, 272.1166, 
    272.4925, 272.6417, 272.764, 272.845, 272.8794, 272.8367, 272.7551, 
    272.7593,
  277.8316, 275.4879, 273.3513, 272.1338, 271.8802, 272.1019, 272.1255, 
    272.5931, 272.7188, 272.7941, 272.8463, 272.8707, 272.815, 272.7453, 
    272.7913,
  276.8305, 275.2286, 273.1208, 272.5558, 272.309, 271.6907, 271.9033, 
    272.3005, 272.4935, 272.6437, 272.8499, 272.778, 272.7229, 272.6348, 
    273.1577,
  274.3991, 273.7768, 275.8335, 274.1709, 274.4199, 275.5328, 272.7982, 
    272.8318, 273.3348, 287.2235, 288.8983, 284.0172, 287.0425, 286.7821, 
    288.6121,
  273.5799, 273.5104, 274.0629, 273.9556, 277.3849, 276.917, 272.9313, 
    272.8776, 272.7687, 276.3467, 287.5812, 281.3407, 280.5276, 287.6961, 
    289.042,
  274.3416, 274.5337, 274.6311, 273.9371, 276.5168, 272.6873, 274.0765, 
    272.9547, 272.9081, 272.9893, 277.2021, 279.2519, 274.9246, 274.0301, 
    281.8031,
  275.6074, 275.1267, 274.4807, 274.5526, 273.9037, 277.2749, 273.2969, 
    274.8865, 272.9611, 272.947, 272.9581, 273.1028, 272.9915, 273.5235, 
    277.2545,
  275.938, 274.7928, 274.3931, 274.1989, 273.1308, 273.0826, 275.8336, 
    273.562, 273.07, 276.0146, 273.1772, 272.8651, 272.8633, 272.8662, 272.802,
  276.3593, 274.9771, 274.0098, 272.955, 272.8395, 272.6412, 272.3556, 
    273.679, 277.0745, 276.105, 275.9076, 272.8138, 272.8429, 272.7956, 
    272.7515,
  277.0752, 275.6185, 273.2352, 272.3586, 272.6649, 272.8029, 272.5037, 
    272.5993, 272.6222, 272.619, 272.6835, 272.8008, 272.8381, 272.7822, 
    272.7308,
  277.7996, 275.9915, 273.3013, 272.4975, 272.5095, 272.8096, 272.2019, 
    272.4072, 272.608, 272.7269, 272.8372, 272.867, 272.8382, 272.7746, 
    272.7998,
  277.741, 275.3373, 273.1165, 272.2536, 271.9516, 272.1458, 272.3232, 
    272.7287, 272.8538, 272.9349, 272.9268, 272.8896, 272.8533, 272.7888, 
    272.9945,
  277.0654, 275.3706, 272.8911, 272.5435, 272.3156, 271.8303, 272.43, 
    272.6624, 272.883, 272.9532, 273.0774, 272.8616, 272.8145, 272.6957, 
    273.2587,
  276.562, 273.8059, 275.2944, 274.1802, 274.0682, 274.4641, 272.7345, 
    272.5078, 272.6722, 281.1562, 287.4497, 283.3395, 284.8742, 285.1127, 
    286.2331,
  273.6652, 273.5172, 274.0293, 274.0123, 275.7304, 275.3548, 272.8163, 
    272.5058, 272.2378, 274.9931, 285.9301, 281.7635, 281.1473, 285.4304, 
    286.7089,
  274.3621, 274.579, 274.6064, 273.9422, 275.5488, 272.8352, 273.8551, 
    272.446, 272.4323, 272.9071, 278.0688, 281.0569, 276.6753, 274.0086, 
    281.0578,
  275.6834, 275.1562, 274.4814, 274.4941, 273.9296, 276.8839, 273.2584, 
    273.8144, 272.541, 272.9075, 272.9967, 273.5543, 273.1227, 273.5124, 
    277.5645,
  275.9427, 274.7999, 274.4421, 274.3439, 273.1577, 273.6251, 276.0678, 
    273.3111, 272.8832, 275.523, 273.1017, 272.7018, 272.8044, 272.8196, 
    272.8649,
  276.3964, 274.9258, 274.022, 273.1808, 273.0231, 273.0077, 272.6931, 
    273.8361, 276.5591, 276.1674, 275.7715, 272.7739, 272.7744, 272.7823, 
    272.7466,
  277.0909, 275.5655, 273.2268, 272.5002, 273.0553, 273.0962, 272.6544, 
    272.4533, 272.5923, 272.7084, 272.7503, 272.7918, 272.8404, 272.8014, 
    272.718,
  277.8438, 275.9167, 273.2798, 272.5245, 272.7034, 273.2038, 272.3452, 
    272.2225, 272.6071, 272.7433, 272.8144, 272.868, 272.8479, 272.7925, 
    272.7405,
  277.8217, 275.402, 273.0925, 272.3175, 272.0656, 272.3594, 272.122, 
    272.7169, 272.9001, 272.9893, 272.9188, 272.8921, 272.8693, 272.8172, 
    273.1926,
  277.3241, 275.6424, 273.108, 272.4545, 272.2977, 271.9115, 272.35, 
    272.6562, 272.9221, 272.9505, 273.1641, 272.8458, 272.8394, 272.6763, 
    273.3712,
  280.3509, 274.7863, 276.7858, 274.2893, 274.1751, 274.2298, 272.8154, 
    272.7716, 272.4754, 277.3114, 281.3319, 282.1646, 284.9293, 285.2046, 
    286.56,
  274.4344, 274.0073, 274.2206, 274.1497, 275.9526, 275.0471, 272.8193, 
    272.7537, 272.2081, 274.2938, 281.0982, 281.7822, 281.5359, 284.6557, 
    286.2341,
  274.9033, 274.8331, 274.6248, 274.06, 275.7155, 273.2813, 273.2283, 
    272.7093, 272.4532, 272.9913, 278.4995, 282.1751, 278.1616, 274.1779, 
    280.1685,
  276.0673, 275.3984, 274.4917, 274.4869, 273.9612, 275.882, 272.5621, 
    274.0278, 272.636, 272.8484, 273.0787, 274.1045, 273.2404, 273.4779, 
    276.8181,
  276.209, 275.06, 274.5861, 274.0182, 273.1576, 273.4848, 275.3623, 
    272.0544, 272.2197, 274.7399, 272.9285, 272.7253, 272.936, 273.045, 
    273.205,
  276.7558, 275.1859, 274.0948, 273.0568, 272.8207, 272.9069, 272.7737, 
    273.7493, 275.0993, 275.7279, 275.0151, 272.5721, 272.5044, 272.5775, 
    272.7536,
  277.3658, 275.6243, 273.2826, 272.5414, 272.8743, 273.026, 272.7472, 
    272.3562, 272.5527, 272.7516, 272.7672, 272.7571, 272.7541, 272.5817, 
    272.5999,
  277.9421, 275.9112, 273.3897, 272.5903, 272.7074, 273.0926, 272.4706, 
    272.209, 272.5201, 272.6702, 272.7561, 272.7911, 272.7448, 272.5406, 
    272.5404,
  277.8169, 275.3797, 273.1129, 272.449, 272.1786, 272.4112, 272.0942, 
    272.6148, 272.8292, 272.8824, 272.8437, 272.7129, 272.5513, 272.4868, 
    272.9633,
  277.203, 275.5735, 273.2179, 272.4599, 272.3949, 272.0152, 272.2073, 
    272.6062, 272.7424, 273.2038, 273.3915, 272.8418, 272.7375, 272.6261, 
    273.4028,
  280.1353, 275.5596, 276.705, 274.669, 274.5348, 273.888, 272.7908, 
    272.8291, 272.9425, 276.8592, 283.168, 283.7115, 286.0356, 286.7682, 
    288.5278,
  275.1132, 274.5292, 275.0169, 274.7505, 276.7535, 275.2752, 272.6274, 
    272.6729, 272.6813, 274.2413, 281.8799, 282.684, 282.2057, 286.7719, 
    288.3548,
  275.2123, 275.1449, 275.3382, 274.759, 276.4623, 273.4781, 273.3521, 
    272.7664, 272.6681, 273.1387, 278.9989, 282.9974, 279.8004, 274.6159, 
    281.0601,
  276.379, 275.6985, 275.0108, 275.1159, 274.5121, 276.5053, 272.7799, 
    273.1957, 272.4135, 272.695, 273.2486, 274.6281, 273.6019, 273.5182, 
    277.2579,
  277.0546, 275.794, 274.9972, 274.3296, 273.4782, 273.7502, 275.4073, 
    272.4896, 271.6346, 273.5755, 272.7585, 272.7357, 273.1579, 273.2191, 
    273.5775,
  277.32, 275.5976, 274.3015, 273.1942, 272.8633, 273.0026, 272.8978, 
    273.7005, 274.6403, 275.2319, 274.306, 272.4744, 272.5725, 272.7379, 
    273.1717,
  277.5314, 275.774, 273.3979, 272.6403, 272.8416, 272.9391, 272.7876, 
    272.2816, 272.5137, 272.7717, 272.7503, 272.4395, 272.4059, 272.5484, 
    272.8509,
  278.0081, 275.9812, 273.5492, 272.6905, 272.7233, 272.9761, 272.5092, 
    272.2305, 272.427, 272.7809, 272.7785, 272.6192, 272.3871, 272.4876, 
    272.7119,
  277.7564, 275.4305, 273.2191, 272.5547, 272.3039, 272.4094, 272.1254, 
    272.4276, 272.8303, 272.7944, 272.7854, 272.539, 272.2715, 272.4447, 
    272.9523,
  276.9515, 275.3599, 273.2441, 272.7621, 272.6375, 272.0728, 272.1749, 
    272.6872, 272.9205, 273.5417, 273.409, 272.6834, 272.1416, 272.4984, 
    273.3936 ;

}
