netcdf atmos.1980-1981.aliq.02 {
dimensions:
	time = UNLIMITED ; // (1 currently)
	pfull = 65 ;
	lat = 18 ;
	lon = 29 ;
	bnds = 2 ;
variables:
	float aliq(time, pfull, lat, lon) ;
		aliq:long_name = "Cloud fraction for large-scale liquid clouds" ;
		aliq:units = "dimensionless" ;
		aliq:_FillValue = -999.f ;
		aliq:missing_value = -999.f ;
		aliq:interp_method = "conserve_order2" ;
		aliq:cell_methods = "time: mean within months time: mean over years" ;
		aliq:time_avg_info = "average_T1,average_T2,average_DT" ;
	double average_DT(time) ;
		average_DT:long_name = "Length of average period" ;
		average_DT:units = "days" ;
	double average_T1(time) ;
		average_T1:long_name = "Start time for average period" ;
		average_T1:units = "days since 1979-01-01 00:00:00" ;
	double average_T2(time) ;
		average_T2:long_name = "End time for average period" ;
		average_T2:units = "days since 1979-01-01 00:00:00" ;
	double climatology_bounds(time, bnds) ;
	double lat(lat) ;
		lat:standard_name = "latitude" ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_N" ;
		lat:axis = "Y" ;
		lat:bounds = "lat_bnds" ;
	double lat_bnds(lat, bnds) ;
	double lon(lon) ;
		lon:standard_name = "longitude" ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_E" ;
		lon:axis = "X" ;
		lon:bounds = "lon_bnds" ;
	double lon_bnds(lon, bnds) ;
	double pfull(pfull) ;
		pfull:standard_name = "air_pressure" ;
		pfull:long_name = "ref full pressure level" ;
		pfull:units = "mb" ;
		pfull:positive = "down" ;
		pfull:axis = "Z" ;
	double time(time) ;
		time:standard_name = "time" ;
		time:long_name = "time" ;
		time:climatology = "climatology_bounds" ;
		time:units = "days since 1979-01-01 00:00:00" ;
		time:calendar = "standard" ;
		time:axis = "T" ;

// global attributes:
		:CDI = "Climate Data Interface version 2.4.4 (https://mpimet.mpg.de/cdi)" ;
		:Conventions = "CF-1.6" ;
		:title = "c96L65_am5f9d8r0_amip" ;
		:associated_files = "area: 19800101.grid_spec.nc" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
		:code_release_version = "2024.05" ;
		:git_hash = "5d306c05d9fe755cab04eedc8fd3de0d3c8355a0" ;
		:creationtime = "Mon Aug 25 14:09:46 2025" ;
		:hostname = "pp050" ;
		:history = "Mon Aug 25 13:32:16 2025: ncks -d lat,,,10 -d lon,,,10 atmos.1980-1981.aliq.02.nc reduced/atmos.1980-1981.aliq.02.nc\n",
			"Mon Aug 25 14:40:31 2025: cdo -O -s -select,month=2 merged_output.nc monthly_nc_files/all_years.2.nc\n",
			"Mon Aug 25 14:40:11 2025: cdo -O -s -mergetime /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/shards/ts/regrid-xy/180_288.conserve_order2/atmos_month/P1M/P1Y/atmos_month.198001-198012.aliq.nc /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/shards/ts/regrid-xy/180_288.conserve_order2/atmos_month/P1M/P1Y/atmos_month.198101-198112.aliq.nc merged_output.nc\n",
			"Mon Aug 25 14:12:17 2025: cdo --history splitname 19800101.atmos_month.nc /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/cycle/19800101T0000Z/split/regrid-xy/180_288.conserve_order2/19800101.atmos_month.\n",
			"fregrid --debug --standard_dimension --input_mosaic C96_mosaic.nc --input_dir /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/cycle/19800101T0000Z/history/native --input_file 19800101.atmos_month --associated_file_dir /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/cycle/19800101T0000Z/history/native --interp_method conserve_order2 --remap_file fregrid_remap_file_288_by_180.nc --nlon 288 --nlat 180 --scalar_field (**please see the field list in this file**) --output_file 19800101.atmos_month.nc" ;
		:CDO = "Climate Data Operators version 2.4.4 (https://mpimet.mpg.de/cdo)" ;
		:comment = "FMS time averaging, version 3.0, precision=double" ;
		:NCO = "netCDF Operators version 5.2.4 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco, Citation = 10.1016/j.envsoft.2008.03.004)" ;
data:

 aliq =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2.705909e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, -1.636048e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.082363e-05, 0, 0.0001027796, 0, 
    9.432776e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, -1.129048e-05, 0, 0, -6.526495e-07, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, -2.705956e-05, 0, 6.186365e-05, 0, -1.498187e-05, 0, 
    -1.064838e-05, 0, 0, 0.0005347569, 0, 0.0003598959, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, -1.677897e-06, 0, 0, 0, 0, 0, 0, 0, -1.894136e-05, 0, 0.0001541694, 
    0, 0.001523186, 0, 0, 0, 0, 0, 0, 0, 0, -3.441667e-06, -1.049463e-05, 
    -1.517001e-05, 0, 0, 0,
  0, 0, 0, 0, 1.309506e-05, 0, 0, 0, 0, -1.680732e-05, 0, 0, -1.880535e-06, 
    0, 0.0006288755, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 1.197376e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, -1.293972e-06, 0, 0, 0,
  0, -1.102099e-05, 3.92292e-06, -6.981099e-05, -3.247878e-05, 0.0001201991, 
    0, 0.001670542, 0, 0.0001530518, 0, -1.873185e-06, 0.000582825, 
    -1.10033e-05, 0.001123685, -7.836831e-06, 0, 0, 0, 0, 0, 0, 0, 0, 
    -4.302812e-05, 0, 0, 0, 0,
  0, 0, -9.149824e-06, 4.725949e-05, -3.570134e-05, 0.000116194, 0, 
    -2.963798e-06, -1.342722e-05, 0, -5.889923e-05, -4.747063e-06, 
    0.000191167, 0, 0.002872409, 0.0002521506, -2.603141e-06, 0, 0, 0, 0, 0, 
    0, 0.0001136147, 0.000286874, -2.90469e-05, 0, 0, 0,
  0, 0, 0, 0, 4.456661e-05, -1.518631e-08, 0, 0, 0, -1.645862e-05, 0, 0, 
    -3.172819e-05, 1.790702e-06, 0.0006174279, 0, 0, 0, 0, 0, 0, 0, 0, 
    -2.265013e-05, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.160752e-05, 0, -4.853643e-06, 0, 0, 0, 0, 
    0, 0.0001033507, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, -9.995935e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0.001183903, 0, 0, 0, 0, 0, 0, -1.632491e-08, 0, -6.599125e-06, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -7.638067e-05, 0, 0, 0,
  0, -1.854171e-05, 2.511038e-05, -8.258962e-05, 0.00036525, 0.0004910757, 0, 
    0.003818728, 0, 0.002123557, 0.0004692226, -2.374704e-05, 0.0009933349, 
    -9.953436e-06, 0.001495595, -9.526268e-05, -6.433327e-05, 0, 0, 0, 0, 0, 
    0, 0, 0.0006558292, 5.810031e-06, 0, 0, 0,
  0, -8.654471e-06, 2.017483e-05, 0.0004098256, -0.0001093507, 0.0001944116, 
    -1.105903e-05, 0.0005502718, -5.90079e-05, -8.829699e-06, -0.0001676939, 
    -1.186766e-05, 0.0007004185, 0, 0.004755169, 0.002936505, -4.882317e-05, 
    -7.568797e-07, 0, 0, 0, 0, 0, 0.0001182349, 0.0009756388, -5.106795e-05, 
    0, 0, 0,
  0, 0, 0, 0, -4.773157e-05, -1.978007e-05, 0, 0.0009699623, 9.111633e-05, 
    5.135531e-05, 0, 0, -3.859495e-07, 0.0001627064, 0.00151093, 
    3.875428e-05, 0, -1.804619e-06, 0, 0, 0, 0, 0, -2.683012e-05, 
    0.0001131635, 0.0001605014, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0004089732, -1.063486e-05, -2.743204e-05, 
    0, 0, 0, 0, 0, 0.0002812898, -3.300919e-05, -1.695767e-05, 0, 0, 0, 0, 0, 
    0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, -4.386038e-06, 0, 0.0003560348, 0, 0, 0, 0, 0, 0, 0, 0, 
    -3.728792e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.765572e-07, 0, 0, 0,
  0, 0, 0, 0, 0.003313332, 0, 0, 0, 0, -2.250412e-05, 0, -3.264982e-08, 0, 
    -1.131894e-05, 0, 0, 5.672832e-05, 0.0002499004, 0.001647102, 
    1.110263e-05, 0, 0, 0, 0, 0, -0.0001737316, -1.750577e-06, 0, 0,
  0, -4.259391e-05, 0.0005254413, 0.0007097205, 0.0009874818, 0.001814467, 
    4.743721e-05, 0.006930246, 0, 0.00430678, 0.001108971, -8.080097e-05, 
    0.002240418, 0.001681189, 0.00133339, -3.446401e-05, 0.0006316685, 
    -4.781069e-06, 0, 0, 0, 0, 0, 0, 0.00402753, 0.0006612433, 0, 0, 0,
  0, 0.0002844951, 0.001447767, 0.001450405, -5.717047e-05, 0.0005771066, 
    -1.935329e-05, 0.00183998, 0.0002327679, 0.0001200012, -0.0002724431, 
    -1.841114e-05, 0.00151042, -0.0001220252, 0.01011875, 0.00384849, 
    -0.0001154128, -1.844258e-05, 0, 0, 0, 0, 0, 0.002541261, 0.001591894, 
    -7.581906e-05, 0, 0, 0,
  0, 0, 0, 0, 0.00244546, -8.251626e-05, -3.8589e-05, 0.00174159, 
    0.0002799148, 0.0006876867, 0, 0, -7.248078e-05, 0.002317995, 
    0.002504987, 4.599304e-05, 0, -1.198909e-05, 0, 0, 0, 0, -1.517708e-07, 
    -3.071973e-05, 0.0001996502, 0.00120284, 0, 0, 0,
  0, 0, 0, 0, -9.090092e-06, 0, 0, 0, 0, 0, 0.002536424, -0.0001324017, 
    0.001123083, 0, 0, 0, -4.619402e-05, 0, 0.0006766719, 0.0004698619, 
    0.000125334, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -8.066397e-11, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, -1.454683e-05, -1.381711e-07, 0.001927259, 0, 0, 0, 0, 
    -9.167945e-06, 0, 0.0001916876, -8.053074e-07, 0.0004802263, 
    -4.899885e-07, 0, 0, 0, 0, 0, 0, 0, 0, 0, -3.827235e-05, -1.35963e-05, 0, 0,
  0, 0, 6.567569e-05, 0, 0.01108415, 0, 0, 0, 0, 0.0001541688, 0, 
    -4.095707e-06, 0, 0.0002272877, 0.001460197, 0, 0.001423076, 
    0.0007482043, 0.006748875, 5.687541e-05, 0, 0, 0, 0, 0, 0.001448818, 
    -1.653045e-05, 0, 0,
  0, -8.183555e-05, 0.001273584, 0.001779506, 0.003782863, 0.002549092, 
    0.000185403, 0.01443958, 0, 0.005937382, 0.004794294, 0.0003883007, 
    0.006297796, 0.005350218, 0.001378563, 0.0009773615, 0.006684646, 
    0.0005063714, 0, -2.15919e-05, 0, 0, 0, 0, 0.006438565, 0.001066474, 0, 
    0, 0,
  0, 0.001150743, 0.005132967, 0.002900098, 0.0004552691, 0.001056722, 
    -6.163715e-07, 0.002593569, 0.001877473, 0.000396631, 0.001196962, 
    0.0001130246, 0.002688008, 0.000175615, 0.0221433, 0.01054386, 
    0.0002228685, -2.999693e-05, 0, 0, 0, 0, 0, 0.003040853, 0.004670689, 
    0.0003778407, 0, 0, 0,
  0, 0, 0, 0, 0.00934066, 0.001074941, 5.216005e-05, 0.003867687, 
    0.001189858, 0.004521663, 0, -3.56682e-06, -7.935265e-05, 0.003596581, 
    0.002807218, 2.104769e-05, 0, 3.147393e-05, -2.572463e-05, -4.75816e-08, 
    0, 0, 1.005744e-05, 1.025354e-05, 0.0002280292, 0.003326153, 0, 0, 0,
  0, 0, 0, 0, -2.181622e-05, 0, 0, -2.215277e-05, 0, -4.747469e-05, 
    0.005348408, -0.0001493671, 0.003947961, -1.021907e-06, -2.979101e-06, 
    0.0003697855, 0.0001301345, 0, 0.002297394, 0.001407882, 0.001345285, 
    -1.748795e-05, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -7.624874e-05, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, -1.866741e-05, -6.174399e-05, 0, 0, 0, 0, 9.361939e-05, 
    0, 0, -7.913734e-08, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, -1.196286e-07, -5.087911e-05, 1.367109e-05, 0.00526863, 0.000311126, 
    0.0004216798, 0, 0, 0.0003157893, -4.556763e-06, 0.001267009, 
    0.0005042986, 0.001725283, 0.0004393672, 4.747791e-06, -1.295494e-06, 
    0.0006776595, -1.255519e-05, 0, 0, 0, 0, 0.0008123562, 0.002229001, 
    5.542921e-06, 0, 0,
  0, 0, 0.0002616344, 0, 0.02614962, -2.369461e-05, 0, 0, 0, 0.0003234054, 0, 
    -5.361823e-05, 0, 0.001887789, 0.003239927, 0, 0.003714009, 0.001470764, 
    0.009721591, 0.0005916963, 0, 0, 0, 0, 3.25471e-05, 0.006362978, 
    0.001122944, 0, 1.586761e-05,
  0, 7.663354e-05, 0.00283963, 0.005681586, 0.01363703, 0.007270776, 
    0.0003530587, 0.02301329, 0, 0.009702591, 0.01291554, 0.001724618, 
    0.0178382, 0.008897105, 0.005217201, 0.004874431, 0.01202608, 
    0.001620758, 0, 0.000554172, 0, 0, 0, -3.405537e-06, 0.01051552, 
    0.002533561, -8.17684e-06, 0, 0,
  0, 0.002347997, 0.01149672, 0.005675265, 0.002773747, 0.003604772, 
    8.260838e-05, 0.003771455, 0.004341213, 0.001710105, 0.005102734, 
    0.0007181698, 0.004316008, 0.001407549, 0.04186069, 0.02224054, 
    0.0003745195, -4.732201e-05, 0, 0, 0, 0, 0, 0.006142808, 0.01008463, 
    0.001022804, 0, 0, 0,
  0, 0, 0, 0, 0.01471123, 0.00679068, 0.002224806, 0.005187211, 0.004643987, 
    0.007872741, -7.004833e-06, 5.441577e-05, 0.0006347364, 0.006368103, 
    0.006189456, 0.001885397, 0, 0.0001057691, -9.628052e-05, -5.517563e-06, 
    0, 0, 3.158277e-05, 0.0001027484, 0.0007609393, 0.007845938, 
    -3.666943e-06, 0, 0,
  0, 0, 0, 0, -3.500576e-05, -3.002231e-06, 0, -9.113194e-05, 0, 
    -8.302325e-05, 0.009084283, 0.00130428, 0.006429766, 0.0003264702, 
    -2.537414e-05, 0.0006000366, 0.00315406, 6.204315e-05, 0.00689445, 
    0.001978534, 0.002062348, -0.0001139289, 0, 0, -1.637161e-07, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -9.670705e-06, 0, 0, 0, 0, 0, 
    -0.0001512158, 0, -2.396255e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, -3.169697e-06, 0, 0, 0, 0, 0, 0, 0, 3.35193e-05, 
    0, 0, 0, 0, 0, 0, 0, -5.988689e-06, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -7.465825e-06, 0, -9.873747e-06, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.956328e-05, 0, 0, 0, 0, 0, 0, 0, 0, -4.275659e-06, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0002345358,
  0, 0, 0, -6.837091e-06, 6.32399e-05, 9.025554e-06, 0.001444159, 
    0.002138574, -1.125628e-05, 0, 0, -2.889463e-06, 0.004753133, 
    -5.037096e-07, -1.54073e-05, 0.0007652466, 0.0002823537, 0, 0, 0, 
    0.0002810462, -5.974045e-06, 0.0006160247, 2.18758e-06, 0, 0.0003447288, 
    0.000570249, 0, -3.397776e-07,
  -1.531816e-05, 0, -2.874568e-06, -0.0001138364, 0.002818848, 0.01343547, 
    0.00269496, 0.0007736267, 0, 0, 0.001810758, 0.00183372, 0.00440787, 
    0.003121911, 0.008983792, 0.004961793, 0.001977066, -5.946582e-05, 
    0.006140395, 0.0009095364, -2.398942e-05, 0, 0, 0, 0.002814076, 
    0.01091608, -0.0002108495, 0.00079232, 0.0001013303,
  0, 0, 0.0009164582, -1.519895e-05, 0.04908048, 0.003996089, 0.0037571, 0, 
    0, 0.0006820772, -3.371215e-05, 0.0004353643, 0, 0.008234042, 
    0.007795211, 1.470196e-06, 0.007356673, 0.005322646, 0.01416126, 
    0.001599633, 0, 0, 0, 0, 0.0002231294, 0.02431218, 0.003440203, 
    0.0005574827, 0.0004125204,
  0, -9.860931e-06, 0.005341482, 0.01101913, 0.0415241, 0.01716684, 
    0.0005854961, 0.03401166, 0, 0.01530186, 0.01833644, 0.004840669, 
    0.02998803, 0.0146379, 0.01330781, 0.01555522, 0.02193911, 0.003089319, 
    0.001841971, 0.0009087413, 0, 0, 0, 0.0003210456, 0.02449383, 
    0.005104381, -0.0001122077, 0, 0,
  0, 0.003011848, 0.02298257, 0.009286834, 0.009608928, 0.01336056, 
    0.002232636, 0.0061625, 0.01146719, 0.003902888, 0.009420566, 
    0.003512637, 0.01121188, 0.01299424, 0.07003881, 0.03355437, 0.00279008, 
    0.0001397496, 6.611073e-09, 9.075566e-06, 0, 0, 0, 0.01391281, 
    0.02563607, 0.001862354, -1.070268e-05, 0, 0,
  0, 0, -1.720165e-06, 0, 0.02618093, 0.01672088, 0.005894753, 0.007721313, 
    0.010417, 0.0139837, 2.963469e-05, 0.0007133319, 0.01063, 0.01352865, 
    0.01560032, 0.002732558, -3.247629e-05, 0.002673132, -0.0001034007, 
    -4.337428e-05, 1.644952e-05, 0, 0.0006585207, 0.002192543, 0.003581958, 
    0.0154322, -1.121631e-05, 0, 0,
  0, 0, 0, 0, -4.90726e-05, -1.591607e-05, -2.225983e-05, 1.92625e-05, 0, 
    -0.0001517891, 0.02582862, 0.006632818, 0.01181327, 0.003225856, 
    -0.0001942483, 0.001114418, 0.007654375, 0.00539556, 0.0157277, 
    0.004172458, 0.00360429, -9.865784e-05, -1.583018e-07, 0, 2.765312e-06, 
    0.0009316398, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0002135721, 7.105841e-05, -4.52085e-08, 0, 
    0, 0, -7.57318e-07, 0.002172984, -1.506675e-06, -7.031441e-05, 
    -7.812295e-06, -3.60731e-11, 0, 0, -3.687996e-07, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, -7.011781e-05, 2.025833e-07, -2.612773e-06, 
    8.507218e-05, 0, -7.944911e-09, 0, 2.690436e-05, 0.004386348, 
    -1.636628e-06, 0, 0, 0, 0, 4.231515e-05, 0, 0.002959311, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.55144e-06, 0, 0, 0, -2.868499e-06, 0, 
    0, -5.108698e-06, 0, 0, 0, -1.284673e-05, 0.001676772, 0.0003954085, 
    0.001004518, 0.0006913315, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4.290527e-05, 0, 0, 0, 
    0, 0, -2.082235e-05, 0, 0, -5.113245e-07, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, -1.491983e-07, 0, 0, 0, 0.0002199464, 0, 3.854968e-05, 0, 0, 0, 0, 
    0, 0, 0.00263276, -0.0001153117, 0.001814128, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0006299565,
  0.000336635, 0.0002343797, -4.505108e-06, 0.001754712, 0.003273813, 
    0.002938466, 0.006359805, 0.006314048, 0.001220909, 0, 0, -6.679567e-05, 
    0.01075295, 0.002517766, -7.857216e-05, 0.01431278, 0.003399687, 
    -3.124116e-06, 0, -2.991878e-08, 0.001531523, -7.590325e-05, 0.002349593, 
    0.0005512371, 0, 0.007276746, 0.002126951, 0.003353781, 0.001238094,
  0.0002349804, -1.841046e-05, 0.0007000676, 0.0008256562, 0.01309241, 
    0.02233464, 0.008941958, 0.00317748, 0, -7.526215e-07, 0.005935864, 
    0.01631838, 0.007353608, 0.01595988, 0.01643996, 0.02247189, 0.006188274, 
    0.002227526, 0.013726, 0.006652614, -0.0001263535, 0, 0, 0, 0.005895807, 
    0.02453544, 0.005520717, 0.003459325, 0.002559583,
  -1.963082e-05, 0, 0.002217478, -6.652906e-05, 0.06838825, 0.009760998, 
    0.01183955, -2.312035e-06, 0.005139633, 0.00111013, 0.001094445, 
    0.001900626, -5.702559e-05, 0.02416542, 0.02747432, 0.001053408, 
    0.01387977, 0.0209007, 0.02624534, 0.00224756, 0, 0, 0, 0, 0.001856267, 
    0.04528399, 0.00965487, 0.00517921, 0.003445577,
  1.943251e-06, 0.005146621, 0.011926, 0.01761701, 0.07896107, 0.03136012, 
    0.00265955, 0.04259906, 5.506047e-06, 0.02558525, 0.03312513, 0.02170077, 
    0.04762623, 0.03250823, 0.04251686, 0.03535925, 0.03218257, 0.007893899, 
    0.003343752, 0.004210412, 0, -9.615113e-10, 0, 0.001783954, 0.05387048, 
    0.01227961, 0.0002175196, 0, 0,
  0, 0.005416088, 0.04506553, 0.02243974, 0.02637277, 0.0222047, 0.007576573, 
    0.01054549, 0.02795324, 0.01037958, 0.01959161, 0.01948646, 0.02980298, 
    0.0791126, 0.1199366, 0.04299139, 0.011953, 0.0005458089, -1.046723e-05, 
    4.186916e-05, 0, 0, 1.564681e-09, 0.06048325, 0.06832609, 0.01003279, 
    0.00015867, 0, 0,
  0, -6.496797e-06, -1.034834e-05, 0.00017772, 0.04321846, 0.03159788, 
    0.01687145, 0.01346153, 0.02927011, 0.02134521, 0.002202786, 0.00346814, 
    0.02811087, 0.04401673, 0.029317, 0.004937334, -0.0001011014, 
    0.006262041, 0.001445705, -0.0001050451, 0.002107344, 0, 0.002711225, 
    0.0139339, 0.01575147, 0.02810684, 0.000724947, 0, 0,
  0, 0, 0, -6.633497e-07, 0.001125791, -4.7744e-05, 3.286454e-05, 
    0.000132562, 1.425438e-06, 3.70896e-05, 0.05412559, 0.01953745, 
    0.01986727, 0.01395126, 0.0007285652, 0.0016237, 0.02001589, 0.01749869, 
    0.02525064, 0.0133537, 0.008560489, 0.004866506, 0.001829096, 0, 
    0.0001643227, 0.003227887, -4.001565e-05, -7.985271e-07, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0001602455, 0.003169782, 0.001069278, 
    0.0001348455, -4.081206e-06, 5.272725e-08, -8.377516e-08, 0.004903212, 
    0.009304799, 0.0007084367, 0.00319779, 0.0008554552, 0.002706196, 0, 0, 
    -7.44627e-05, -5.746066e-08, 0, 1.897993e-06, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, -0.0001567419, 1.274854e-05, 0.0003075614, 
    0.0003741768, 0.0001171895, 0.000212919, -7.704782e-06, 0.000934797, 
    0.01591155, 7.895593e-05, -1.975901e-08, -4.223795e-06, 0.0003403044, 
    0.001638686, 0.006452517, 6.29059e-05, 0.008949078, -1.32246e-08, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.002521419, -5.350763e-07, 0.001358772, 0, 
    0, -3.463356e-05, -2.91111e-05, -8.270772e-07, -9.932154e-06, 
    -3.116135e-05, 0, -1.033797e-05, 0.001895456, 0.007438816, 0.00595132, 
    0.004056196, 0.004088432, 0, 0,
  -3.755468e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2.947955e-05, 0, 0, 0, 0, 0, -4.949469e-05, -2.874619e-05, 0.0004391618, 
    0.0001531941, 0.0008669837, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  -1.444221e-05, 0, 0, -1.108663e-05, 0.0003096772, -7.496168e-07, 0, 
    0.0009208738, 0.0009572044, 0.0007114056, 0, 0, 0, -2.997431e-06, 
    1.691827e-05, -5.809824e-06, 0.005487234, 0.003996763, 0.005175048, 0, 0, 
    0, 0, 0, 0, 0, -1.115772e-06, -1.069464e-06, 0.001415802,
  0.002900735, 0.002443856, 0.0003498947, 0.00681199, 0.01214954, 0.01249237, 
    0.01395047, 0.01713581, 0.004951125, 0.001503557, 0.000229672, 
    0.0005441248, 0.01831478, 0.01169143, 0.002960031, 0.0249393, 
    0.006234739, 0.0006284838, -2.52193e-05, 0.0002598802, 0.005957415, 
    0.009101236, 0.00788765, 0.001742866, -2.256175e-05, 0.01526742, 
    0.005216493, 0.0116046, 0.006758687,
  0.005886977, 0.0007179244, 0.001938681, 0.007522382, 0.02520277, 
    0.03597369, 0.01284031, 0.008095955, 5.89014e-08, 0.000231593, 
    0.02013691, 0.03281756, 0.01308837, 0.03246696, 0.03860691, 0.06819069, 
    0.01368517, 0.01288928, 0.02875025, 0.02378815, 0.004420205, 
    0.0003824363, 0.0006272406, 7.050756e-08, 0.01032475, 0.03565359, 
    0.02321542, 0.01411866, 0.008423901,
  -0.0001019697, -7.169994e-07, 0.01164365, 0.005168422, 0.1006598, 
    0.04489516, 0.02421996, 0.000698751, 0.01502733, 0.001955329, 0.01646988, 
    0.01843537, 0.003837255, 0.05929628, 0.07787388, 0.01204295, 0.03101542, 
    0.04687348, 0.04397767, 0.003994867, -4.764717e-05, 3.802677e-05, 
    1.374658e-10, 0, 0.01369255, 0.09656402, 0.01651503, 0.007674302, 
    0.01000521,
  0.0002823143, 0.0335873, 0.03811097, 0.06631474, 0.1769367, 0.07246286, 
    0.009721467, 0.05467599, 0.0009516153, 0.07165661, 0.1565668, 0.1238779, 
    0.1245259, 0.08302689, 0.1515059, 0.1044058, 0.08463567, 0.03581092, 
    0.006999371, 0.009034394, 6.355277e-06, -3.956871e-05, -1.30208e-05, 
    0.007087761, 0.2328496, 0.03401357, 0.004686056, -1.944504e-12, 
    -1.55819e-07,
  1.183342e-07, 0.01395721, 0.1068773, 0.07025205, 0.06402668, 0.06532887, 
    0.0333472, 0.05361259, 0.0774244, 0.1268071, 0.1029722, 0.1897317, 
    0.2185294, 0.3156835, 0.3262307, 0.1073214, 0.05708491, 0.02026558, 
    0.0001947797, 0.002666614, 0.0005777919, -4.680263e-09, 0.01708061, 
    0.1932828, 0.2533574, 0.04158471, 0.001659798, 1.505872e-05, 0,
  -9.628722e-10, 0.0009845787, 2.133309e-05, 0.000837235, 0.06504928, 
    0.06163283, 0.06937367, 0.03865109, 0.09319404, 0.06136182, 0.05390777, 
    0.07042958, 0.1585415, 0.2543817, 0.09374598, 0.02145585, 0.005841017, 
    0.01632345, 0.009434089, 0.003359699, 0.004235359, 1.967817e-09, 
    0.00418393, 0.06748998, 0.0694347, 0.06328756, 0.001877589, 0.0006470042, 0,
  2.461289e-05, 0, -1.132698e-08, -8.238177e-06, 0.007817479, 0.000376592, 
    0.000317551, 0.008170359, -2.992784e-05, 0.0009012511, 0.1088532, 
    0.08253603, 0.06109682, 0.04727827, 0.0193693, 0.003604252, 0.04250322, 
    0.02881365, 0.03850433, 0.02774323, 0.01264918, 0.01351114, 0.004562375, 
    1.960419e-05, 0.000336874, 0.007242674, 0.000195934, -2.004974e-05, 
    9.280538e-06,
  -1.519884e-06, 0, 0, 1.449178e-08, 6.660235e-08, 2.096211e-08, 
    -4.498309e-06, 0, 0, 0.0003209072, 0.00690372, 0.002020005, 0.00131213, 
    -1.427216e-05, 0.0001925635, -1.879838e-06, 0.01666835, 0.0256538, 
    0.01795968, 0.01168178, 0.006981174, 0.0114979, -2.159676e-05, 
    -7.997683e-08, -0.0004505308, -3.564758e-06, -1.376761e-09, 0.001296373, 
    2.314418e-05,
  0, 0, 0, 0, -2.343606e-07, 7.000125e-07, -1.064996e-09, 0, 0, 0.002703426, 
    0.003457398, 0.003158808, 0.004424176, 0.002651021, 0.006430039, 
    0.004328564, 0.006741662, 0.0414649, 0.003485892, -3.894473e-05, 
    -7.430732e-05, 0.002703601, 0.004337495, 0.01013622, 0.004309162, 
    0.01526257, 0.0002667761, 0.001313007, 0,
  5.034953e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.006130937, -4.755484e-05, 
    0.005019878, 0.0009493285, -6.043496e-06, 0.00828755, -0.0001679451, 
    0.01087573, 0.0007955974, 0.001930616, 0, -5.112329e-05, 0.008028113, 
    0.01713364, 0.01292377, 0.009241605, 0.01248093, 0.002068053, 7.668415e-06,
  -2.035268e-05, 0.0004899903, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -9.10263e-06, 0, 
    0, 0, 0.0003337176, 0.001722525, 0.000426225, -4.563415e-06, 0, 
    -1.695807e-05, -1.529113e-05, 0.0003127585, 0.0002677238, 0.00362319, 
    0.002701612, 0.004124544, 0.0007088249,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.0006486729, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -4.191977e-06, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0.0004940704, -1.362273e-08, -5.645397e-09, -1.301563e-05, 0.00123512, 
    0.001877536, 0.0002436888, 0.003394053, 0.002168723, 0.001433215, 
    -8.108493e-06, 0.001399115, -6.195533e-06, 3.216824e-05, 0.004206372, 
    0.002609312, 0.01407906, 0.008527359, 0.009053306, -2.236082e-05, 0, 0, 
    0.0005975948, 0.000130033, -1.368767e-05, -0.0001611423, 0.0002523215, 
    0.0009560414, 0.00204147,
  0.01015896, 0.008970466, 0.002981373, 0.0145406, 0.02052665, 0.03046934, 
    0.02329888, 0.02599112, 0.01539012, 0.005243952, 0.002196174, 
    0.002913098, 0.02876772, 0.02727632, 0.01586038, 0.03744537, 0.01758788, 
    0.007439528, 0.002365412, 0.00390492, 0.01131624, 0.025436, 0.01797052, 
    0.007527811, 8.737561e-05, 0.02330176, 0.02106915, 0.03015797, 0.02210782,
  0.02849647, 0.008398283, 0.004107007, 0.02125126, 0.05644798, 0.1086387, 
    0.05513325, 0.02354775, 0.002482238, 0.004666857, 0.03365146, 0.05838758, 
    0.03207828, 0.05713468, 0.08513625, 0.1373229, 0.06012727, 0.05130231, 
    0.05270698, 0.05101683, 0.02795832, 0.004878258, 0.002634413, 
    0.001712847, 0.02334042, 0.07364506, 0.100288, 0.06303123, 0.03495404,
  -0.0001748401, 4.027249e-06, 0.08374282, 0.02951898, 0.1397817, 0.1394282, 
    0.1122071, 0.04681712, 0.06240322, 0.01390401, 0.03857644, 0.03773436, 
    0.01916873, 0.150152, 0.1656404, 0.08192413, 0.1270812, 0.1710847, 
    0.1767152, 0.04402181, 0.000845441, 0.0259697, 0.003551813, 
    -2.712917e-05, 0.08069277, 0.2389809, 0.1501783, 0.0615503, 0.02495223,
  0.004320382, 0.1388111, 0.1574747, 0.05863912, 0.1830132, 0.09995991, 
    0.01719022, 0.06645782, 0.0009150201, 0.05613707, 0.1406715, 0.1216465, 
    0.1133012, 0.07650761, 0.128236, 0.1341505, 0.1848605, 0.1887199, 
    0.09969181, 0.07474854, 0.00144481, 0.02441927, 0.01059208, 0.009047274, 
    0.2405078, 0.160697, 0.09706166, 0.009713298, -8.10446e-05,
  0.002287844, 0.08930105, 0.4990917, 0.2771019, 0.1197851, 0.1248561, 
    0.08248568, 0.06562023, 0.09277258, 0.1340339, 0.1111672, 0.1642278, 
    0.1727452, 0.2499341, 0.2915675, 0.1146683, 0.07739979, 0.04695228, 
    0.02775143, 0.01020694, 0.01612632, 7.301003e-07, 0.06739774, 0.4246916, 
    0.3891182, 0.2271498, 0.1628569, 0.03877104, 7.993533e-07,
  9.594554e-06, 0.04641776, 0.1332625, 0.08177485, 0.1284656, 0.232127, 
    0.1557948, 0.1722953, 0.3064005, 0.2453499, 0.08512964, 0.1200397, 
    0.1594304, 0.2163483, 0.06513214, 0.01021672, 0.004513186, 0.02741356, 
    0.01572787, 0.01397915, 0.01293549, 2.164219e-06, 0.009142788, 0.297601, 
    0.3101045, 0.1989243, 0.1219507, 0.01532487, 3.621392e-07,
  0.0001137318, 5.466281e-06, 0.0001840624, 4.200204e-05, 0.04416269, 
    0.01678012, 0.02101646, 0.01691417, 0.002774152, 0.03177161, 0.1408966, 
    0.07894816, 0.04631645, 0.03206722, 0.01506794, 0.003549607, 0.05379373, 
    0.06295623, 0.1223657, 0.1225738, 0.1268836, 0.04106414, 0.00765017, 
    4.509102e-06, 0.005946493, 0.06194941, 0.05745209, 0.0907105, 0.000283921,
  0.0002340096, 3.288626e-05, -5.56148e-09, 7.031974e-06, 3.508973e-05, 
    6.961056e-05, 9.368747e-05, 2.03716e-05, 1.780754e-07, 5.378757e-05, 
    0.01640858, 0.002878728, 0.006872234, 0.001257281, 0.004789446, 
    -1.488471e-05, 0.03297583, 0.05527817, 0.06612545, 0.06874356, 0.1056312, 
    0.04949781, 0.007995061, 0.001269927, 0.001129301, -6.064482e-05, 
    0.0004347466, 0.0299279, 0.002913826,
  -2.797692e-06, -7.686882e-06, 0.0002147388, 0, 0.0001528218, 0.0007951912, 
    9.331322e-05, 0, 0, 0.009596888, 0.01328875, 0.02161194, 0.01289262, 
    0.01165447, 0.01675492, 0.01665458, 0.04089119, 0.08211744, 0.02045456, 
    0.003669956, 0.0009419642, 0.01955493, 0.01703615, 0.02065704, 0.0120039, 
    0.02150633, 0.004679071, 0.003247123, -5.118047e-07,
  0.0110362, -4.592892e-10, 1.399774e-07, 0, 0.0003055212, 0, 0, 0, 0, 
    -1.243021e-06, 0.008661953, 0.003712617, 0.007868643, 0.003996318, 
    0.002125264, 0.02507953, 0.007427855, 0.03437084, 0.01046991, 0.01086985, 
    -6.926874e-06, -8.941276e-05, 0.01495485, 0.04746722, 0.03254031, 
    0.02542416, 0.02254883, 0.006795683, 0.005145603,
  0.001558259, 0.001830962, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001204422, 
    -2.238204e-05, 0, 0, 0.001748581, 0.004689316, 0.001828669, 
    -1.318929e-05, 0, -2.918153e-05, -9.347345e-05, 0.001720778, 0.002061646, 
    0.007483245, 0.0119431, 0.01163649, 0.00251274,
  3.174235e-05, -1.323295e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, -1.514426e-05, 0.001627874, -8.112007e-06, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.032114e-08, 0, -6.908213e-05, 
    -2.496079e-05, 0.0007062772, -5.199444e-05, -3.676315e-07, -2.147276e-08, 
    0, 0, 0, -7.495229e-06, 0, 0, 0, 0, 0,
  0.001846784, 0.0001479768, 0.0007421268, 2.252514e-05, 0.00308982, 
    0.005052751, 0.0002011699, 0.004504285, 0.00450571, 0.001694524, 
    0.001252824, 0.00574512, -0.0001197168, 0.004643109, 0.02672868, 
    0.03503745, 0.04092495, 0.02810294, 0.01615606, -3.623344e-05, 
    -1.058754e-08, -7.207512e-06, 0.002333765, 0.002767992, 0.004726023, 
    0.002981311, 0.00649938, 0.006584173, 0.005010914,
  0.042302, 0.04525863, 0.04067521, 0.05589642, 0.05670925, 0.08439231, 
    0.0953251, 0.05520756, 0.04494748, 0.03044227, 0.04446954, 0.05327721, 
    0.07010676, 0.06152518, 0.07145953, 0.121632, 0.1302658, 0.0680948, 
    0.03756317, 0.02441949, 0.02825254, 0.07279769, 0.06003129, 0.02202459, 
    0.01026737, 0.04562494, 0.03713514, 0.07730414, 0.07799281,
  0.1099838, 0.05916596, 0.03263076, 0.05515428, 0.08649706, 0.1504372, 
    0.09962722, 0.08872022, 0.0394059, 0.07139587, 0.07750024, 0.1001732, 
    0.05455366, 0.07501309, 0.1144508, 0.1833615, 0.1347859, 0.1302561, 
    0.1228495, 0.1497625, 0.1095939, 0.06428026, 0.02459792, 0.006556286, 
    0.06992304, 0.1187986, 0.1447331, 0.1255976, 0.0947217,
  -0.0002374622, 7.282811e-06, 0.1124998, 0.02839937, 0.1293624, 0.1386934, 
    0.1222491, 0.05617607, 0.05846152, 0.0107435, 0.05090926, 0.03681355, 
    0.02565433, 0.1375908, 0.1611452, 0.09205425, 0.1781185, 0.2054999, 
    0.2239926, 0.1548896, 0.06763658, 0.01053041, 0.0008130734, 9.133061e-05, 
    0.09389393, 0.2273381, 0.1403017, 0.07795183, 0.06082729,
  0.00048927, 0.1031038, 0.1253794, 0.04834514, 0.1541904, 0.0872644, 
    0.009489976, 0.07172761, 0.001204199, 0.03875742, 0.1368926, 0.09176117, 
    0.1013152, 0.06865285, 0.112817, 0.1196741, 0.1588876, 0.1378557, 
    0.09356366, 0.08931834, 0.01630279, 0.01647673, 0.004122423, 0.009353455, 
    0.1904052, 0.1474883, 0.09210047, 0.002727518, -3.102347e-06,
  0.001287257, 0.0582952, 0.4694574, 0.2447848, 0.08784029, 0.08737655, 
    0.06081199, 0.0490967, 0.08331814, 0.1062734, 0.0905562, 0.1327809, 
    0.1268916, 0.199477, 0.2470466, 0.08818745, 0.05156069, 0.03437809, 
    0.0172454, 0.007470273, 0.01814834, 1.242543e-07, 0.0320227, 0.378228, 
    0.3388429, 0.1965751, 0.1283709, 0.01284714, 1.486122e-07,
  5.766817e-06, 0.02250591, 0.04930754, 0.07067034, 0.1018994, 0.173766, 
    0.1145027, 0.1213882, 0.2386068, 0.1939978, 0.05047807, 0.08265488, 
    0.116942, 0.1727444, 0.06298284, 0.00665928, 0.004722674, 0.01731356, 
    0.00632744, 0.006159502, 0.01053497, 1.044077e-06, 0.003428843, 
    0.1550064, 0.2693241, 0.1565903, 0.08181284, 0.009014995, 2.35873e-06,
  3.620599e-05, 3.928716e-06, 0.0001790038, 0.001085779, 0.02417988, 
    0.01218458, 0.008214924, 0.01034858, 0.001231604, 0.02035665, 0.134851, 
    0.06713292, 0.03518276, 0.02978342, 0.006515201, 0.003209686, 0.04524046, 
    0.0653953, 0.1046175, 0.07830173, 0.08590855, 0.03085711, 0.008306146, 
    -1.272678e-05, 0.001632702, 0.03625212, 0.04647175, 0.07850194, 0.02149743,
  0.1039875, 0.004893897, -1.593999e-06, 1.566438e-06, 6.279754e-06, 
    2.454064e-05, 6.617098e-06, 1.619827e-05, 1.256931e-07, 5.950125e-05, 
    0.01565926, 0.007369591, 0.0113589, 0.0005110955, 0.006773728, 
    0.0001419131, 0.03022859, 0.06165468, 0.09388594, 0.07486303, 0.09242785, 
    0.05381671, 0.01932453, 0.01669143, 0.007865705, 9.415053e-06, 
    0.00281255, 0.04475355, 0.1226215,
  0.004956037, 0.001756849, 0.002824914, -6.130015e-11, 0.001715643, 
    0.003096165, 0.005684472, 0, -5.127349e-14, 0.03133266, 0.02404227, 
    0.04206619, 0.03050108, 0.02775559, 0.03522647, 0.06135174, 0.06684079, 
    0.1429329, 0.1200646, 0.04075705, 0.008519285, 0.07947765, 0.1070013, 
    0.07352132, 0.07605571, 0.0644654, 0.02811813, 0.01003282, -0.0002299527,
  0.03571051, 0.0001642495, 3.225335e-05, 0, 0.0006597501, 0, -5.094264e-06, 
    0, 0, -1.040576e-05, 0.01287133, 0.0166909, 0.01754213, 0.01906574, 
    0.01174308, 0.04143089, 0.03069223, 0.06675559, 0.02953179, 0.02721427, 
    0.0006946882, 0.00976667, 0.03666356, 0.1154479, 0.09375536, 0.08241966, 
    0.06420946, 0.0272022, 0.0249029,
  0.007703144, 0.00273511, -1.113944e-06, 0, 3.820187e-06, 0, 0, 0, 0, 0, 0, 
    -2.491797e-05, 0.006123343, 0.0006179846, 0.0002147575, 0.002053342, 
    0.005661078, 0.009042653, 0.008401988, 0.0002877824, -6.976227e-10, 
    0.0002880565, 0.0001809663, 0.00456463, 0.006653453, 0.01590078, 
    0.02952839, 0.0309726, 0.008665836,
  0.00105154, 0.0002410715, -2.11847e-05, 8.164209e-05, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, -4.020143e-05, 0, 0, 0, 0, 0, 0, 0, 0.0007386389, 
    0.003934659, 0.001964537, 0.001173544,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 8.028651e-05, 3.124892e-06,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  -3.033003e-05, 0, 0, 0, -6.053036e-06, 0, -7.060225e-07, -3.876358e-05, 
    -5.630121e-05, -8.694356e-06, 0, 0, -6.70785e-08, 4.245507e-07, 
    0.0007532686, 0.002502698, 0.006106541, 0.003903762, 2.995978e-05, 
    -9.111258e-06, 0, 0, 7.590625e-07, 0.0007033853, 0, 0, 0, 0, -2.087745e-05,
  0.01634221, 0.02324029, 0.02457476, 0.005069041, 0.03747144, 0.03850536, 
    0.04104137, 0.02062833, 0.03038538, 0.02362654, 0.02474292, 0.0214432, 
    0.01289759, 0.04417208, 0.08987622, 0.107632, 0.1028283, 0.08119398, 
    0.05449836, 0.006881807, 0.000230515, -2.485973e-06, 0.002785972, 
    0.01961575, 0.0348841, 0.02086773, 0.03697249, 0.04039289, 0.02355538,
  0.09979989, 0.08814291, 0.1035666, 0.1413529, 0.1721497, 0.1750165, 
    0.1370178, 0.1571413, 0.1086098, 0.08799266, 0.1082026, 0.1516499, 
    0.1588256, 0.1158073, 0.1013578, 0.1691847, 0.1604463, 0.1064973, 
    0.09833187, 0.1017755, 0.1220816, 0.1815591, 0.1510098, 0.05682464, 
    0.09905528, 0.1367426, 0.09269731, 0.1408253, 0.1447675,
  0.09826447, 0.06706921, 0.03074344, 0.05298153, 0.07048093, 0.1416432, 
    0.08628826, 0.1024683, 0.03390364, 0.06493649, 0.070635, 0.1042578, 
    0.05508529, 0.07359245, 0.1258661, 0.1999002, 0.1242976, 0.1102822, 
    0.1195577, 0.1478258, 0.1182083, 0.06062584, 0.01585647, 0.01540208, 
    0.07012814, 0.1099112, 0.1251885, 0.1316535, 0.1006192,
  -0.0002204508, 1.074032e-05, 0.1145665, 0.02190797, 0.1073672, 0.150766, 
    0.1158769, 0.05253775, 0.0506817, 0.01578134, 0.05409845, 0.03724267, 
    0.02037159, 0.1275804, 0.1446445, 0.0729334, 0.1645106, 0.1847506, 
    0.2010142, 0.1216509, 0.05364409, 0.00327288, 0.0001661171, 0.0004566582, 
    0.07605084, 0.2048697, 0.1286761, 0.06443538, 0.05434049,
  0.0002076483, 0.08220863, 0.1015208, 0.04564767, 0.1378684, 0.07776333, 
    0.009230837, 0.0570591, 4.30823e-05, 0.0338709, 0.1437685, 0.0720399, 
    0.08826139, 0.07055408, 0.1116816, 0.1106051, 0.1609407, 0.1144476, 
    0.07345211, 0.06602744, 0.01510235, 0.007769217, 7.747026e-05, 
    0.008026881, 0.15849, 0.1389551, 0.08594956, 0.002024772, 1.090969e-05,
  0.0004527936, 0.03970858, 0.4245879, 0.2289236, 0.07781976, 0.07071619, 
    0.05261046, 0.04123713, 0.08017445, 0.09591255, 0.07953694, 0.1200461, 
    0.09408057, 0.1627638, 0.2240316, 0.08926567, 0.04742227, 0.0135216, 
    0.008188149, 0.006081246, 0.01048246, 4.364574e-08, 0.01188943, 0.349486, 
    0.3265312, 0.1718347, 0.07931762, 0.002654725, 4.55019e-08,
  7.511737e-06, 0.01388368, 0.01155215, 0.02964976, 0.08746058, 0.1401086, 
    0.1094893, 0.100423, 0.2008799, 0.1726815, 0.03665195, 0.05923114, 
    0.0972169, 0.1530715, 0.06379706, 0.004787668, 0.008653034, 0.02211115, 
    0.004816966, 0.004040641, 0.01119551, 6.967809e-09, 0.002162252, 
    0.08676035, 0.2176545, 0.1482015, 0.0601079, 0.005204671, 5.858582e-07,
  4.647417e-06, 1.737406e-06, 4.330678e-05, 0.0003994081, 0.01966968, 
    0.01009459, 0.005427483, 0.007122809, 0.001530385, 0.01447115, 0.1360717, 
    0.06494507, 0.03512705, 0.02830501, 0.004721782, 0.005517041, 0.0448099, 
    0.06743564, 0.09783866, 0.06735451, 0.06614216, 0.01757056, 0.008860166, 
    0.0002041283, 0.001862864, 0.02338633, 0.04473776, 0.04394805, 0.01993624,
  0.09241663, 0.00504729, -2.779495e-06, 1.506888e-07, 2.12923e-06, 
    1.133275e-05, 2.214154e-06, 8.003752e-06, 1.673725e-07, 0.000230999, 
    0.01309731, 0.01429482, 0.01540505, 0.002236532, 0.0117098, 0.0006378485, 
    0.02422815, 0.06064726, 0.08884398, 0.04790368, 0.06183817, 0.03911392, 
    0.01411457, 0.01642043, 0.008770383, 0.0006351814, 0.01187612, 0.0629761, 
    0.1814814,
  0.04972105, 0.03132145, 0.005916904, 1.484467e-05, 0.002784649, 0.01194927, 
    0.01453979, 0, 3.065868e-11, 0.06852396, 0.05137044, 0.06311402, 
    0.05895582, 0.05579849, 0.08295503, 0.1252484, 0.13171, 0.2189178, 
    0.1967097, 0.09013403, 0.03011641, 0.1110776, 0.1498228, 0.0992912, 
    0.1071746, 0.06812783, 0.08086175, 0.06373959, 0.01742657,
  0.07458379, 0.02133536, 0.0008753266, 0.001310973, 0.004070414, 
    0.002680193, -9.45956e-06, 0, 0, -2.796926e-05, 0.02320533, 0.02401472, 
    0.03256284, 0.04134368, 0.03091546, 0.0930372, 0.09328131, 0.1952641, 
    0.1097025, 0.06155146, 0.002776591, 0.02847545, 0.09901468, 0.185152, 
    0.1942337, 0.1697456, 0.1248073, 0.05380109, 0.0491933,
  0.04105491, 0.006505239, 0.0005871847, 1.458631e-05, 0.000873555, 0, 0, 0, 
    0, 0, 0, -6.097851e-05, 0.01279459, 0.00526247, 0.0007070057, 
    0.005837382, 0.01129707, 0.03459832, 0.0485386, 0.01090479, 2.618716e-05, 
    0.002903398, 0.004829445, 0.00870976, 0.01471661, 0.02924319, 0.05942302, 
    0.04867807, 0.0428834,
  0.007627334, 0.002536654, 0.001784539, 0.001453768, 0.0003960566, 0, 0, 0, 
    0, 0, 0, 0, -7.794454e-06, -1.205e-06, 0, 0, -8.658988e-06, 0.003181254, 
    0.0002847681, -1.57107e-05, 6.367983e-11, 0, 0, 0, -6.203366e-06, 
    0.00283114, 0.01838826, 0.01142059, 0.005982121,
  -2.808312e-05, 1.949733e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, -2.812367e-06, 0.0005943917, 0.00137695,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0.007771883, 0.01200579, 0.01482662, 0.002049395, -6.199459e-05, 
    -0.0001449713, 0.001790024, 0.00117558, -1.264622e-05, -0.0009079898, 
    -2.255367e-05, -1.111559e-07, -0.0001807226, -0.0004358545, 0.03134069, 
    0.04581322, 0.04469068, 0.02704356, 0.01593483, 0.006525125, 
    -0.0002056825, 0.003333765, 0.007657141, 0.006809706, 0.008877059, 
    0.01021473, 0.005856161, 0.002781288, 0.008865846,
  0.0558879, 0.06435267, 0.04040974, 0.06137302, 0.06564121, 0.07069184, 
    0.08903979, 0.07815816, 0.09472682, 0.09163956, 0.07977113, 0.090863, 
    0.09853921, 0.1569487, 0.1507683, 0.1415771, 0.1403227, 0.113526, 
    0.08877848, 0.05380337, 0.03232509, 0.02421012, 0.02631365, 0.05431974, 
    0.08669703, 0.09172612, 0.1110982, 0.1035546, 0.05232852,
  0.1413544, 0.1438787, 0.1570743, 0.1924208, 0.2038628, 0.1779091, 
    0.1541847, 0.1626158, 0.154211, 0.151331, 0.1416068, 0.1885232, 
    0.1779135, 0.1315302, 0.09677599, 0.162039, 0.1468037, 0.1159197, 
    0.1145036, 0.129907, 0.158917, 0.2107995, 0.178924, 0.09955859, 
    0.1214947, 0.1675474, 0.1166349, 0.1509592, 0.1658047,
  0.08081166, 0.0590045, 0.02902993, 0.04712334, 0.06519487, 0.1370874, 
    0.08073467, 0.1006183, 0.02222054, 0.05594581, 0.05513975, 0.0983509, 
    0.05757583, 0.06079642, 0.1199052, 0.1719414, 0.1194523, 0.08899309, 
    0.1144819, 0.1460699, 0.1064176, 0.04720598, 0.0163283, 0.01538275, 
    0.07232937, 0.09076849, 0.1035903, 0.1236622, 0.08365421,
  -0.0001021565, 7.694872e-05, 0.1106463, 0.03046197, 0.09617403, 0.1510906, 
    0.1106539, 0.03464802, 0.04971273, 0.01356045, 0.04954549, 0.03296758, 
    0.01848679, 0.1233899, 0.1262302, 0.05640014, 0.1476805, 0.1744238, 
    0.1784919, 0.1192471, 0.03741665, 0.002252215, 1.814966e-05, 
    0.0004039012, 0.05457816, 0.1883163, 0.1362595, 0.0664925, 0.04576234,
  0.0001625472, 0.06773701, 0.07889503, 0.0378396, 0.1417252, 0.06513787, 
    0.007392675, 0.05822311, 1.820028e-05, 0.03068333, 0.1533276, 0.05777361, 
    0.08115707, 0.07132129, 0.1221742, 0.1063891, 0.1605874, 0.09829301, 
    0.0571161, 0.05996341, 0.003899866, 0.01239668, 3.460393e-05, 
    0.005904887, 0.1225638, 0.146314, 0.0829962, 0.01013984, 0.0008739922,
  1.169127e-05, 0.0326772, 0.389859, 0.2001703, 0.06810222, 0.05532035, 
    0.04891402, 0.03577064, 0.07472833, 0.08425929, 0.06942134, 0.1104026, 
    0.07143132, 0.1278748, 0.2123515, 0.08643351, 0.04494022, 0.008427801, 
    0.007028859, 0.00591339, 0.0001650777, 2.892177e-08, 0.007605747, 
    0.2857105, 0.306015, 0.1436021, 0.04178659, 0.0001274922, 2.770431e-09,
  2.068368e-06, 0.008245391, 0.004571859, 0.01482418, 0.07670297, 0.1132076, 
    0.09003136, 0.08290836, 0.1580061, 0.1412012, 0.02442375, 0.04623888, 
    0.08193781, 0.1270799, 0.06742524, 0.006045073, 0.01081505, 0.01363431, 
    0.01233906, 0.006526456, 0.01359074, 7.484236e-08, 0.002164217, 0.044827, 
    0.1680524, 0.155884, 0.05013205, 0.003898209, 4.579065e-07,
  1.507476e-06, 4.629869e-07, 8.744533e-06, 0.0003029451, 0.01713881, 
    0.006322789, 0.002295653, 0.005563241, 0.001545222, 0.0128522, 0.1371614, 
    0.05925928, 0.03291297, 0.02665272, 0.003560264, 0.008340293, 0.05111299, 
    0.07364964, 0.07780892, 0.0658865, 0.05491931, 0.002154016, 0.01280402, 
    0.001437374, 0.002942709, 0.02186247, 0.04033465, 0.04602633, 0.006624764,
  0.1026888, 0.002875114, -1.891409e-06, 3.460867e-08, 1.33798e-06, 
    2.441382e-05, -4.98247e-06, 2.020164e-06, 1.847467e-07, 0.0001462551, 
    0.01572119, 0.01099875, 0.00662909, 0.005374253, 0.01765491, 0.000600785, 
    0.02529504, 0.06206091, 0.07957971, 0.05135837, 0.04876908, 0.03078838, 
    0.009868779, 0.01723218, 0.007707718, 0.001889601, 0.0298315, 0.04866043, 
    0.1638582,
  0.06611606, 0.05383089, 0.01752905, 0.005699601, 0.004496687, 0.03647564, 
    0.01884329, -9.196175e-10, -7.547851e-06, 0.1203918, 0.08475615, 
    0.06606643, 0.07028047, 0.07030236, 0.1233106, 0.1449697, 0.1423395, 
    0.215355, 0.1422366, 0.05784554, 0.05625844, 0.09639058, 0.1450417, 
    0.07133303, 0.06924438, 0.05903926, 0.06817432, 0.081819, 0.04677259,
  0.114094, 0.04066971, 0.0189427, 0.00945829, 0.005430052, 0.005791703, 
    0.0002032491, -1.581193e-05, 0.002182008, -1.052791e-05, 0.02955581, 
    0.04529487, 0.07099926, 0.07186213, 0.06522621, 0.1461572, 0.1732597, 
    0.2369568, 0.1531663, 0.09209812, 0.008831032, 0.08597933, 0.1579698, 
    0.2214851, 0.2031318, 0.210646, 0.2024618, 0.1376509, 0.1404276,
  0.07500732, 0.02920642, 0.02232447, 0.007490906, 0.002942219, 0, 0, 0, 0, 
    0, 0, 0.0002078091, 0.01657541, 0.01469073, 0.01564129, 0.01307435, 
    0.03241746, 0.1008731, 0.1579232, 0.02925167, 0.005433429, 0.02156411, 
    0.032326, 0.02406262, 0.0588097, 0.07516085, 0.1303868, 0.1174642, 
    0.07379629,
  0.04288492, 0.02284101, 0.01044109, 0.006482448, 0.0008990005, 
    -2.602732e-06, 0, 0, 0, 0, 0, -1.589229e-06, -8.973845e-05, 0.003881419, 
    0.003612584, 4.053206e-08, -0.0001393599, 0.01852736, 0.003684155, 
    0.002244669, 0.0007700893, 0, 1.594209e-07, -8.601229e-09, 0.001116778, 
    0.00841555, 0.04514835, 0.03881482, 0.03610683,
  0.005579875, 0.003849061, 0.0007313861, -1.715833e-05, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, -7.619605e-06, 0.002439532, 0, 0, 0, 0, 0, 0, 0, 
    1.640381e-05, 0.003198756, 0.006138767,
  -9.299694e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.0002592868,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0.0006926763, -0.0003605429, 
    0.002005627, -4.819438e-06, 0, 0, 0, 0, 0.0001145009, -1.171818e-05, 
    -2.055948e-07, 0, 0, 0,
  0.03902423, 0.04143805, 0.03621709, 0.02278561, 0.0006440808, 0.001693444, 
    0.02141832, 0.001677708, 0.004938369, 0.005947994, 0.003106165, 
    -9.759374e-05, 0.0005881491, 0.0348179, 0.09025863, 0.1177963, 0.1497829, 
    0.1078279, 0.09142917, 0.0580392, 0.06276578, 0.03293984, 0.02030835, 
    0.01693711, 0.06298266, 0.05955896, 0.02636255, 0.04756861, 0.01728825,
  0.1089282, 0.09009624, 0.0592311, 0.1200826, 0.1278727, 0.1135577, 
    0.1499013, 0.1377231, 0.1408305, 0.1356078, 0.1627366, 0.1506795, 
    0.1801542, 0.2146438, 0.1805971, 0.1484649, 0.1438636, 0.1302897, 
    0.1203937, 0.09156929, 0.0775156, 0.06357536, 0.09914477, 0.1399931, 
    0.1788225, 0.1459954, 0.1874802, 0.1549469, 0.1154882,
  0.155615, 0.1886477, 0.1868252, 0.1817802, 0.193509, 0.1620378, 0.1420332, 
    0.1557018, 0.1755354, 0.1909833, 0.1492226, 0.1784169, 0.1886001, 
    0.1482639, 0.09036337, 0.1624854, 0.1319482, 0.120757, 0.1251247, 
    0.1390622, 0.1555929, 0.2010193, 0.1768084, 0.09896396, 0.119863, 
    0.1693335, 0.1206783, 0.1422193, 0.169346,
  0.06824467, 0.05705575, 0.03072175, 0.05099846, 0.05828434, 0.1302889, 
    0.07797545, 0.08465579, 0.01961501, 0.04282299, 0.04850267, 0.09383342, 
    0.0553444, 0.05569585, 0.118616, 0.1565842, 0.1003305, 0.07329778, 
    0.1090569, 0.1519893, 0.1013891, 0.05441613, 0.01496612, 0.01008936, 
    0.0654782, 0.07762133, 0.08519144, 0.1104039, 0.06592193,
  0.0008772774, 1.602633e-07, 0.1099097, 0.01739925, 0.08491553, 0.1571776, 
    0.1012206, 0.02626183, 0.02840311, 0.01962657, 0.04975464, 0.01953327, 
    0.01425634, 0.1168336, 0.1326391, 0.02968507, 0.1463235, 0.1570101, 
    0.1632228, 0.1195999, 0.02525289, 0.002615189, 5.706873e-07, 
    6.168303e-05, 0.04143155, 0.1611751, 0.107941, 0.05945044, 0.04132325,
  0.0002325458, 0.06056897, 0.05805808, 0.03226499, 0.1416456, 0.0580169, 
    0.004343156, 0.05829334, 3.925951e-05, 0.02638417, 0.1274851, 0.04300769, 
    0.07420935, 0.06627137, 0.1174768, 0.1013175, 0.1484075, 0.07660349, 
    0.04193493, 0.04675511, 0.001434805, 0.006323929, 2.369293e-05, 
    0.005602697, 0.09838714, 0.1372552, 0.07549108, 0.01398007, 0.0004067672,
  6.93739e-06, 0.02476555, 0.3432639, 0.1672617, 0.05075674, 0.0421863, 
    0.0392506, 0.03126801, 0.06584676, 0.07188152, 0.05626095, 0.09326765, 
    0.05780663, 0.09062503, 0.2033117, 0.077936, 0.03620311, 0.007198105, 
    0.005008196, 0.006094251, 3.614344e-06, -8.081374e-09, 0.004533949, 
    0.2209881, 0.2834556, 0.1261849, 0.02691768, 4.388632e-05, -5.786092e-09,
  -1.439861e-06, 0.007256665, 0.004091651, 0.009436593, 0.08628914, 
    0.08011273, 0.06905082, 0.06181027, 0.1148076, 0.1172051, 0.01745403, 
    0.02891145, 0.06343879, 0.08958632, 0.0670106, 0.005495645, 0.007256564, 
    0.008207224, 0.01117152, 0.01102579, 0.01349624, -1.517072e-07, 
    0.01368451, 0.02779751, 0.115733, 0.1636934, 0.03166062, 0.003382801, 
    5.087924e-07,
  4.470916e-07, 1.778271e-07, 5.803159e-06, 0.0005370519, 0.01745692, 
    0.004850458, 0.00256151, 0.002585316, 0.001398665, 0.01366689, 0.131384, 
    0.05376641, 0.038036, 0.02592488, 0.003652104, 0.009223562, 0.0605977, 
    0.07208391, 0.07501837, 0.06675382, 0.04782689, 0.00249419, 0.004902416, 
    0.0007555523, 0.004165251, 0.02008829, 0.03653534, 0.08584136, 0.00161332,
  0.08464159, 0.0007766609, 0.0001888277, -6.447634e-07, 1.986779e-06, 
    0.001240768, -6.911117e-05, 7.554139e-07, 2.301822e-07, 8.704744e-05, 
    0.02184512, 0.02649547, 0.007932548, 0.02058913, 0.01423721, 0.003134368, 
    0.02745359, 0.06684692, 0.05720483, 0.05016105, 0.04282608, 0.02849759, 
    0.004212415, 0.01833064, 0.006986396, 0.003492352, 0.01904487, 
    0.04208947, 0.1362896,
  0.0502792, 0.04374574, 0.01743589, 0.01352009, 0.007445599, 0.04041538, 
    0.01759228, -1.358608e-08, 0.0004936357, 0.1482902, 0.1060363, 
    0.08695779, 0.07124411, 0.07980555, 0.1322718, 0.1512465, 0.1316261, 
    0.1470237, 0.1034116, 0.04104029, 0.05869141, 0.08258958, 0.1234168, 
    0.05621428, 0.05625269, 0.04949258, 0.06119346, 0.05909404, 0.04332445,
  0.1490624, 0.08365303, 0.06024437, 0.03734027, 0.02762622, 0.02593245, 
    0.002423357, 0.02494763, 0.006008015, 0.007549062, 0.0486802, 0.09777449, 
    0.09589916, 0.1124533, 0.1226964, 0.1754612, 0.2075324, 0.2365287, 
    0.1359651, 0.1362996, 0.03354938, 0.1206583, 0.1830957, 0.2130259, 
    0.2098016, 0.2023267, 0.1965844, 0.1424883, 0.163721,
  0.1694974, 0.1004722, 0.07544179, 0.04784893, 0.0437429, 0.00601919, 
    7.759956e-05, -5.067998e-06, 0, 0, 0.004738105, 0.002975343, 0.05762513, 
    0.03640502, 0.05190663, 0.0624171, 0.08578499, 0.1282392, 0.2067286, 
    0.09623429, 0.0423323, 0.04750306, 0.07900257, 0.07127514, 0.1179234, 
    0.1203676, 0.1623672, 0.1435969, 0.1306173,
  0.1021981, 0.08534481, 0.05018456, 0.04403451, 0.005790699, 0.002863178, 
    -8.004114e-05, -2.719095e-09, 0, 0, 0, -6.356918e-06, 0.001246678, 
    0.009471454, 0.007806181, 0.02116394, 0.01879255, 0.04385049, 0.01625967, 
    0.01553095, 0.02164558, 0.01272523, 0.01255943, 0.0006930448, 
    0.008059754, 0.03047308, 0.0827769, 0.1186809, 0.09986968,
  0.02627171, 0.02917846, 0.00572504, 0.005149259, -8.096615e-06, 
    -2.59473e-05, -1.766061e-05, 0.001383875, 0, 0, 0, 0, -1.634777e-05, 
    0.01142659, 0.02931729, 0.01569657, 0.01756976, 0.009856528, 0.0128648, 
    0.01230934, 0.004141814, -3.721847e-08, 0, 0, 0, 7.454703e-06, 
    -3.668207e-06, 0.01951005, 0.02891599,
  -0.0001236701, 0.000166633, -1.379632e-07, -5.595229e-06, -2.281575e-06, 0, 
    0, 0, 0, 0, 0, 0, 1.139456e-06, 1.895389e-06, 5.949364e-09, 1.775386e-07, 
    -5.485198e-08, 4.880545e-07, 7.697406e-06, -4.102232e-09, 0, 0, 0, 0, 0, 
    0, 0, -6.798932e-05, 0.0003292223,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4.439429e-06, 0.0006311615, 
    0.01464317, 0.0619413, 0.04134853, 0.00242641, -1.424117e-05, 
    -2.185093e-06, 0, 0.00383306, 0.02270907, 0.0110929, 0.02546076, 
    0.01577564, -0.0001843927, 0,
  0.1534262, 0.1184341, 0.1359174, 0.07221896, 0.001159013, 0.009591414, 
    0.06499965, 0.00229435, 0.02227789, 0.03511689, 0.01660413, 
    -0.0002509286, 0.003384974, 0.1295657, 0.1560197, 0.1716461, 0.1899081, 
    0.1527924, 0.1634355, 0.1450349, 0.0866427, 0.065331, 0.115033, 0.145499, 
    0.1920562, 0.1341264, 0.06161075, 0.1278418, 0.1420388,
  0.1762182, 0.158328, 0.1386911, 0.1876848, 0.188705, 0.1457876, 0.1972421, 
    0.2120607, 0.1945879, 0.2133559, 0.2155511, 0.2014982, 0.2020731, 
    0.221599, 0.1633945, 0.1406106, 0.1504175, 0.1626466, 0.1554571, 
    0.1757436, 0.1526646, 0.1378387, 0.1755818, 0.2234862, 0.2540041, 
    0.1950355, 0.236334, 0.1845238, 0.180235,
  0.1735497, 0.1927886, 0.1919249, 0.1787427, 0.1816181, 0.1481202, 
    0.1237471, 0.1494514, 0.1706167, 0.1841726, 0.1713034, 0.1633081, 
    0.1725749, 0.1492599, 0.0870693, 0.1552898, 0.1226022, 0.1259648, 
    0.1220508, 0.1347558, 0.1531989, 0.1911526, 0.1736536, 0.09816504, 
    0.09492093, 0.1644192, 0.1198692, 0.1456952, 0.1696984,
  0.06351329, 0.04621909, 0.03105989, 0.05404909, 0.04941129, 0.1234316, 
    0.08309107, 0.08428477, 0.01124682, 0.02824183, 0.03404858, 0.07829623, 
    0.05529594, 0.05157031, 0.1142627, 0.1491286, 0.07386933, 0.06168931, 
    0.1125425, 0.1354096, 0.09017701, 0.05641758, 0.01533361, 0.006881739, 
    0.05514056, 0.07047758, 0.07596245, 0.1006564, 0.06202126,
  0.002071025, 5.899858e-07, 0.1035411, 0.01557222, 0.0790686, 0.1431122, 
    0.09102872, 0.02103793, 0.0202049, 0.02110837, 0.05085652, 0.01774375, 
    0.01172687, 0.1096561, 0.1468421, 0.02146333, 0.1467414, 0.145033, 
    0.137298, 0.09231055, 0.01037331, 0.00171197, 1.371392e-07, 
    -3.748496e-05, 0.03432211, 0.1528363, 0.07583811, 0.05788349, 0.03651833,
  1.019767e-05, 0.05278797, 0.04425398, 0.03601192, 0.1606937, 0.05391096, 
    0.004099852, 0.0597152, 9.124907e-05, 0.01924753, 0.1073398, 0.0310562, 
    0.06696977, 0.05681404, 0.1166049, 0.09600825, 0.1250585, 0.06205754, 
    0.0291836, 0.03838558, 0.0003533011, 0.001451697, 3.014988e-06, 
    0.006606923, 0.08108567, 0.141594, 0.04790935, 0.002201381, -8.026086e-06,
  1.336411e-05, 0.02193348, 0.2849877, 0.1257205, 0.03800473, 0.02972687, 
    0.03826947, 0.0300587, 0.05091377, 0.05760003, 0.04720197, 0.07726643, 
    0.05438747, 0.07559723, 0.1984057, 0.06626347, 0.02916116, 0.006503641, 
    0.003756813, 0.003272675, 9.356245e-07, 3.613681e-08, 0.002879006, 
    0.1676989, 0.2745785, 0.1109501, 0.01324832, 4.036286e-05, -1.348465e-07,
  1.650089e-05, 0.006946331, 0.004298443, 0.006952039, 0.08838219, 
    0.07464781, 0.07060204, 0.04831662, 0.09340508, 0.09771966, 0.01396655, 
    0.01764645, 0.04877193, 0.06522308, 0.0657002, 0.007525533, 0.01084366, 
    0.006634981, 0.01189153, 0.01881734, 0.0114575, -5.782138e-07, 0.0215799, 
    0.02387932, 0.07637862, 0.1726044, 0.01752068, 0.002251312, 2.109014e-06,
  9.334958e-08, 4.980901e-08, 1.375256e-06, 0.0008077263, 0.0107765, 
    0.007826242, 0.00109587, 0.001433137, 0.001177784, 0.01609677, 0.1331244, 
    0.04803077, 0.03821517, 0.02430384, 0.01907637, 0.008361721, 0.07436425, 
    0.06929101, 0.07532591, 0.0601015, 0.04861763, 0.0009969871, 0.001373599, 
    0.0006038367, 0.009806721, 0.01972214, 0.01717166, 0.03242071, 
    0.0001442557,
  0.04810046, 2.262459e-06, 1.338723e-05, -1.785244e-06, 2.090703e-06, 
    0.00370819, -5.184659e-05, 2.160049e-07, 6.850701e-08, 0.0001061934, 
    0.03635353, 0.03794612, 0.0046676, 0.02705537, 0.01777238, 0.01394057, 
    0.01892122, 0.06237221, 0.04091909, 0.04615759, 0.03221669, 0.02356857, 
    0.002259576, 0.01011476, 0.006150724, 0.003923804, 0.005540664, 
    0.03466066, 0.089513,
  0.03570985, 0.03203127, 0.01865226, 0.01761622, 0.01118944, 0.04095609, 
    0.01934913, 3.237935e-06, 0.004268331, 0.1712039, 0.1294817, 0.09089283, 
    0.07412681, 0.08915167, 0.1346253, 0.1522377, 0.1150925, 0.1141618, 
    0.08229473, 0.0357701, 0.05135875, 0.07504942, 0.1005126, 0.04239289, 
    0.05182423, 0.04308415, 0.05193216, 0.04695321, 0.04084884,
  0.1509664, 0.08998787, 0.07063144, 0.05174216, 0.1016103, 0.08324637, 
    0.01049473, 0.08345445, 0.04843246, 0.03285933, 0.08572295, 0.1257797, 
    0.1255807, 0.1381399, 0.1281846, 0.1837924, 0.2373676, 0.237299, 
    0.1353101, 0.1462037, 0.1031928, 0.138463, 0.1782238, 0.2129076, 
    0.2011752, 0.1947097, 0.1943326, 0.136516, 0.1532804,
  0.1685132, 0.1608459, 0.1337597, 0.1241888, 0.1633935, 0.1316118, 
    0.05453969, -3.405163e-05, 0.0001173392, -0.0002769723, 0.01146543, 
    0.002411277, 0.09350547, 0.08101275, 0.123542, 0.09902481, 0.1413641, 
    0.1508197, 0.216407, 0.1712435, 0.08315355, 0.08568788, 0.1252236, 
    0.1083581, 0.1520696, 0.1404343, 0.1732645, 0.1612951, 0.1458467,
  0.1656129, 0.1529838, 0.1105159, 0.1088902, 0.07934888, 0.02487697, 
    0.02228128, 0.00619798, 0.005427156, 0.001171185, 0, 4.471211e-05, 
    0.007636532, 0.0525178, 0.02630625, 0.07449984, 0.04715165, 0.06953818, 
    0.04132694, 0.04405182, 0.03999465, 0.05729005, 0.0396077, 0.02629001, 
    0.02894394, 0.06096324, 0.1389215, 0.1641891, 0.1216905,
  0.08980283, 0.08253218, 0.02634044, 0.02801715, 0.01689196, 0.01390343, 
    0.008218837, 0.003228339, 0, 0, -1.43298e-07, -3.320641e-05, 0.01507429, 
    0.05839086, 0.05020027, 0.03507506, 0.08726609, 0.07990457, 0.02781865, 
    0.02920247, 0.01432332, -0.0001168417, -5.555095e-08, -1.343419e-07, 
    0.001579988, 0.001576872, -0.0001931031, 0.05654197, 0.0779997,
  0.006267896, 0.00118321, 0.0003091479, 0.0005585229, 0.00083019, 
    -4.558781e-07, 0, 0, 0, 0, 0, -2.301385e-05, 0.001106163, -6.83419e-05, 
    1.311301e-05, 0.000154635, 0.0003955732, 0.001446502, 6.155554e-05, 
    -1.244118e-05, 4.534602e-07, -7.009169e-06, -1.160569e-05, -4.509025e-06, 
    -5.268419e-05, 1.545571e-05, -5.804306e-05, -0.001421674, 0.01297429,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001930239, 0.03408608, 0.1275216, 
    0.2070957, 0.2160432, 0.0913081, 0.005221148, -0.0003584632, 
    -0.0004661703, 0.01792372, 0.06525484, 0.05151429, 0.07261354, 0.1360433, 
    -0.002439856, 0,
  0.2060618, 0.2222278, 0.2395065, 0.1941703, 0.01028255, 0.02008904, 
    0.09972949, 0.006535805, 0.04567517, 0.05022066, 0.03925691, 0.009194433, 
    0.07272829, 0.2421659, 0.1981515, 0.2020586, 0.2111507, 0.1969524, 
    0.2029102, 0.1572263, 0.09489837, 0.1468688, 0.2823591, 0.2285278, 
    0.3020601, 0.1675355, 0.1012668, 0.1873437, 0.1726722,
  0.2020888, 0.1886021, 0.1862085, 0.2309826, 0.2161816, 0.1596139, 0.206679, 
    0.2251974, 0.2394426, 0.2498057, 0.2349074, 0.2444255, 0.2157485, 
    0.2207297, 0.167353, 0.1432286, 0.1520647, 0.1903323, 0.1712817, 
    0.2208744, 0.2147768, 0.2126236, 0.2088832, 0.2343596, 0.2678794, 
    0.2135452, 0.2617064, 0.2059129, 0.2154507,
  0.1770246, 0.1866553, 0.1950479, 0.1785391, 0.1701755, 0.1571735, 
    0.1171167, 0.1449691, 0.1651454, 0.181272, 0.1733263, 0.1576924, 
    0.1520671, 0.1390792, 0.09108061, 0.1535693, 0.1231615, 0.1212315, 
    0.113497, 0.1281452, 0.1471886, 0.1721883, 0.1809346, 0.09867568, 
    0.09272981, 0.1625109, 0.1142594, 0.1474742, 0.1813084,
  0.05795681, 0.04404665, 0.02709325, 0.06503675, 0.04883144, 0.1096864, 
    0.07611102, 0.07404715, 0.01272363, 0.02132588, 0.03152647, 0.06944363, 
    0.05279738, 0.04495157, 0.1126429, 0.1480031, 0.06679463, 0.04766234, 
    0.09399965, 0.1106592, 0.08631481, 0.05414714, 0.009367866, 0.006902021, 
    0.05314928, 0.06902531, 0.07175022, 0.09316805, 0.0524027,
  0.002085275, 1.667239e-06, 0.09092337, 0.009967767, 0.08034501, 0.1189139, 
    0.07774181, 0.01572469, 0.009706841, 0.02153346, 0.05279307, 0.02075383, 
    0.01537608, 0.1045768, 0.1545101, 0.01336165, 0.132547, 0.1447281, 
    0.1355534, 0.07274947, 0.007511319, 0.000141318, 4.786848e-08, 
    -7.835817e-05, 0.03175182, 0.1661562, 0.0564243, 0.03686932, 0.03492964,
  0.001191663, 0.03931789, 0.03373345, 0.03035016, 0.1689063, 0.05138106, 
    0.003993001, 0.05849679, 0.0007466189, 0.01612298, 0.09659941, 
    0.02538559, 0.05664095, 0.05341933, 0.122895, 0.09028364, 0.1038325, 
    0.06086582, 0.0244961, 0.03252563, 0.0001524231, 0.0007351431, 
    9.692294e-08, 0.00698936, 0.07682774, 0.1497958, 0.02551226, 0.002525234, 
    -9.019677e-05,
  6.671243e-06, 0.02723737, 0.246556, 0.1085451, 0.03499789, 0.02941967, 
    0.03972698, 0.0311822, 0.03729338, 0.04470835, 0.0391285, 0.0725936, 
    0.06109442, 0.07762706, 0.1888225, 0.05480413, 0.02462906, 0.007181376, 
    0.003467353, 0.0007701411, 5.965451e-08, 3.568456e-08, 0.002553942, 
    0.1427473, 0.2913593, 0.1127189, 0.01168967, 0.0002500079, -2.687101e-07,
  0.0001687902, 0.006789234, 0.004952865, 0.005135894, 0.08590338, 
    0.06830543, 0.0763033, 0.05445419, 0.08561061, 0.0876029, 0.01746943, 
    0.01201871, 0.03478679, 0.04798976, 0.06265634, 0.007518599, 0.005035112, 
    0.007029757, 0.01163752, 0.0187626, 0.008567739, 4.822012e-05, 
    0.02243973, 0.0241522, 0.06503975, 0.1823504, 0.01628016, 0.002808307, 
    2.042897e-05,
  -2.483526e-07, 1.744497e-07, 1.132761e-06, 0.001817115, 0.01268978, 
    0.003834021, 0.0006126569, 0.0005420885, 0.001073748, 0.01605017, 
    0.130422, 0.0495497, 0.0439212, 0.03095439, 0.02324908, 0.01159379, 
    0.08296448, 0.06903706, 0.07939475, 0.05394975, 0.05597726, 0.001497625, 
    0.001564323, 0.0007015126, 0.02324855, 0.02540644, 0.02069747, 
    0.01307263, 0.002206796,
  0.01054247, -3.897109e-05, 1.295527e-07, -9.625649e-08, 1.598712e-06, 
    0.00111923, 0.0001071778, 1.300175e-07, 9.302591e-08, 0.000402173, 
    0.04679317, 0.05503323, 0.001131462, 0.02237225, 0.01582876, 0.01408694, 
    0.01511269, 0.04603125, 0.02046694, 0.04114766, 0.02076993, 0.02179344, 
    0.003117513, 0.006921842, 0.007364499, 0.005763409, 0.0005663198, 
    0.03072645, 0.06761616,
  0.02884846, 0.02279182, 0.01635019, 0.01608378, 0.01317161, 0.0422532, 
    0.01861949, 0.0003941256, 0.01661732, 0.200017, 0.1537173, 0.09643944, 
    0.07934254, 0.09625643, 0.1149969, 0.1283637, 0.09378932, 0.114126, 
    0.06911073, 0.02332989, 0.04147832, 0.06979828, 0.08792973, 0.04111941, 
    0.04969459, 0.04133147, 0.042709, 0.051137, 0.04195996,
  0.1397726, 0.08152819, 0.06780376, 0.07513537, 0.09110678, 0.1077452, 
    0.0298565, 0.1428771, 0.08244285, 0.07254484, 0.1080583, 0.1467831, 
    0.1429262, 0.137399, 0.1344468, 0.202523, 0.2408624, 0.2367511, 
    0.1440653, 0.1449491, 0.1369492, 0.1531983, 0.1717302, 0.2156219, 
    0.1810147, 0.2057399, 0.1869678, 0.1229987, 0.153251,
  0.1638245, 0.192191, 0.1229231, 0.1390615, 0.182947, 0.1574497, 0.1673901, 
    0.00118646, 0.0003303649, 0.01805491, 0.02799272, 0.04426061, 0.1267307, 
    0.1424667, 0.2299387, 0.144357, 0.1678707, 0.1701266, 0.2095193, 
    0.1978299, 0.1019578, 0.1159342, 0.1732102, 0.1362449, 0.2036449, 
    0.1704626, 0.1960026, 0.1840185, 0.1628501,
  0.1898097, 0.1901738, 0.1675479, 0.1606664, 0.1762851, 0.1374169, 0.103235, 
    0.1298191, 0.0524403, 0.02952919, 0.003275491, 2.682737e-05, 0.01841701, 
    0.1111308, 0.1165273, 0.1070271, 0.06670066, 0.1109845, 0.06027624, 
    0.09255205, 0.07001543, 0.1052556, 0.0518498, 0.04967064, 0.04476938, 
    0.1140485, 0.196767, 0.2341453, 0.1828864,
  0.164274, 0.1127305, 0.06067882, 0.08142285, 0.07204995, 0.06329852, 
    0.04684932, 0.04986758, 0.006479973, -7.246969e-07, -8.491411e-07, 
    0.004434423, 0.02991968, 0.06002648, 0.06215543, 0.06463081, 0.1127454, 
    0.1043825, 0.04567926, 0.04966283, 0.01810171, 0.003324375, 
    -0.0001292158, -0.0001370106, 0.02833358, 0.008269871, 0.005502163, 
    0.1272842, 0.1469443,
  0.05742806, 0.04416455, 0.03370805, 0.02134502, 0.01529648, 0.001267702, 
    0.002245897, 0.002696595, 0.0005206882, 9.268631e-05, -4.089097e-07, 
    0.0007555897, 0.01223847, 0.01126946, 0.01119411, 0.01534398, 
    0.007934386, 0.02028227, 0.02673428, 0.0154008, 0.009853949, 0.007191568, 
    4.408173e-05, -0.0003976754, 0.001025895, -1.450133e-05, -0.001663457, 
    0.0171747, 0.05775772,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, -8.788774e-09, 0, 0, 0, 0, 0, 0, 0, 0, -1.716951e-07, -7.066027e-07, 
    3.981664e-05, 0.05242685, 0.07766518, 0.2000858, 0.2248446, 0.2801746, 
    0.1925065, 0.09709121, 0.04616995, 0.008765001, 0.0945446, 0.06007354, 
    0.08222957, 0.1019456, 0.1707223, 0.1313384, 0.001020209,
  0.2230891, 0.2943419, 0.3064008, 0.258143, 0.04695129, 0.07855329, 
    0.1158163, 0.02989842, 0.05710024, 0.06389468, 0.05669342, 0.0239595, 
    0.1800342, 0.2290302, 0.2203283, 0.2135009, 0.2138483, 0.2014515, 
    0.240591, 0.1668492, 0.09339938, 0.1915575, 0.3124254, 0.2433016, 
    0.2986298, 0.1668703, 0.1131666, 0.2085096, 0.2023786,
  0.2111514, 0.2001915, 0.1886544, 0.2384966, 0.2335168, 0.1741951, 
    0.2012205, 0.2451352, 0.2595764, 0.2649724, 0.2261766, 0.2565715, 
    0.2250749, 0.2232207, 0.1714404, 0.1343004, 0.1520929, 0.19525, 
    0.1831062, 0.2408512, 0.2331116, 0.244784, 0.2095497, 0.2390858, 
    0.2615341, 0.2244914, 0.2561385, 0.2056336, 0.2407834,
  0.1739439, 0.1819479, 0.1835139, 0.1856771, 0.1617354, 0.1437085, 
    0.1066315, 0.1428829, 0.1570392, 0.1885792, 0.1658704, 0.1568567, 
    0.1474529, 0.1343644, 0.0969574, 0.1399629, 0.1253932, 0.1037929, 
    0.09567429, 0.1263564, 0.1389207, 0.1658211, 0.1589268, 0.09224759, 
    0.08587502, 0.1607537, 0.1093298, 0.1487712, 0.1883052,
  0.05286421, 0.03312124, 0.02135304, 0.0756868, 0.0397326, 0.1073752, 
    0.07072283, 0.06231781, 0.01737122, 0.01719099, 0.03657232, 0.06964932, 
    0.05570763, 0.04440195, 0.1100744, 0.1408168, 0.05592227, 0.04118066, 
    0.08448499, 0.1030133, 0.0801929, 0.05810564, 0.01386486, 0.005779536, 
    0.05039653, 0.06954479, 0.06465953, 0.09225669, 0.04546696,
  0.003467956, 3.13064e-06, 0.08214413, 0.007846261, 0.0793929, 0.1033864, 
    0.06418436, 0.0167992, 0.007808391, 0.01729996, 0.07233377, 0.04026678, 
    0.01469814, 0.1116772, 0.1495472, 0.007951138, 0.1303593, 0.1355684, 
    0.1243044, 0.05374528, 0.005591245, 0.0001408716, 2.079615e-10, 
    -4.0036e-05, 0.03053259, 0.1636989, 0.03943701, 0.02420381, 0.03468985,
  0.000390384, 0.03463623, 0.02962372, 0.03758749, 0.1618715, 0.05474177, 
    0.004935553, 0.05528563, 0.001466714, 0.01313091, 0.09965833, 0.02464224, 
    0.04497587, 0.05554983, 0.1236405, 0.08382068, 0.09035129, 0.06685663, 
    0.02578331, 0.02829969, -3.446628e-06, 0.000349066, 5.84654e-06, 
    0.006161551, 0.07552307, 0.1633354, 0.009755415, 0.0005265338, 
    -3.755209e-05,
  0.0008331239, 0.03931483, 0.2290157, 0.1023094, 0.03698992, 0.03311611, 
    0.04675579, 0.03125906, 0.03449728, 0.04112139, 0.04873792, 0.06421038, 
    0.07636034, 0.07374038, 0.1780178, 0.04621034, 0.02334383, 0.008711999, 
    0.003549056, 0.0002341117, 3.801785e-09, 5.62461e-08, 0.002316395, 
    0.1287612, 0.2970333, 0.1160083, 0.01028754, 0.0002492846, 2.266988e-05,
  0.0193981, 0.01423702, 0.004950304, 0.006928351, 0.07977123, 0.055249, 
    0.07381298, 0.06282545, 0.07762634, 0.09413753, 0.02296423, 0.009647169, 
    0.02284561, 0.03919943, 0.05469793, 0.005570477, 0.00237714, 0.002890708, 
    0.02267917, 0.01792745, 0.007715769, 0.00742919, 0.03262508, 0.02703858, 
    0.05229048, 0.1845625, 0.01736361, 0.005072529, 0.0005429352,
  4.310241e-07, 7.221696e-07, 1.011494e-06, 0.0015173, 0.01394668, 
    0.001944555, 0.0005509983, 0.0001331535, 0.0007913839, 0.01868625, 
    0.1376254, 0.0587376, 0.04372791, 0.03689521, 0.02946811, 0.02234603, 
    0.08766323, 0.06936068, 0.07108655, 0.05943662, 0.05661402, 0.005636015, 
    0.0009156981, 0.0009460637, 0.0329124, 0.02217643, 0.01940851, 
    0.006047044, 0.00100551,
  0.002552878, -1.30078e-06, 1.345683e-07, 8.574672e-09, 1.447302e-06, 
    0.0001714863, 0.0006623869, 2.324837e-07, 7.85226e-08, 0.003100234, 
    0.05864961, 0.05374973, 0.001344299, 0.02025223, 0.01597261, 0.01415597, 
    0.02276164, 0.03805255, 0.02103361, 0.03825759, 0.01188715, 0.02210127, 
    0.003674827, 0.002762686, 0.006385046, 0.00957167, 0.0004009538, 
    0.0311803, 0.04431163,
  0.02100813, 0.0169177, 0.01464287, 0.02269029, 0.01764552, 0.04565268, 
    0.0182381, 0.001142849, 0.04228983, 0.2312192, 0.1752096, 0.08454082, 
    0.07853658, 0.08500902, 0.1146391, 0.103713, 0.08163655, 0.1014429, 
    0.06653917, 0.0117187, 0.03424999, 0.07300492, 0.0724006, 0.03466032, 
    0.04343271, 0.03952901, 0.03667567, 0.05271176, 0.04166208,
  0.1290663, 0.07585588, 0.06499389, 0.09869504, 0.08426169, 0.09528831, 
    0.06624635, 0.1507023, 0.0938565, 0.08051015, 0.114106, 0.1387696, 
    0.1370715, 0.1435017, 0.1565514, 0.2075901, 0.2255049, 0.2432035, 
    0.14894, 0.1396857, 0.1402178, 0.146054, 0.1690126, 0.2114547, 0.1601191, 
    0.1909706, 0.1551245, 0.1054945, 0.1325114,
  0.15662, 0.1813366, 0.1162899, 0.1318716, 0.184265, 0.1658827, 0.2316564, 
    0.0169174, 0.02133735, 0.04864988, 0.0775625, 0.0747842, 0.1615133, 
    0.2044436, 0.2599328, 0.1684341, 0.1762748, 0.1729569, 0.2111934, 
    0.2253036, 0.1191391, 0.1366143, 0.198566, 0.180087, 0.2398216, 0.206332, 
    0.213902, 0.1976153, 0.1600294,
  0.2216404, 0.2081161, 0.2025495, 0.2437281, 0.2787981, 0.2188647, 
    0.1899889, 0.1915743, 0.1405932, 0.1187962, 0.09594724, 0.009165434, 
    0.03113527, 0.1643041, 0.1802889, 0.1676943, 0.1128983, 0.1775073, 
    0.1147538, 0.1365188, 0.1232492, 0.1292137, 0.08470768, 0.06650712, 
    0.1065502, 0.1930222, 0.2501287, 0.2848831, 0.2247715,
  0.2125205, 0.174252, 0.1367583, 0.1919458, 0.1604692, 0.1283813, 
    0.08379856, 0.08827733, 0.04129095, 0.02535884, 0.01398622, 0.02823933, 
    0.05283729, 0.08208062, 0.1106794, 0.1036334, 0.1524853, 0.1571941, 
    0.09720016, 0.06952355, 0.03206267, 0.008618236, 0.01495711, 
    -0.001103141, 0.0676451, 0.02645944, 0.01161698, 0.2070124, 0.2032147,
  0.08419845, 0.08529226, 0.06656706, 0.0528087, 0.04455451, 0.02447699, 
    0.02224307, 0.02804575, 0.03735143, 0.02692476, 0.02836693, 0.02947763, 
    0.0294109, 0.0275972, 0.03557991, 0.06619446, 0.0787669, 0.07274043, 
    0.05859194, 0.05583419, 0.03741981, 0.01892641, 0.006969049, 
    -0.0003266095, 0.005106764, 0.001493777, 0.001396509, 0.04883231, 
    0.1076102,
  7.75249e-06, 2.520815e-06, -2.71086e-06, -7.942534e-06, -1.317421e-05, 
    -1.840588e-05, -2.363756e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -8.080056e-05, -7.556888e-05, -7.033721e-05, -6.510553e-05, 
    -5.987386e-05, -5.464218e-05, -4.94105e-05, 1.193783e-05,
  0.001915041, -9.769019e-05, 0, 0, 0, -5.000024e-05, 0, 0, 0, 0.0001098891, 
    0.000407086, 0.001540173, 0.0005202476, 0.1153923, 0.1054924, 0.2249554, 
    0.205785, 0.2730326, 0.2041428, 0.1601193, 0.1068371, 0.08368233, 
    0.1181803, 0.07040638, 0.09108516, 0.1145724, 0.1791189, 0.1631402, 
    0.05296697,
  0.2567706, 0.3113299, 0.2732869, 0.2544065, 0.1245637, 0.1639177, 
    0.1339491, 0.08446646, 0.08512209, 0.1177075, 0.1067637, 0.06203649, 
    0.24629, 0.1907315, 0.2211521, 0.2127005, 0.2085268, 0.2052453, 
    0.2562844, 0.1428781, 0.09724661, 0.2370836, 0.3236538, 0.2468818, 
    0.2836798, 0.1513017, 0.1361764, 0.2136052, 0.210762,
  0.2296179, 0.2194758, 0.1963085, 0.2432705, 0.2497097, 0.1946547, 
    0.1969226, 0.2448733, 0.2733169, 0.2616619, 0.232547, 0.2479766, 
    0.2341093, 0.2377155, 0.1849972, 0.1421589, 0.1496886, 0.1965729, 
    0.1857544, 0.2593259, 0.256312, 0.272421, 0.2268002, 0.2565153, 
    0.2688631, 0.2228388, 0.2562338, 0.2197052, 0.2604953,
  0.1875121, 0.1760541, 0.1858336, 0.1731296, 0.1605127, 0.1401136, 
    0.1268076, 0.1448961, 0.1562859, 0.1932459, 0.1703542, 0.1452521, 
    0.1448902, 0.134623, 0.1059714, 0.1293807, 0.1238472, 0.1008377, 
    0.09721048, 0.1239303, 0.132467, 0.1692811, 0.176952, 0.0825661, 
    0.08332193, 0.1544467, 0.1176085, 0.1441322, 0.1827333,
  0.05019152, 0.03481495, 0.01919527, 0.09445731, 0.0323003, 0.1015494, 
    0.05572125, 0.05715578, 0.02563731, 0.01855127, 0.04267518, 0.06227855, 
    0.05600444, 0.03886739, 0.1126891, 0.13094, 0.05778198, 0.04138279, 
    0.07593061, 0.09183972, 0.08653328, 0.05367787, 0.005327095, 0.004846812, 
    0.05189839, 0.060816, 0.06235999, 0.0824228, 0.04288857,
  0.005431564, 4.064205e-06, 0.07902893, 0.007799602, 0.07512393, 0.09706667, 
    0.04786456, 0.00941672, 0.004744964, 0.01271019, 0.09999031, 0.06307112, 
    0.02057547, 0.1162719, 0.1400096, 0.01158319, 0.1281582, 0.1248087, 
    0.1148943, 0.0475122, 0.006822255, 0.0001094925, -3.625244e-08, 
    0.0001195057, 0.03055927, 0.1676393, 0.02634347, 0.02131501, 0.0342293,
  0.001140323, 0.039667, 0.03407488, 0.04907115, 0.1629289, 0.05953569, 
    0.007963421, 0.05420969, 0.001123494, 0.01934036, 0.1097326, 0.02362831, 
    0.04296109, 0.06111208, 0.1396215, 0.08526712, 0.08226445, 0.07188923, 
    0.02853426, 0.02692284, 1.4601e-07, -7.421156e-06, 1.178264e-05, 
    0.01037554, 0.08373508, 0.1631606, 0.004757612, 5.110191e-05, 
    -1.629396e-06,
  0.007086505, 0.05612723, 0.2290567, 0.1173894, 0.03658593, 0.03530212, 
    0.05136209, 0.02742959, 0.03557532, 0.05056793, 0.0746682, 0.06835772, 
    0.1074691, 0.0746107, 0.1784417, 0.04067124, 0.02412176, 0.009362347, 
    0.003497829, 0.0002500548, -4.613571e-08, -5.21326e-05, 0.004958996, 
    0.1416083, 0.3176089, 0.1172584, 0.009477045, 0.0001868126, 0.001491102,
  0.08626761, 0.02717864, 0.02505641, 0.00790113, 0.07246835, 0.05814819, 
    0.08450749, 0.06483193, 0.07188341, 0.1105421, 0.03769892, 0.009465137, 
    0.0202075, 0.0405913, 0.048209, 0.005254194, 0.002456439, 0.001457866, 
    0.01643356, 0.01223172, 0.008284502, 0.01747336, 0.05132306, 0.03605868, 
    0.05689184, 0.1865287, 0.02050437, 0.004282911, 0.03089831,
  1.636123e-05, 1.088265e-06, 1.407098e-06, 0.001511915, 0.01798292, 
    0.00106119, 0.0007810573, 5.292999e-05, 0.0011688, 0.02324082, 0.1410557, 
    0.05492418, 0.0490447, 0.04764862, 0.02680197, 0.03730596, 0.08192784, 
    0.08978437, 0.07484286, 0.06517646, 0.05723159, 0.006969599, 0.002242228, 
    0.001366677, 0.03567367, 0.03684989, 0.02444367, 0.00103275, 0.0003051811,
  0.001010238, 2.216731e-07, 6.904635e-08, 1.759219e-08, 1.154e-06, 
    0.0002040856, 4.758842e-05, -7.58091e-07, 4.362336e-08, 0.004164334, 
    0.05270399, 0.03980566, 0.0007471274, 0.01568632, 0.01960146, 0.00649885, 
    0.03744756, 0.03584651, 0.02081602, 0.03053914, 0.009159314, 0.0265442, 
    0.007428984, 0.001822192, 0.005148656, 0.01658141, 0.0001884598, 
    0.02074748, 0.04649427,
  0.01161933, 0.01227438, 0.01366062, 0.02448181, 0.02668804, 0.05112224, 
    0.02205933, 0.001506567, 0.07699631, 0.2441446, 0.1847734, 0.07833187, 
    0.06897795, 0.09217383, 0.09646589, 0.08821017, 0.05977287, 0.0890324, 
    0.06388418, 0.008797864, 0.02430129, 0.07233835, 0.06579984, 0.03108791, 
    0.03704099, 0.0391145, 0.03548168, 0.04951512, 0.03401827,
  0.1172194, 0.06855625, 0.05657554, 0.09850277, 0.08658566, 0.07895985, 
    0.1162941, 0.136952, 0.09107369, 0.07814649, 0.1081794, 0.1362206, 
    0.133305, 0.1509063, 0.1699595, 0.2175603, 0.2244473, 0.2257378, 
    0.1362334, 0.1385227, 0.1513635, 0.1308612, 0.1630481, 0.1980799, 
    0.1532484, 0.1744554, 0.1372337, 0.10874, 0.1197114,
  0.1458124, 0.1523442, 0.1031928, 0.1149052, 0.181326, 0.1759141, 0.2483359, 
    0.07478033, 0.0659896, 0.07106398, 0.07939659, 0.1086947, 0.1885766, 
    0.2372235, 0.2821854, 0.1666859, 0.1692967, 0.1720389, 0.2274554, 
    0.244172, 0.1609122, 0.1529371, 0.2193606, 0.1853849, 0.2427218, 
    0.2144613, 0.2260774, 0.1996686, 0.1543152,
  0.2127171, 0.2133146, 0.2075506, 0.2640748, 0.3029033, 0.2793585, 0.271237, 
    0.3133848, 0.2130541, 0.190762, 0.1628657, 0.07614422, 0.09822071, 
    0.2092354, 0.2222899, 0.1853493, 0.1347811, 0.2020544, 0.1291293, 
    0.2351417, 0.1781778, 0.1602283, 0.1280859, 0.1261138, 0.1813319, 
    0.2686328, 0.2770151, 0.2984843, 0.210806,
  0.2276008, 0.2318456, 0.2587474, 0.2977778, 0.236067, 0.1616738, 0.1262953, 
    0.1639849, 0.1165688, 0.09503211, 0.05324043, 0.07149846, 0.08974291, 
    0.09642524, 0.1719104, 0.1439528, 0.2031612, 0.2015356, 0.1323775, 
    0.08641133, 0.05308891, 0.03929047, 0.04205683, 0.004174648, 0.1135016, 
    0.04022565, 0.03002941, 0.2483782, 0.223231,
  0.09363627, 0.1109546, 0.1099034, 0.09695207, 0.09330089, 0.09898798, 
    0.1117583, 0.1442815, 0.1552894, 0.08812318, 0.06789394, 0.06171868, 
    0.07130059, 0.09268516, 0.1238105, 0.1210234, 0.1044714, 0.08070718, 
    0.08329293, 0.06975323, 0.05439215, 0.0434289, 0.02187462, -0.001160899, 
    0.02440487, 0.009186093, 0.02078856, 0.1024396, 0.1299537,
  0.00481344, 0.004111921, 0.003410402, 0.002708882, 0.002007363, 
    0.001305844, 0.0006043243, 0.002220706, 0.002281747, 0.002342787, 
    0.002403828, 0.002464869, 0.00252591, 0.00258695, 0.006181938, 
    0.007049856, 0.007917775, 0.008785693, 0.009653613, 0.01052153, 
    0.01138945, 0.01128366, 0.01105622, 0.01082878, 0.01060134, 0.0103739, 
    0.01014646, 0.009919016, 0.005374656,
  0.04959956, 0.001794936, -0.0001214653, 0, -0.0001006459, 0.0007143399, 
    0.0005869545, 0.002220551, 0.006211421, 0.003383511, 0.004953875, 
    0.007645709, 0.004335499, 0.1441282, 0.09888919, 0.1987381, 0.2112893, 
    0.2508308, 0.2057544, 0.1853303, 0.1780566, 0.1567513, 0.1454007, 
    0.0951346, 0.1139098, 0.1152399, 0.1818949, 0.1582706, 0.1094899,
  0.2736006, 0.3114718, 0.2632992, 0.2610527, 0.2247355, 0.1914391, 
    0.1269581, 0.1760581, 0.1549485, 0.2030765, 0.1684455, 0.1552032, 
    0.2520928, 0.1728497, 0.2331603, 0.2171565, 0.2187734, 0.2123361, 
    0.2509512, 0.1376651, 0.1407673, 0.2732879, 0.3393484, 0.2989482, 
    0.2930339, 0.1454798, 0.1807475, 0.2180178, 0.2348642,
  0.2464211, 0.2319957, 0.2388359, 0.2809908, 0.2697346, 0.2160367, 
    0.2275217, 0.27242, 0.2951443, 0.2685502, 0.2321407, 0.2578646, 
    0.2613943, 0.2320783, 0.1965152, 0.1394874, 0.1670876, 0.2082164, 
    0.1925962, 0.2752922, 0.2784936, 0.3187499, 0.2425976, 0.2707676, 
    0.2872708, 0.2340871, 0.2561585, 0.2366465, 0.2786546,
  0.1868201, 0.1558455, 0.1778326, 0.1652613, 0.14913, 0.1290251, 0.1361811, 
    0.138096, 0.1525137, 0.165435, 0.1741372, 0.153013, 0.1519943, 0.1352134, 
    0.09774509, 0.1211244, 0.1311263, 0.1023268, 0.08486056, 0.142004, 
    0.1287721, 0.1553347, 0.1477054, 0.08099226, 0.08507663, 0.1566672, 
    0.1185593, 0.1351555, 0.1962691,
  0.04604068, 0.03711671, 0.01697129, 0.09531775, 0.03168959, 0.1009326, 
    0.055571, 0.06024759, 0.02239591, 0.02652068, 0.03634297, 0.06086653, 
    0.05696996, 0.04051645, 0.1053975, 0.121827, 0.05740912, 0.04729009, 
    0.07513648, 0.08462243, 0.08454359, 0.04916135, 0.006038821, 0.003913755, 
    0.06125102, 0.06250492, 0.06584062, 0.08504585, 0.04359084,
  0.0084362, -6.116659e-07, 0.08606531, 0.009758068, 0.07197394, 0.09177247, 
    0.03594498, 0.007658951, 0.005128921, 0.01425315, 0.1095365, 0.08011854, 
    0.01929809, 0.118046, 0.1504547, 0.02241673, 0.1426731, 0.1092942, 
    0.1074678, 0.04967884, 0.01472448, 0.0001108537, -1.383329e-08, 
    0.0006255719, 0.02739093, 0.18456, 0.02490653, 0.0195644, 0.03773857,
  0.0004079675, 0.06055764, 0.04796698, 0.06174971, 0.1907607, 0.07292902, 
    0.009757323, 0.05764107, 0.001756752, 0.02525722, 0.1326637, 0.03416315, 
    0.04356889, 0.05813672, 0.1580893, 0.08792809, 0.09134797, 0.09336919, 
    0.03753779, 0.03102515, 5.563538e-07, 3.315784e-06, 6.020958e-06, 
    0.01098204, 0.1012534, 0.164986, 0.002822291, 6.633611e-05, -8.456878e-06,
  0.005115087, 0.07041773, 0.2518165, 0.1421579, 0.0444063, 0.04991037, 
    0.0588438, 0.0330998, 0.04391981, 0.07140585, 0.1139213, 0.08262023, 
    0.1559138, 0.1041526, 0.1931085, 0.04481163, 0.02576684, 0.009801446, 
    0.004534085, 0.0005583002, 5.172585e-08, 0.001900777, 0.004995291, 
    0.1717486, 0.3529414, 0.1330718, 0.0131687, 0.0001982172, 0.01666569,
  0.178578, 0.0439504, 0.04395741, 0.01254381, 0.07113308, 0.06430423, 
    0.09320278, 0.07719812, 0.09538276, 0.1394293, 0.05086127, 0.017192, 
    0.02720898, 0.04472622, 0.05224527, 0.007026001, 0.005639427, 
    0.002241807, 0.008316392, 0.00624834, 0.01956295, 0.03876843, 0.07746153, 
    0.05765361, 0.07990491, 0.2129204, 0.02656056, 0.005018051, 0.06557956,
  0.0001167052, 1.294323e-06, 7.730629e-05, 0.01452805, 0.01019877, 
    0.001307732, 0.001406714, 0.00045971, 0.001509934, 0.02308355, 0.1615921, 
    0.06236673, 0.06479845, 0.06222602, 0.03207786, 0.03842334, 0.09209663, 
    0.1040761, 0.08331661, 0.06451718, 0.06285628, 0.006029209, 0.004373412, 
    0.001925986, 0.03651201, 0.04693962, 0.02691115, 0.001242215, 0.0007214381,
  -1.428175e-07, 1.464579e-06, 2.525084e-08, 7.9114e-10, 3.853979e-05, 
    0.0004185669, -7.844783e-06, 9.653297e-08, 2.742838e-08, 0.008059436, 
    0.05274612, 0.03820202, 6.868264e-05, 0.01149629, 0.03074098, 
    0.0005561037, 0.04213841, 0.03360186, 0.01153691, 0.02791788, 
    0.005647704, 0.03634864, 0.01583197, 0.003453203, 0.004527868, 
    0.02438821, 0.000417026, 0.04047278, 0.03758383,
  0.009146748, 0.01160375, 0.0142154, 0.02313685, 0.03600984, 0.05837297, 
    0.02192215, 0.002045634, 0.1128869, 0.2704416, 0.1868987, 0.07728967, 
    0.05597311, 0.09019536, 0.0735912, 0.07167579, 0.04829836, 0.08660558, 
    0.0491483, 0.008658865, 0.02058575, 0.0663592, 0.06530353, 0.03024676, 
    0.03560643, 0.04229348, 0.03021226, 0.04820378, 0.03980592,
  0.09842145, 0.0604788, 0.05147108, 0.09313985, 0.08502412, 0.08295631, 
    0.1813863, 0.1045377, 0.08338577, 0.0707385, 0.1018922, 0.1232598, 
    0.1357782, 0.1606697, 0.1706091, 0.2195047, 0.2160583, 0.2148684, 
    0.1234931, 0.1406953, 0.165616, 0.1300427, 0.158467, 0.1914549, 0.145895, 
    0.1567125, 0.1284572, 0.09582617, 0.1132771,
  0.1415569, 0.1321675, 0.09800757, 0.1297267, 0.179494, 0.1782389, 
    0.2269023, 0.1400561, 0.103671, 0.08933081, 0.07708994, 0.09638683, 
    0.1793698, 0.2759375, 0.2812459, 0.1532438, 0.1455342, 0.1544826, 
    0.2301694, 0.2722096, 0.1881779, 0.1513744, 0.2175981, 0.1943659, 
    0.2645898, 0.231395, 0.2374401, 0.1882069, 0.1532124,
  0.1986197, 0.2083263, 0.2006701, 0.2674253, 0.3369696, 0.3013399, 
    0.3177338, 0.3637029, 0.301037, 0.2586621, 0.2036111, 0.1403783, 
    0.217061, 0.2258467, 0.2142231, 0.190398, 0.1476713, 0.1979161, 
    0.1729712, 0.28415, 0.1806442, 0.1811672, 0.1682292, 0.1803998, 
    0.2082341, 0.3125814, 0.2617009, 0.2969015, 0.1832143,
  0.2172055, 0.2079944, 0.2702539, 0.3087641, 0.2282762, 0.1974623, 
    0.1652446, 0.2621543, 0.215567, 0.178322, 0.1065945, 0.1375026, 
    0.1793288, 0.1931894, 0.2057926, 0.2012108, 0.2378674, 0.2053619, 
    0.123674, 0.1201693, 0.08981849, 0.06611606, 0.1225172, 0.03649947, 
    0.1560807, 0.09294388, 0.04910352, 0.2528934, 0.2204458,
  0.1000473, 0.1670968, 0.2088677, 0.2359529, 0.2203982, 0.1706561, 
    0.1845467, 0.2275015, 0.2548655, 0.1831198, 0.1366954, 0.1476174, 
    0.1971284, 0.185497, 0.1786124, 0.1558458, 0.1257859, 0.1102125, 
    0.09538373, 0.07104438, 0.06686694, 0.07471915, 0.0312463, -0.003433376, 
    0.05105214, 0.0189996, 0.05430525, 0.1082886, 0.1299494,
  0.02724427, 0.02612538, 0.02500649, 0.02388761, 0.02276872, 0.02164983, 
    0.02053095, 0.03281726, 0.03407464, 0.03533202, 0.03658941, 0.03784679, 
    0.03910416, 0.04036155, 0.0320925, 0.03377928, 0.03546606, 0.03715284, 
    0.03883962, 0.0405264, 0.04221318, 0.03821925, 0.03639397, 0.0345687, 
    0.03274343, 0.03091816, 0.02909288, 0.02726761, 0.02813938,
  0.09301814, 0.03263973, 0.0141618, 0.00775505, -0.0003862894, 0.006547232, 
    0.01019307, 0.01497733, 0.009885846, 0.008291327, 0.01270079, 0.01263938, 
    0.07786369, 0.1500502, 0.1014694, 0.1826974, 0.2152861, 0.2570546, 
    0.1857178, 0.1728386, 0.2286038, 0.2265991, 0.1653902, 0.1204683, 
    0.1800746, 0.132872, 0.1739141, 0.127113, 0.113629,
  0.3011969, 0.3101723, 0.2825701, 0.2844252, 0.2570318, 0.2006911, 
    0.1522064, 0.2421974, 0.2084968, 0.2688161, 0.2289055, 0.265878, 
    0.2430695, 0.1767196, 0.2543102, 0.213107, 0.2105729, 0.2332719, 
    0.2822112, 0.1508449, 0.1706427, 0.2835493, 0.3288228, 0.3895383, 
    0.3077812, 0.1805383, 0.2328803, 0.2315181, 0.2628951,
  0.242894, 0.2380612, 0.2712786, 0.293689, 0.2797558, 0.2414273, 0.2542526, 
    0.2774314, 0.2911064, 0.2964873, 0.2395444, 0.3008501, 0.271274, 
    0.2397268, 0.2157509, 0.1474029, 0.187275, 0.2110346, 0.2310978, 
    0.3031744, 0.332406, 0.3069549, 0.2623557, 0.2742139, 0.2884788, 
    0.2334208, 0.2564681, 0.2538597, 0.2956857,
  0.2059563, 0.1654802, 0.1970473, 0.1586358, 0.1600449, 0.1443677, 
    0.1285655, 0.1498094, 0.1625844, 0.1767827, 0.1624634, 0.1439661, 
    0.1549632, 0.1315698, 0.1031799, 0.1194493, 0.1198261, 0.09728334, 
    0.07997271, 0.1527153, 0.137044, 0.1513577, 0.1472233, 0.07856591, 
    0.08951336, 0.1510624, 0.1201033, 0.1449577, 0.1876883,
  0.04553302, 0.03937338, 0.01667256, 0.09863759, 0.03148033, 0.1036515, 
    0.05745991, 0.06563754, 0.02426834, 0.03122559, 0.03342743, 0.05484571, 
    0.06745024, 0.04554665, 0.115081, 0.1262913, 0.05772319, 0.04914571, 
    0.08613802, 0.09204611, 0.08772841, 0.04844134, 0.005913612, 0.005538394, 
    0.06015151, 0.05754248, 0.08543268, 0.09064293, 0.0492286,
  0.016347, -1.539085e-05, 0.0868711, 0.01247839, 0.07876807, 0.1108668, 
    0.03171232, 0.0053729, 0.009397263, 0.01519211, 0.1101312, 0.07054041, 
    0.02464233, 0.1234559, 0.1684856, 0.02613582, 0.1523514, 0.1015071, 
    0.1086864, 0.05901663, 0.02764232, 0.000644686, 1.322327e-07, 
    0.001671354, 0.02746873, 0.2119766, 0.02796265, 0.01890511, 0.04087101,
  0.0004068639, 0.09406825, 0.07052944, 0.06722718, 0.1995008, 0.08321069, 
    0.01381525, 0.05971022, 0.001390744, 0.03628617, 0.1528003, 0.04062957, 
    0.05253712, 0.05843536, 0.1746879, 0.09315215, 0.1097129, 0.1103323, 
    0.04863921, 0.03970191, 8.986881e-06, 2.582088e-06, 5.683689e-06, 
    0.006780767, 0.1310533, 0.179219, 0.004021353, 9.66575e-05, 5.981854e-06,
  0.003982325, 0.07759403, 0.3019968, 0.1793505, 0.05694968, 0.06006528, 
    0.06029607, 0.03636876, 0.05673721, 0.0837054, 0.1332287, 0.0872923, 
    0.1898583, 0.1162732, 0.2110744, 0.04979955, 0.03171773, 0.0132687, 
    0.01032318, 0.001275516, 1.537902e-06, 0.01223706, 0.004937928, 
    0.2019313, 0.3743451, 0.1605864, 0.0140503, 0.0004931861, 0.005657848,
  0.1745157, 0.05208634, 0.04782999, 0.02445471, 0.0725547, 0.07238465, 
    0.1074671, 0.09181843, 0.1224149, 0.1749503, 0.06183939, 0.02224249, 
    0.03230973, 0.05891339, 0.05542277, 0.0102759, 0.00392015, 0.003417232, 
    0.01883519, 0.01720915, 0.04225225, 0.04459165, 0.1026457, 0.09040175, 
    0.1124234, 0.2212203, 0.02512001, 0.004124991, 0.05697905,
  4.882372e-05, 5.709568e-06, 0.004090463, 0.05256438, 0.01059408, 
    0.001820466, 0.002559718, 0.001340569, 0.001563942, 0.02425318, 
    0.1795405, 0.07670973, 0.07562833, 0.0667935, 0.032943, 0.03647101, 
    0.08556988, 0.1115507, 0.08648247, 0.06656255, 0.06875652, 0.005511562, 
    0.008234967, 0.003426272, 0.04171783, 0.03450691, 0.01507304, 0.00439423, 
    0.008246265,
  -5.696254e-07, 1.726057e-06, 1.707531e-07, 2.490124e-08, 0.001099199, 
    0.0001240029, -9.633061e-06, 7.283482e-05, 9.855884e-08, 0.0101973, 
    0.05523198, 0.04231076, 5.696565e-05, 0.02187178, 0.03042531, 
    0.0007056777, 0.04260117, 0.03203826, 0.01185892, 0.04337218, 0.00541442, 
    0.05193512, 0.01769855, 0.004977727, 0.006017701, 0.02469391, 
    0.0008724498, 0.02158967, 0.01470677,
  0.008741641, 0.01526237, 0.01324084, 0.02509492, 0.04520068, 0.06036333, 
    0.02543294, 0.007760854, 0.1399114, 0.2767065, 0.1786885, 0.07246336, 
    0.05877443, 0.08495349, 0.07291333, 0.07305133, 0.04421028, 0.08529522, 
    0.03847055, 0.009308755, 0.01985455, 0.05790621, 0.06616861, 0.03112628, 
    0.03812826, 0.04497518, 0.02365729, 0.03308699, 0.02890363,
  0.0904812, 0.05519515, 0.04627933, 0.08811393, 0.07543164, 0.07101969, 
    0.2044532, 0.0603874, 0.07276734, 0.06314468, 0.09771693, 0.1114892, 
    0.1337206, 0.1805282, 0.1834827, 0.2212202, 0.2031032, 0.1983417, 
    0.117947, 0.14298, 0.181332, 0.1426771, 0.1492529, 0.1876173, 0.1337333, 
    0.1346567, 0.1381015, 0.09879535, 0.1142589,
  0.1391191, 0.1240796, 0.09979726, 0.1195048, 0.1744636, 0.174428, 
    0.2147229, 0.1665419, 0.1170066, 0.08525781, 0.06971651, 0.09046128, 
    0.1743588, 0.2771876, 0.2758346, 0.1383745, 0.1282395, 0.1434079, 
    0.2228814, 0.2991445, 0.1880344, 0.1465998, 0.2286389, 0.1923244, 
    0.2688414, 0.2295342, 0.2336939, 0.2027184, 0.1605648,
  0.1862922, 0.2057769, 0.2003917, 0.2669448, 0.3288675, 0.2894252, 
    0.3178734, 0.352609, 0.3185231, 0.2707841, 0.2588903, 0.1505563, 
    0.2538199, 0.2451845, 0.1898936, 0.1883659, 0.1565337, 0.1917274, 
    0.1942782, 0.2937894, 0.1782786, 0.1969339, 0.1830023, 0.1960302, 
    0.2149895, 0.3430719, 0.2594988, 0.2943204, 0.1960928,
  0.2099786, 0.2160482, 0.2875977, 0.2993603, 0.2376887, 0.220828, 0.1800361, 
    0.3304556, 0.3256584, 0.2572147, 0.1402567, 0.2030573, 0.2334412, 
    0.1840663, 0.2187701, 0.1927632, 0.2311244, 0.2076418, 0.119494, 
    0.1234903, 0.09907846, 0.07400818, 0.1116647, 0.08242489, 0.1633905, 
    0.1480953, 0.09260923, 0.2347506, 0.2261533,
  0.1065998, 0.1988685, 0.2066511, 0.2466483, 0.2515803, 0.2085383, 
    0.2119712, 0.2504981, 0.2782916, 0.2320853, 0.1573955, 0.202024, 
    0.2431621, 0.2261743, 0.1757968, 0.1512275, 0.127152, 0.1234908, 
    0.1060037, 0.1089075, 0.1094592, 0.112381, 0.07813279, 0.01717786, 
    0.05375461, 0.02964262, 0.08099056, 0.1047002, 0.1275296,
  0.1008114, 0.09478155, 0.0887517, 0.08272187, 0.07669202, 0.07066218, 
    0.06463234, 0.06664799, 0.07184572, 0.07704344, 0.08224116, 0.08743888, 
    0.09263661, 0.09783433, 0.08079353, 0.08591528, 0.09103704, 0.0961588, 
    0.1012806, 0.1064023, 0.1115241, 0.1414156, 0.137126, 0.1328363, 
    0.1285467, 0.1242571, 0.1199674, 0.1156778, 0.1056353,
  0.09905592, 0.08490454, 0.05452631, 0.0247951, 0.02389254, 0.02076882, 
    0.0219565, 0.01984833, 0.01433607, 0.007411429, 0.007954906, 0.1071372, 
    0.1994262, 0.178446, 0.102117, 0.2095526, 0.210937, 0.2421119, 0.1673959, 
    0.146428, 0.2165809, 0.2406492, 0.1850063, 0.1097985, 0.1727388, 
    0.1416153, 0.1587435, 0.1217222, 0.1006967,
  0.3124442, 0.3228245, 0.3058805, 0.3076741, 0.2518571, 0.1894537, 0.203111, 
    0.2748747, 0.259745, 0.3194672, 0.2763629, 0.2830043, 0.2162874, 
    0.1630789, 0.2630509, 0.2344904, 0.2445496, 0.240802, 0.2885354, 
    0.1933162, 0.2667103, 0.3892543, 0.3571928, 0.3355226, 0.3017241, 
    0.2035859, 0.229402, 0.2780929, 0.293846,
  0.292807, 0.26855, 0.3021977, 0.334518, 0.3360958, 0.2748782, 0.3102134, 
    0.3656082, 0.3713186, 0.3264778, 0.250734, 0.2765241, 0.2735112, 
    0.245249, 0.2107616, 0.1498845, 0.1798814, 0.2322824, 0.2331729, 
    0.3480989, 0.3297604, 0.3267395, 0.2769932, 0.3156343, 0.2884748, 
    0.2544232, 0.2893163, 0.2796043, 0.3396983,
  0.2176937, 0.1779957, 0.2035272, 0.1704869, 0.18332, 0.1288852, 0.1445182, 
    0.1685968, 0.1593716, 0.1816586, 0.184292, 0.152091, 0.1589482, 
    0.1276733, 0.09468679, 0.131272, 0.1202514, 0.1043779, 0.1049194, 
    0.1689628, 0.1478883, 0.1511398, 0.146705, 0.08374407, 0.09771562, 
    0.1429588, 0.1247395, 0.1345188, 0.2005482,
  0.05598001, 0.04442252, 0.01226245, 0.09899732, 0.0355961, 0.1153284, 
    0.06142581, 0.06602004, 0.03733891, 0.03550073, 0.03768443, 0.05542466, 
    0.06738259, 0.05058669, 0.1297105, 0.1293003, 0.06618156, 0.05707593, 
    0.09139542, 0.09606391, 0.09663709, 0.05805593, 0.009676209, 0.004185994, 
    0.05443831, 0.06145042, 0.1049246, 0.0998293, 0.05655706,
  0.01476082, -1.359522e-06, 0.09507436, 0.009981577, 0.07860905, 0.1237836, 
    0.02959133, 0.004815521, 0.01287109, 0.0088876, 0.08800759, 0.03656679, 
    0.03666652, 0.1297756, 0.1524935, 0.03910409, 0.1714848, 0.1120849, 
    0.1158356, 0.06703068, 0.03689483, 0.002465206, 1.664616e-07, 
    0.001215923, 0.03407807, 0.2284349, 0.03389963, 0.02216993, 0.04363164,
  0.0002971548, 0.1037845, 0.08814146, 0.06518668, 0.1726362, 0.07801022, 
    0.02396385, 0.05753875, 0.001494275, 0.02787206, 0.1453163, 0.03942052, 
    0.04250652, 0.05577157, 0.1379249, 0.09069389, 0.1037177, 0.1030836, 
    0.05003317, 0.04213232, 0.0008685606, 1.124067e-06, 3.324473e-06, 
    0.001383677, 0.126062, 0.2105713, 0.006474369, 3.405235e-07, 5.682782e-07,
  8.109084e-05, 0.05996313, 0.3479705, 0.1856688, 0.04361574, 0.05441065, 
    0.05342674, 0.03503946, 0.04932518, 0.06464285, 0.1118478, 0.06216753, 
    0.1693342, 0.08551356, 0.167808, 0.04177859, 0.02651708, 0.01963925, 
    0.01232695, 0.001852263, 4.079015e-05, 0.02053113, 0.0006395759, 
    0.2245924, 0.3483744, 0.1883263, 0.01419917, 0.0002168526, 0.0001671452,
  0.08475684, 0.05295902, 0.05505874, 0.02915673, 0.06701046, 0.06872693, 
    0.1021629, 0.1011326, 0.1363869, 0.2003553, 0.0636511, 0.01905401, 
    0.02014786, 0.04730131, 0.04764879, 0.01802107, 0.004696974, 0.01054022, 
    0.03375913, 0.01247946, 0.03087742, 0.02699734, 0.1382379, 0.09969794, 
    0.147805, 0.2212785, 0.02875163, 0.005935516, 0.01445839,
  -0.0001706467, 4.638856e-06, 0.001811682, 0.1271299, 0.008255095, 
    0.00652462, 0.003235026, 0.001444721, 0.00338031, 0.02069689, 0.1883963, 
    0.07448791, 0.06418692, 0.05826284, 0.03168627, 0.04055283, 0.08279598, 
    0.1098738, 0.0943075, 0.0719454, 0.07747313, 0.007100163, 0.008227208, 
    0.005060748, 0.03775311, 0.03650701, 0.008511379, 0.004647348, 0.01127783,
  2.018869e-06, 7.764358e-07, 5.357035e-07, 1.28137e-07, 0.00300887, 
    7.472068e-06, -1.29951e-06, 5.419973e-05, 8.558867e-07, 0.007995226, 
    0.07203174, 0.04203819, 0.003590279, 0.02265472, 0.0291285, 0.001494032, 
    0.05421109, 0.03552264, 0.01518792, 0.02980823, 0.003169748, 0.06898914, 
    0.01836556, 0.007393795, 0.009937446, 0.03209538, 0.002168196, 
    0.01177344, 0.001510044,
  0.008849616, 0.01718961, 0.009673556, 0.02934531, 0.05653324, 0.05801027, 
    0.02689382, 0.01329379, 0.1563097, 0.2701609, 0.1830143, 0.07614808, 
    0.06332605, 0.08149755, 0.08591804, 0.07746832, 0.04472205, 0.09283903, 
    0.03163752, 0.01419231, 0.02497172, 0.05561223, 0.06904052, 0.03226959, 
    0.04564378, 0.04576553, 0.02649673, 0.02958084, 0.01841807,
  0.07646427, 0.0471184, 0.03918013, 0.08965196, 0.06122278, 0.06291427, 
    0.2137627, 0.03186825, 0.05449125, 0.06605566, 0.09235749, 0.1021413, 
    0.1273249, 0.1833925, 0.1950361, 0.2159457, 0.1926222, 0.1946353, 
    0.1221971, 0.1441159, 0.1968695, 0.1299495, 0.1429137, 0.1864287, 
    0.1256049, 0.1368447, 0.1451996, 0.0993543, 0.1232901,
  0.1309159, 0.108955, 0.09408481, 0.1190433, 0.1592163, 0.1653314, 
    0.1843753, 0.1822049, 0.1081064, 0.08532556, 0.07078695, 0.08613973, 
    0.1667766, 0.2713705, 0.2996373, 0.1232264, 0.1231631, 0.1568532, 
    0.230287, 0.2867983, 0.1938338, 0.1500479, 0.2386548, 0.2021589, 
    0.2747431, 0.220429, 0.2442409, 0.204837, 0.1586191,
  0.1696771, 0.2116362, 0.2106076, 0.2795767, 0.3527115, 0.2836719, 
    0.3311878, 0.3793893, 0.3158619, 0.2613905, 0.2969898, 0.1554253, 
    0.276228, 0.2605728, 0.1695265, 0.1756776, 0.158545, 0.1955964, 
    0.2132261, 0.275109, 0.1811647, 0.2176654, 0.1934336, 0.2067896, 
    0.2132691, 0.3314691, 0.2559236, 0.2838558, 0.2066544,
  0.210077, 0.2212573, 0.2981486, 0.3285398, 0.2547231, 0.2205613, 0.2186792, 
    0.357241, 0.3462096, 0.3138054, 0.1752945, 0.2238667, 0.2049451, 
    0.1689771, 0.2339728, 0.2095549, 0.2308143, 0.2151869, 0.1194698, 
    0.1283887, 0.1121936, 0.07677191, 0.1147369, 0.1027093, 0.1494142, 
    0.1993225, 0.1718734, 0.2251629, 0.2170385,
  0.1294897, 0.2004186, 0.1959076, 0.2621083, 0.2453681, 0.204086, 0.2036953, 
    0.2623389, 0.302451, 0.2737285, 0.2052528, 0.2318241, 0.2225479, 
    0.2313114, 0.1900016, 0.1573832, 0.1236098, 0.1503151, 0.151413, 
    0.1696297, 0.1548191, 0.1625616, 0.1136862, 0.05691607, 0.06176864, 
    0.04208981, 0.08774204, 0.09870079, 0.1314513,
  0.1676785, 0.1657333, 0.163788, 0.1618427, 0.1598975, 0.1579522, 0.1560069, 
    0.1463156, 0.1540446, 0.1617735, 0.1695025, 0.1772315, 0.1849604, 
    0.1926894, 0.2004943, 0.1998763, 0.1992583, 0.1986403, 0.1980222, 
    0.1974042, 0.1967862, 0.1995052, 0.1943396, 0.1891739, 0.1840083, 
    0.1788426, 0.1736769, 0.1685113, 0.1692348,
  0.10292, 0.09203213, 0.1195052, 0.04466872, 0.04938931, 0.05752005, 
    0.0556667, 0.03749003, 0.02077091, 0.007119037, 0.04725532, 0.1810979, 
    0.2326391, 0.2120711, 0.140119, 0.2636357, 0.2612145, 0.2452908, 
    0.1888968, 0.1863132, 0.2471626, 0.2886763, 0.1991669, 0.1581142, 
    0.1755784, 0.155019, 0.1520516, 0.12277, 0.08929881,
  0.3371108, 0.3395544, 0.300754, 0.3500569, 0.2663145, 0.18685, 0.2609376, 
    0.2918361, 0.2854531, 0.3308845, 0.2753934, 0.2733243, 0.2072572, 
    0.175466, 0.278513, 0.2971583, 0.2554456, 0.2803805, 0.3527459, 
    0.2230816, 0.3092793, 0.3726049, 0.3551026, 0.3649643, 0.2773937, 
    0.1711243, 0.2041035, 0.300713, 0.391556,
  0.2845515, 0.3293489, 0.3218725, 0.2850049, 0.3065093, 0.2705475, 
    0.3103419, 0.3341926, 0.3424475, 0.310816, 0.2564827, 0.3293346, 
    0.2714118, 0.2307551, 0.2091447, 0.1683641, 0.1763258, 0.2383768, 
    0.2599168, 0.337061, 0.321989, 0.2826866, 0.2800208, 0.2968683, 
    0.2794935, 0.2633546, 0.3116359, 0.2925555, 0.3722558,
  0.2262591, 0.1938701, 0.2056173, 0.1728779, 0.174041, 0.1469464, 0.1463964, 
    0.1715909, 0.1720177, 0.184414, 0.1816548, 0.1595796, 0.1731904, 
    0.1304986, 0.1096932, 0.1320337, 0.1122079, 0.110621, 0.1104259, 
    0.1775871, 0.1587689, 0.1648294, 0.1647359, 0.09625645, 0.09383282, 
    0.1401057, 0.1193668, 0.1315004, 0.2177396,
  0.05865524, 0.05965878, 0.01218128, 0.0981323, 0.04818422, 0.1249932, 
    0.07268877, 0.06796378, 0.05204386, 0.03190485, 0.04099948, 0.05111365, 
    0.05956678, 0.05005884, 0.1492458, 0.1238313, 0.07968247, 0.06616429, 
    0.09437255, 0.1007905, 0.1001906, 0.05946937, 0.01722451, 0.00389758, 
    0.0439067, 0.06047388, 0.1283296, 0.10708, 0.06015623,
  0.01374761, -7.881246e-06, 0.1176942, 0.01262528, 0.06361642, 0.1235436, 
    0.02635434, 0.004253452, 0.0134504, 0.01154908, 0.04744096, 0.01776849, 
    0.05016124, 0.1092812, 0.1255772, 0.04927587, 0.1577042, 0.1108474, 
    0.1008066, 0.067622, 0.04155488, 0.003683374, -8.933112e-07, 
    0.0006360685, 0.02990449, 0.1869117, 0.03633904, 0.02456264, 0.04327241,
  0.001275856, 0.08744884, 0.08970998, 0.06674785, 0.1415899, 0.07259543, 
    0.03479698, 0.05217389, 0.0006925181, 0.01330109, 0.1229235, 0.03105798, 
    0.03162873, 0.04986347, 0.1059474, 0.07327966, 0.08219047, 0.07969101, 
    0.04739891, 0.04360312, 0.008085988, 4.665446e-07, 2.178735e-06, 
    0.0003251733, 0.110324, 0.2219059, 0.01321757, 0.000996538, 1.595383e-05,
  8.803838e-05, 0.02518415, 0.3788609, 0.119302, 0.03172092, 0.04664897, 
    0.04678443, 0.03419636, 0.04014302, 0.04758292, 0.09069853, 0.04547638, 
    0.151977, 0.07298061, 0.1392567, 0.03803599, 0.02554725, 0.01862304, 
    0.01794786, 0.003776921, 0.0002156626, 0.006836445, 0.000372072, 
    0.1631181, 0.2373492, 0.1583088, 0.01593197, 0.0007742461, 5.143719e-06,
  0.02338091, 0.04116008, 0.03375852, 0.04342563, 0.05875214, 0.06508075, 
    0.0973575, 0.09983149, 0.1243898, 0.1869876, 0.05957507, 0.01640102, 
    0.01360923, 0.03549935, 0.04235915, 0.02520453, 0.004840803, 0.009544805, 
    0.02926451, 0.01326853, 0.02428607, 0.0196712, 0.156668, 0.09566654, 
    0.1403784, 0.2114082, 0.03388447, 0.008951705, 0.001315214,
  -8.699333e-05, 2.565627e-06, 0.0001584416, 0.2177455, 0.00962574, 
    0.01747826, 0.003888133, 0.001945803, 0.007038458, 0.02707396, 0.191315, 
    0.07432104, 0.05141269, 0.05015128, 0.03053706, 0.042078, 0.06961773, 
    0.100737, 0.0828919, 0.07451741, 0.07965979, 0.007202705, 0.01131262, 
    0.009872602, 0.02956959, 0.01747139, 0.002058449, 0.001195004, 0.002410239,
  1.869344e-06, 4.49701e-07, 1.8346e-07, 7.027129e-06, 0.007217078, 
    9.550629e-06, -8.731226e-07, 0.0003925974, 3.619403e-05, 0.009617076, 
    0.1361576, 0.02955134, 0.007779559, 0.01756744, 0.0278023, 0.002867265, 
    0.06904366, 0.03554798, 0.01100421, 0.01500285, 0.0007584852, 0.08405166, 
    0.01905368, 0.01688325, 0.01454272, 0.04355557, 0.004959908, 0.00381896, 
    0.0008920514,
  0.003410585, 0.02039103, 0.01077758, 0.0321633, 0.06622869, 0.05505402, 
    0.02959043, 0.01593366, 0.1605225, 0.2571114, 0.1576658, 0.07649127, 
    0.08036891, 0.0895125, 0.0925246, 0.08911209, 0.05590896, 0.1053279, 
    0.03458585, 0.01927249, 0.02753823, 0.05962904, 0.07006866, 0.03838957, 
    0.05858049, 0.04847686, 0.03528871, 0.02025205, 0.00465995,
  0.07462157, 0.04334373, 0.03616388, 0.09701706, 0.05983765, 0.05976702, 
    0.2196, 0.0203198, 0.0392985, 0.07653475, 0.09215851, 0.0995858, 
    0.1251196, 0.2105483, 0.1876178, 0.209442, 0.1864179, 0.1894675, 
    0.1352034, 0.1491138, 0.1997368, 0.1273783, 0.1507779, 0.185759, 
    0.127744, 0.1383832, 0.1556629, 0.1027345, 0.1366367,
  0.1301746, 0.1015028, 0.09577876, 0.1295733, 0.1531334, 0.1803152, 
    0.183256, 0.200162, 0.1000052, 0.07430781, 0.06647841, 0.08647116, 
    0.1604588, 0.2816396, 0.3308163, 0.1132783, 0.118341, 0.1531446, 
    0.245392, 0.2870536, 0.1928776, 0.1549344, 0.2400668, 0.1937487, 
    0.2866933, 0.2195717, 0.2466099, 0.2158061, 0.1598861,
  0.1668607, 0.2199432, 0.240083, 0.2898679, 0.3612912, 0.3060749, 0.3509378, 
    0.395799, 0.2954351, 0.2713922, 0.3071451, 0.152539, 0.2877972, 0.284131, 
    0.1818047, 0.1829829, 0.1717439, 0.1950332, 0.2273645, 0.2619005, 
    0.2043048, 0.2270978, 0.2017027, 0.2097303, 0.2040827, 0.3304883, 
    0.2545359, 0.2902061, 0.2007704,
  0.2190419, 0.2279159, 0.3255684, 0.3460167, 0.2799055, 0.23073, 0.2374208, 
    0.3760686, 0.3552866, 0.3319428, 0.1829699, 0.2234907, 0.1958607, 
    0.1827489, 0.237466, 0.2132481, 0.2546686, 0.2299791, 0.1207642, 0.1291, 
    0.1227632, 0.1033374, 0.1281289, 0.1211484, 0.1349585, 0.3040266, 
    0.2637348, 0.2409388, 0.2290153,
  0.134411, 0.2148667, 0.2088657, 0.2734603, 0.2409749, 0.2167502, 0.2053973, 
    0.259568, 0.3031209, 0.2882547, 0.2096755, 0.2391182, 0.2201862, 
    0.2338927, 0.217221, 0.1821224, 0.1567461, 0.1820141, 0.1772688, 
    0.215969, 0.1734822, 0.1886178, 0.1465418, 0.07586724, 0.06987528, 
    0.04668071, 0.0911348, 0.09008123, 0.1353263,
  0.1693149, 0.1695054, 0.1696959, 0.1698863, 0.1700768, 0.1702673, 
    0.1704577, 0.1716127, 0.180393, 0.1891734, 0.1979537, 0.2067341, 
    0.2155144, 0.2242948, 0.2328371, 0.2285156, 0.224194, 0.2198725, 
    0.2155509, 0.2112294, 0.2069079, 0.1961189, 0.1914696, 0.1868203, 
    0.1821711, 0.1775218, 0.1728725, 0.1682232, 0.1691626,
  0.1071582, 0.09924354, 0.1471616, 0.1406231, 0.1042327, 0.1383648, 
    0.1081229, 0.06446987, 0.01941042, 0.01094219, 0.1395079, 0.2124499, 
    0.2349432, 0.23957, 0.1237361, 0.2374197, 0.2169189, 0.2208537, 
    0.1824396, 0.1758993, 0.2872382, 0.3080582, 0.1988677, 0.1221899, 
    0.1493928, 0.135861, 0.1231392, 0.1377397, 0.08392166,
  0.3517995, 0.3723667, 0.3374555, 0.4239787, 0.2975188, 0.2021704, 
    0.2720383, 0.336106, 0.2959795, 0.3318118, 0.2897985, 0.2522107, 
    0.1970869, 0.1965195, 0.3184868, 0.367556, 0.2994811, 0.2766952, 
    0.4110193, 0.2611093, 0.3214484, 0.3541768, 0.3762417, 0.3878842, 
    0.2443219, 0.1681952, 0.2662061, 0.3848321, 0.4597878,
  0.3015884, 0.3747337, 0.3721571, 0.3366806, 0.3511771, 0.3195075, 
    0.3581817, 0.407142, 0.3866438, 0.3457979, 0.2975084, 0.3341874, 
    0.2793837, 0.2235831, 0.2297048, 0.1830762, 0.1955381, 0.282432, 
    0.311424, 0.360797, 0.342517, 0.2752864, 0.2663184, 0.3015116, 0.2949476, 
    0.2986946, 0.3028299, 0.2808886, 0.3368741,
  0.2241708, 0.1927198, 0.2246393, 0.1940362, 0.1756292, 0.1505565, 
    0.1713637, 0.1759928, 0.1812641, 0.2048276, 0.2158016, 0.158718, 
    0.1699954, 0.1408797, 0.1263364, 0.1420766, 0.116185, 0.1198957, 
    0.1383909, 0.1862063, 0.1726449, 0.1817453, 0.1659772, 0.1173978, 
    0.09228605, 0.1588354, 0.1171357, 0.1472871, 0.2145549,
  0.06890556, 0.05950484, 0.0207912, 0.1016889, 0.04683067, 0.1321613, 
    0.07176993, 0.0858428, 0.07174772, 0.04131129, 0.03333939, 0.05083562, 
    0.05539586, 0.0532826, 0.1726711, 0.1092428, 0.07555205, 0.06320974, 
    0.08521628, 0.09650309, 0.1004571, 0.06680193, 0.02055727, 0.003728554, 
    0.03320112, 0.05897936, 0.114914, 0.1075159, 0.05286299,
  0.01996988, -6.673333e-06, 0.1168855, 0.01928711, 0.05394322, 0.1201389, 
    0.02264553, 0.002180688, 0.01089968, 0.02469033, 0.02998561, 0.008817664, 
    0.04669901, 0.08524162, 0.1164012, 0.05916433, 0.1481231, 0.09692828, 
    0.07495105, 0.06657183, 0.0450038, 0.00398816, -6.349863e-06, 
    0.0003645565, 0.02010725, 0.1723761, 0.02981273, 0.03063808, 0.04302415,
  0.001350317, 0.0755422, 0.07887275, 0.07027565, 0.122618, 0.06841844, 
    0.03583674, 0.058144, 0.0009946248, 0.009497101, 0.1095759, 0.03055805, 
    0.03061716, 0.04048177, 0.09230787, 0.06367489, 0.06822477, 0.06319766, 
    0.05027739, 0.05655638, 0.02851317, 4.104633e-05, 1.586034e-06, 
    3.619342e-05, 0.1119066, 0.2007925, 0.02362931, 0.008061121, 0.001099704,
  2.851869e-06, 0.006592555, 0.2627721, 0.08365003, 0.02614592, 0.04092944, 
    0.05020192, 0.03314069, 0.03676412, 0.03899019, 0.07960767, 0.03539139, 
    0.1215672, 0.06372206, 0.1255099, 0.04215033, 0.04036448, 0.01800247, 
    0.0203453, 0.01469495, 0.0003483722, 0.001834045, 0.0002238087, 
    0.1547684, 0.1943539, 0.1354249, 0.02171429, 0.001859251, 1.525255e-06,
  0.006848336, 0.02773246, 0.01652535, 0.07363932, 0.0571185, 0.06517769, 
    0.09086919, 0.1051724, 0.1306008, 0.1979336, 0.05093197, 0.01468261, 
    0.01290479, 0.0368275, 0.04741509, 0.04556289, 0.004845676, 0.01299837, 
    0.03059321, 0.01017958, 0.02125599, 0.02103414, 0.1452761, 0.0918977, 
    0.1386354, 0.195055, 0.04476106, 0.0120312, 0.001236055,
  -1.081691e-05, 9.462683e-07, 7.77878e-06, 0.258495, 0.01358089, 0.02224452, 
    0.004847812, 0.002787316, 0.01819376, 0.03848168, 0.2029288, 0.0764317, 
    0.0481444, 0.04723793, 0.03736156, 0.04951169, 0.06684904, 0.09028587, 
    0.07819151, 0.07958224, 0.0784793, 0.009177541, 0.02551908, 0.01922212, 
    0.03266529, 0.008060837, -3.296304e-05, 1.15173e-05, 6.093962e-05,
  1.458807e-06, 2.921901e-07, 9.348556e-08, 0.0005397688, 0.009484353, 
    9.748192e-06, -4.110815e-06, 0.001233345, 0.003496371, 0.0172793, 
    0.1653951, 0.0286518, 0.01262944, 0.02795191, 0.02770351, 0.005463805, 
    0.07890633, 0.03120937, 0.007462921, 0.007445018, 0.0001521808, 
    0.09634909, 0.02006077, 0.0230132, 0.02177859, 0.04732509, 0.01099456, 
    0.002775691, 0.0006825489,
  0.006407327, 0.0160538, 0.02865817, 0.03410799, 0.0781469, 0.05723093, 
    0.0202059, 0.01663357, 0.1558023, 0.2470475, 0.1604691, 0.07708864, 
    0.08868378, 0.09913917, 0.1052857, 0.107976, 0.08302457, 0.1262951, 
    0.04382083, 0.02512069, 0.03449665, 0.07214418, 0.06941689, 0.04940604, 
    0.06188401, 0.04902441, 0.04080181, 0.02353062, 0.001636379,
  0.07466142, 0.03844171, 0.03736507, 0.1178097, 0.06899767, 0.07764781, 
    0.2234396, 0.01264229, 0.02651563, 0.07889201, 0.09633108, 0.105101, 
    0.1415295, 0.2465869, 0.1866003, 0.2066005, 0.1776437, 0.1886644, 
    0.1506085, 0.152813, 0.2151621, 0.1102119, 0.150555, 0.1758099, 
    0.1417693, 0.1502466, 0.1685763, 0.1421117, 0.1558092,
  0.140235, 0.08962356, 0.1095867, 0.16269, 0.191187, 0.2084651, 0.1822506, 
    0.2085749, 0.08542633, 0.06542783, 0.06014142, 0.09343905, 0.1670603, 
    0.3108028, 0.3373655, 0.1270385, 0.1206276, 0.1814322, 0.255078, 
    0.2997032, 0.1939268, 0.140468, 0.2077536, 0.2067251, 0.2926421, 
    0.2233626, 0.2771036, 0.2156366, 0.1624135,
  0.1756676, 0.212389, 0.2402002, 0.3459284, 0.4217348, 0.3312824, 0.3708764, 
    0.4357609, 0.30409, 0.2909722, 0.3044378, 0.1479408, 0.2914592, 
    0.3216541, 0.1907823, 0.2223983, 0.1724281, 0.2033854, 0.2347513, 
    0.2578747, 0.2067246, 0.2266194, 0.1900555, 0.2076155, 0.1903952, 
    0.3341766, 0.2719997, 0.2972764, 0.2033937,
  0.2308591, 0.2389098, 0.3368942, 0.3610806, 0.2823232, 0.2263535, 
    0.2767922, 0.4030108, 0.3707032, 0.3342835, 0.1922248, 0.2283563, 
    0.1830257, 0.1973939, 0.2401424, 0.2185894, 0.2842364, 0.2342621, 
    0.1260867, 0.1493251, 0.1402785, 0.1400984, 0.1316018, 0.109753, 
    0.1203326, 0.3777849, 0.3108191, 0.2536495, 0.2365302,
  0.1543795, 0.2523473, 0.2327149, 0.2743475, 0.248639, 0.2354967, 0.2233211, 
    0.2815939, 0.317842, 0.3035447, 0.2435644, 0.262109, 0.2260016, 
    0.2253143, 0.2124072, 0.1780185, 0.1647869, 0.172144, 0.1808518, 
    0.2321926, 0.1834509, 0.1971232, 0.1569842, 0.1028584, 0.07586631, 
    0.04222728, 0.1008721, 0.1068754, 0.1598893,
  0.1760083, 0.1774321, 0.1788559, 0.1802796, 0.1817034, 0.1831272, 0.184551, 
    0.178435, 0.1877867, 0.1971384, 0.2064901, 0.2158418, 0.2251935, 
    0.2345452, 0.2450214, 0.2387643, 0.2325073, 0.2262502, 0.2199932, 
    0.2137361, 0.207479, 0.1987687, 0.1942503, 0.1897319, 0.1852135, 
    0.1806951, 0.1761767, 0.1716582, 0.1748692,
  0.1221607, 0.1196064, 0.1527011, 0.233933, 0.1645073, 0.2037706, 0.1254239, 
    0.05907262, 0.02351676, 0.1083462, 0.1734637, 0.2226774, 0.2473239, 
    0.2422644, 0.1844774, 0.2451516, 0.1806948, 0.1946422, 0.1788433, 
    0.1782825, 0.2959976, 0.3346127, 0.1934941, 0.0989123, 0.1276679, 
    0.1250483, 0.09568319, 0.1346912, 0.1256239,
  0.333072, 0.3731117, 0.3240893, 0.3786148, 0.3249915, 0.2215552, 0.2735221, 
    0.3754343, 0.3134118, 0.3528859, 0.2855099, 0.2272401, 0.1718939, 
    0.2021299, 0.319575, 0.3779858, 0.3288021, 0.3352707, 0.4095984, 
    0.1898492, 0.2752485, 0.3412299, 0.3880885, 0.3869091, 0.2212934, 
    0.1458098, 0.2162169, 0.3341829, 0.388237,
  0.2864866, 0.3499463, 0.3678471, 0.3334471, 0.3527687, 0.2973816, 
    0.3376519, 0.348889, 0.3709383, 0.3383651, 0.2766887, 0.3409792, 
    0.2848384, 0.2492956, 0.2397517, 0.1893929, 0.2053915, 0.2916879, 
    0.3485646, 0.3717336, 0.3111893, 0.2788627, 0.2853127, 0.2866473, 
    0.3385271, 0.3122362, 0.3057794, 0.2940711, 0.3010384,
  0.2478257, 0.2237785, 0.2397263, 0.2061474, 0.1811986, 0.1724138, 0.178724, 
    0.1846035, 0.1934313, 0.2488052, 0.2247386, 0.1813269, 0.1898877, 
    0.1485212, 0.1331782, 0.1366547, 0.1136832, 0.1219164, 0.1619388, 
    0.2089927, 0.2073845, 0.1996951, 0.1765013, 0.1465466, 0.07818864, 
    0.1316493, 0.1168234, 0.1735712, 0.2175517,
  0.066744, 0.06891022, 0.03220502, 0.1182571, 0.05043673, 0.1269731, 
    0.06213812, 0.1053783, 0.0833139, 0.05332204, 0.02763098, 0.05406917, 
    0.06564554, 0.05624654, 0.1717525, 0.1019353, 0.06072484, 0.06770015, 
    0.07941064, 0.09228328, 0.1075996, 0.07792133, 0.03310334, 0.003777812, 
    0.01773822, 0.06088357, 0.1082149, 0.08661767, 0.05216081,
  0.02279018, -2.831054e-05, 0.09818682, 0.02455025, 0.05848323, 0.1129742, 
    0.03290387, 0.004408347, 0.007724534, 0.01724356, 0.01611704, 
    0.006657435, 0.04313367, 0.06786512, 0.1271926, 0.06306583, 0.1536338, 
    0.1092947, 0.08585958, 0.06205507, 0.04911302, 0.009728868, 
    -3.186241e-05, 0.0001993428, 0.01906194, 0.164216, 0.02864249, 
    0.03936545, 0.05045385,
  0.006396739, 0.04836263, 0.09258398, 0.07083189, 0.1176315, 0.06135612, 
    0.04530349, 0.05979659, 0.006203666, 0.01017951, 0.09456626, 0.02345856, 
    0.03761432, 0.03980083, 0.08239206, 0.05747545, 0.06019139, 0.05107303, 
    0.05129041, 0.06085413, 0.07100776, 0.006473081, 7.618353e-07, 
    -2.054476e-05, 0.1179296, 0.1874839, 0.03384653, 0.02799235, 0.0116858,
  1.260371e-06, 0.001086111, 0.2098849, 0.06360886, 0.02354621, 0.03541186, 
    0.05199394, 0.03221636, 0.03470375, 0.03757445, 0.07599805, 0.03010051, 
    0.1029346, 0.05398937, 0.1139746, 0.04326609, 0.04869941, 0.02208797, 
    0.02312453, 0.02340559, 0.003858834, 0.001747999, 0.0003111504, 
    0.1481981, 0.1606881, 0.1070545, 0.02940447, 0.001625599, -2.006352e-06,
  0.001652286, 0.01433604, 0.009176201, 0.05846147, 0.05716722, 0.06114792, 
    0.08530729, 0.1044748, 0.1517708, 0.1937166, 0.04459249, 0.01506251, 
    0.01345978, 0.03883314, 0.04856379, 0.04955168, 0.00690691, 0.01606974, 
    0.03127085, 0.0174211, 0.02673372, 0.02909141, 0.1127126, 0.08042783, 
    0.1343706, 0.1790991, 0.04281453, 0.01636397, 0.00130251,
  -3.935466e-06, 1.975927e-07, 1.241544e-06, 0.1493004, 0.01958396, 
    0.0265364, 0.008626243, 0.003527922, 0.02540965, 0.04510904, 0.2174031, 
    0.07553273, 0.0515472, 0.04740182, 0.03564149, 0.05219905, 0.06065886, 
    0.08834541, 0.0777158, 0.08312993, 0.07947643, 0.01172668, 0.04253845, 
    0.03796929, 0.04496112, 0.008204097, 6.368668e-05, 9.600607e-07, 
    -2.213051e-05,
  1.111839e-06, 1.25969e-07, 5.709395e-08, 0.001396363, 0.005321173, 
    1.109761e-05, 0.0009865934, 0.001248672, 0.01893227, 0.01979201, 
    0.1515112, 0.04327958, 0.02243945, 0.02909829, 0.0351503, 0.01215223, 
    0.0765972, 0.02816422, 0.007151276, 0.010862, 0.0001676884, 0.10795, 
    0.02385544, 0.02490772, 0.02417079, 0.04207984, 0.02218615, 0.002251491, 
    7.745614e-05,
  0.00815081, 0.01147876, 0.07986538, 0.05361351, 0.08105016, 0.05118403, 
    0.008097881, 0.01725704, 0.1409527, 0.2276627, 0.1662795, 0.08185475, 
    0.1064272, 0.1230646, 0.1322647, 0.1227063, 0.08667265, 0.1393578, 
    0.05761707, 0.02773762, 0.03160618, 0.09396382, 0.08958484, 0.05718818, 
    0.06390597, 0.05384525, 0.04399328, 0.03948161, 0.001335437,
  0.07314686, 0.03826935, 0.04249108, 0.1509289, 0.0692457, 0.06119636, 
    0.2239965, 0.007901911, 0.01681602, 0.07771786, 0.08060393, 0.1225273, 
    0.1708328, 0.2615319, 0.1886942, 0.2033139, 0.2161537, 0.1960033, 
    0.160387, 0.1688492, 0.2079011, 0.09469108, 0.1553858, 0.1715167, 
    0.1548923, 0.174506, 0.178967, 0.153606, 0.1646544,
  0.1374434, 0.09597762, 0.1219655, 0.1842736, 0.1879178, 0.2213134, 
    0.1797173, 0.2053777, 0.0759986, 0.05486276, 0.05640024, 0.09149261, 
    0.1622455, 0.3497336, 0.3630072, 0.1260671, 0.1340652, 0.1903284, 
    0.2753078, 0.3058141, 0.1855626, 0.1162609, 0.2029622, 0.2352506, 
    0.2793255, 0.2441172, 0.2912352, 0.2386021, 0.1503875,
  0.1734015, 0.1956604, 0.2363965, 0.3432834, 0.4324775, 0.3564125, 
    0.3988144, 0.4470743, 0.3038332, 0.2939387, 0.3113325, 0.1475237, 
    0.2844807, 0.3264601, 0.2057396, 0.268615, 0.1773062, 0.2076817, 
    0.2681493, 0.2652843, 0.1890991, 0.2022806, 0.1703574, 0.2253494, 
    0.1713701, 0.3406718, 0.2941863, 0.302976, 0.2130504,
  0.2418391, 0.25867, 0.3374869, 0.3739021, 0.287597, 0.219713, 0.27728, 
    0.4232784, 0.3710748, 0.334244, 0.2068515, 0.23743, 0.170772, 0.2414934, 
    0.2649598, 0.2139453, 0.2833968, 0.2649371, 0.1167665, 0.1515553, 
    0.1477053, 0.1379838, 0.1267151, 0.07564735, 0.1048257, 0.4266103, 
    0.3357446, 0.2851625, 0.2577819,
  0.2168252, 0.2621666, 0.2534651, 0.2622187, 0.2459686, 0.2504503, 
    0.2618489, 0.3210958, 0.341526, 0.303158, 0.2638629, 0.2726699, 
    0.2355194, 0.2160985, 0.2021094, 0.1754349, 0.1512703, 0.1719756, 
    0.1957209, 0.2419931, 0.1954056, 0.2036372, 0.1677299, 0.1023321, 
    0.07260007, 0.04573574, 0.1007853, 0.1306753, 0.1812336,
  0.1780684, 0.1802385, 0.1824087, 0.1845788, 0.1867489, 0.188919, 0.1910892, 
    0.1839513, 0.192758, 0.2015647, 0.2103714, 0.2191781, 0.2279848, 
    0.2367915, 0.2447473, 0.2380949, 0.2314425, 0.2247901, 0.2181377, 
    0.2114853, 0.204833, 0.1977354, 0.1934109, 0.1890865, 0.1847621, 
    0.1804376, 0.1761132, 0.1717888, 0.1763323,
  0.1342222, 0.1343382, 0.1682979, 0.265137, 0.1966722, 0.2236016, 0.14979, 
    0.09353268, 0.1108131, 0.140964, 0.1738771, 0.2204999, 0.2634408, 
    0.1938155, 0.1569099, 0.1750952, 0.1624603, 0.1649034, 0.1481507, 
    0.2164971, 0.3160044, 0.3427888, 0.1852279, 0.06454062, 0.1466409, 
    0.1361998, 0.1608026, 0.1292342, 0.122473,
  0.2788541, 0.3449442, 0.2802011, 0.3086194, 0.3099188, 0.2538457, 
    0.2390655, 0.3918294, 0.3274756, 0.3509045, 0.2961255, 0.2094372, 
    0.1696533, 0.1984642, 0.2981815, 0.3556679, 0.3409753, 0.3035729, 
    0.3269112, 0.2406881, 0.2456094, 0.2978657, 0.2996594, 0.331304, 
    0.2243982, 0.1605147, 0.2436567, 0.2952309, 0.2814938,
  0.3158978, 0.3320053, 0.3228939, 0.3200315, 0.3097441, 0.2649171, 
    0.3077126, 0.2978683, 0.3262649, 0.3169838, 0.2739096, 0.2889541, 
    0.2683591, 0.2404127, 0.2804007, 0.2188754, 0.1999834, 0.2906263, 
    0.3494521, 0.3635594, 0.3048401, 0.2643998, 0.2654976, 0.3039395, 
    0.3226536, 0.2706814, 0.28645, 0.2864743, 0.2745438,
  0.2486, 0.229007, 0.2486245, 0.2102217, 0.1898455, 0.1822283, 0.180344, 
    0.1808538, 0.1884521, 0.2716172, 0.2448724, 0.1981892, 0.2136888, 
    0.1611779, 0.1326818, 0.1411343, 0.1201199, 0.1271567, 0.1854452, 
    0.2410894, 0.2362696, 0.2129765, 0.1824121, 0.1652089, 0.05460896, 
    0.09627114, 0.136278, 0.1574671, 0.2162033,
  0.07021748, 0.09210318, 0.03736925, 0.1284071, 0.06256147, 0.1305114, 
    0.06838962, 0.1301124, 0.0823947, 0.04454565, 0.03705415, 0.06346589, 
    0.07209015, 0.05801211, 0.1657497, 0.1063878, 0.05285895, 0.07204045, 
    0.08403312, 0.1017361, 0.1307647, 0.07983845, 0.03912055, 0.005272408, 
    0.007179583, 0.06450386, 0.1010209, 0.08399544, 0.05620628,
  0.03745357, 1.706128e-05, 0.1042226, 0.03046817, 0.09049654, 0.1055891, 
    0.04423991, 0.01685863, 0.009113152, 0.01769497, 0.01362419, 0.005335634, 
    0.02911565, 0.07061466, 0.1364016, 0.0675291, 0.1541237, 0.1232078, 
    0.08869719, 0.05983572, 0.05412669, 0.02268011, 0.0002178352, 
    9.060114e-05, 0.0158833, 0.1553845, 0.03011977, 0.04518631, 0.08109483,
  0.007557689, 0.03134653, 0.09792627, 0.06447886, 0.104771, 0.05124839, 
    0.04769336, 0.07784705, 0.006834467, 0.01597226, 0.08730505, 0.02308678, 
    0.03942867, 0.03517289, 0.07201509, 0.05523299, 0.05040879, 0.03986366, 
    0.04206247, 0.04705034, 0.09173647, 0.05281902, 1.777487e-05, 
    3.519067e-05, 0.1160119, 0.1743381, 0.03314304, 0.06197026, 0.0394218,
  -6.555986e-06, 0.003416628, 0.1728719, 0.05534795, 0.02060982, 0.03028395, 
    0.04408975, 0.02926454, 0.03359779, 0.03756291, 0.07064891, 0.02530554, 
    0.08607584, 0.0427176, 0.09072518, 0.0365653, 0.038217, 0.0229593, 
    0.0247411, 0.02314989, 0.005264005, 0.003748736, 0.0008468644, 0.1362699, 
    0.1410626, 0.08476871, 0.03411739, 0.00340892, 0.0009755947,
  0.001054929, 0.009205291, 0.005487865, 0.03402223, 0.05881526, 0.05640866, 
    0.07639828, 0.1011846, 0.1603782, 0.2057536, 0.03906163, 0.01617426, 
    0.01430469, 0.03613062, 0.04711298, 0.04830097, 0.01304425, 0.02148182, 
    0.03854839, 0.02843527, 0.03550871, 0.03714137, 0.095482, 0.07051513, 
    0.1317307, 0.1581119, 0.03772398, 0.01693582, 0.00201712,
  -1.243036e-06, 4.910883e-08, 1.973806e-07, 0.05927078, 0.02772482, 
    0.02958622, 0.01120812, 0.007343144, 0.03265978, 0.05011597, 0.2034333, 
    0.06694158, 0.04932284, 0.0454357, 0.04127533, 0.05155345, 0.05778734, 
    0.08390167, 0.08085619, 0.08344354, 0.07533511, 0.01352993, 0.05624483, 
    0.0567644, 0.04640976, 0.01005145, 0.0003012345, 1.458303e-07, 
    1.396469e-05,
  8.611628e-07, 6.012633e-08, 2.925791e-08, 0.007513577, 0.0006191681, 
    3.916695e-05, 0.001912853, 0.003078077, 0.03284147, 0.03375594, 
    0.1451255, 0.07139494, 0.02690258, 0.03607969, 0.05378847, 0.0184721, 
    0.07397239, 0.03317128, 0.01852787, 0.01850831, 0.0002367695, 0.1204461, 
    0.02279573, 0.02839386, 0.02818263, 0.04187945, 0.03472187, 0.00109553, 
    5.48967e-06,
  0.008394836, 0.02217072, 0.09244065, 0.03149331, 0.08166976, 0.0438023, 
    0.0007143129, 0.010118, 0.1212895, 0.2087106, 0.1793193, 0.1149513, 
    0.1301308, 0.1355048, 0.1440008, 0.1350565, 0.09201044, 0.141038, 
    0.07245088, 0.02773808, 0.02741969, 0.1015765, 0.09316888, 0.0689104, 
    0.06097925, 0.05870235, 0.051096, 0.05159817, 0.0001214593,
  0.0727368, 0.04232673, 0.04814396, 0.1740977, 0.06856401, 0.05232615, 
    0.2221734, 0.004020031, 0.01364064, 0.08506737, 0.06644326, 0.1790634, 
    0.214389, 0.2896905, 0.2041585, 0.2251014, 0.2592297, 0.2077748, 
    0.1742897, 0.1800019, 0.1937096, 0.08947203, 0.1682844, 0.1687128, 
    0.195443, 0.1945946, 0.1937816, 0.1535566, 0.179641,
  0.1344978, 0.1102693, 0.1198036, 0.1718405, 0.1550872, 0.238171, 0.175074, 
    0.1971691, 0.06186418, 0.04225338, 0.0538111, 0.08650278, 0.1549454, 
    0.3422877, 0.3642392, 0.1430971, 0.1590669, 0.2177751, 0.2904098, 
    0.3276163, 0.1794824, 0.1055965, 0.2125324, 0.2478839, 0.2776244, 
    0.3042893, 0.308818, 0.2516728, 0.1562582,
  0.1865498, 0.1789653, 0.2538637, 0.3367428, 0.4326749, 0.350399, 0.4462757, 
    0.4494516, 0.3242824, 0.2919064, 0.2741169, 0.1432563, 0.2742844, 
    0.3769595, 0.2747182, 0.236109, 0.191643, 0.2077942, 0.2773952, 
    0.2808291, 0.1703077, 0.1821507, 0.1505317, 0.2254252, 0.1662107, 
    0.3630058, 0.3026859, 0.3094129, 0.2278347,
  0.2473198, 0.2681151, 0.3396567, 0.3683017, 0.2599999, 0.1765195, 
    0.2567286, 0.4343899, 0.3586668, 0.3342646, 0.2234673, 0.2413779, 
    0.1729767, 0.2600689, 0.2876633, 0.2251958, 0.3003948, 0.2798705, 
    0.1193237, 0.1602232, 0.150277, 0.1387636, 0.1481604, 0.04867469, 
    0.07729357, 0.4405239, 0.3394955, 0.2746085, 0.2728966,
  0.1903589, 0.2271825, 0.2487225, 0.2581985, 0.2289331, 0.2470897, 
    0.2806015, 0.3248069, 0.3670603, 0.3391537, 0.2887142, 0.287452, 
    0.2518539, 0.2173983, 0.202052, 0.1992109, 0.1708232, 0.2015865, 
    0.226971, 0.2674913, 0.2276632, 0.2039913, 0.1725393, 0.1056696, 
    0.06781064, 0.05129334, 0.09909879, 0.1577019, 0.2386538,
  0.1760776, 0.1780888, 0.1801, 0.1821112, 0.1841224, 0.1861336, 0.1881447, 
    0.184544, 0.1935308, 0.2025176, 0.2115043, 0.2204911, 0.2294779, 
    0.2384647, 0.2426757, 0.2364714, 0.2302671, 0.2240628, 0.2178584, 
    0.2116541, 0.2054498, 0.2056757, 0.2008821, 0.1960884, 0.1912948, 
    0.1865011, 0.1817075, 0.1769138, 0.1744687,
  0.147202, 0.1407095, 0.2007303, 0.2964897, 0.2239634, 0.250065, 0.1931499, 
    0.1178017, 0.145337, 0.175843, 0.1747135, 0.2169951, 0.2988385, 
    0.1214618, 0.09676326, 0.1390972, 0.1580369, 0.1397023, 0.1066086, 
    0.1819569, 0.3425395, 0.3275997, 0.1675303, 0.04823862, 0.1262435, 
    0.1918142, 0.1764475, 0.115575, 0.141291,
  0.2716333, 0.324853, 0.2870238, 0.2837218, 0.3079265, 0.2251124, 0.2226646, 
    0.3818561, 0.3573143, 0.3468321, 0.2902946, 0.1644938, 0.1534, 0.234877, 
    0.3874177, 0.3945093, 0.3768382, 0.3422382, 0.3757827, 0.2636122, 
    0.2769429, 0.3069559, 0.3109998, 0.3289468, 0.2634582, 0.234273, 
    0.2444208, 0.3116135, 0.3471092,
  0.3651997, 0.3388646, 0.2954913, 0.3481017, 0.3182544, 0.3075367, 
    0.3126355, 0.3097042, 0.3521595, 0.365448, 0.2916558, 0.3319822, 
    0.2863511, 0.2898245, 0.3080466, 0.2457712, 0.2514098, 0.3041436, 
    0.3611389, 0.3895914, 0.3243643, 0.2647095, 0.2917128, 0.3425731, 
    0.2981868, 0.2942912, 0.3004499, 0.3314331, 0.3447787,
  0.2659954, 0.2506498, 0.2749904, 0.23371, 0.2061055, 0.2051907, 0.1978376, 
    0.217602, 0.2319722, 0.3114879, 0.2703323, 0.2402582, 0.2359489, 
    0.1749211, 0.1531648, 0.1563371, 0.1364442, 0.1619335, 0.2484961, 
    0.3021609, 0.2586043, 0.2592159, 0.2265834, 0.1653831, 0.04199558, 
    0.08494221, 0.1493625, 0.1602974, 0.2422625,
  0.092359, 0.1185014, 0.09057777, 0.1458613, 0.1065091, 0.1553668, 
    0.08796286, 0.1485598, 0.1343376, 0.07914032, 0.09769517, 0.1040986, 
    0.07755176, 0.07819659, 0.1654074, 0.1352056, 0.07292629, 0.08264953, 
    0.1113043, 0.1183526, 0.1608094, 0.127318, 0.06598473, 0.007782527, 
    0.01281431, 0.08069965, 0.1062201, 0.09551305, 0.08322704,
  0.05728864, 0.001003668, 0.1015098, 0.05922897, 0.09878707, 0.1005207, 
    0.05489922, 0.06717603, 0.01185994, 0.01742116, 0.01860609, 0.004830776, 
    0.01571168, 0.1008192, 0.150692, 0.08233963, 0.1656546, 0.1479096, 
    0.06847954, 0.06095353, 0.05179769, 0.04028745, 0.00645656, 7.559919e-05, 
    0.01420313, 0.148938, 0.03107858, 0.04971472, 0.09818541,
  0.01212345, 0.02196238, 0.08997263, 0.05953482, 0.08188729, 0.0416556, 
    0.0395086, 0.0862906, 0.01311546, 0.018488, 0.07776212, 0.02429157, 
    0.03695171, 0.03630419, 0.06297392, 0.05264945, 0.0439296, 0.03267545, 
    0.03301707, 0.03221308, 0.06340222, 0.1149542, 0.004902036, 0.0001524797, 
    0.1126846, 0.1664008, 0.02726634, 0.04478915, 0.07767452,
  0.002298605, 0.002318896, 0.1457399, 0.05322212, 0.02000559, 0.02819326, 
    0.0384049, 0.0303066, 0.03969248, 0.03122973, 0.06297237, 0.02062678, 
    0.07350147, 0.03299734, 0.07225086, 0.03288253, 0.03247558, 0.02327776, 
    0.02526302, 0.03106378, 0.009509313, 0.008903669, 0.0107191, 0.119529, 
    0.1178044, 0.06902538, 0.03711066, 0.0217847, 0.01354012,
  0.001292822, 0.01008661, 0.003582717, 0.02211323, 0.06094595, 0.06356439, 
    0.0624348, 0.08988668, 0.1536246, 0.21841, 0.0325253, 0.0172144, 
    0.0169438, 0.0324524, 0.04300281, 0.03772033, 0.01695629, 0.02466078, 
    0.04803202, 0.0395974, 0.05189643, 0.03730212, 0.0784017, 0.06439574, 
    0.120732, 0.1279973, 0.03176054, 0.01725317, 0.001838149,
  -8.866825e-08, 1.324957e-08, 2.773267e-08, 0.02882586, 0.05440769, 
    0.02855586, 0.01252196, 0.01222098, 0.02757744, 0.05180359, 0.1913218, 
    0.05978575, 0.04875019, 0.04161799, 0.04346504, 0.04522285, 0.05526297, 
    0.08232819, 0.08625069, 0.07460865, 0.06085514, 0.01444719, 0.06950854, 
    0.06415284, 0.0417272, 0.01199366, 0.0051944, 5.667202e-08, 1.54638e-05,
  5.068844e-07, 3.467137e-08, 1.625181e-08, 0.0229352, 4.77892e-05, 
    0.0006983427, 0.0002853755, 0.004540418, 0.01187377, 0.09425273, 
    0.1576878, 0.08073759, 0.04468141, 0.05876609, 0.07764223, 0.02977654, 
    0.07277585, 0.03961833, 0.0292857, 0.02373708, -1.296505e-05, 0.1619197, 
    0.02989269, 0.03244266, 0.04933107, 0.0554328, 0.04611034, -4.801419e-06, 
    2.018476e-06,
  0.007213081, 0.04432862, 0.1051809, 0.0335145, 0.0738534, 0.03817953, 
    -0.001498902, 0.003403302, 0.1071007, 0.186943, 0.1935083, 0.2098679, 
    0.182896, 0.1861207, 0.1839783, 0.1544196, 0.1237486, 0.1509781, 
    0.1086526, 0.03493045, 0.03462102, 0.1089202, 0.1108412, 0.1036894, 
    0.06818189, 0.07022834, 0.07095402, 0.06733774, 0.001911658,
  0.08829785, 0.04059012, 0.0701203, 0.2071577, 0.09111968, 0.06148374, 
    0.2147461, 0.001731082, 0.01496648, 0.08557104, 0.06360193, 0.2458553, 
    0.3061365, 0.2688636, 0.2511411, 0.2523983, 0.2787127, 0.248896, 
    0.2186991, 0.201598, 0.1974628, 0.08147527, 0.1817966, 0.1803522, 
    0.2646092, 0.2419112, 0.237125, 0.184607, 0.214716,
  0.1449251, 0.1340307, 0.112881, 0.1890194, 0.1702041, 0.2431524, 0.1743014, 
    0.1955743, 0.04690054, 0.0309641, 0.03846467, 0.08142093, 0.1869409, 
    0.3341797, 0.3620271, 0.1804353, 0.2033775, 0.2726921, 0.2766077, 
    0.3711154, 0.1702573, 0.09070686, 0.242859, 0.2650772, 0.2821853, 
    0.3926358, 0.3040377, 0.2430455, 0.158794,
  0.2059605, 0.1907653, 0.2681437, 0.2911507, 0.4424839, 0.3354417, 
    0.4221098, 0.4901053, 0.3588495, 0.3082241, 0.2916338, 0.1421163, 
    0.2627161, 0.4034176, 0.291803, 0.2133703, 0.2288093, 0.2085912, 
    0.281077, 0.2899749, 0.1707495, 0.1855009, 0.1615349, 0.2295489, 
    0.2112306, 0.3503926, 0.2955038, 0.3145871, 0.2751226,
  0.2876239, 0.2697419, 0.3355943, 0.3851547, 0.24268, 0.193711, 0.293186, 
    0.4479768, 0.3495136, 0.3392792, 0.2552094, 0.2446796, 0.1792581, 
    0.2652269, 0.2991959, 0.2220643, 0.2804484, 0.2638623, 0.1180668, 
    0.1814157, 0.1720126, 0.1532223, 0.1528249, 0.03486055, 0.06405293, 
    0.4400927, 0.3466476, 0.2637841, 0.3008345,
  0.1473466, 0.2222023, 0.253957, 0.2567783, 0.2048689, 0.2472851, 0.2892417, 
    0.3247331, 0.3954988, 0.3675381, 0.3158148, 0.3004389, 0.265454, 
    0.2346101, 0.2033626, 0.2114397, 0.2166966, 0.2307302, 0.2435801, 
    0.2826963, 0.2416038, 0.2197014, 0.1712151, 0.1003547, 0.07453348, 
    0.0463902, 0.09603653, 0.1794052, 0.2371902,
  0.174702, 0.1771754, 0.1796488, 0.1821222, 0.1845957, 0.1870691, 0.1895425, 
    0.1868735, 0.1958825, 0.2048914, 0.2139004, 0.2229093, 0.2319182, 
    0.2409272, 0.2471633, 0.2422357, 0.2373081, 0.2323805, 0.2274529, 
    0.2225253, 0.2175977, 0.2122356, 0.2056808, 0.1991261, 0.1925713, 
    0.1860166, 0.1794618, 0.1729071, 0.1727233,
  0.158749, 0.1447772, 0.2111688, 0.3253312, 0.2389597, 0.2460824, 0.2311058, 
    0.1718126, 0.1960601, 0.2094832, 0.2041764, 0.2425322, 0.3151486, 
    0.07318197, 0.1075664, 0.09822696, 0.1677845, 0.1240462, 0.1020825, 
    0.162859, 0.3590238, 0.3289166, 0.1645503, 0.05827722, 0.104826, 
    0.1762991, 0.1587908, 0.09101493, 0.1337813,
  0.3346524, 0.3384781, 0.2841801, 0.2663498, 0.2794449, 0.2197081, 
    0.2011008, 0.3797984, 0.3678622, 0.3405583, 0.2777183, 0.1246378, 
    0.1443575, 0.2426315, 0.4478413, 0.4430691, 0.4185151, 0.4581448, 
    0.412323, 0.358647, 0.3159925, 0.3795148, 0.3717578, 0.3483629, 
    0.3142953, 0.3849083, 0.3526988, 0.4161435, 0.4769868,
  0.3905968, 0.3627344, 0.3489692, 0.3772142, 0.3807271, 0.3918085, 
    0.4064489, 0.3554559, 0.3884109, 0.4115262, 0.3086566, 0.3893987, 
    0.3781653, 0.3934491, 0.3757339, 0.2911341, 0.3057221, 0.3409326, 
    0.3996481, 0.4006979, 0.3596236, 0.2960882, 0.3512772, 0.4241486, 
    0.3244819, 0.3938322, 0.404378, 0.4253024, 0.4345553,
  0.3585407, 0.3099765, 0.3063866, 0.277526, 0.2390816, 0.2438699, 0.2241724, 
    0.2559358, 0.2660652, 0.3687345, 0.3321931, 0.3031145, 0.2783389, 
    0.1991358, 0.1779349, 0.2091142, 0.1897629, 0.2219177, 0.3071346, 
    0.3359316, 0.2929381, 0.3008912, 0.2671562, 0.1772376, 0.02532705, 
    0.1040314, 0.1716966, 0.2098169, 0.3159123,
  0.1711752, 0.20565, 0.2075077, 0.1815874, 0.1579983, 0.2025548, 0.1566199, 
    0.1953814, 0.1820784, 0.1489178, 0.1645187, 0.1642466, 0.1261442, 
    0.1021384, 0.1977933, 0.1710048, 0.1096731, 0.1448139, 0.1633254, 
    0.2029432, 0.2068221, 0.1646105, 0.1438012, 0.01191921, 0.01844431, 
    0.1181291, 0.1301379, 0.1173568, 0.1502185,
  0.1023504, 0.0108739, 0.09358928, 0.0862163, 0.09537095, 0.1004987, 
    0.05600167, 0.1004284, 0.07986579, 0.02215272, 0.01724542, 0.006103139, 
    0.006803042, 0.1236619, 0.1696959, 0.09827895, 0.164565, 0.1603669, 
    0.06195439, 0.07012941, 0.04758048, 0.08053653, 0.05833708, 0.0001660293, 
    0.01498639, 0.1521533, 0.03132232, 0.04974872, 0.1057876,
  0.0723468, 0.01942881, 0.06535441, 0.06034952, 0.06724525, 0.03787524, 
    0.04742277, 0.09473586, 0.03732707, 0.01785662, 0.06892804, 0.01810666, 
    0.04167381, 0.04348507, 0.04696954, 0.04639044, 0.0413585, 0.03100371, 
    0.03038502, 0.03177636, 0.04553907, 0.1852974, 0.05802375, 0.000119332, 
    0.1001812, 0.1681944, 0.02917213, 0.04119513, 0.08838436,
  0.02206658, 0.003835391, 0.1162006, 0.06038791, 0.02279511, 0.02842047, 
    0.03796604, 0.03465964, 0.05084166, 0.02829955, 0.05558047, 0.01962428, 
    0.0647921, 0.0309763, 0.06279429, 0.03439723, 0.03194384, 0.02573699, 
    0.02776131, 0.03171334, 0.02519253, 0.01550309, 0.04592852, 0.1037635, 
    0.09741404, 0.0587561, 0.04398777, 0.04158902, 0.05329943,
  0.002565622, 0.01164035, 0.001715713, 0.01691517, 0.06145608, 0.05233323, 
    0.05850318, 0.0742237, 0.1448949, 0.2064595, 0.02805157, 0.02071233, 
    0.02175162, 0.03261391, 0.04316109, 0.03130329, 0.0158908, 0.02412284, 
    0.04207389, 0.03554061, 0.05486428, 0.03065307, 0.06723306, 0.05758299, 
    0.1123255, 0.09519273, 0.02922478, 0.02227797, 0.003010847,
  -5.839981e-08, 3.889545e-09, 7.173255e-09, 0.01081039, 0.09474533, 
    0.03390606, 0.01500197, 0.02900327, 0.01691866, 0.05740371, 0.1662332, 
    0.05652183, 0.05255272, 0.05368453, 0.04899141, 0.04841164, 0.05548877, 
    0.08002711, 0.1017246, 0.0863526, 0.04983708, 0.01925458, 0.09807579, 
    0.08400137, 0.0448738, 0.02163994, 0.01173555, 1.012473e-07, 1.427063e-05,
  2.16536e-07, 2.707833e-08, -3.402021e-07, 0.004582884, 1.748437e-05, 
    0.02473929, 7.027302e-05, 0.007832409, 0.005755618, 0.1240423, 0.1720744, 
    0.1285972, 0.06998908, 0.1173447, 0.1131476, 0.05138085, 0.08713252, 
    0.0513375, 0.07089444, 0.04813636, 0.007061532, 0.200968, 0.03468759, 
    0.02483756, 0.0641045, 0.09556408, 0.09056804, 0.02206263, 9.334256e-07,
  0.001792723, 0.04962005, 0.1353598, 0.03202659, 0.06731391, 0.03328693, 
    -0.001935069, 0.001251202, 0.1044216, 0.168181, 0.2545797, 0.2426023, 
    0.188874, 0.1907267, 0.1725069, 0.1899906, 0.1585229, 0.1720633, 
    0.1625242, 0.03900802, 0.03794004, 0.1410828, 0.1122811, 0.1448493, 
    0.09317021, 0.1122961, 0.1077955, 0.0746557, 0.005326019,
  0.1061234, 0.04963314, 0.08663776, 0.2500967, 0.1354056, 0.05752005, 
    0.1972452, 0.000292442, 0.01767191, 0.08031914, 0.05568181, 0.2812251, 
    0.403819, 0.2694127, 0.2460947, 0.2757991, 0.3374124, 0.308803, 
    0.2255973, 0.2201006, 0.2112258, 0.08054358, 0.1963025, 0.2016861, 
    0.3738996, 0.3188824, 0.2665056, 0.2028485, 0.2137482,
  0.1473055, 0.1437367, 0.138782, 0.2111726, 0.2221125, 0.2709911, 0.1977228, 
    0.202683, 0.03803561, 0.02409612, 0.03213334, 0.07859711, 0.2587108, 
    0.3870093, 0.3740563, 0.2807404, 0.2881465, 0.3269736, 0.2806115, 
    0.3945296, 0.1537805, 0.1016054, 0.2569592, 0.286301, 0.3036788, 
    0.4532354, 0.2797396, 0.2266601, 0.1580088,
  0.2253467, 0.2226405, 0.2505394, 0.3210912, 0.4353592, 0.3747256, 
    0.4686378, 0.5038189, 0.402603, 0.3853797, 0.3247948, 0.1499657, 
    0.2295127, 0.4569327, 0.3471153, 0.2413848, 0.2388644, 0.2142633, 
    0.2974864, 0.2717766, 0.1885992, 0.2131251, 0.1852539, 0.2376525, 
    0.3603033, 0.3301662, 0.2448092, 0.3088619, 0.2636025,
  0.3951156, 0.2493563, 0.3547193, 0.4420049, 0.2773438, 0.2258554, 
    0.3213049, 0.4578169, 0.3589986, 0.3527664, 0.3041354, 0.2479028, 
    0.1950792, 0.2931703, 0.3133923, 0.2276224, 0.3126683, 0.2736523, 
    0.1343812, 0.2168115, 0.1990703, 0.1865191, 0.1658473, 0.03447808, 
    0.05530617, 0.4316154, 0.3625301, 0.2711732, 0.3461527,
  0.1513051, 0.2071297, 0.2685127, 0.2474339, 0.1868778, 0.2787305, 
    0.3144193, 0.3609465, 0.4313138, 0.4096555, 0.362067, 0.3117278, 
    0.2916436, 0.2638911, 0.220193, 0.2363982, 0.2478583, 0.2751282, 
    0.2637928, 0.291138, 0.2584282, 0.2368406, 0.1761796, 0.1041624, 
    0.07537279, 0.04447719, 0.09575871, 0.1931351, 0.2232443,
  0.1772873, 0.1800762, 0.182865, 0.1856539, 0.1884428, 0.1912317, 0.1940206, 
    0.1996081, 0.2092738, 0.2189394, 0.228605, 0.2382706, 0.2479362, 
    0.2576019, 0.2698688, 0.2649002, 0.2599317, 0.2549632, 0.2499946, 
    0.2450261, 0.2400575, 0.2215168, 0.2140308, 0.2065449, 0.1990589, 
    0.191573, 0.184087, 0.1766011, 0.1750562,
  0.1713431, 0.1576829, 0.2115994, 0.3419101, 0.2601482, 0.2555977, 
    0.2553347, 0.2059861, 0.2411436, 0.2320804, 0.2128963, 0.2581657, 
    0.3434444, 0.05834168, 0.12123, 0.0900989, 0.1047302, 0.12927, 0.1382655, 
    0.1488054, 0.3397064, 0.3158655, 0.1524187, 0.1118942, 0.1733439, 
    0.2591021, 0.121995, 0.1029142, 0.1742212,
  0.3524147, 0.3341598, 0.3146088, 0.2406033, 0.2473337, 0.2168283, 
    0.1789933, 0.3816491, 0.3627763, 0.3398317, 0.2529078, 0.1014329, 
    0.1353802, 0.2218674, 0.4044511, 0.410846, 0.3552669, 0.4372334, 
    0.4701498, 0.4141834, 0.3723544, 0.459015, 0.3984134, 0.3679386, 
    0.3551768, 0.4365516, 0.4345207, 0.4615044, 0.518958,
  0.4165664, 0.4031247, 0.4170028, 0.4352254, 0.435951, 0.4409446, 0.4698615, 
    0.4449233, 0.4369366, 0.4226585, 0.3475349, 0.4378045, 0.4751284, 
    0.4736807, 0.452315, 0.387524, 0.3660832, 0.4362602, 0.4535971, 
    0.3822383, 0.3598362, 0.3083697, 0.3744225, 0.4514486, 0.4085135, 
    0.5149578, 0.4648813, 0.4878076, 0.4974751,
  0.4063131, 0.3609424, 0.3619741, 0.316703, 0.2910626, 0.3027575, 0.2761267, 
    0.3325603, 0.3715099, 0.4137321, 0.3738195, 0.3636566, 0.3294745, 
    0.265798, 0.2985823, 0.2917644, 0.3415629, 0.3489213, 0.3358571, 
    0.3569444, 0.2835035, 0.2867281, 0.3142206, 0.1891948, 0.01666898, 
    0.135573, 0.2382704, 0.2968793, 0.387913,
  0.2391402, 0.287694, 0.247006, 0.2770811, 0.2494531, 0.30378, 0.2080564, 
    0.2689427, 0.3338574, 0.2416367, 0.2207122, 0.2636332, 0.12994, 
    0.1463152, 0.2118714, 0.2454484, 0.2020664, 0.2967947, 0.2878701, 
    0.2300581, 0.2057391, 0.1818875, 0.2211379, 0.01491018, 0.03515094, 
    0.1498383, 0.1758718, 0.1793593, 0.2567693,
  0.172911, 0.06414834, 0.08964302, 0.1242414, 0.09334899, 0.107752, 
    0.06931872, 0.140073, 0.248872, 0.02105894, 0.0167683, 0.005302512, 
    0.003504686, 0.1471109, 0.1870005, 0.1184647, 0.1600741, 0.1933309, 
    0.06481997, 0.08958977, 0.05266163, 0.163554, 0.2103775, 0.0003306605, 
    0.01497472, 0.1516211, 0.05043909, 0.063943, 0.1305816,
  0.2023013, 0.02245236, 0.04582101, 0.07030087, 0.06124524, 0.044929, 
    0.06336078, 0.1051928, 0.1081728, 0.02921512, 0.05763038, 0.01263548, 
    0.04600054, 0.05896421, 0.04274013, 0.05542099, 0.04800079, 0.03181887, 
    0.04982321, 0.04286139, 0.04883338, 0.1732046, 0.2728288, 0.0005142387, 
    0.07546144, 0.1619577, 0.0568904, 0.0444192, 0.1023527,
  0.07681379, 0.01174509, 0.09045213, 0.06412284, 0.0292352, 0.03412784, 
    0.04180155, 0.05541731, 0.06654968, 0.02895678, 0.05340222, 0.02258251, 
    0.05646361, 0.03466074, 0.05578446, 0.03950863, 0.04231831, 0.04157462, 
    0.05406924, 0.04816442, 0.05998486, 0.05198144, 0.09067802, 0.08955421, 
    0.07823543, 0.03899654, 0.06029222, 0.05674955, 0.08820109,
  0.004065648, 0.00957316, 0.0008594268, 0.01572965, 0.06436626, 0.05010129, 
    0.06178243, 0.06999291, 0.1536282, 0.1751698, 0.03129262, 0.02775983, 
    0.02816786, 0.04058155, 0.05307455, 0.03420098, 0.01616578, 0.01798096, 
    0.03651622, 0.02858582, 0.0447553, 0.03340463, 0.05802851, 0.04029349, 
    0.09668015, 0.07129013, 0.03221329, 0.03435687, 0.00757046,
  -4.256728e-08, 1.549549e-09, 1.476582e-09, 0.001936628, 0.09394284, 
    0.1506947, 0.009455739, 0.09857564, 0.01203959, 0.08637363, 0.1573734, 
    0.05934234, 0.0731549, 0.07453395, 0.0607644, 0.0614804, 0.06300826, 
    0.08952519, 0.1039403, 0.0885843, 0.04875009, 0.03308076, 0.1183897, 
    0.08137607, 0.06335589, 0.116641, 0.04013422, 1.0106e-07, 8.337783e-06,
  7.406757e-08, 1.812733e-08, -4.442707e-06, 0.005537944, -1.496527e-06, 
    0.01802153, 3.666252e-05, 0.008436032, 0.003802861, 0.1984835, 0.2173527, 
    0.1694563, 0.1251898, 0.1464952, 0.1889791, 0.10567, 0.1266638, 
    0.07080086, 0.1466632, 0.2081611, 0.008074163, 0.2451442, 0.04135729, 
    0.02688439, 0.05903009, 0.09620282, 0.08096275, 0.02715571, 4.433148e-07,
  0.0001350955, 0.04043571, 0.08200958, 0.0322258, 0.06329293, 0.02972811, 
    -0.002104412, 0.0005295128, 0.09245961, 0.1702815, 0.238511, 0.1471445, 
    0.1255589, 0.1401419, 0.1562353, 0.1807729, 0.1982964, 0.1928666, 
    0.2120961, 0.04808237, 0.04077107, 0.191498, 0.1210379, 0.1546445, 
    0.09577344, 0.1528427, 0.1302129, 0.1269679, 0.00329059,
  0.1300784, 0.05801067, 0.09238801, 0.2802418, 0.1299328, 0.05425447, 
    0.1814691, -0.000139123, 0.02181982, 0.07315378, 0.05858842, 0.2242521, 
    0.3307772, 0.1978291, 0.2025301, 0.2692083, 0.377078, 0.3109521, 
    0.2208077, 0.224765, 0.223095, 0.1109441, 0.2167388, 0.2345094, 
    0.3516716, 0.2760698, 0.2503754, 0.21173, 0.2146147,
  0.1870732, 0.1613921, 0.1614133, 0.2279236, 0.3012979, 0.3058037, 
    0.2346727, 0.2105932, 0.03100927, 0.02256939, 0.02768112, 0.07736664, 
    0.2981478, 0.4039094, 0.4343557, 0.3215969, 0.300824, 0.2566865, 
    0.2342632, 0.4330483, 0.1526686, 0.1512214, 0.2872266, 0.3132826, 
    0.3442912, 0.396067, 0.2191225, 0.232677, 0.159934,
  0.2363079, 0.1952273, 0.2799276, 0.3868482, 0.516845, 0.3982199, 0.4916035, 
    0.542146, 0.4198652, 0.475169, 0.3535045, 0.1749764, 0.2285015, 
    0.4272746, 0.487214, 0.2337666, 0.2656171, 0.2234846, 0.3055883, 
    0.2665545, 0.2104037, 0.2325199, 0.2007982, 0.2538955, 0.6160147, 
    0.2558415, 0.1823834, 0.2570903, 0.2421868,
  0.3327157, 0.2316149, 0.3393949, 0.4703144, 0.3005858, 0.2588072, 
    0.3453027, 0.4936554, 0.3764588, 0.3779202, 0.3721724, 0.2655944, 
    0.2015337, 0.3071854, 0.3488883, 0.2650547, 0.3419076, 0.3083428, 
    0.1540684, 0.2292953, 0.2133732, 0.2185281, 0.1862397, 0.03874956, 
    0.05139354, 0.3979619, 0.3678027, 0.2557662, 0.4214158,
  0.1636024, 0.2037111, 0.2698779, 0.2396627, 0.2235518, 0.3253517, 
    0.3989976, 0.3978201, 0.4775258, 0.4490657, 0.396033, 0.3437648, 
    0.3272519, 0.3105235, 0.2634331, 0.2944216, 0.2851112, 0.3119218, 
    0.288345, 0.3223749, 0.2818917, 0.2613462, 0.190493, 0.09760953, 
    0.07485995, 0.04773012, 0.09331728, 0.1989931, 0.2243953,
  0.2137329, 0.2146626, 0.2155923, 0.2165219, 0.2174516, 0.2183813, 0.219311, 
    0.216273, 0.2249576, 0.2336421, 0.2423266, 0.2510111, 0.2596956, 
    0.2683801, 0.2760611, 0.2714767, 0.2668924, 0.262308, 0.2577237, 
    0.2531393, 0.248555, 0.2424747, 0.2374448, 0.232415, 0.2273851, 
    0.2223553, 0.2173255, 0.2122956, 0.2129892,
  0.2201871, 0.1910039, 0.2164541, 0.3746551, 0.2819608, 0.2649441, 
    0.2609999, 0.2370318, 0.2736914, 0.260484, 0.2292774, 0.25668, 0.334896, 
    0.04146233, 0.1167254, 0.09699911, 0.1101126, 0.1595928, 0.1664041, 
    0.146928, 0.3588821, 0.3271769, 0.1574291, 0.150683, 0.2254653, 
    0.2947528, 0.1122406, 0.115284, 0.1911054,
  0.3599111, 0.3212604, 0.2898379, 0.1671827, 0.2172007, 0.2001433, 0.138348, 
    0.3852051, 0.3998961, 0.360161, 0.2482264, 0.07542764, 0.1134021, 
    0.1891098, 0.3081765, 0.3741327, 0.342492, 0.4182391, 0.4686556, 
    0.4521005, 0.4184477, 0.4590414, 0.4597757, 0.3856432, 0.3368225, 
    0.4146191, 0.391113, 0.4261981, 0.4256611,
  0.4428849, 0.40322, 0.4106534, 0.4808181, 0.4858466, 0.4476914, 0.4631266, 
    0.4498747, 0.4577881, 0.3933306, 0.3931017, 0.4928379, 0.5133356, 
    0.5119003, 0.4445272, 0.4362686, 0.445547, 0.5171956, 0.45186, 0.3529769, 
    0.3374759, 0.3207799, 0.3869036, 0.4407073, 0.4696913, 0.4748712, 
    0.4933234, 0.4788173, 0.4849135,
  0.404659, 0.3934537, 0.4120802, 0.3604748, 0.3296093, 0.3636429, 0.3601723, 
    0.3448131, 0.3620925, 0.408168, 0.3520487, 0.4851964, 0.4043398, 
    0.337204, 0.3333242, 0.4179758, 0.4097601, 0.461542, 0.3389565, 0.328104, 
    0.2572623, 0.3026376, 0.2863903, 0.1993617, 0.01203097, 0.1392893, 
    0.3147004, 0.4007233, 0.4128573,
  0.3064471, 0.2886068, 0.2389448, 0.3170679, 0.2871163, 0.2639123, 
    0.2268202, 0.2912212, 0.3755516, 0.336591, 0.3301434, 0.2367302, 
    0.08362389, 0.1878017, 0.2347255, 0.3336609, 0.3083005, 0.3143246, 
    0.3316227, 0.268045, 0.2456702, 0.1929728, 0.274555, 0.01840587, 
    0.02639263, 0.1887848, 0.2045228, 0.2475177, 0.2729163,
  0.1559728, 0.1179136, 0.07466379, 0.1199248, 0.1330924, 0.1177474, 
    0.09052648, 0.1714354, 0.232256, 0.02035414, 0.02504143, 0.007557584, 
    0.0007518844, 0.103477, 0.2132128, 0.115858, 0.1702826, 0.2317119, 
    0.1324198, 0.08700387, 0.1227734, 0.1706197, 0.3235874, 0.0006346975, 
    0.01567438, 0.1585943, 0.08425903, 0.08640094, 0.155745,
  0.2668386, 0.02969886, 0.02700784, 0.1072741, 0.05658951, 0.06401362, 
    0.06482878, 0.08467019, 0.1770155, 0.07410952, 0.04301101, 0.00612391, 
    0.04541411, 0.1062867, 0.1069512, 0.07902721, 0.06589558, 0.06851597, 
    0.0428457, 0.0420969, 0.04571863, 0.1058222, 0.374663, 0.007554469, 
    0.05642287, 0.1542338, 0.04696689, 0.05194853, 0.08061263,
  0.1588415, 0.06300066, 0.05896857, 0.05926128, 0.05578795, 0.08463525, 
    0.09883849, 0.06837626, 0.1144157, 0.04675806, 0.05162232, 0.0357184, 
    0.05195797, 0.07388224, 0.08989261, 0.07650384, 0.05071476, 0.06959966, 
    0.0706526, 0.09488387, 0.1480998, 0.1612891, 0.1542203, 0.05842816, 
    0.05697614, 0.02438754, 0.07409588, 0.1168884, 0.1344685,
  0.03402497, 0.005502729, 0.0003333723, 0.01139442, 0.07840277, 0.06720649, 
    0.09990046, 0.06310323, 0.1247092, 0.1414309, 0.05153045, 0.0686359, 
    0.0886005, 0.05779179, 0.09717378, 0.06638175, 0.02552259, 0.0171334, 
    0.03929362, 0.02803065, 0.05179637, 0.05047352, 0.04869173, 0.01887987, 
    0.05980311, 0.08095533, 0.04184658, 0.09634096, 0.05739862,
  -2.332465e-08, 8.845001e-10, 4.392898e-10, -0.001512694, 0.1149403, 
    0.1230373, 0.006009783, 0.09890893, 0.01401399, 0.1230187, 0.1577519, 
    0.05383008, 0.04769947, 0.06246433, 0.08644149, 0.0893679, 0.1115162, 
    0.0875192, 0.1012148, 0.08823849, 0.05865776, 0.06688462, 0.2049455, 
    0.09390405, 0.04089117, 0.06171774, 0.1966093, -8.085022e-05, 3.818802e-06,
  3.998217e-08, 1.124066e-08, -2.513431e-06, 0.0008868483, -1.935767e-07, 
    0.02108464, -3.05299e-07, 0.007159789, 0.002686795, 0.3033271, 0.2010862, 
    0.1307098, 0.09305948, 0.1249678, 0.141659, 0.08015344, 0.1409832, 
    0.1061124, 0.1195445, 0.2142476, 0.01280609, 0.2587419, 0.06466587, 
    0.02210091, 0.02536767, 0.0461885, 0.07839179, 0.005590778, 2.940087e-07,
  -5.057085e-05, 0.03844419, 0.03414019, 0.03368667, 0.05845356, 0.02083888, 
    -0.002071818, 0.0002277263, 0.06810173, 0.1619436, 0.1802989, 0.09261842, 
    0.1016852, 0.1049575, 0.1596547, 0.1462503, 0.1788759, 0.2124998, 
    0.1582035, 0.08271796, 0.05019798, 0.2220042, 0.1287657, 0.1659549, 
    0.1789533, 0.1720668, 0.07115982, 0.1071272, 0.001592829,
  0.1240364, 0.0489939, 0.08743791, 0.3000549, 0.07455126, 0.03186103, 
    0.1700156, -0.0001706459, 0.01524812, 0.05641093, 0.07109457, 0.139452, 
    0.2304746, 0.1657772, 0.1531015, 0.2367455, 0.353082, 0.2808246, 
    0.1809793, 0.2401657, 0.2243724, 0.134845, 0.2421049, 0.2512789, 
    0.2805173, 0.2452083, 0.2206039, 0.2259107, 0.2133086,
  0.2353861, 0.1964625, 0.1890789, 0.2603166, 0.454196, 0.3519894, 0.2102918, 
    0.2134359, 0.02890329, 0.02325383, 0.02536055, 0.0813892, 0.3001151, 
    0.3347844, 0.4289336, 0.2845924, 0.2328846, 0.2179585, 0.2042506, 
    0.4761126, 0.1423261, 0.2208856, 0.2943507, 0.3369861, 0.3702587, 
    0.2851712, 0.1743294, 0.1889098, 0.2377919,
  0.2520787, 0.2149488, 0.3622518, 0.5023961, 0.607686, 0.3925255, 0.5146642, 
    0.5737761, 0.4331524, 0.4908352, 0.3721706, 0.2166166, 0.2307708, 
    0.3691364, 0.479821, 0.2245349, 0.2834832, 0.2351349, 0.307536, 
    0.2857983, 0.2483083, 0.2404935, 0.2139493, 0.2492106, 0.7741309, 
    0.1771584, 0.1399632, 0.2245972, 0.2047534,
  0.2425417, 0.1764276, 0.3375964, 0.4119892, 0.3155079, 0.2975336, 
    0.3830101, 0.5041116, 0.3894807, 0.4204658, 0.4248962, 0.2624349, 
    0.2045383, 0.3362, 0.3878402, 0.2788094, 0.4113594, 0.3285512, 0.1772934, 
    0.2746469, 0.2061988, 0.2621394, 0.2096115, 0.04350674, 0.05149603, 
    0.3629186, 0.3706769, 0.2490879, 0.401705,
  0.1973867, 0.2232805, 0.2555453, 0.2270647, 0.2560999, 0.3762469, 
    0.4531952, 0.4487457, 0.5395094, 0.4784707, 0.4437782, 0.3600214, 
    0.3698128, 0.3734284, 0.3034801, 0.3518832, 0.326066, 0.3451561, 
    0.3384294, 0.3741011, 0.330731, 0.2774691, 0.197684, 0.08132957, 
    0.07821773, 0.05465924, 0.08770791, 0.2050179, 0.2384105,
  0.2843591, 0.2860836, 0.2878081, 0.2895326, 0.2912571, 0.2929816, 
    0.2947061, 0.3003111, 0.3074334, 0.3145557, 0.321678, 0.3288003, 
    0.3359226, 0.3430449, 0.3412363, 0.3355381, 0.3298398, 0.3241416, 
    0.3184433, 0.3127451, 0.3070469, 0.3175291, 0.3143806, 0.311232, 
    0.3080834, 0.3049349, 0.3017863, 0.2986377, 0.2829795,
  0.2259782, 0.2310189, 0.2609324, 0.4154013, 0.3123224, 0.2714005, 
    0.2895287, 0.2807321, 0.3136407, 0.2909812, 0.2728997, 0.2702756, 
    0.3582722, 0.03232784, 0.1186683, 0.1476738, 0.1652296, 0.1809503, 
    0.1603083, 0.1381824, 0.4049187, 0.3472483, 0.1748277, 0.1700433, 
    0.221807, 0.3004754, 0.07173514, 0.1087713, 0.160517,
  0.3247109, 0.2405262, 0.2477636, 0.1120462, 0.1633456, 0.1887084, 
    0.09278839, 0.3245101, 0.3899846, 0.3494474, 0.232519, 0.06797729, 
    0.09141549, 0.1239956, 0.2510346, 0.3570991, 0.3291489, 0.3871374, 
    0.4604256, 0.3218366, 0.4101423, 0.3811728, 0.4266016, 0.3520898, 
    0.2904033, 0.3136715, 0.3213805, 0.3141577, 0.3271687,
  0.4277282, 0.4194194, 0.3804266, 0.4841323, 0.4797004, 0.439597, 0.4806349, 
    0.4296095, 0.4404294, 0.3435405, 0.3997063, 0.4924576, 0.5261393, 
    0.5079587, 0.4222767, 0.4326079, 0.4494405, 0.5192612, 0.4066342, 
    0.3072233, 0.2806024, 0.3184215, 0.3418144, 0.4051892, 0.4607053, 
    0.4574991, 0.5031583, 0.4483001, 0.4610914,
  0.4016294, 0.3925599, 0.4574749, 0.4052837, 0.3702387, 0.3765186, 
    0.3720794, 0.3438245, 0.3353123, 0.3549027, 0.2797484, 0.3931484, 
    0.3279347, 0.3061563, 0.3337896, 0.4089125, 0.382987, 0.4075595, 
    0.3362378, 0.2868506, 0.2285327, 0.304028, 0.2915505, 0.1941886, 
    0.01044243, 0.1524138, 0.3552338, 0.3924336, 0.4181046,
  0.2321881, 0.2485312, 0.1891991, 0.2693272, 0.2357821, 0.2957698, 
    0.2453817, 0.2606371, 0.3364885, 0.2626156, 0.2083169, 0.1238091, 
    0.04304824, 0.1690305, 0.2670032, 0.2594745, 0.2227877, 0.2902318, 
    0.3097325, 0.1777858, 0.2271147, 0.2245481, 0.2579224, 0.02089649, 
    0.02929563, 0.2474596, 0.2407275, 0.2476931, 0.2292946,
  0.1159009, 0.1224923, 0.06344298, 0.07987054, 0.1044127, 0.1092393, 
    0.06177361, 0.09345195, 0.1868453, 0.01457897, 0.02216368, 0.009251143, 
    0.001282461, 0.06553623, 0.1896706, 0.1140345, 0.1691711, 0.1839561, 
    0.1551837, 0.05215552, 0.09865277, 0.04437745, 0.1612759, 0.003907493, 
    0.0208515, 0.1375885, 0.05988832, 0.05561119, 0.07977931,
  0.105712, 0.04952812, 0.01273943, 0.03689428, 0.04638042, 0.01971019, 
    0.05149952, 0.04096362, 0.1139731, 0.06454848, 0.03203248, 0.002273844, 
    0.05966589, 0.03256734, 0.04178622, 0.05970268, 0.07836351, 0.03597417, 
    0.01803029, 0.007989811, 0.009647466, 0.04582363, 0.1966324, 0.2807275, 
    0.04303424, 0.1518831, 0.02412883, 0.01589729, 0.02245518,
  0.2993072, 0.1549788, 0.04117372, 0.05324569, 0.07504918, 0.07143648, 
    0.03427671, 0.02139799, 0.04315296, 0.05858426, 0.04002761, 0.0638976, 
    0.03438224, 0.02801992, 0.05670661, 0.02267412, 0.01715224, 0.01797803, 
    0.01901363, 0.02551993, 0.0385774, 0.07658437, 0.1448907, 0.03528622, 
    0.04706386, 0.0151679, 0.02341902, 0.05213242, 0.1342521,
  0.03863107, 0.004018488, 0.0001725134, 0.006967997, 0.06877439, 0.06169595, 
    0.05748824, 0.05236663, 0.07697855, 0.1095243, 0.03806381, 0.09650028, 
    0.02660193, 0.0352899, 0.03918224, 0.03823781, 0.0405714, 0.02646254, 
    0.03877135, 0.03390183, 0.07027049, 0.1760052, 0.06705849, 0.007424938, 
    0.03102873, 0.06958403, 0.02842074, 0.03873467, 0.1186891,
  -8.544729e-09, 6.655125e-10, 2.822799e-10, -0.001625888, 0.1268519, 
    0.03503823, 0.002633499, 0.03558488, 0.0119242, 0.09641086, 0.1493454, 
    0.03181332, 0.01782469, 0.04042165, 0.03055277, 0.03682069, 0.05578414, 
    0.07856804, 0.08137313, 0.05741117, 0.03768186, 0.03686525, 0.3934948, 
    0.1301109, 0.01543272, 0.02091697, 0.07919718, 0.003033202, -6.079352e-07,
  3.30346e-08, 7.858913e-09, -2.358785e-06, 0.0002338676, -5.239919e-08, 
    0.01243545, 5.256631e-08, 0.0108793, 0.002750858, 0.2904739, 0.1460856, 
    0.08292918, 0.04262619, 0.0617561, 0.0717448, 0.03990435, 0.09204684, 
    0.09335994, 0.0689095, 0.1450938, 0.007148375, 0.2290488, 0.01821514, 
    0.01007905, 0.005128361, 0.01005072, 0.03877317, 0.001317284, 2.513893e-07,
  -1.648607e-05, 0.03682198, 0.01204627, 0.0265296, 0.05100562, 0.01754739, 
    -0.001970922, 0.0001045042, 0.04783041, 0.1893297, 0.1464459, 0.05933242, 
    0.0720047, 0.09562777, 0.1366788, 0.1251018, 0.1502127, 0.1544767, 
    0.0951029, 0.07568338, 0.04944191, 0.2299409, 0.1208161, 0.1666521, 
    0.1738534, 0.1121335, 0.07827312, 0.07691897, 0.00107852,
  0.1016396, 0.01494788, 0.0519207, 0.3193334, 0.03255715, 0.04228303, 
    0.1640007, -0.0001051928, 0.007776179, 0.05650138, 0.08439439, 
    0.09646232, 0.178673, 0.1471855, 0.1338372, 0.1922987, 0.3381439, 
    0.2876249, 0.1676581, 0.2545131, 0.2119872, 0.1595084, 0.2515766, 
    0.2388825, 0.2675251, 0.2071473, 0.204679, 0.1579642, 0.2031513,
  0.2384256, 0.2139231, 0.2219549, 0.3169526, 0.4501317, 0.35454, 0.1827479, 
    0.2155108, 0.0241991, 0.02445399, 0.01527008, 0.07980199, 0.2261115, 
    0.2914219, 0.3428443, 0.1825598, 0.1953599, 0.1990592, 0.1975639, 
    0.481346, 0.1379838, 0.2255874, 0.2538688, 0.3717995, 0.358537, 
    0.1989265, 0.1526398, 0.1705576, 0.2032913,
  0.2382548, 0.2438712, 0.4003673, 0.5956396, 0.6143922, 0.3780578, 
    0.5338041, 0.563181, 0.4168293, 0.4694257, 0.3915245, 0.2691207, 
    0.2352014, 0.3361669, 0.3992784, 0.1903036, 0.3002982, 0.2261517, 
    0.3236862, 0.2982849, 0.3133982, 0.2707095, 0.2216311, 0.2052324, 
    0.7734303, 0.1212787, 0.0982326, 0.2126579, 0.1728215,
  0.1876999, 0.1318067, 0.2996403, 0.3209566, 0.3396352, 0.3233704, 
    0.4451223, 0.5472445, 0.4017666, 0.4440593, 0.4559898, 0.2727142, 
    0.2325092, 0.3556623, 0.4130078, 0.2647389, 0.4846776, 0.3636253, 
    0.2067488, 0.3513462, 0.2067784, 0.3191627, 0.2227536, 0.04112088, 
    0.04953981, 0.3316883, 0.3728947, 0.2492132, 0.3314006,
  0.2206738, 0.3068187, 0.2771748, 0.2385905, 0.2856067, 0.4124877, 
    0.5032447, 0.5077435, 0.5672544, 0.5208822, 0.4729731, 0.4224855, 
    0.4056357, 0.4238416, 0.3565375, 0.4138024, 0.3769037, 0.3815679, 
    0.3748145, 0.4268104, 0.3882862, 0.2894027, 0.2077733, 0.07823623, 
    0.08599246, 0.06386133, 0.06838887, 0.2240233, 0.2716671,
  0.3721125, 0.375854, 0.3795955, 0.3833369, 0.3870784, 0.3908198, 0.3945613, 
    0.4049536, 0.4089568, 0.4129599, 0.4169631, 0.4209663, 0.4249694, 
    0.4289726, 0.4179829, 0.4113497, 0.4047164, 0.3980831, 0.3914498, 
    0.3848165, 0.3781833, 0.3797188, 0.3786075, 0.3774961, 0.3763847, 
    0.3752734, 0.374162, 0.3730506, 0.3691193,
  0.2345239, 0.2649868, 0.3338204, 0.4599279, 0.3441388, 0.2995712, 
    0.3130752, 0.34321, 0.3345089, 0.3524049, 0.3260777, 0.2552454, 
    0.3627951, 0.02037186, 0.1766273, 0.2151313, 0.2664791, 0.1777484, 
    0.1065693, 0.1431667, 0.3907687, 0.3768919, 0.1739551, 0.1659637, 
    0.2316608, 0.2294081, 0.0824948, 0.09070171, 0.130235,
  0.2299009, 0.1942046, 0.2120439, 0.06879978, 0.08821577, 0.1646763, 
    0.07058784, 0.233706, 0.3189546, 0.2991963, 0.2070977, 0.06970023, 
    0.06808387, 0.09001068, 0.2170456, 0.3524304, 0.3202506, 0.368158, 
    0.4261789, 0.2387067, 0.3598948, 0.3599318, 0.4440778, 0.3274193, 
    0.296108, 0.2465457, 0.2552096, 0.2276657, 0.2607139,
  0.4118091, 0.4071546, 0.3384678, 0.4290846, 0.45984, 0.4168008, 0.4730794, 
    0.4021166, 0.3994428, 0.30541, 0.3670443, 0.4681396, 0.5174716, 0.474625, 
    0.4066302, 0.4207653, 0.4420167, 0.507015, 0.3580199, 0.2480976, 
    0.2453507, 0.2919503, 0.3054228, 0.3945388, 0.4244915, 0.4759516, 
    0.5026699, 0.4266812, 0.4185089,
  0.404833, 0.3957711, 0.4804543, 0.4215859, 0.3905229, 0.3629539, 0.3770914, 
    0.3233953, 0.3255283, 0.3216957, 0.2076657, 0.2781423, 0.2697713, 
    0.2575095, 0.2946168, 0.3490181, 0.3296017, 0.3116955, 0.2847274, 
    0.2499842, 0.2018003, 0.2779489, 0.2944063, 0.1769025, 0.01257873, 
    0.2187752, 0.3468497, 0.4022905, 0.417609,
  0.168541, 0.1771055, 0.1151388, 0.2254902, 0.2167826, 0.265915, 0.1973602, 
    0.2401921, 0.2753454, 0.1722946, 0.1021354, 0.06752058, 0.02875664, 
    0.123338, 0.2868395, 0.2293407, 0.162205, 0.2036633, 0.2164203, 
    0.1623278, 0.2173204, 0.2082821, 0.1844501, 0.03048059, 0.03760393, 
    0.2309088, 0.2905726, 0.2252246, 0.1627636,
  0.07173853, 0.06503075, 0.05619697, 0.02592111, 0.1101787, 0.0826513, 
    0.02080253, 0.04246923, 0.1214125, 0.005999436, 0.01270452, 0.004978551, 
    0.0007789053, 0.04035594, 0.1423102, 0.07399528, 0.1552783, 0.1636257, 
    0.08068886, 0.03283341, 0.03833658, 0.01222284, 0.05365457, 0.04200441, 
    0.02434966, 0.1031251, 0.01937273, 0.01299106, 0.04391059,
  0.02805322, 0.09602135, 0.0102229, 0.01505221, 0.01896564, 0.004996104, 
    0.0126314, 0.02247828, 0.0477195, 0.04828374, 0.0248586, 0.0007289548, 
    0.02136273, 0.01051764, 0.01724903, 0.03080485, 0.02695319, 0.01106741, 
    0.002724059, 0.0005688067, 0.0003989363, 0.01033128, 0.05601868, 
    0.1672083, 0.03164357, 0.1400616, 0.004841706, 0.005039797, 0.003809772,
  0.07169886, 0.0788484, 0.03240637, 0.04110837, 0.01568408, 0.01079125, 
    0.01108105, 0.002699225, 0.01373472, 0.01131136, 0.02029347, 0.008887857, 
    0.01870057, 0.007499149, 0.04354761, 0.006280402, 0.00177946, 
    0.003935487, 0.002692578, 0.004636053, 0.00866155, 0.01579557, 
    0.02715901, 0.02590173, 0.03898527, 0.01127317, 0.00105367, 0.007907483, 
    0.02404628,
  0.004873529, 0.004175114, 0.00019897, 0.004350679, 0.04618199, 0.0189489, 
    0.02026491, 0.03438172, 0.04608187, 0.08017179, 0.01366751, 0.02589997, 
    0.005741829, 0.009785929, 0.01401682, 0.009371002, 0.01408395, 
    0.02683353, 0.02879432, 0.02695557, 0.05984621, 0.1930034, 0.1452083, 
    0.003299221, 0.01982679, 0.04795974, 0.008160152, 0.005240241, 0.02083966,
  -1.876255e-09, 5.847514e-10, 2.24658e-10, -0.0008172507, 0.09376364, 
    0.009278772, -0.0004130986, 0.006774984, 0.003036186, 0.04981699, 
    0.1019467, 0.01322936, 0.004506973, 0.01297448, 0.005481532, 0.0107868, 
    0.02781859, 0.05331215, 0.04928174, 0.0419713, 0.01641289, 0.005599997, 
    0.4053682, 0.1263741, 0.003413965, 0.006565718, 0.02811425, 0.0004893638, 
    -2.546712e-06,
  3.039193e-08, 6.292574e-09, -9.321319e-07, 8.414065e-05, -6.893833e-08, 
    0.002624829, 3.728476e-08, 0.006506934, 0.001463056, 0.2331302, 
    0.09972364, 0.04134213, 0.00981966, 0.02064014, 0.03367829, 0.00976552, 
    0.05642237, 0.04367166, 0.02194318, 0.06631532, 0.008205583, 0.1940655, 
    0.004219009, 0.001232926, 0.001364046, 0.004849102, 0.01329833, 
    0.0005014535, 2.315265e-07,
  -6.41552e-06, 0.0182265, 0.006255202, 0.01436144, 0.04462612, 0.01490972, 
    -0.001778274, 6.559139e-05, 0.0309644, 0.2038361, 0.1165673, 0.04129469, 
    0.05496408, 0.08011821, 0.1142032, 0.1933755, 0.1171056, 0.1296146, 
    0.06019511, 0.04190237, 0.04186787, 0.2208557, 0.1194685, 0.2087972, 
    0.08687156, 0.05316687, 0.04077668, 0.03461947, 0.001341953,
  0.07459497, 0.005393597, 0.02648692, 0.3145961, 0.01546224, 0.07756259, 
    0.1597404, -6.66312e-05, 0.006576931, 0.04963364, 0.08646842, 0.07267345, 
    0.1484721, 0.1363631, 0.1097763, 0.1715074, 0.3290754, 0.2708057, 
    0.1479594, 0.2540298, 0.207519, 0.1395693, 0.241442, 0.2041421, 
    0.2131148, 0.1656112, 0.167652, 0.1052491, 0.1632134,
  0.2124915, 0.1856475, 0.2684057, 0.404521, 0.4022476, 0.3641745, 0.1497212, 
    0.1953112, 0.01913006, 0.02224981, 0.007816829, 0.07063497, 0.1812507, 
    0.2711613, 0.2705297, 0.1230771, 0.1588354, 0.1959337, 0.1915971, 
    0.4762107, 0.1346909, 0.2044035, 0.2162298, 0.4153842, 0.3097646, 
    0.1523955, 0.1274335, 0.144439, 0.1748474,
  0.1935165, 0.2768376, 0.4016069, 0.6333668, 0.5694357, 0.3462326, 
    0.5327321, 0.5539646, 0.4263644, 0.4531955, 0.4142762, 0.3353817, 
    0.2311409, 0.3137314, 0.3118467, 0.1924588, 0.3185559, 0.2064771, 
    0.3426719, 0.3126962, 0.3637612, 0.2941756, 0.2454378, 0.1799276, 
    0.7334301, 0.08477136, 0.08086973, 0.179959, 0.139402,
  0.1566678, 0.09638677, 0.2708564, 0.2486961, 0.3770902, 0.3859188, 
    0.534509, 0.5848176, 0.3493167, 0.4578457, 0.5165533, 0.3238165, 
    0.2707302, 0.4029234, 0.4151357, 0.2978481, 0.5318081, 0.36629, 
    0.2538204, 0.4111108, 0.1916598, 0.3511583, 0.2305174, 0.05805274, 
    0.05569354, 0.3040144, 0.3768481, 0.2144568, 0.2828435,
  0.2673992, 0.3671347, 0.3195871, 0.2669946, 0.2966795, 0.4443767, 
    0.5771127, 0.5706401, 0.6135285, 0.5870509, 0.5043485, 0.4813525, 
    0.4664398, 0.4951192, 0.4246193, 0.48524, 0.4317845, 0.4263196, 
    0.4089651, 0.4943221, 0.4361439, 0.2943171, 0.2331353, 0.1060107, 
    0.115063, 0.08023477, 0.0687089, 0.2424668, 0.3239299,
  0.4509113, 0.4582232, 0.4655349, 0.4728467, 0.4801585, 0.4874703, 
    0.4947821, 0.4854176, 0.4891508, 0.4928841, 0.4966173, 0.5003505, 
    0.5040838, 0.507817, 0.4895454, 0.4792064, 0.4688672, 0.4585281, 
    0.448189, 0.4378499, 0.4275108, 0.4321793, 0.4314734, 0.4307675, 
    0.4300616, 0.4293556, 0.4286497, 0.4279438, 0.4450619,
  0.2192344, 0.2967325, 0.4021227, 0.4799689, 0.3707142, 0.3074282, 
    0.3407631, 0.4057552, 0.3664534, 0.3725099, 0.2817661, 0.2141372, 
    0.3387486, 0.01313214, 0.2158997, 0.2111327, 0.3606288, 0.1955106, 
    0.08661009, 0.1404513, 0.3756703, 0.3875699, 0.161363, 0.1462334, 
    0.2218666, 0.1916067, 0.07754007, 0.07097164, 0.1075491,
  0.1570158, 0.1193061, 0.1479727, 0.04311201, 0.04669952, 0.1402501, 
    0.04439515, 0.153087, 0.2424316, 0.2348825, 0.1683168, 0.06681297, 
    0.04579045, 0.06715706, 0.1850047, 0.3172673, 0.294091, 0.3034771, 
    0.3580565, 0.2029553, 0.3019127, 0.3382265, 0.4377194, 0.2778071, 
    0.2582483, 0.2126847, 0.2346666, 0.1804285, 0.2056337,
  0.3547701, 0.3464182, 0.2816942, 0.3677568, 0.4177732, 0.3750495, 
    0.4339062, 0.3428361, 0.3433115, 0.277979, 0.3225152, 0.4377717, 
    0.4969774, 0.447749, 0.359663, 0.3968174, 0.4185474, 0.467798, 0.3221259, 
    0.2087532, 0.2148121, 0.2375282, 0.2529178, 0.3406275, 0.386356, 
    0.4601495, 0.4847601, 0.3865862, 0.3692537,
  0.3702717, 0.3573735, 0.4169765, 0.3586429, 0.3718166, 0.364863, 0.3735399, 
    0.2775267, 0.2943678, 0.2775972, 0.1677224, 0.2070315, 0.2301492, 
    0.2310681, 0.2621957, 0.2917749, 0.2528204, 0.2242624, 0.2390002, 
    0.2064613, 0.1661466, 0.2297715, 0.2584591, 0.1452577, 0.03713202, 
    0.2333849, 0.3092551, 0.3742462, 0.4034648,
  0.1311311, 0.1098071, 0.06329883, 0.181199, 0.1652898, 0.2264875, 
    0.1618606, 0.2186981, 0.2086549, 0.117464, 0.05615452, 0.03616866, 
    0.02411973, 0.08489722, 0.2843689, 0.1852973, 0.1046038, 0.1634464, 
    0.1548217, 0.1334508, 0.1791961, 0.1538485, 0.1112216, 0.04115107, 
    0.0343663, 0.1917889, 0.2813818, 0.1813388, 0.1158259,
  0.03239731, 0.02753979, 0.04781349, 0.009165134, 0.06950317, 0.05789459, 
    0.004841577, 0.01442982, 0.04651359, 0.006177319, 0.006700705, 
    0.002794882, 0.001983079, 0.02882804, 0.08732726, 0.0429299, 0.13366, 
    0.1310333, 0.0515978, 0.01704263, 0.01128819, 0.00444514, 0.01878184, 
    0.06134234, 0.0202191, 0.06129938, 0.005659156, 0.002103854, 0.02075845,
  0.008257125, 0.1205115, 0.006171202, 0.004982451, 0.004719146, 0.001540626, 
    0.004315166, 0.01308528, 0.01515099, 0.03144608, 0.01826829, 
    0.0001606983, 0.006190439, 0.004273996, 0.006814799, 0.01256892, 
    0.01082482, 0.004766707, 0.0002407294, 0.0001083607, 8.177891e-05, 
    0.002960745, 0.01885885, 0.0571052, 0.02320529, 0.1258792, 0.001704609, 
    0.0005808336, 0.000928989,
  0.02593285, 0.02266107, 0.02871101, 0.03370046, 0.003668922, 0.002356307, 
    0.00593212, 0.0005370444, 0.003463767, 0.0009688449, 0.008663838, 
    0.002260669, 0.003724312, 0.0007068586, 0.02533841, 0.002872443, 
    0.0002429366, 0.001063067, 0.0007620162, 0.001158316, 0.002955905, 
    0.005196531, 0.008982833, 0.02510933, 0.03552381, 0.00572564, 
    -0.0006476067, 0.002542143, 0.008021557,
  0.001042055, 0.004167917, 0.0001694416, 0.003949851, 0.02378988, 
    0.009131146, 0.01590523, 0.01967504, 0.02931184, 0.06732449, 0.001717711, 
    0.004542173, 0.000927515, 0.004497709, 0.009856279, 0.002066337, 
    0.001360672, 0.004550336, 0.008574903, 0.00557078, 0.01551787, 
    0.04032652, 0.0481381, 0.001507843, 0.01303014, 0.02462843, 0.001377809, 
    0.001433152, 0.005155993,
  -4.552027e-09, 5.581292e-10, 1.89192e-10, -0.0004574187, 0.04769286, 
    0.003023584, -0.001380549, 0.00248642, 0.0004012456, 0.01610612, 
    0.05242104, 0.004093464, 0.001119817, 0.003534026, 0.000680915, 
    0.003678063, 0.01236087, 0.021027, 0.02219854, 0.01459678, 0.006225037, 
    0.001299242, 0.3000228, 0.1084761, 0.0009678272, 0.00270363, 0.01294312, 
    0.0001275145, -1.653629e-05,
  2.868836e-08, 5.531254e-09, -2.716599e-07, 5.408712e-05, -5.261548e-08, 
    0.0009221014, 2.662963e-08, 0.003173083, 0.001013278, 0.1672005, 
    0.0554003, 0.01814036, 0.004076119, 0.007268979, 0.0123289, 0.003136931, 
    0.03211055, 0.0160328, 0.008517123, 0.03187725, 0.01208932, 0.1512725, 
    0.001170397, -0.001027689, 0.0006017475, 0.002719977, 0.0066072, 
    0.0002503977, 2.1384e-07,
  -8.250969e-06, 0.009883731, 0.003141273, 0.006791511, 0.03975612, 
    0.0116177, -0.00153964, 0.0001017801, 0.0220309, 0.1883923, 0.09317333, 
    0.03007267, 0.03518656, 0.06103112, 0.09181914, 0.1709788, 0.07718848, 
    0.1048057, 0.04529849, 0.02236397, 0.03237705, 0.1916215, 0.09889149, 
    0.1482464, 0.04580246, 0.02514143, 0.01830719, 0.01550611, 0.0009563366,
  0.05498819, 0.001995619, 0.0162509, 0.2981558, 0.007857027, 0.07047135, 
    0.1527274, -3.006805e-05, 0.006554928, 0.03322436, 0.08180238, 
    0.05622279, 0.1194268, 0.1170715, 0.08359624, 0.1456355, 0.2809401, 
    0.2240175, 0.1131335, 0.245003, 0.1884645, 0.1102628, 0.2047478, 
    0.1918648, 0.1573308, 0.1118451, 0.1107523, 0.06237546, 0.1295326,
  0.1560815, 0.158854, 0.243433, 0.4090328, 0.3719476, 0.3112379, 0.1097545, 
    0.16615, 0.01853339, 0.02047309, 0.003651233, 0.0683047, 0.1651489, 
    0.2326247, 0.2194067, 0.0921976, 0.125944, 0.1756156, 0.1666238, 
    0.4569818, 0.1216349, 0.1703317, 0.1831741, 0.4056268, 0.2625331, 
    0.1220792, 0.1022836, 0.1140362, 0.1255936,
  0.1434326, 0.3223909, 0.4005887, 0.5978842, 0.5307878, 0.3529395, 
    0.4904151, 0.4917396, 0.41079, 0.4170637, 0.4037313, 0.3846622, 
    0.2154539, 0.2858456, 0.2483818, 0.2167043, 0.3308569, 0.2056959, 
    0.3405411, 0.2979965, 0.3851094, 0.2552377, 0.2723879, 0.1686188, 
    0.6997297, 0.0611369, 0.06929592, 0.1392178, 0.0985543,
  0.1296908, 0.07084277, 0.2606985, 0.1736754, 0.4563186, 0.4482527, 
    0.6249803, 0.5382048, 0.3180059, 0.4975719, 0.5805702, 0.3583233, 
    0.3303837, 0.4549277, 0.4001573, 0.3787003, 0.5263046, 0.341866, 
    0.2794315, 0.4450802, 0.1809679, 0.3975889, 0.2481343, 0.1080351, 
    0.06695037, 0.2754186, 0.3805444, 0.1802006, 0.2338087,
  0.3545144, 0.4354071, 0.3687741, 0.2990654, 0.2781829, 0.4826212, 
    0.6083332, 0.6245704, 0.6786662, 0.6472104, 0.6199117, 0.5890805, 
    0.5761176, 0.599991, 0.5612314, 0.5629439, 0.5197514, 0.5092425, 
    0.5344599, 0.5581849, 0.5288039, 0.3060342, 0.235912, 0.1619374, 
    0.139804, 0.1031601, 0.04939, 0.2777615, 0.4236092,
  0.4762921, 0.4842118, 0.4921315, 0.5000511, 0.5079708, 0.5158905, 
    0.5238101, 0.477221, 0.4855211, 0.4938213, 0.5021214, 0.5104215, 
    0.5187216, 0.5270218, 0.5808916, 0.5681472, 0.5554029, 0.5426586, 
    0.5299142, 0.5171699, 0.5044255, 0.4933129, 0.4898374, 0.486362, 
    0.4828865, 0.479411, 0.4759356, 0.4724601, 0.4699564,
  0.1979804, 0.2901727, 0.3671052, 0.5139803, 0.4331201, 0.28971, 0.351121, 
    0.4574244, 0.2705048, 0.2666203, 0.2255228, 0.1722456, 0.270982, 
    0.006369411, 0.2124331, 0.3078359, 0.3156955, 0.2128007, 0.06319396, 
    0.1796651, 0.3514475, 0.3939229, 0.1248845, 0.09568384, 0.1873153, 
    0.1838584, 0.09005646, 0.05400863, 0.08745623,
  0.1065015, 0.0752386, 0.09436469, 0.02686879, 0.02522016, 0.1143943, 
    0.03027568, 0.09370831, 0.1716937, 0.1786489, 0.1181113, 0.06656957, 
    0.02979674, 0.05014564, 0.1549114, 0.2738333, 0.2356485, 0.2359693, 
    0.2879882, 0.1643013, 0.2539349, 0.2958225, 0.4265231, 0.2142619, 
    0.206626, 0.1882778, 0.1802798, 0.1289228, 0.1572607,
  0.2638648, 0.2712947, 0.2263346, 0.3108345, 0.3398099, 0.3046148, 0.342139, 
    0.2719027, 0.2893219, 0.2444168, 0.2795782, 0.3843209, 0.4461286, 
    0.3839906, 0.2974471, 0.3328201, 0.3596463, 0.4011527, 0.2769171, 
    0.1658762, 0.1763826, 0.1871097, 0.1838599, 0.270676, 0.3427838, 
    0.4235094, 0.4386097, 0.3319006, 0.3080081,
  0.2902571, 0.2710596, 0.3234742, 0.2771297, 0.3013002, 0.3181707, 
    0.3176809, 0.2236303, 0.2292568, 0.2190038, 0.1213067, 0.1467503, 
    0.1785362, 0.1892319, 0.2383071, 0.262016, 0.2205399, 0.1678205, 
    0.1745123, 0.1552421, 0.1176972, 0.1711105, 0.1973566, 0.1134339, 
    0.04402521, 0.2090481, 0.275132, 0.3091928, 0.3377145,
  0.09402421, 0.06781942, 0.0405977, 0.1375767, 0.1184378, 0.1847442, 
    0.1132861, 0.190588, 0.1595323, 0.08498853, 0.0339166, 0.0194691, 
    0.01772108, 0.05622378, 0.252025, 0.1380583, 0.08538566, 0.1408452, 
    0.1250397, 0.09430926, 0.1300013, 0.09428765, 0.06729382, 0.04639122, 
    0.04023235, 0.1416452, 0.2225335, 0.133677, 0.07839164,
  0.01642555, 0.0128583, 0.03753067, 0.003710715, 0.03037873, 0.03590931, 
    0.001823499, 0.006772751, 0.0217141, 0.001653656, 0.002929963, 
    0.001475236, 0.0008950492, 0.01935857, 0.0535771, 0.02927585, 0.1040916, 
    0.111875, 0.03907221, 0.008433993, 0.005086142, 0.002420675, 0.009722706, 
    0.04746881, 0.01538798, 0.02933096, 0.002111099, 0.000697517, 0.006937139,
  0.003882163, 0.1130395, 0.003327826, 0.001910903, 0.000674889, 
    0.0005379381, 0.001801442, 0.006477697, 0.007158445, 0.01495465, 
    0.0131187, 8.253415e-05, 0.002007366, 0.001802298, 0.002827129, 
    0.005616699, 0.005771524, 0.001397313, 6.619156e-05, 3.057296e-05, 
    3.486295e-05, 0.001238025, 0.008918381, 0.03037296, 0.01647757, 
    0.1077426, 0.0009453965, 0.000235748, 0.0004425063,
  0.01369942, 0.008341706, 0.02846764, 0.02714977, 0.001392483, 0.001136872, 
    0.005243241, 0.000216568, 0.001767878, -0.0001923525, 0.003737895, 
    0.001038254, 0.0008673671, 0.0001212578, 0.01482876, 0.001359441, 
    0.0001043928, 0.0005787646, 0.0003831653, 0.0006053813, 0.001666199, 
    0.002675749, 0.00465659, 0.02804019, 0.03621506, 0.004334503, 
    -0.0002618168, 0.001351694, 0.004268633,
  0.000483881, 0.002940093, 0.0001802342, 0.004917193, 0.01262953, 
    0.006077123, 0.01281684, 0.01022284, 0.02746522, 0.0619684, 0.0006490532, 
    0.001766574, 0.0003289087, 0.003703007, 0.01054107, 0.0005696168, 
    0.0004197598, 0.0004089182, 0.003399189, 0.0007179807, 0.00453674, 
    0.01275284, 0.01451018, 0.0006203548, 0.008642379, 0.009549115, 
    0.0003163496, 0.0007962394, 0.002608876,
  1.451475e-10, 5.482352e-10, 1.720608e-10, 0.001041468, 0.02548494, 
    0.001501716, -0.001655437, 0.001431961, 0.0001585702, 0.006925384, 
    0.0230346, 0.0008388418, 0.0003825524, 0.001050251, 0.0003580655, 
    0.001464223, 0.004704332, 0.01118028, 0.008941432, 0.005346743, 
    0.0021207, 0.0006364553, 0.2031998, 0.08537063, 0.0002342853, 0.00147661, 
    0.007247447, 5.042519e-05, -6.008645e-05,
  2.679925e-08, 5.224309e-09, -1.092829e-07, 3.825914e-05, -3.913712e-08, 
    0.0005193492, 1.971082e-08, 0.001067798, 0.0008283467, 0.1059559, 
    0.02750586, 0.008712399, 0.002663281, 0.003372655, 0.004468806, 
    0.001759911, 0.01850569, 0.007467382, 0.004701493, 0.01802183, 
    0.005983361, 0.1201058, 0.0005500272, -0.0008944634, 0.0001993242, 
    0.001251298, 0.003998199, 0.0001504626, 2.027425e-07,
  -4.437545e-06, 0.005870233, 0.001659933, 0.003431433, 0.03483315, 
    0.008370182, -0.001332513, 0.000257384, 0.01712882, 0.1536256, 
    0.06861506, 0.01575647, 0.02113882, 0.04024668, 0.0664956, 0.09131376, 
    0.05033306, 0.07898821, 0.02834613, 0.01242365, 0.02582436, 0.1505708, 
    0.07311013, 0.06010049, 0.02571267, 0.0134553, 0.00960137, 0.007133916, 
    0.001101234,
  0.04090454, 0.001075306, 0.01404783, 0.2762342, 0.004831324, 0.05461416, 
    0.1434538, -1.691641e-05, 0.006198934, 0.02782389, 0.07441714, 
    0.04285038, 0.09336114, 0.09885053, 0.06182222, 0.1135485, 0.2102858, 
    0.1719348, 0.07518855, 0.2260259, 0.1601138, 0.08781147, 0.1634307, 
    0.1688076, 0.1109571, 0.07405125, 0.06609204, 0.03507151, 0.09306216,
  0.1350358, 0.1423799, 0.2100642, 0.3779926, 0.3050067, 0.2430371, 
    0.07901645, 0.1440323, 0.02042069, 0.02369911, 0.002291554, 0.06827685, 
    0.1586159, 0.1852122, 0.1824428, 0.07140516, 0.1051991, 0.1468537, 
    0.1314161, 0.4341263, 0.09805301, 0.1253311, 0.1491216, 0.3858114, 
    0.2100293, 0.1009705, 0.07997082, 0.07759973, 0.0873166,
  0.1010027, 0.3362389, 0.3571648, 0.5302272, 0.4746698, 0.3556476, 0.422371, 
    0.4021084, 0.364633, 0.3488105, 0.378931, 0.4397457, 0.196037, 0.2666883, 
    0.2111535, 0.2199586, 0.3556004, 0.1912407, 0.3028086, 0.3067268, 
    0.3807851, 0.2071667, 0.2699026, 0.1391584, 0.6764414, 0.04509303, 
    0.05870022, 0.0989143, 0.06447938,
  0.1019758, 0.05146838, 0.2558339, 0.1239532, 0.5115471, 0.4402061, 
    0.7081858, 0.5282651, 0.3323679, 0.5321852, 0.6601213, 0.3521423, 
    0.5057646, 0.4487954, 0.403329, 0.4159747, 0.4728377, 0.3036006, 
    0.3276974, 0.4244354, 0.2603273, 0.5202664, 0.3041613, 0.1734233, 
    0.09177853, 0.2351777, 0.3885637, 0.1473107, 0.1941044,
  0.4605963, 0.4337806, 0.4861775, 0.3516136, 0.3453415, 0.58187, 0.6661489, 
    0.6249152, 0.6250718, 0.6711715, 0.6798408, 0.6153797, 0.5919825, 
    0.6298006, 0.5844802, 0.6485673, 0.6172345, 0.6413789, 0.5812573, 
    0.580682, 0.6032213, 0.2640893, 0.2412727, 0.2190996, 0.1184305, 
    0.1201763, 0.04056093, 0.2785147, 0.4818441,
  0.419843, 0.4275108, 0.4351785, 0.4428463, 0.450514, 0.4581818, 0.4658496, 
    0.4028049, 0.4161991, 0.4295933, 0.4429875, 0.4563817, 0.4697759, 
    0.4831702, 0.6095927, 0.5939652, 0.5783377, 0.5627102, 0.5470827, 
    0.5314551, 0.5158276, 0.4674947, 0.4620602, 0.4566258, 0.4511913, 
    0.4457568, 0.4403224, 0.4348879, 0.4137088,
  0.1765084, 0.2393865, 0.2944548, 0.4872611, 0.4934442, 0.2445586, 
    0.3136608, 0.4096809, 0.2224359, 0.1803663, 0.1442727, 0.1222489, 
    0.1847959, 0.004507977, 0.2107945, 0.3038504, 0.2430915, 0.2006798, 
    0.06109885, 0.2036714, 0.3193674, 0.3670902, 0.09761033, 0.07102807, 
    0.1537842, 0.1716166, 0.113139, 0.03782993, 0.07348779,
  0.07007163, 0.05474846, 0.06197003, 0.01941335, 0.01618016, 0.09624344, 
    0.02139976, 0.06104506, 0.1333768, 0.1410157, 0.09102358, 0.06474767, 
    0.01883283, 0.03267557, 0.1223197, 0.2157125, 0.1751909, 0.1800458, 
    0.2251061, 0.1278231, 0.1937182, 0.2399161, 0.3723406, 0.1680222, 
    0.1741213, 0.1540281, 0.1386865, 0.08443211, 0.1090099,
  0.1819645, 0.19694, 0.1706901, 0.24428, 0.2607728, 0.2210449, 0.2461347, 
    0.2045501, 0.2247664, 0.1889133, 0.2135153, 0.2886083, 0.3528108, 
    0.2930708, 0.2276956, 0.2559909, 0.2867036, 0.3332524, 0.2227613, 
    0.1237116, 0.1236349, 0.1286802, 0.1188512, 0.1928786, 0.2804741, 
    0.3663332, 0.3605928, 0.2551907, 0.2260255,
  0.2060118, 0.1907873, 0.2404376, 0.2067589, 0.2360222, 0.2557449, 
    0.2493924, 0.1650171, 0.161184, 0.1511636, 0.07778629, 0.09384182, 
    0.1235253, 0.1331101, 0.2046639, 0.21384, 0.1645726, 0.1213728, 
    0.1189022, 0.1016771, 0.07638488, 0.1184411, 0.1352874, 0.08867141, 
    0.03996219, 0.1674207, 0.2329459, 0.2385732, 0.260224,
  0.06130784, 0.04420653, 0.02739671, 0.09355716, 0.08471207, 0.1230519, 
    0.07995883, 0.1542513, 0.114703, 0.05492426, 0.02155844, 0.01102025, 
    0.01082174, 0.03214849, 0.2133703, 0.08488785, 0.06119706, 0.1113143, 
    0.09357952, 0.0592288, 0.08985232, 0.05345518, 0.03146303, 0.05200291, 
    0.03052748, 0.09276158, 0.1642453, 0.08406125, 0.04891744,
  0.007643622, 0.006239424, 0.02506888, 0.001637912, 0.0167177, 0.0211341, 
    0.001122824, 0.004221191, 0.0134042, 0.0007771869, 0.00147397, 
    0.0008017518, -0.0001431107, 0.008575028, 0.02814789, 0.01651551, 
    0.06798755, 0.07848635, 0.02860299, 0.004549127, 0.003075387, 
    0.001619377, 0.006234117, 0.02826987, 0.01108135, 0.009427797, 
    0.001150864, 0.0003940153, 0.00232391,
  0.002357987, 0.08483809, 0.001167459, 0.0007725898, -0.0005936432, 
    0.0002489182, 0.001052053, 0.002530639, 0.004363109, 0.008324286, 
    0.008027561, -1.811946e-05, 0.0008462337, 0.0009034655, 0.00136957, 
    0.002813229, 0.003064972, 0.0005583105, 3.653741e-05, 1.433656e-05, 
    2.05523e-05, 0.0006760357, 0.00528627, 0.02015647, 0.01113682, 
    0.08122299, 0.0006248502, 0.0001459475, 0.000268891,
  0.008892361, 0.004519145, 0.02592176, 0.0232325, 0.000773291, 0.0007052928, 
    0.003330494, 0.0001345711, 0.0008216772, -8.983174e-05, 0.001104676, 
    0.000605773, 0.0002515298, 7.311342e-05, 0.006804935, 0.000653467, 
    6.837286e-05, 0.0003873713, 0.0002365112, 0.0003840283, 0.001113067, 
    0.00169808, 0.002982441, 0.02091471, 0.03846994, 0.003545929, 
    -8.190505e-05, 0.0008766559, 0.002778959,
  0.0002864463, 0.002880264, 0.0001816175, 0.004338889, 0.005603223, 
    0.003376832, 0.007545541, 0.004659566, 0.02857598, 0.06552779, 
    0.0003489465, 0.001034174, 0.0001983713, 0.002049546, 0.006613838, 
    0.0002890205, 0.0002535547, 0.0001391594, 0.001106463, 0.0002715179, 
    0.001997678, 0.006476757, 0.006570654, 0.0007411534, 0.004797912, 
    0.003719145, 0.0001163421, 0.000535989, 0.001652798,
  4.780574e-10, 5.433145e-10, 1.605144e-10, 0.001307977, 0.01551048, 
    0.0009887951, -0.001290254, 0.0009806361, 8.206148e-05, 0.003223738, 
    0.009583334, 0.0002397973, 0.0001828003, 0.0005652565, 0.0002588488, 
    0.0007076895, 0.00206137, 0.005694333, 0.003343304, 0.00201638, 
    0.0007328936, 0.0003926918, 0.1655898, 0.06344478, 5.233421e-05, 
    0.0009034429, 0.004754003, 2.872732e-05, -0.0002174434,
  2.595908e-08, 5.118376e-09, -6.338415e-08, 2.878994e-05, -3.971844e-08, 
    0.0003595329, 1.6882e-08, 0.0003891708, 0.000347531, 0.06015353, 
    0.01150853, 0.00406094, 0.001910998, 0.002138221, 0.002268889, 
    0.001209429, 0.009218162, 0.00406463, 0.003124054, 0.01189794, 
    0.002922205, 0.09823605, 0.0003355207, -0.0007942365, 9.268981e-05, 
    0.0006660213, 0.002816786, 0.0001031825, 1.959874e-07,
  -2.335623e-06, 0.004381191, 0.001063815, 0.002438441, 0.02909327, 
    0.005604361, -0.001153607, 0.001520987, 0.01598335, 0.1141722, 
    0.05155224, 0.009510074, 0.01166433, 0.02473339, 0.03881066, 0.05331768, 
    0.03089506, 0.05554689, 0.01521112, 0.00600663, 0.0203397, 0.1136234, 
    0.05279775, 0.02956815, 0.01400512, 0.008204577, 0.005371912, 
    0.004199076, 0.001190746,
  0.02933468, 0.0005426722, 0.0116651, 0.259627, 0.003557541, 0.04302893, 
    0.1335785, -1.049362e-05, 0.005544919, 0.02956193, 0.0608618, 0.03419825, 
    0.07234072, 0.07600426, 0.04014975, 0.07990433, 0.1465498, 0.1169038, 
    0.04257027, 0.2048585, 0.1346422, 0.06778668, 0.1354555, 0.1493195, 
    0.08013958, 0.04764558, 0.0380698, 0.01844534, 0.06179189,
  0.1094875, 0.1270737, 0.1741552, 0.33284, 0.2376796, 0.1813371, 0.05911141, 
    0.1263773, 0.02906473, 0.02834147, 0.002593242, 0.07475104, 0.1477084, 
    0.1418842, 0.1488415, 0.05626817, 0.08437885, 0.1099418, 0.08980494, 
    0.4023613, 0.07669772, 0.09151418, 0.1091465, 0.3526087, 0.172844, 
    0.08586995, 0.05940254, 0.05018716, 0.06177799,
  0.07601494, 0.3244647, 0.3024166, 0.4624096, 0.4113944, 0.3115414, 
    0.3486106, 0.3414164, 0.3029987, 0.2911101, 0.3312855, 0.4814755, 
    0.2127017, 0.2360232, 0.1860542, 0.2135095, 0.3822103, 0.1830729, 
    0.2807761, 0.3088745, 0.3749661, 0.2225851, 0.2294061, 0.150335, 
    0.6596532, 0.03520935, 0.04797477, 0.07015291, 0.04192853,
  0.07717779, 0.0371908, 0.2576098, 0.0955766, 0.4853028, 0.4147561, 
    0.6971544, 0.4876836, 0.396776, 0.5918276, 0.6712739, 0.3557444, 
    0.6846224, 0.3384481, 0.3672777, 0.4046895, 0.4350114, 0.2604521, 
    0.380157, 0.3733575, 0.271414, 0.5583488, 0.4430289, 0.2486759, 
    0.1055882, 0.1822838, 0.4017856, 0.1237928, 0.1558849,
  0.544834, 0.4793344, 0.5339175, 0.3585035, 0.3964221, 0.605009, 0.6091037, 
    0.5829172, 0.598263, 0.5360218, 0.5907986, 0.5650085, 0.5328221, 
    0.5194927, 0.5538989, 0.5536578, 0.5883325, 0.5889397, 0.5298798, 
    0.5521792, 0.5510452, 0.2479393, 0.2342892, 0.2821897, 0.1031266, 
    0.0920203, 0.03569971, 0.2579195, 0.4610005,
  0.3043083, 0.309477, 0.3146457, 0.3198144, 0.3249832, 0.3301519, 0.3353206, 
    0.2958811, 0.3070386, 0.318196, 0.3293535, 0.3405109, 0.3516684, 
    0.3628258, 0.4772877, 0.4678198, 0.4583519, 0.4488841, 0.4394162, 
    0.4299483, 0.4204804, 0.3570853, 0.350227, 0.3433686, 0.3365104, 
    0.3296521, 0.3227938, 0.3159355, 0.3001733,
  0.156468, 0.1878448, 0.2280992, 0.406122, 0.4352266, 0.212728, 0.2437721, 
    0.3032909, 0.1702685, 0.1074253, 0.08828159, 0.09485377, 0.1368496, 
    0.001853151, 0.205339, 0.2814031, 0.2059685, 0.1676745, 0.04542178, 
    0.2042069, 0.2709998, 0.3405356, 0.0802184, 0.06183476, 0.129738, 
    0.1632224, 0.1367622, 0.03126356, 0.07202077,
  0.05618785, 0.03984843, 0.04738729, 0.01422584, 0.01300285, 0.08446408, 
    0.0174868, 0.04746772, 0.1116492, 0.1222508, 0.08050847, 0.06204309, 
    0.01530364, 0.02161661, 0.09038328, 0.1709197, 0.1347927, 0.1425067, 
    0.1740034, 0.1038531, 0.1469462, 0.1867637, 0.3126043, 0.1357882, 
    0.1484025, 0.123478, 0.1118235, 0.06000181, 0.07946694,
  0.1408628, 0.1554224, 0.1317726, 0.2041852, 0.2063182, 0.1728954, 0.192431, 
    0.1597562, 0.178929, 0.1530729, 0.1605734, 0.2169677, 0.2745731, 
    0.2302814, 0.1779364, 0.2005764, 0.2338807, 0.279018, 0.1831549, 
    0.09716383, 0.08918548, 0.08808471, 0.08071552, 0.1343437, 0.2226443, 
    0.2933896, 0.2938591, 0.2045287, 0.1776238,
  0.1565817, 0.1445766, 0.1877688, 0.1637498, 0.1903861, 0.2093133, 
    0.1960836, 0.1276387, 0.1191218, 0.109041, 0.05337073, 0.06152921, 
    0.08070789, 0.09516545, 0.16975, 0.1580232, 0.1133907, 0.088504, 
    0.08505917, 0.07054021, 0.05250093, 0.08735803, 0.1004431, 0.07498044, 
    0.03238941, 0.1265281, 0.1985569, 0.1907454, 0.2094424,
  0.04093284, 0.02975396, 0.01804713, 0.05869479, 0.06022095, 0.07757856, 
    0.05695889, 0.1183019, 0.0737128, 0.03471997, 0.01452349, 0.007145096, 
    0.007563422, 0.01844393, 0.1814705, 0.05317132, 0.03627673, 0.08274025, 
    0.0644238, 0.03894361, 0.05827405, 0.03311624, 0.01564427, 0.05701226, 
    0.02099153, 0.06184975, 0.1126769, 0.05451946, 0.03188264,
  0.004423083, 0.003487368, 0.01648849, 0.001137976, 0.009753566, 0.01146219, 
    0.0008499504, 0.003102529, 0.009803778, 0.0004831044, 0.0007853063, 
    0.0005226224, 0.0001442258, 0.004802988, 0.01552045, 0.009575431, 
    0.03986786, 0.04791948, 0.02041347, 0.002628872, 0.002236035, 
    0.001221615, 0.004583814, 0.02077476, 0.008655287, 0.004065606, 
    0.0008005531, 0.0002788435, 0.00125749,
  0.001662165, 0.06262996, 0.0005870964, 0.0004434224, -0.0007054717, 
    0.000161453, 0.0007389284, 0.001183752, 0.003112862, 0.005506219, 
    0.004390279, 2.867649e-05, 0.0005591454, 0.0005695336, 0.0006530193, 
    0.001594072, 0.001748834, 0.0003234875, 2.648787e-05, 1.011776e-05, 
    1.443601e-05, 0.0004435328, 0.003682198, 0.01519391, 0.007187103, 
    0.05930882, 0.0004640266, 0.0001055026, 0.0001902931,
  0.006564, 0.003106167, 0.02912633, 0.03105311, 0.0005298102, 0.0004957163, 
    0.00178454, 0.000100812, 0.0005507801, 6.773876e-05, 0.0005089276, 
    0.000429997, 0.0001062191, 5.116526e-05, 0.00311851, 0.0003734837, 
    5.085423e-05, 0.0002916543, 0.0001876876, 0.0002787494, 0.0008371663, 
    0.001236397, 0.002183607, 0.01729569, 0.03122282, 0.005336431, 
    -3.972533e-05, 0.0006470479, 0.002055614,
  0.0001992724, 0.01224785, 0.0004370474, 0.004646512, 0.002506088, 
    0.001652427, 0.003911417, 0.002302782, 0.03312358, 0.06682374, 
    0.0002308766, 0.0007228857, 0.000152283, 0.001117046, 0.003157576, 
    0.000179708, 0.0001838646, 7.874364e-05, 0.0004885248, 0.0001302927, 
    0.001020923, 0.004210918, 0.003877259, 0.003091085, 0.0031769, 
    0.001647233, 6.632982e-05, 0.0004063716, 0.001200574,
  5.200849e-10, 5.392831e-10, 1.505937e-10, 0.002425899, 0.01010763, 
    0.0007363809, -0.000911574, 0.0007409949, 1.019834e-05, 0.001661777, 
    0.00429945, 0.0001221967, 0.0001268244, 0.000385129, 0.0001943227, 
    0.0004380321, 0.0009756802, 0.00293219, 0.001509434, 0.0009727831, 
    0.0003286675, 0.0002800748, 0.1222898, 0.04390734, 3.094222e-05, 
    0.0006331784, 0.003525894, 1.960418e-05, -0.0003400941,
  2.528918e-08, 5.091563e-09, -4.417841e-08, 2.396639e-05, -3.275905e-08, 
    0.0002792352, 1.498976e-08, 0.0002219112, 0.0002131064, 0.03677936, 
    0.005967762, 0.002254612, 0.001388153, 0.001590302, 0.001550155, 
    0.0009340993, 0.004402291, 0.002772391, 0.002350298, 0.008885888, 
    0.001714024, 0.0821947, 0.0002477908, -0.000745612, 6.438365e-05, 
    0.000467173, 0.002192776, 7.911817e-05, 1.93376e-07,
  -1.744722e-06, 0.003911971, 0.0009206774, 0.001977181, 0.02490947, 
    0.003585326, -0.001030608, 0.01545419, 0.01677314, 0.08776157, 
    0.03790526, 0.006098268, 0.006289402, 0.01573558, 0.02311482, 0.02991821, 
    0.01883574, 0.03381482, 0.008220262, 0.00317185, 0.01641126, 0.08824624, 
    0.04290134, 0.01760623, 0.008353812, 0.005761916, 0.003902384, 
    0.002923013, 0.0007725056,
  0.02049607, 0.0003179436, 0.01019334, 0.240939, 0.00290384, 0.03654461, 
    0.1283889, -6.328173e-06, 0.003603611, 0.03527464, 0.05341191, 
    0.02995251, 0.05704307, 0.05869859, 0.02631128, 0.05467435, 0.106069, 
    0.08256003, 0.02472341, 0.1857678, 0.1254289, 0.05770793, 0.1184996, 
    0.1357324, 0.06006964, 0.03252653, 0.02310207, 0.01092068, 0.04328438,
  0.09334114, 0.114787, 0.1552362, 0.3023342, 0.2057333, 0.1680324, 
    0.05108472, 0.1327502, 0.05627616, 0.02985726, 0.004692679, 0.08205387, 
    0.1386075, 0.1177236, 0.1252472, 0.0463348, 0.06871431, 0.08387014, 
    0.0665729, 0.3798369, 0.06634545, 0.07202373, 0.09073028, 0.3070695, 
    0.1510457, 0.07426784, 0.04616454, 0.03582754, 0.0476069,
  0.06224651, 0.3244811, 0.2696152, 0.4228882, 0.3648157, 0.2688351, 
    0.2913696, 0.2984504, 0.2491203, 0.2477913, 0.3039692, 0.5435202, 
    0.2679485, 0.2226279, 0.1700566, 0.2123212, 0.4024499, 0.22183, 
    0.3070359, 0.291237, 0.3464482, 0.2446336, 0.1352284, 0.1596893, 
    0.6476743, 0.03137168, 0.03951918, 0.05416327, 0.03064235,
  0.06268141, 0.02902455, 0.2594167, 0.0784395, 0.4739292, 0.323662, 
    0.6167271, 0.4856276, 0.47966, 0.6017166, 0.663808, 0.3877892, 0.6666335, 
    0.2405462, 0.2784105, 0.3362122, 0.4241396, 0.2231172, 0.3675476, 
    0.2462054, 0.285464, 0.4477758, 0.3176811, 0.2846608, 0.1132537, 
    0.1480004, 0.4515244, 0.11163, 0.1330632,
  0.5202895, 0.4783695, 0.5111322, 0.2912812, 0.3571323, 0.4582016, 
    0.4551691, 0.4131322, 0.4555469, 0.3953592, 0.4058218, 0.408956, 
    0.3429179, 0.3242839, 0.3815167, 0.4315896, 0.4399793, 0.4027672, 
    0.358427, 0.3735499, 0.3633735, 0.2572092, 0.2263299, 0.3641087, 
    0.09960489, 0.05943592, 0.04003475, 0.255415, 0.3548836,
  0.2123475, 0.2151578, 0.217968, 0.2207782, 0.2235885, 0.2263987, 0.229209, 
    0.1909586, 0.2019855, 0.2130123, 0.2240392, 0.235066, 0.2460929, 
    0.2571197, 0.3576828, 0.3513137, 0.3449445, 0.3385755, 0.3322064, 
    0.3258373, 0.3194682, 0.277472, 0.270004, 0.262536, 0.2550681, 0.2476001, 
    0.2401321, 0.2326641, 0.2100993,
  0.1560873, 0.1795674, 0.1916587, 0.3078817, 0.353343, 0.1939584, 0.1999942, 
    0.2518348, 0.1406608, 0.07794933, 0.06751838, 0.07843629, 0.1091367, 
    0.001340345, 0.2158734, 0.2712507, 0.1900499, 0.1626318, 0.03872195, 
    0.1977586, 0.2389969, 0.3266635, 0.07607935, 0.06548578, 0.1138008, 
    0.1629749, 0.1416238, 0.03545288, 0.07026018,
  0.0484015, 0.0339126, 0.03990227, 0.01258352, 0.01631446, 0.07733018, 
    0.01500348, 0.04030991, 0.102802, 0.1187092, 0.08030969, 0.06331221, 
    0.01503158, 0.01746953, 0.0722326, 0.1405701, 0.111151, 0.1177937, 
    0.1397245, 0.08872291, 0.1216004, 0.1567376, 0.2724858, 0.1193276, 
    0.1361013, 0.1045896, 0.09556075, 0.04881584, 0.06669307,
  0.1182199, 0.1314127, 0.1106518, 0.1799666, 0.1767855, 0.1478257, 
    0.1614484, 0.1339494, 0.1526382, 0.1230563, 0.1274908, 0.1743168, 
    0.2272533, 0.1847451, 0.1438267, 0.1693301, 0.1982718, 0.2404149, 
    0.1520567, 0.08240567, 0.07236556, 0.0684672, 0.06212813, 0.1054349, 
    0.1706563, 0.2296866, 0.2439147, 0.1703796, 0.1522356,
  0.1306199, 0.1216771, 0.1530664, 0.1384594, 0.1571384, 0.1747669, 
    0.1638255, 0.1070208, 0.09816088, 0.08840123, 0.04232628, 0.04516917, 
    0.0579445, 0.07269216, 0.1339755, 0.1198298, 0.08643487, 0.06812643, 
    0.06572814, 0.05453654, 0.03969261, 0.06993781, 0.08212856, 0.07888361, 
    0.02666394, 0.1003622, 0.1646919, 0.1600581, 0.1775442,
  0.03002381, 0.02106605, 0.01201019, 0.03941786, 0.04344747, 0.05360848, 
    0.04088253, 0.08922412, 0.05240373, 0.02417137, 0.01125296, 0.005578711, 
    0.006072524, 0.01208837, 0.1794012, 0.03505732, 0.02271379, 0.06103928, 
    0.04386044, 0.02717894, 0.04187617, 0.02328314, 0.0101323, 0.06275823, 
    0.01656445, 0.04436207, 0.08095554, 0.03852326, 0.02383501,
  0.003245526, 0.002564661, 0.016853, 0.0009147755, 0.005760003, 0.007154576, 
    0.0007056079, 0.002559502, 0.008080839, 0.0003774189, 0.0005688972, 
    0.000390557, 0.00474776, 0.003431872, 0.008474577, 0.004716212, 
    0.02423224, 0.02885854, 0.0127887, 0.001829691, 0.001805061, 0.0010178, 
    0.00380427, 0.01712818, 0.01289591, 0.002619337, 0.0006535688, 
    0.0002248668, 0.0009495197,
  0.001359729, 0.04977167, 0.00382741, 0.0003317342, -0.0008033491, 
    0.0001321212, 0.0005966314, 0.0008232553, 0.002541821, 0.004266356, 
    0.005344456, 0.0004994966, 0.0004465906, 0.0004380796, 0.0004366176, 
    0.001103708, 0.001217437, 0.0002511172, 2.225876e-05, 8.566107e-06, 
    1.177596e-05, 0.0003430962, 0.002957932, 0.01241389, 0.01520716, 
    0.07446006, 0.0003828885, 8.571999e-05, 0.0001529398,
  0.005381922, 0.002367712, 0.06685261, 0.1366045, 0.0004239877, 
    0.0003946503, 0.001159187, 8.439669e-05, 0.0004391214, 6.964335e-05, 
    0.0003653269, 0.0003489521, 6.864028e-05, 4.032838e-05, 0.001976187, 
    0.0002670908, 4.103423e-05, 0.0002431365, 0.000162694, 0.0002292035, 
    0.0007033748, 0.001014231, 0.001789797, 0.1019188, 0.05006916, 
    0.03357964, -0.0001054085, 0.0005354547, 0.00169274,
  0.0001577882, 0.06452537, 0.001501647, 0.004282579, 0.001468581, 
    0.001092625, 0.002426279, 0.001524131, 0.05366059, 0.09931245, 
    0.0001841446, 0.0005777621, 0.0001275889, 0.000761355, 0.00184759, 
    0.0001389809, 0.0001516446, 5.770999e-05, 0.0002841971, 8.585204e-05, 
    0.000664451, 0.00326751, 0.002858127, 0.06531611, 0.03160036, 
    0.001068304, 4.738699e-05, 0.0003403264, 0.0009757576,
  5.732909e-10, 5.365947e-10, 1.433529e-10, 0.003808534, 0.007402718, 
    0.0006393171, -0.0006935392, 0.0006276803, -0.0005203154, 0.001111129, 
    0.002655633, 8.701284e-05, 0.0001061714, 0.000314319, 0.0001628273, 
    0.0003501725, 0.0006384281, 0.001833717, 0.0009375044, 0.0006921542, 
    0.0002199697, 0.0002302489, 0.1442656, 0.03903014, 2.370957e-05, 
    0.0005322771, 0.002948158, 1.582133e-05, -0.00072444,
  2.512304e-08, 5.083061e-09, -3.289628e-08, 2.161717e-05, -2.505507e-08, 
    0.0002390483, 1.398356e-08, 0.000158161, 0.0003196546, 0.02356928, 
    0.003741294, 0.001562401, 0.001132707, 0.001331089, 0.001272998, 
    0.0007973582, 0.002674584, 0.002244154, 0.001976462, 0.007384616, 
    0.001228475, 0.07426924, 0.0002073306, -0.001087784, 5.372998e-05, 
    0.000379439, 0.001874139, 6.863607e-05, 1.946455e-07,
  -2.637094e-06, 0.003463896, 0.001179869, 0.001729866, 0.02351549, 
    0.002675725, -0.001040348, 0.0646078, 0.02513833, 0.07964804, 0.02630326, 
    0.004771011, 0.003984522, 0.01101222, 0.0154216, 0.0190777, 0.01281078, 
    0.02273048, 0.005194176, 0.002184776, 0.01447765, 0.08145819, 0.04779169, 
    0.0119191, 0.006260216, 0.00469116, 0.003218874, 0.002371749, 0.0006477026,
  0.01656227, 0.0001877568, 0.01040692, 0.2378972, 0.002496526, 0.03230303, 
    0.1450469, -4.693681e-06, 0.002910157, 0.0378847, 0.05558977, 0.02508077, 
    0.04945886, 0.04807829, 0.0197322, 0.03899636, 0.08420452, 0.06273519, 
    0.01706228, 0.1798761, 0.1236163, 0.05688788, 0.1227488, 0.1196979, 
    0.05037131, 0.02484965, 0.01600415, 0.007892076, 0.03635539,
  0.08407253, 0.1089293, 0.1510379, 0.3070327, 0.1920107, 0.1649241, 
    0.05145838, 0.1942451, 0.1602083, 0.04139311, 0.01758898, 0.1326875, 
    0.1333559, 0.1043939, 0.1084049, 0.04076767, 0.05696721, 0.06791193, 
    0.05392718, 0.3896907, 0.06642695, 0.07171926, 0.1062109, 0.3035549, 
    0.1428082, 0.06721406, 0.03963302, 0.02918806, 0.0403682,
  0.05562409, 0.4008203, 0.2831789, 0.4184378, 0.3656228, 0.2837025, 
    0.2822459, 0.2909983, 0.26412, 0.2652032, 0.3364422, 0.6599336, 
    0.3472852, 0.2256225, 0.1625178, 0.2028041, 0.4543903, 0.244487, 
    0.3621415, 0.3232124, 0.368188, 0.2773089, 0.1054406, 0.19642, 0.6442151, 
    0.03336206, 0.03532673, 0.04705824, 0.02539312,
  0.05350851, 0.02494476, 0.3120021, 0.06888708, 0.4681234, 0.2810536, 
    0.493327, 0.4523565, 0.5285131, 0.5816624, 0.6911382, 0.5401253, 
    0.5069911, 0.2289624, 0.2428823, 0.2873643, 0.4560698, 0.2476785, 
    0.3262658, 0.1900907, 0.2665766, 0.3641545, 0.2399426, 0.3326486, 
    0.1088031, 0.1406712, 0.5471841, 0.1080237, 0.1227593,
  0.5004803, 0.4881263, 0.4600914, 0.2613734, 0.2816322, 0.3629329, 0.34878, 
    0.3076749, 0.3683794, 0.3120129, 0.320803, 0.2875353, 0.2553217, 
    0.2341018, 0.2733694, 0.3053757, 0.2956488, 0.2783793, 0.2751173, 
    0.282182, 0.2648836, 0.256533, 0.2639455, 0.4459879, 0.102018, 0.0295193, 
    0.05022892, 0.2575523, 0.2794023 ;

 average_DT = 731 ;

 average_T1 = 45 ;

 average_T2 = 776 ;

 climatology_bounds =
  45, 776 ;

 lat = -89.5, -79.5, -69.5, -59.5, -49.5, -39.5, -29.5, -19.5, -9.5, 0.5, 
    10.5, 20.5, 30.5, 40.5, 50.5, 60.5, 70.5, 80.5 ;

 lat_bnds =
  -90, -89,
  -80, -79,
  -70, -69,
  -60, -59,
  -50, -49,
  -40, -39,
  -30, -29,
  -20, -19,
  -10, -9,
  0, 1,
  10, 11,
  20, 21,
  30, 31,
  40, 41,
  50, 51,
  60, 61,
  70, 71,
  80, 81 ;

 lon = 0.625, 13.125, 25.625, 38.125, 50.625, 63.125, 75.625, 88.125, 
    100.625, 113.125, 125.625, 138.125, 150.625, 163.125, 175.625, 188.125, 
    200.625, 213.125, 225.625, 238.125, 250.625, 263.125, 275.625, 288.125, 
    300.625, 313.125, 325.625, 338.125, 350.625 ;

 lon_bnds =
  0, 1.25,
  12.5, 13.75,
  25, 26.25,
  37.5, 38.75,
  50, 51.25,
  62.5, 63.75,
  75, 76.25,
  87.5, 88.75,
  100, 101.25,
  112.5, 113.75,
  125, 126.25,
  137.5, 138.75,
  150, 151.25,
  162.5, 163.75,
  175, 176.25,
  187.5, 188.75,
  200, 201.25,
  212.5, 213.75,
  225, 226.25,
  237.5, 238.75,
  250, 251.25,
  262.5, 263.75,
  275, 276.25,
  287.5, 288.75,
  300, 301.25,
  312.5, 313.75,
  325, 326.25,
  337.5, 338.75,
  350, 351.25 ;

 pfull = 0.0252729048206747, 0.0885404738757409, 0.213072411383256, 
    0.41190537807884, 0.671080828691593, 0.987471468515016, 1.36790961365676, 
    1.82562112064242, 2.38097588033244, 3.06218961364243, 3.90121721567151, 
    4.9296281825995, 6.18008131929323, 7.68875807563375, 9.49537809361575, 
    11.643153995098, 14.1786857151188, 17.1517875598959, 20.6152476986609, 
    24.6245259348741, 29.237386591333, 34.5134757786445, 40.5138467378254, 
    47.3004421634272, 54.9355325495126, 63.4811392623337, 72.9984371159701, 
    83.5471442618119, 95.1849171805989, 107.966767294215, 121.944503506415, 
    137.166169497631, 153.675572970355, 171.511834307961, 190.708985325578, 
    211.295632932361, 233.294677858721, 256.723099608772, 281.591803639405, 
    307.905555737256, 335.66293113824, 364.856338389786, 395.47216160598, 
    427.490864234311, 460.887168786725, 495.630391513078, 531.761718445649, 
    569.289185351388, 607.768705103107, 646.445374671436, 684.792067788697, 
    722.468679913451, 759.124006783627, 794.401045766566, 827.769968639223, 
    858.597822486016, 886.389109609622, 910.841030891388, 931.860653469283, 
    949.549679924174, 964.159924710431, 976.012345333387, 985.470174132691, 
    992.77226220014, 997.948601287575 ;

 time = 0 ;
}
