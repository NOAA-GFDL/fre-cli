netcdf tracer_level.0002-0002.scale_salt_emis {
dimensions:
	bnds = 2 ;
	lat = 18 ;
	lon = 29 ;
	time = UNLIMITED ; // (1 currently)
variables:
	double bnds(bnds) ;
		bnds:long_name = "vertex number" ;
	double lat(lat) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_N" ;
		lat:axis = "Y" ;
		lat:bounds = "lat_bnds" ;
	double lat_bnds(lat, bnds) ;
		lat_bnds:long_name = "latitude bounds" ;
		lat_bnds:units = "degrees_N" ;
		lat_bnds:axis = "Y" ;
	double lon(lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_E" ;
		lon:axis = "X" ;
		lon:bounds = "lon_bnds" ;
	double lon_bnds(lon, bnds) ;
		lon_bnds:long_name = "longitude bounds" ;
		lon_bnds:units = "degrees_E" ;
		lon_bnds:axis = "X" ;
	float scale_salt_emis(time, lat, lon) ;
		scale_salt_emis:_FillValue = 1.e+20f ;
		scale_salt_emis:missing_value = 1.e+20f ;
		scale_salt_emis:units = "unitless" ;
		scale_salt_emis:long_name = "scale salt emis" ;
		scale_salt_emis:interp_method = "conserve_order1" ;
		scale_salt_emis:cell_methods = "time: mean" ;
	double time(time) ;
		time:units = "days since 0001-01-01 00:00:00" ;
		time:long_name = "time" ;
		time:axis = "T" ;
		time:calendar_type = "NOLEAP" ;
		time:calendar = "noleap" ;
		time:bounds = "time_bnds" ;
	double time_bnds(time, bnds) ;
		time_bnds:units = "days since 0001-01-01 00:00:00" ;
		time_bnds:long_name = "time axis boundaries" ;

// global attributes:
		:title = "cm5_c96_am5f7c1r0_b06_piC_galb_noiceinit_alb" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
		:code_release_version = "2024.02" ;
		:git_hash = "b86d27037f755a82c586e55073dd575245c144b1" ;
		:creationtime = "Fri Dec  6 17:15:31 2024" ;
		:hostname = "pp329" ;
		:history = "Tue Aug 12 16:31:58 2025: ncks -d lat,,,10 -d lon,,,10 tracer_level.0002-0002.scale_salt_emis.nc reduced/tracer_level.0002-0002.scale_salt_emis.nc\n",
			"fregrid --standard_dimension --input_mosaic C96_mosaic.nc --input_file 00020101.atmos_tracer --interp_method conserve_order1 --remap_file .fregrid_remap_file_288_by_180.nc --nlon 288 --nlat 180 --scalar_field bk,pk,radon,ssalt1_emis,ssalt2_emis,ssalt3_emis,ssalt4_emis,ssalt5_emis,ssalt1_setl,ssalt2_setl,ssalt3_setl,ssalt4_setl,ssalt5_setl,ssalt1_wet_dep,ssalt2_wet_dep,ssalt3_wet_dep,ssalt4_wet_dep,ssalt5_wet_dep,ssalt1_dvel,ssalt2_dvel,ssalt3_dvel,ssalt4_dvel,ssalt5_dvel,ssalt1_ddep,ssalt2_ddep,ssalt3_ddep,ssalt4_ddep,ssalt5_ddep,scale_salt_emis,time_bnds --output_file out.nc" ;
		:comment = "FMS time averaging, version 3.0, precision=double" ;
		:NCO = "netCDF Operators version 5.2.4 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco, Citation = 10.1016/j.envsoft.2008.03.004)" ;
data:

 bnds = 1, 2 ;

 lat = -89.5, -79.5, -69.5, -59.5, -49.5, -39.5, -29.5, -19.5, -9.5, 0.5, 
    10.5, 20.5, 30.5, 40.5, 50.5, 60.5, 70.5, 80.5 ;

 lat_bnds =
  -90, -89,
  -80, -79,
  -70, -69,
  -60, -59,
  -50, -49,
  -40, -39,
  -30, -29,
  -20, -19,
  -10, -9,
  0, 1,
  10, 11,
  20, 21,
  30, 31,
  40, 41,
  50, 51,
  60, 61,
  70, 71,
  80, 81 ;

 lon = 0.625, 13.125, 25.625, 38.125, 50.625, 63.125, 75.625, 88.125, 
    100.625, 113.125, 125.625, 138.125, 150.625, 163.125, 175.625, 188.125, 
    200.625, 213.125, 225.625, 238.125, 250.625, 263.125, 275.625, 288.125, 
    300.625, 313.125, 325.625, 338.125, 350.625 ;

 lon_bnds =
  0, 1.25,
  12.5, 13.75,
  25, 26.25,
  37.5, 38.75,
  50, 51.25,
  62.5, 63.75,
  75, 76.25,
  87.5, 88.75,
  100, 101.25,
  112.5, 113.75,
  125, 126.25,
  137.5, 138.75,
  150, 151.25,
  162.5, 163.75,
  175, 176.25,
  187.5, 188.75,
  200, 201.25,
  212.5, 213.75,
  225, 226.25,
  237.5, 238.75,
  250, 251.25,
  262.5, 263.75,
  275, 276.25,
  287.5, 288.75,
  300, 301.25,
  312.5, 313.75,
  325, 326.25,
  337.5, 338.75,
  350, 351.25 ;

 scale_salt_emis =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9102186, 0.8604528, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1,
  0.3296477, 0.3290002, 0.3290007, 0.3309282, 1, 1, 0.3314292, 1, 1, 1, 1, 1, 
    0.6211897, 0.3302617, 0.329, 0.329, 0.329, 0.3290168, 0.3290002, 
    0.3290001, 0.329119, 0.3297966, 0.3369154, 0.3331891, 0.3295439, 0.329, 
    0.329, 0.329, 0.3295651,
  0.3371729, 0.3386994, 0.3408951, 0.3395075, 0.3470881, 0.3722999, 
    0.3518886, 0.3952325, 0.348536, 0.3448845, 0.3701847, 0.397248, 
    0.3910242, 0.5976994, 0.6396083, 0.5569168, 0.4495965, 0.4010386, 
    0.511073, 0.514978, 0.5259352, 0.5797572, 0.60065, 0.6067469, 0.39921, 
    0.4114034, 0.3989161, 0.3748124, 0.3432934,
  0.6298555, 0.6027915, 0.5656114, 0.588512, 0.5961135, 0.60136, 0.5706596, 
    0.6861383, 0.634931, 0.6396075, 0.6895247, 0.6879635, 0.7093733, 
    0.7184394, 0.704713, 0.7305059, 0.7294949, 0.7221748, 0.700253, 
    0.6811001, 0.681775, 0.6758776, 0.6821724, 1, 0.6879607, 0.6614476, 
    0.6307729, 0.6351866, 0.5826361,
  0.7520998, 0.750919, 0.7993714, 0.8148194, 0.8029634, 0.7861974, 0.7851042, 
    0.7608019, 0.7430172, 0.742758, 0.7490817, 0.7782386, 0.817667, 
    0.8027568, 0.9636984, 0.8060386, 0.7921332, 0.7768064, 0.7630197, 
    0.7614706, 0.7661467, 0.7651634, 0.7690724, 1, 0.7952487, 0.7929625, 
    0.7891757, 0.7733648, 0.7630287,
  0.8797275, 0.8449149, 1, 1.153171, 1.093907, 1.068495, 0.9878888, 
    0.9260218, 0.8675792, 1.085712, 1, 1, 1, 1.033729, 1.043196, 1.043852, 
    1.041912, 1.04601, 1.071271, 1.08346, 1.095675, 1.024644, 0.8937485, 
    0.9138233, 1, 1.058399, 1.004075, 0.9895277, 0.9382431,
  0.9863473, 1.238238, 1, 1.62324, 1.484143, 1.367136, 1.224457, 1.170952, 
    1.188306, 1.454394, 1, 1, 1.451664, 1.463599, 1.534147, 1.515187, 
    1.486369, 1.423484, 1.359231, 1.249717, 1.108656, 0.9777949, 0.9129261, 
    1.059994, 1, 1, 1.264084, 1.087481, 0.9913942,
  1.503706, 1.680604, 1, 1, 1.620708, 1.654683, 1.621423, 1.671825, 1.785053, 
    1.868382, 1.746655, 1.812026, 1.839639, 1.977715, 1.911868, 1.82181, 
    1.731165, 1.609439, 1.49022, 1.380854, 1.283819, 1.201916, 1.210948, 1, 
    1, 1, 1.479333, 1.507641, 1.479214,
  1.857402, 1, 1, 1, 1.640938, 1.911062, 1.907253, 1.91518, 1.056642, 1, 
    2.069844, 2.067556, 2.0059, 1.884957, 1.717608, 1.591674, 1.49585, 
    1.401825, 1.270026, 1.172125, 1.104888, 1.175035, 1.450881, 1, 1, 
    1.631075, 1.57507, 1.647949, 1.758816,
  1, 1, 1, 1, 1.528613, 1.727899, 1.706319, 1.799111, 1.799193, 1.79817, 
    1.80352, 1.859412, 1.845677, 1.773694, 1.694453, 1.658343, 1.624091, 
    1.634069, 1.669537, 1.672654, 1.67479, 1.668777, 1.088935, 1.501016, 
    1.65305, 1.599206, 1.544332, 1.524576, 1,
  1, 1, 1, 1.729381, 1, 1.396547, 1, 1.696521, 1, 1.570495, 1.548481, 
    1.538056, 1.566143, 1.503188, 1.442366, 1.391122, 1.370778, 1.194978, 
    1.117747, 1.209273, 1.619209, 1.372711, 1.687163, 1.585171, 1.437394, 
    1.310064, 1.20201, 1.141775, 1,
  1, 1, 1.046025, 1, 1.146102, 1, 1, 1, 1, 1, 1.045999, 1.188558, 1.093168, 
    1.04286, 1.011154, 0.9655874, 0.9502635, 0.9372212, 0.8859323, 0.8466945, 
    1, 1, 1.084712, 1.277099, 1.22488, 1.187116, 1.041395, 0.9524601, 1.163123,
  0.96485, 0.9695348, 0.918228, 0.9037478, 1, 1, 1, 1, 1, 1, 1, 0.8554919, 
    0.8092672, 0.7816681, 0.7716753, 0.7676703, 0.7876042, 0.7910683, 
    0.7699994, 1, 1, 1, 1, 0.8339392, 0.9305618, 0.8820788, 0.8601742, 
    0.8206283, 0.8196361,
  0.7452157, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9946604, 0.5294534, 0.569612, 
    0.615425, 0.6288385, 0.6414759, 0.6605721, 0.7047323, 1, 1, 1, 1, 1, 
    0.6390572, 0.6848722, 0.7314101, 0.7470665, 0.7431206,
  0.7034169, 1, 0.5765121, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.6503509, 0.4700027, 
    0.5122825, 0.4229538, 1, 0.4874792, 1, 1, 1, 0.9688244, 0.4324096, 
    0.9528526, 0.5369457, 0.5754016, 0.6870786, 0.7125688, 0.7134482,
  0.5586247, 0.6111827, 0.4210862, 0.4291934, 0.3743742, 0.333806, 0.3961508, 
    1, 1, 1, 1, 0.9392857, 0.7811477, 0.3662757, 0.358023, 0.3834543, 
    0.4382198, 0.4172753, 0.4246714, 0.3971203, 1, 0.3623618, 0.4200918, 
    0.6465928, 0.4138302, 0.9794093, 1, 0.3438256, 0.3906454,
  0.329, 0.329, 0.3307337, 0.329, 0.3299954, 0.3304242, 0.329, 0.3442636, 
    0.3349507, 0.3309646, 0.3306479, 0.3300624, 0.3311481, 0.336798, 
    0.340131, 0.3430622, 0.3490393, 0.3432007, 0.3361313, 0.3332506, 
    0.3327981, 0.3455813, 0.3500048, 0.329956, 0.6671661, 0.9717175, 1, 
    0.4145629, 0.329 ;

 time = 547.5 ;

 time_bnds =
  365, 730 ;
}
