netcdf tracer_level.0003-0003.radon {
dimensions:
	bnds = 2 ;
	lat = 18 ;
	lon = 29 ;
	pfull = 65 ;
	time = UNLIMITED ; // (1 currently)
variables:
	double bnds(bnds) ;
		bnds:long_name = "vertex number" ;
	double lat(lat) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_N" ;
		lat:axis = "Y" ;
		lat:bounds = "lat_bnds" ;
	double lat_bnds(lat, bnds) ;
		lat_bnds:long_name = "latitude bounds" ;
		lat_bnds:units = "degrees_N" ;
		lat_bnds:axis = "Y" ;
	double lon(lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_E" ;
		lon:axis = "X" ;
		lon:bounds = "lon_bnds" ;
	double lon_bnds(lon, bnds) ;
		lon_bnds:long_name = "longitude bounds" ;
		lon_bnds:units = "degrees_E" ;
		lon_bnds:axis = "X" ;
	double pfull(pfull) ;
		pfull:units = "mb" ;
		pfull:long_name = "ref full pressure level" ;
		pfull:axis = "Z" ;
		pfull:positive = "down" ;
	float radon(time, pfull, lat, lon) ;
		radon:_FillValue = -1.e+10f ;
		radon:missing_value = -1.e+10f ;
		radon:units = "vmr*1e21" ;
		radon:long_name = "radon-222" ;
		radon:interp_method = "conserve_order1" ;
		radon:cell_methods = "time: mean" ;
	double time(time) ;
		time:units = "days since 0001-01-01 00:00:00" ;
		time:long_name = "time" ;
		time:axis = "T" ;
		time:calendar_type = "NOLEAP" ;
		time:calendar = "noleap" ;
		time:bounds = "time_bnds" ;
	double time_bnds(time, bnds) ;
		time_bnds:units = "days since 0001-01-01 00:00:00" ;
		time_bnds:long_name = "time axis boundaries" ;

// global attributes:
		:title = "cm5_c96_am5f7c1r0_b06_piC_galb_noiceinit_alb" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
		:code_release_version = "2024.02" ;
		:git_hash = "b86d27037f755a82c586e55073dd575245c144b1" ;
		:creationtime = "Fri Dec  6 16:33:51 2024" ;
		:hostname = "pp211" ;
		:history = "Tue Aug 12 16:38:49 2025: ncks -d lat,,,10 -d lon,,,10 tracer_level.0003-0003.radon.nc reduced/tracer_level.0003-0003.radon.nc\n",
			"fregrid --standard_dimension --input_mosaic C96_mosaic.nc --input_file 00030101.atmos_tracer --interp_method conserve_order1 --remap_file .fregrid_remap_file_288_by_180.nc --nlon 288 --nlat 180 --scalar_field bk,pk,radon,ssalt1_emis,ssalt2_emis,ssalt3_emis,ssalt4_emis,ssalt5_emis,ssalt1_setl,ssalt2_setl,ssalt3_setl,ssalt4_setl,ssalt5_setl,ssalt1_wet_dep,ssalt2_wet_dep,ssalt3_wet_dep,ssalt4_wet_dep,ssalt5_wet_dep,ssalt1_dvel,ssalt2_dvel,ssalt3_dvel,ssalt4_dvel,ssalt5_dvel,ssalt1_ddep,ssalt2_ddep,ssalt3_ddep,ssalt4_ddep,ssalt5_ddep,scale_salt_emis,time_bnds --output_file out.nc" ;
		:comment = "FMS time averaging, version 3.0, precision=double" ;
		:NCO = "netCDF Operators version 5.2.4 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco, Citation = 10.1016/j.envsoft.2008.03.004)" ;
data:

 bnds = 1, 2 ;

 lat = -89.5, -79.5, -69.5, -59.5, -49.5, -39.5, -29.5, -19.5, -9.5, 0.5, 
    10.5, 20.5, 30.5, 40.5, 50.5, 60.5, 70.5, 80.5 ;

 lat_bnds =
  -90, -89,
  -80, -79,
  -70, -69,
  -60, -59,
  -50, -49,
  -40, -39,
  -30, -29,
  -20, -19,
  -10, -9,
  0, 1,
  10, 11,
  20, 21,
  30, 31,
  40, 41,
  50, 51,
  60, 61,
  70, 71,
  80, 81 ;

 lon = 0.625, 13.125, 25.625, 38.125, 50.625, 63.125, 75.625, 88.125, 
    100.625, 113.125, 125.625, 138.125, 150.625, 163.125, 175.625, 188.125, 
    200.625, 213.125, 225.625, 238.125, 250.625, 263.125, 275.625, 288.125, 
    300.625, 313.125, 325.625, 338.125, 350.625 ;

 lon_bnds =
  0, 1.25,
  12.5, 13.75,
  25, 26.25,
  37.5, 38.75,
  50, 51.25,
  62.5, 63.75,
  75, 76.25,
  87.5, 88.75,
  100, 101.25,
  112.5, 113.75,
  125, 126.25,
  137.5, 138.75,
  150, 151.25,
  162.5, 163.75,
  175, 176.25,
  187.5, 188.75,
  200, 201.25,
  212.5, 213.75,
  225, 226.25,
  237.5, 238.75,
  250, 251.25,
  262.5, 263.75,
  275, 276.25,
  287.5, 288.75,
  300, 301.25,
  312.5, 313.75,
  325, 326.25,
  337.5, 338.75,
  350, 351.25 ;

 pfull = 0.0252729048206747, 0.0885404738757409, 0.213072411383256, 
    0.41190537807884, 0.671080828691593, 0.987471468515016, 1.36790961365676, 
    1.82562112064242, 2.38097588033244, 3.06218961364243, 3.90121721567151, 
    4.9296281825995, 6.18008131929323, 7.68875807563375, 9.49537809361575, 
    11.643153995098, 14.1786857151188, 17.1517875598959, 20.6152476986609, 
    24.6245259348741, 29.237386591333, 34.5134757786445, 40.5138467378254, 
    47.3004421634272, 54.9355325495126, 63.4811392623337, 72.9984371159701, 
    83.5471442618119, 95.1849171805989, 107.966767294215, 121.944503506415, 
    137.166169497631, 153.675572970355, 171.511834307961, 190.708985325578, 
    211.295632932361, 233.294677858721, 256.723099608772, 281.591803639405, 
    307.905555737256, 335.66293113824, 364.856338389786, 395.47216160598, 
    427.490864234311, 460.887168786725, 495.630391513078, 531.761718445649, 
    569.289185351388, 607.768705103107, 646.445374671436, 684.792067788697, 
    722.468679913451, 759.124006783627, 794.401045766566, 827.769968639223, 
    858.597822486016, 886.389109609622, 910.841030891388, 931.860653469283, 
    949.549679924174, 964.159924710431, 976.012345333387, 985.470174132691, 
    992.77226220014, 997.948601287575 ;

 radon =
  1.529905e-20, 1.529905e-20, 1.529905e-20, 1.529905e-20, 1.529905e-20, 
    1.529905e-20, 1.529905e-20, 1.570424e-20, 1.570424e-20, 1.570424e-20, 
    1.570424e-20, 1.570424e-20, 1.570424e-20, 1.570424e-20, 1.461861e-20, 
    1.461861e-20, 1.461861e-20, 1.461861e-20, 1.461861e-20, 1.461861e-20, 
    1.461861e-20, 1.417031e-20, 1.417031e-20, 1.417031e-20, 1.417031e-20, 
    1.417031e-20, 1.417031e-20, 1.417031e-20, 1.529905e-20,
  2.792644e-20, 2.94163e-20, 2.990711e-20, 3.043833e-20, 3.104231e-20, 
    3.198042e-20, 3.219991e-20, 3.186235e-20, 3.133002e-20, 3.069218e-20, 
    2.994387e-20, 2.861837e-20, 2.740331e-20, 2.62316e-20, 2.509186e-20, 
    2.377209e-20, 2.223065e-20, 2.093378e-20, 1.976975e-20, 1.846463e-20, 
    1.737695e-20, 1.687829e-20, 1.683034e-20, 1.692227e-20, 1.87837e-20, 
    2.191543e-20, 2.380868e-20, 2.531372e-20, 2.744932e-20,
  6.291285e-20, 6.356922e-20, 6.209972e-20, 6.370077e-20, 6.515402e-20, 
    6.613891e-20, 6.609035e-20, 6.591663e-20, 6.583151e-20, 6.240656e-20, 
    5.902473e-20, 5.541319e-20, 5.273494e-20, 5.033542e-20, 4.591586e-20, 
    4.304027e-20, 4.009911e-20, 3.783607e-20, 3.612019e-20, 3.450833e-20, 
    3.465537e-20, 3.655801e-20, 4.173054e-20, 4.590905e-20, 4.863177e-20, 
    4.851119e-20, 5.317074e-20, 5.845196e-20, 6.134737e-20,
  1.339326e-19, 1.378785e-19, 1.383572e-19, 1.421069e-19, 1.374414e-19, 
    1.37718e-19, 1.335003e-19, 1.293423e-19, 1.270034e-19, 1.222106e-19, 
    1.140254e-19, 1.102128e-19, 1.055618e-19, 1.024667e-19, 9.996735e-20, 
    9.522275e-20, 9.232591e-20, 9.927119e-20, 1.014957e-19, 9.952638e-20, 
    1.001275e-19, 1.002523e-19, 1.049665e-19, 1.143355e-19, 1.209165e-19, 
    1.222613e-19, 1.27011e-19, 1.239263e-19, 1.322282e-19,
  3.687176e-19, 3.766959e-19, 3.598953e-19, 3.500167e-19, 3.499452e-19, 
    3.427155e-19, 3.251263e-19, 3.174702e-19, 2.994454e-19, 3.065455e-19, 
    3.207701e-19, 3.097657e-19, 3.103803e-19, 3.25053e-19, 3.261128e-19, 
    3.368267e-19, 3.452066e-19, 3.253044e-19, 3.100357e-19, 3.204692e-19, 
    3.431552e-19, 3.491795e-19, 3.548529e-19, 3.545652e-19, 3.408539e-19, 
    3.546602e-19, 3.641355e-19, 3.590176e-19, 3.558187e-19,
  6.836935e-19, 6.758511e-19, 6.600581e-19, 6.567139e-19, 6.534449e-19, 
    6.506283e-19, 6.249643e-19, 6.435146e-19, 6.456624e-19, 6.100797e-19, 
    6.00116e-19, 5.920137e-19, 5.970792e-19, 6.048863e-19, 6.218084e-19, 
    6.24877e-19, 6.436755e-19, 6.517679e-19, 6.574299e-19, 6.866661e-19, 
    6.717213e-19, 6.578521e-19, 6.568273e-19, 6.697756e-19, 6.582734e-19, 
    6.796152e-19, 6.943658e-19, 7.123142e-19, 6.913157e-19,
  8.410984e-19, 8.393758e-19, 8.282354e-19, 8.16854e-19, 8.158556e-19, 
    8.45247e-19, 8.794888e-19, 8.677967e-19, 8.20273e-19, 8.003768e-19, 
    7.99527e-19, 7.813897e-19, 7.617919e-19, 7.634965e-19, 7.518716e-19, 
    7.795946e-19, 8.067737e-19, 8.102195e-19, 8.161774e-19, 8.570868e-19, 
    8.820782e-19, 8.83071e-19, 8.279955e-19, 8.472959e-19, 8.474791e-19, 
    8.85373e-19, 9.104047e-19, 8.963234e-19, 8.629073e-19,
  1.529364e-18, 1.441613e-18, 1.389551e-18, 1.481377e-18, 1.518948e-18, 
    1.609079e-18, 1.595011e-18, 1.612517e-18, 1.598066e-18, 1.428549e-18, 
    1.40217e-18, 1.277455e-18, 1.280097e-18, 1.266934e-18, 1.195355e-18, 
    1.247625e-18, 1.244335e-18, 1.180211e-18, 1.176883e-18, 1.259094e-18, 
    1.286865e-18, 1.303127e-18, 1.412689e-18, 1.383588e-18, 1.399291e-18, 
    1.411239e-18, 1.450886e-18, 1.489284e-18, 1.481969e-18,
  2.309859e-18, 2.260571e-18, 2.247057e-18, 2.342657e-18, 2.496715e-18, 
    2.516091e-18, 2.431865e-18, 2.238618e-18, 2.177682e-18, 2.092994e-18, 
    1.948004e-18, 1.809427e-18, 1.775756e-18, 1.799602e-18, 1.722921e-18, 
    1.733008e-18, 1.675467e-18, 1.723339e-18, 1.74219e-18, 1.782298e-18, 
    1.899084e-18, 2.015597e-18, 2.008239e-18, 2.127551e-18, 2.04813e-18, 
    2.190875e-18, 2.306886e-18, 2.327837e-18, 2.322991e-18,
  2.48718e-18, 2.555999e-18, 2.678844e-18, 2.407835e-18, 2.509911e-18, 
    2.512623e-18, 2.477395e-18, 2.462777e-18, 2.34766e-18, 2.17152e-18, 
    2.087229e-18, 1.947183e-18, 1.887236e-18, 1.830724e-18, 1.787617e-18, 
    1.83408e-18, 1.849676e-18, 1.749673e-18, 1.850597e-18, 1.865563e-18, 
    2.038324e-18, 2.192424e-18, 2.30774e-18, 2.46194e-18, 2.448611e-18, 
    2.43753e-18, 2.357872e-18, 2.557602e-18, 2.585383e-18,
  2.248639e-18, 2.271656e-18, 2.229075e-18, 2.133042e-18, 2.248369e-18, 
    2.265566e-18, 2.176944e-18, 2.160566e-18, 2.025706e-18, 1.934781e-18, 
    1.855758e-18, 1.75437e-18, 1.639255e-18, 1.577406e-18, 1.552321e-18, 
    1.534864e-18, 1.566428e-18, 1.673451e-18, 1.619866e-18, 1.652293e-18, 
    1.835637e-18, 1.867994e-18, 1.967927e-18, 2.076814e-18, 2.074902e-18, 
    2.015617e-18, 1.920688e-18, 2.076585e-18, 2.150319e-18,
  1.297626e-18, 1.258914e-18, 1.278968e-18, 1.328942e-18, 1.462818e-18, 
    1.518581e-18, 1.467145e-18, 1.397982e-18, 1.422046e-18, 1.324788e-18, 
    1.336662e-18, 1.360683e-18, 1.321881e-18, 1.306421e-18, 1.277498e-18, 
    1.210434e-18, 1.165711e-18, 1.16792e-18, 1.169802e-18, 1.215448e-18, 
    1.267507e-18, 1.299639e-18, 1.28498e-18, 1.230338e-18, 1.214607e-18, 
    1.248382e-18, 1.26301e-18, 1.286118e-18, 1.302682e-18,
  6.755676e-19, 6.448173e-19, 6.644589e-19, 6.597928e-19, 6.930701e-19, 
    7.088545e-19, 7.203643e-19, 7.247768e-19, 6.993435e-19, 6.890466e-19, 
    6.879142e-19, 7.113188e-19, 7.371714e-19, 7.250285e-19, 7.371592e-19, 
    7.392653e-19, 7.48707e-19, 7.618746e-19, 7.625732e-19, 7.536131e-19, 
    7.539401e-19, 7.445632e-19, 7.374904e-19, 7.459634e-19, 7.735216e-19, 
    7.872748e-19, 7.682547e-19, 7.352931e-19, 7.010524e-19,
  4.231602e-19, 3.964815e-19, 3.782945e-19, 3.911071e-19, 3.641974e-19, 
    3.665488e-19, 3.669822e-19, 3.597399e-19, 3.726893e-19, 3.803257e-19, 
    3.712741e-19, 3.700621e-19, 3.54276e-19, 3.492298e-19, 3.46752e-19, 
    3.61374e-19, 3.769701e-19, 3.989339e-19, 4.259599e-19, 4.343806e-19, 
    4.342421e-19, 4.330312e-19, 4.265806e-19, 4.226742e-19, 4.305164e-19, 
    4.457013e-19, 4.673632e-19, 4.760536e-19, 4.558912e-19,
  2.554122e-19, 2.398996e-19, 2.517105e-19, 2.530264e-19, 2.487636e-19, 
    2.411612e-19, 2.43711e-19, 2.44708e-19, 2.487262e-19, 2.344839e-19, 
    2.23615e-19, 2.052627e-19, 1.962553e-19, 1.96636e-19, 1.779718e-19, 
    1.716171e-19, 1.694708e-19, 1.742272e-19, 1.776125e-19, 1.878437e-19, 
    1.963663e-19, 2.107088e-19, 2.343268e-19, 2.539544e-19, 2.693412e-19, 
    2.641719e-19, 2.631631e-19, 2.764146e-19, 2.651537e-19,
  1.881961e-19, 1.805493e-19, 1.758531e-19, 1.803266e-19, 1.754786e-19, 
    1.695378e-19, 1.809524e-19, 1.787327e-19, 1.909773e-19, 1.794786e-19, 
    1.746284e-19, 1.628943e-19, 1.464135e-19, 1.345534e-19, 1.245071e-19, 
    1.121896e-19, 1.050615e-19, 9.581917e-20, 9.085416e-20, 9.25267e-20, 
    9.556695e-20, 9.973583e-20, 1.104445e-19, 1.288537e-19, 1.496264e-19, 
    1.597224e-19, 1.750007e-19, 1.809875e-19, 1.841693e-19,
  1.464375e-19, 1.484765e-19, 1.494066e-19, 1.510798e-19, 1.53043e-19, 
    1.491743e-19, 1.476378e-19, 1.471888e-19, 1.483093e-19, 1.469853e-19, 
    1.384596e-19, 1.308295e-19, 1.184412e-19, 1.120846e-19, 1.066391e-19, 
    1.004659e-19, 9.559956e-20, 8.801264e-20, 8.399971e-20, 8.177865e-20, 
    8.303892e-20, 8.287016e-20, 8.265304e-20, 8.74223e-20, 8.968954e-20, 
    9.262664e-20, 1.067183e-19, 1.279745e-19, 1.390544e-19,
  1.156813e-19, 1.257387e-19, 1.321264e-19, 1.337644e-19, 1.388633e-19, 
    1.438769e-19, 1.4638e-19, 1.448198e-19, 1.40311e-19, 1.344297e-19, 
    1.281878e-19, 1.213302e-19, 1.143174e-19, 1.049721e-19, 9.748716e-20, 
    9.114474e-20, 8.617404e-20, 8.262527e-20, 7.843981e-20, 7.572658e-20, 
    7.401408e-20, 7.149407e-20, 6.991637e-20, 6.876957e-20, 7.078766e-20, 
    7.636585e-20, 8.317334e-20, 9.625048e-20, 1.117353e-19,
  3.242325e-20, 3.242325e-20, 3.242325e-20, 3.242325e-20, 3.242325e-20, 
    3.242325e-20, 3.242325e-20, 3.257049e-20, 3.257049e-20, 3.257049e-20, 
    3.257049e-20, 3.257049e-20, 3.257049e-20, 3.257049e-20, 3.021871e-20, 
    3.021871e-20, 3.021871e-20, 3.021871e-20, 3.021871e-20, 3.021871e-20, 
    3.021871e-20, 2.993235e-20, 2.993235e-20, 2.993235e-20, 2.993235e-20, 
    2.993235e-20, 2.993235e-20, 2.993235e-20, 3.242325e-20,
  7.029581e-20, 8.047592e-20, 8.559827e-20, 8.615599e-20, 8.906016e-20, 
    8.875024e-20, 8.809855e-20, 8.625731e-20, 8.323346e-20, 7.964006e-20, 
    8.035555e-20, 7.90436e-20, 7.728811e-20, 7.420181e-20, 6.923716e-20, 
    6.231781e-20, 5.459115e-20, 4.925065e-20, 4.354375e-20, 3.929421e-20, 
    3.530195e-20, 3.38593e-20, 3.209246e-20, 3.286094e-20, 3.713715e-20, 
    4.438604e-20, 4.974586e-20, 5.557107e-20, 6.629825e-20,
  2.044447e-19, 2.232688e-19, 2.286154e-19, 2.339311e-19, 2.404307e-19, 
    2.484625e-19, 2.58791e-19, 2.672724e-19, 2.686793e-19, 2.596689e-19, 
    2.41781e-19, 2.252732e-19, 2.139905e-19, 2.010314e-19, 1.865359e-19, 
    1.756465e-19, 1.612269e-19, 1.508166e-19, 1.363264e-19, 1.201255e-19, 
    1.113628e-19, 1.133402e-19, 1.200546e-19, 1.37325e-19, 1.487299e-19, 
    1.571939e-19, 1.649308e-19, 1.796239e-19, 1.923439e-19,
  6.562758e-19, 7.03591e-19, 6.944993e-19, 7.088025e-19, 7.008139e-19, 
    6.944805e-19, 6.772162e-19, 6.30426e-19, 6.105944e-19, 6.129472e-19, 
    5.966587e-19, 5.562945e-19, 5.374058e-19, 5.149737e-19, 4.74243e-19, 
    4.444378e-19, 4.132849e-19, 3.972794e-19, 4.229769e-19, 4.424964e-19, 
    4.505754e-19, 4.468304e-19, 4.554868e-19, 4.686821e-19, 4.735915e-19, 
    5.07778e-19, 5.186342e-19, 5.622863e-19, 6.040552e-19,
  1.618024e-18, 1.600177e-18, 1.554625e-18, 1.470625e-18, 1.441288e-18, 
    1.45021e-18, 1.427806e-18, 1.415244e-18, 1.362932e-18, 1.354966e-18, 
    1.350921e-18, 1.274714e-18, 1.272936e-18, 1.289551e-18, 1.286411e-18, 
    1.29888e-18, 1.295458e-18, 1.243505e-18, 1.208698e-18, 1.297857e-18, 
    1.344362e-18, 1.334767e-18, 1.367928e-18, 1.398355e-18, 1.44659e-18, 
    1.527619e-18, 1.653101e-18, 1.671746e-18, 1.628738e-18,
  3.18729e-18, 3.081124e-18, 3.022619e-18, 2.949331e-18, 2.819096e-18, 
    2.767871e-18, 2.85794e-18, 2.757101e-18, 2.740142e-18, 2.669628e-18, 
    2.642566e-18, 2.645462e-18, 2.623457e-18, 2.578216e-18, 2.673928e-18, 
    2.609192e-18, 2.609101e-18, 2.716304e-18, 2.830178e-18, 2.945804e-18, 
    3.040861e-18, 3.066788e-18, 3.138506e-18, 3.273527e-18, 3.35741e-18, 
    3.448541e-18, 3.295491e-18, 3.242759e-18, 3.333775e-18,
  3.899575e-18, 3.864113e-18, 3.768397e-18, 3.868997e-18, 3.847597e-18, 
    3.983579e-18, 4.070398e-18, 3.859339e-18, 3.864676e-18, 3.921135e-18, 
    3.904773e-18, 3.88134e-18, 3.744028e-18, 3.747635e-18, 3.725756e-18, 
    3.891378e-18, 4.038157e-18, 3.976294e-18, 4.057749e-18, 4.196298e-18, 
    4.246421e-18, 4.163313e-18, 4.322499e-18, 4.171851e-18, 4.154108e-18, 
    4.065848e-18, 4.093697e-18, 4.009769e-18, 3.944097e-18,
  6.185096e-18, 6.285208e-18, 6.062397e-18, 6.309337e-18, 6.356195e-18, 
    6.930695e-18, 6.716457e-18, 6.738121e-18, 6.958568e-18, 6.380307e-18, 
    6.010909e-18, 5.810158e-18, 5.649354e-18, 5.828608e-18, 5.503446e-18, 
    5.559872e-18, 5.454155e-18, 5.234663e-18, 5.545034e-18, 5.557592e-18, 
    5.69623e-18, 6.066342e-18, 6.263001e-18, 6.23517e-18, 6.455788e-18, 
    6.220098e-18, 6.185148e-18, 5.9627e-18, 6.071808e-18,
  9.433826e-18, 9.217257e-18, 9.562544e-18, 1.004435e-17, 9.29685e-18, 
    9.872941e-18, 1.024477e-17, 1.021597e-17, 1.016537e-17, 9.022554e-18, 
    9.275801e-18, 8.865059e-18, 7.943717e-18, 7.78021e-18, 7.721445e-18, 
    7.583722e-18, 7.419064e-18, 7.275571e-18, 7.675491e-18, 7.982647e-18, 
    8.08515e-18, 8.822335e-18, 9.262451e-18, 9.466358e-18, 9.543417e-18, 
    9.71374e-18, 9.55481e-18, 9.548698e-18, 9.513427e-18,
  1.017767e-17, 9.901928e-18, 1.06116e-17, 1.049977e-17, 9.947212e-18, 
    1.000357e-17, 1.010459e-17, 1.029783e-17, 9.611855e-18, 9.198451e-18, 
    8.771393e-18, 8.211079e-18, 8.119172e-18, 7.791127e-18, 7.79037e-18, 
    8.014176e-18, 7.947424e-18, 8.144726e-18, 7.871806e-18, 8.050958e-18, 
    8.719962e-18, 9.414026e-18, 9.918099e-18, 1.032557e-17, 1.036977e-17, 
    1.033016e-17, 1.067939e-17, 1.080624e-17, 1.073229e-17,
  8.856326e-18, 8.822737e-18, 9.192097e-18, 9.129006e-18, 9.288254e-18, 
    9.279236e-18, 9.078872e-18, 8.702548e-18, 8.477793e-18, 8.047588e-18, 
    7.755339e-18, 7.443301e-18, 7.138093e-18, 6.808658e-18, 6.62688e-18, 
    6.498078e-18, 6.738067e-18, 7.140456e-18, 7.255137e-18, 7.264073e-18, 
    7.641978e-18, 8.091423e-18, 8.515925e-18, 8.512875e-18, 8.708808e-18, 
    8.810704e-18, 8.670078e-18, 8.909088e-18, 9.050466e-18,
  5.805357e-18, 5.86775e-18, 5.769914e-18, 5.980266e-18, 6.283358e-18, 
    6.381583e-18, 6.060596e-18, 5.872539e-18, 5.662115e-18, 5.677145e-18, 
    5.692037e-18, 5.673929e-18, 5.613959e-18, 5.38921e-18, 5.201506e-18, 
    4.981702e-18, 4.90008e-18, 4.931942e-18, 5.032516e-18, 5.186048e-18, 
    5.418617e-18, 5.646916e-18, 5.724858e-18, 5.541123e-18, 5.648706e-18, 
    5.834053e-18, 5.798137e-18, 5.738119e-18, 5.849169e-18,
  3.328421e-18, 3.290345e-18, 3.335255e-18, 3.444658e-18, 3.599759e-18, 
    3.67817e-18, 3.686349e-18, 3.586024e-18, 3.431103e-18, 3.345855e-18, 
    3.222203e-18, 3.245846e-18, 3.257964e-18, 3.26227e-18, 3.290304e-18, 
    3.281655e-18, 3.370318e-18, 3.389905e-18, 3.291865e-18, 3.313524e-18, 
    3.460797e-18, 3.578121e-18, 3.611899e-18, 3.730753e-18, 3.681278e-18, 
    3.646911e-18, 3.457343e-18, 3.375221e-18, 3.357063e-18,
  2.252428e-18, 2.233232e-18, 2.149543e-18, 2.209388e-18, 2.260287e-18, 
    2.282651e-18, 2.227822e-18, 2.123999e-18, 2.092289e-18, 2.040883e-18, 
    1.989161e-18, 1.951502e-18, 1.881841e-18, 1.795531e-18, 1.758878e-18, 
    1.694124e-18, 1.664642e-18, 1.670671e-18, 1.727097e-18, 1.790647e-18, 
    1.938364e-18, 2.107028e-18, 2.218511e-18, 2.265122e-18, 2.400018e-18, 
    2.453733e-18, 2.437233e-18, 2.420937e-18, 2.375716e-18,
  1.275335e-18, 1.315067e-18, 1.365863e-18, 1.380446e-18, 1.508995e-18, 
    1.630455e-18, 1.809213e-18, 1.741367e-18, 1.609068e-18, 1.449787e-18, 
    1.314828e-18, 1.179775e-18, 1.105425e-18, 1.009371e-18, 9.002402e-19, 
    8.139616e-19, 7.819452e-19, 7.347181e-19, 7.166871e-19, 6.949077e-19, 
    7.042017e-19, 7.754284e-19, 9.053389e-19, 9.754969e-19, 1.124961e-18, 
    1.189196e-18, 1.27889e-18, 1.332191e-18, 1.346479e-18,
  7.297035e-19, 7.232628e-19, 7.754188e-19, 8.703986e-19, 9.416114e-19, 
    1.016757e-18, 1.112574e-18, 1.222495e-18, 1.285005e-18, 1.159595e-18, 
    1.003369e-18, 8.764517e-19, 7.633253e-19, 6.910962e-19, 6.280154e-19, 
    5.779921e-19, 5.343221e-19, 4.712265e-19, 4.144207e-19, 3.862302e-19, 
    3.727035e-19, 3.532103e-19, 3.660703e-19, 4.293083e-19, 4.891665e-19, 
    5.195818e-19, 5.353863e-19, 5.927518e-19, 6.548237e-19,
  3.856631e-19, 4.524316e-19, 5.17615e-19, 5.557725e-19, 6.200509e-19, 
    6.622243e-19, 6.75621e-19, 7.326402e-19, 8.222814e-19, 8.17167e-19, 
    7.940709e-19, 7.191267e-19, 6.371172e-19, 5.893461e-19, 5.433711e-19, 
    5.051215e-19, 4.805239e-19, 4.362337e-19, 3.525428e-19, 3.203061e-19, 
    2.923649e-19, 2.594215e-19, 2.440137e-19, 2.413154e-19, 2.598589e-19, 
    2.659854e-19, 2.613845e-19, 2.878961e-19, 3.45867e-19,
  2.898945e-19, 3.195323e-19, 3.749056e-19, 4.082873e-19, 4.396809e-19, 
    4.879304e-19, 5.038373e-19, 5.171666e-19, 5.429365e-19, 5.596609e-19, 
    5.650533e-19, 5.575887e-19, 5.55936e-19, 5.475022e-19, 5.290081e-19, 
    4.727192e-19, 4.042734e-19, 3.58999e-19, 3.353387e-19, 3.031073e-19, 
    2.688815e-19, 2.448446e-19, 2.326755e-19, 2.31612e-19, 2.433072e-19, 
    2.45376e-19, 2.446238e-19, 2.571236e-19, 2.777883e-19,
  6.112494e-20, 6.112494e-20, 6.112494e-20, 6.112494e-20, 6.112494e-20, 
    6.112494e-20, 6.112494e-20, 6.236226e-20, 6.236226e-20, 6.236226e-20, 
    6.236226e-20, 6.236226e-20, 6.236226e-20, 6.236226e-20, 5.756621e-20, 
    5.756621e-20, 5.756621e-20, 5.756621e-20, 5.756621e-20, 5.756621e-20, 
    5.756621e-20, 5.646822e-20, 5.646822e-20, 5.646822e-20, 5.646822e-20, 
    5.646822e-20, 5.646822e-20, 5.646822e-20, 6.112494e-20,
  1.626581e-19, 1.928468e-19, 2.207442e-19, 2.367029e-19, 2.61319e-19, 
    2.65637e-19, 2.62481e-19, 2.515832e-19, 2.355403e-19, 2.233594e-19, 
    2.140054e-19, 1.930589e-19, 1.7685e-19, 1.643728e-19, 1.48688e-19, 
    1.331004e-19, 1.215216e-19, 1.112045e-19, 9.713811e-20, 8.606236e-20, 
    7.719029e-20, 7.125107e-20, 7.195401e-20, 7.765164e-20, 8.234734e-20, 
    9.183363e-20, 1.057524e-19, 1.234391e-19, 1.513517e-19,
  7.645142e-19, 8.242957e-19, 8.786997e-19, 8.990231e-19, 9.30723e-19, 
    9.470894e-19, 9.73505e-19, 9.755315e-19, 9.671617e-19, 9.196267e-19, 
    8.565632e-19, 7.744088e-19, 7.213221e-19, 6.804226e-19, 6.44499e-19, 
    6.172175e-19, 5.765678e-19, 5.245054e-19, 4.677461e-19, 4.22335e-19, 
    3.818529e-19, 3.683765e-19, 3.519592e-19, 5.013088e-19, 5.293777e-19, 
    5.814367e-19, 6.327831e-19, 6.876941e-19, 7.35204e-19,
  3.044912e-18, 3.173055e-18, 3.183955e-18, 3.321957e-18, 3.363808e-18, 
    3.309506e-18, 3.20165e-18, 3.012913e-18, 2.866162e-18, 2.742941e-18, 
    2.588487e-18, 2.421178e-18, 2.373955e-18, 2.354949e-18, 2.2322e-18, 
    2.098062e-18, 2.015503e-18, 1.916023e-18, 1.865674e-18, 2.028064e-18, 
    2.293095e-18, 2.476965e-18, 2.382531e-18, 2.213106e-18, 2.192546e-18, 
    2.27588e-18, 2.340323e-18, 2.565857e-18, 2.844722e-18,
  7.523482e-18, 7.112064e-18, 6.806023e-18, 6.704989e-18, 6.564148e-18, 
    6.467144e-18, 6.493238e-18, 6.406231e-18, 6.28094e-18, 6.22488e-18, 
    6.445141e-18, 6.587706e-18, 6.48831e-18, 6.265461e-18, 6.437482e-18, 
    6.595322e-18, 6.598947e-18, 6.494454e-18, 6.193495e-18, 6.203788e-18, 
    6.530537e-18, 6.542816e-18, 6.649819e-18, 7.045345e-18, 7.45595e-18, 
    7.341457e-18, 7.518295e-18, 7.732288e-18, 7.454684e-18,
  1.664108e-17, 1.569898e-17, 1.486063e-17, 1.45215e-17, 1.442691e-17, 
    1.39543e-17, 1.440192e-17, 1.425604e-17, 1.444891e-17, 1.447679e-17, 
    1.444421e-17, 1.442431e-17, 1.467162e-17, 1.414215e-17, 1.402401e-17, 
    1.394296e-17, 1.4053e-17, 1.408447e-17, 1.466965e-17, 1.53107e-17, 
    1.577757e-17, 1.632022e-17, 1.702419e-17, 1.742578e-17, 1.735737e-17, 
    1.721096e-17, 1.662754e-17, 1.674827e-17, 1.69421e-17,
  2.367196e-17, 2.37269e-17, 2.336516e-17, 2.427363e-17, 2.491568e-17, 
    2.524846e-17, 2.4719e-17, 2.315555e-17, 2.384038e-17, 2.336454e-17, 
    2.393202e-17, 2.360594e-17, 2.304761e-17, 2.288398e-17, 2.28995e-17, 
    2.306385e-17, 2.46759e-17, 2.482307e-17, 2.450299e-17, 2.494919e-17, 
    2.572784e-17, 2.573072e-17, 2.60261e-17, 2.523013e-17, 2.515154e-17, 
    2.484066e-17, 2.445574e-17, 2.418321e-17, 2.400043e-17,
  3.139806e-17, 3.42724e-17, 3.424835e-17, 3.28291e-17, 3.50522e-17, 
    3.624508e-17, 3.615791e-17, 3.723224e-17, 3.751321e-17, 3.388355e-17, 
    3.432689e-17, 3.285153e-17, 3.368191e-17, 3.243543e-17, 3.275453e-17, 
    3.328891e-17, 3.292122e-17, 3.304474e-17, 3.250974e-17, 3.184649e-17, 
    3.197734e-17, 3.255488e-17, 3.29605e-17, 3.346158e-17, 3.443501e-17, 
    3.316509e-17, 3.227477e-17, 3.331256e-17, 3.243012e-17,
  5.104998e-17, 4.91873e-17, 5.115426e-17, 5.179897e-17, 5.156395e-17, 
    5.288479e-17, 5.464574e-17, 5.411195e-17, 5.39852e-17, 5.075914e-17, 
    4.807899e-17, 4.653867e-17, 4.405032e-17, 4.353702e-17, 4.334721e-17, 
    4.541258e-17, 4.355763e-17, 4.189293e-17, 4.290899e-17, 4.44646e-17, 
    4.408426e-17, 4.734303e-17, 5.0812e-17, 5.003158e-17, 5.169061e-17, 
    5.138232e-17, 5.129099e-17, 5.062849e-17, 5.216546e-17,
  5.484931e-17, 5.377593e-17, 5.350345e-17, 5.367153e-17, 5.423013e-17, 
    5.289255e-17, 5.112727e-17, 4.952001e-17, 4.753368e-17, 4.604277e-17, 
    4.468909e-17, 4.39126e-17, 4.214769e-17, 4.154939e-17, 4.221515e-17, 
    4.159245e-17, 4.087607e-17, 4.073141e-17, 4.199738e-17, 4.390461e-17, 
    4.641038e-17, 4.776722e-17, 4.788598e-17, 5.172723e-17, 5.224924e-17, 
    5.174633e-17, 5.336741e-17, 5.469684e-17, 5.387476e-17,
  4.683722e-17, 4.740986e-17, 4.792071e-17, 5.042334e-17, 4.751986e-17, 
    5.047276e-17, 4.816343e-17, 4.56867e-17, 4.568087e-17, 4.403369e-17, 
    4.294138e-17, 4.182808e-17, 3.848028e-17, 3.846106e-17, 3.836582e-17, 
    3.784473e-17, 3.921498e-17, 3.746197e-17, 4.019166e-17, 4.015143e-17, 
    4.03692e-17, 4.108266e-17, 4.254115e-17, 4.378779e-17, 4.582816e-17, 
    4.560005e-17, 4.655987e-17, 4.648535e-17, 4.835561e-17,
  3.570619e-17, 3.629757e-17, 3.591264e-17, 3.629365e-17, 3.726121e-17, 
    3.603898e-17, 3.401864e-17, 3.445019e-17, 3.327743e-17, 3.298572e-17, 
    3.315192e-17, 3.307473e-17, 3.317647e-17, 3.102274e-17, 3.053187e-17, 
    2.947388e-17, 2.86861e-17, 2.9564e-17, 3.131473e-17, 3.123277e-17, 
    3.150979e-17, 3.247116e-17, 3.40042e-17, 3.322636e-17, 3.465379e-17, 
    3.527143e-17, 3.531356e-17, 3.481173e-17, 3.638109e-17,
  2.475624e-17, 2.493589e-17, 2.615915e-17, 2.616324e-17, 2.540718e-17, 
    2.508084e-17, 2.419733e-17, 2.31183e-17, 2.085994e-17, 2.088511e-17, 
    2.061425e-17, 2.067261e-17, 2.078427e-17, 1.976926e-17, 1.979522e-17, 
    1.895898e-17, 1.979081e-17, 2.04431e-17, 2.045295e-17, 2.147699e-17, 
    2.279193e-17, 2.40897e-17, 2.479874e-17, 2.566599e-17, 2.511508e-17, 
    2.541837e-17, 2.528303e-17, 2.531257e-17, 2.501958e-17,
  1.825896e-17, 1.827711e-17, 1.758178e-17, 1.710428e-17, 1.622817e-17, 
    1.580218e-17, 1.543724e-17, 1.461729e-17, 1.350395e-17, 1.285084e-17, 
    1.29653e-17, 1.190689e-17, 1.174572e-17, 1.108134e-17, 1.0479e-17, 
    9.578628e-18, 9.126705e-18, 8.711521e-18, 9.02568e-18, 9.558518e-18, 
    1.061625e-17, 1.251769e-17, 1.381434e-17, 1.503895e-17, 1.585948e-17, 
    1.677784e-17, 1.656083e-17, 1.717023e-17, 1.776088e-17,
  8.688053e-18, 8.646608e-18, 8.66592e-18, 9.039977e-18, 9.194718e-18, 
    1.04694e-17, 1.194626e-17, 1.136212e-17, 1.028161e-17, 9.214655e-18, 
    7.925516e-18, 6.776549e-18, 5.863913e-18, 5.65932e-18, 5.264546e-18, 
    4.975622e-18, 4.508893e-18, 4.10088e-18, 3.738048e-18, 3.581021e-18, 
    3.501638e-18, 3.419511e-18, 3.713668e-18, 4.408887e-18, 5.363157e-18, 
    6.325192e-18, 7.169269e-18, 8.114088e-18, 8.483899e-18,
  2.947679e-18, 3.171073e-18, 3.840174e-18, 3.962778e-18, 4.589684e-18, 
    5.266767e-18, 7.092642e-18, 8.192525e-18, 8.311279e-18, 6.867759e-18, 
    5.846666e-18, 5.154062e-18, 4.660218e-18, 4.53007e-18, 4.14221e-18, 
    3.733351e-18, 3.299989e-18, 3.019645e-18, 2.565334e-18, 1.987641e-18, 
    1.716672e-18, 1.562788e-18, 1.458107e-18, 1.422754e-18, 1.597083e-18, 
    1.794278e-18, 2.009504e-18, 2.199453e-18, 2.427831e-18,
  1.165692e-18, 1.477867e-18, 1.881795e-18, 2.436759e-18, 2.796458e-18, 
    3.40826e-18, 4.132795e-18, 5.086024e-18, 5.149978e-18, 5.14455e-18, 
    5.017042e-18, 4.7851e-18, 4.660682e-18, 4.267579e-18, 3.997289e-18, 
    3.602641e-18, 3.097272e-18, 2.499992e-18, 1.956089e-18, 1.457687e-18, 
    1.217356e-18, 1.170574e-18, 1.032151e-18, 8.54683e-19, 7.344313e-19, 
    7.126125e-19, 7.834199e-19, 8.629106e-19, 9.941743e-19,
  9.299219e-19, 1.031231e-18, 1.253755e-18, 1.49131e-18, 1.832101e-18, 
    2.127719e-18, 2.338539e-18, 2.653864e-18, 2.995652e-18, 3.180016e-18, 
    3.252579e-18, 3.242834e-18, 3.216224e-18, 3.060987e-18, 2.785877e-18, 
    2.500204e-18, 2.15762e-18, 1.792709e-18, 1.601444e-18, 1.410711e-18, 
    1.277108e-18, 1.145361e-18, 1.027038e-18, 9.237148e-19, 8.803068e-19, 
    8.145993e-19, 7.893254e-19, 8.008312e-19, 8.930503e-19,
  1.096101e-19, 1.096101e-19, 1.096101e-19, 1.096101e-19, 1.096101e-19, 
    1.096101e-19, 1.096101e-19, 1.116613e-19, 1.116613e-19, 1.116613e-19, 
    1.116613e-19, 1.116613e-19, 1.116613e-19, 1.116613e-19, 1.073396e-19, 
    1.073396e-19, 1.073396e-19, 1.073396e-19, 1.073396e-19, 1.073396e-19, 
    1.073396e-19, 1.054433e-19, 1.054433e-19, 1.054433e-19, 1.054433e-19, 
    1.054433e-19, 1.054433e-19, 1.054433e-19, 1.096101e-19,
  2.749104e-19, 3.449383e-19, 4.178221e-19, 4.751709e-19, 5.756601e-19, 
    6.140596e-19, 6.114308e-19, 5.862263e-19, 5.247349e-19, 4.615378e-19, 
    4.220895e-19, 3.710078e-19, 3.289759e-19, 2.914486e-19, 2.624829e-19, 
    2.373526e-19, 2.15823e-19, 1.97405e-19, 1.726332e-19, 1.585687e-19, 
    1.496388e-19, 1.406598e-19, 1.345211e-19, 1.359625e-19, 1.42808e-19, 
    1.70081e-19, 1.942016e-19, 2.22735e-19, 2.536156e-19,
  2.382392e-18, 2.638433e-18, 2.749642e-18, 2.905979e-18, 2.965543e-18, 
    2.9957e-18, 3.029488e-18, 3.034502e-18, 3.011245e-18, 2.916302e-18, 
    2.854419e-18, 2.495935e-18, 2.206496e-18, 1.900582e-18, 1.62729e-18, 
    1.373079e-18, 1.2491e-18, 1.081671e-18, 9.297976e-19, 8.339075e-19, 
    7.587267e-19, 7.023828e-19, 6.977462e-19, 7.555292e-19, 9.994634e-19, 
    1.744251e-18, 2.06719e-18, 2.134097e-18, 2.378762e-18,
  9.680448e-18, 1.013353e-17, 1.017459e-17, 1.019568e-17, 1.106327e-17, 
    1.140933e-17, 1.184011e-17, 1.161251e-17, 1.113272e-17, 1.055587e-17, 
    9.947746e-18, 8.974623e-18, 8.613554e-18, 8.260056e-18, 7.876362e-18, 
    7.592866e-18, 7.092041e-18, 6.945706e-18, 6.547694e-18, 6.51294e-18, 
    6.432921e-18, 7.39466e-18, 8.979114e-18, 9.681664e-18, 1.019946e-17, 
    7.953909e-18, 8.17718e-18, 8.709436e-18, 9.284374e-18,
  3.466571e-17, 3.299785e-17, 3.084031e-17, 2.999608e-17, 2.935709e-17, 
    2.938191e-17, 2.890123e-17, 2.870471e-17, 2.852499e-17, 2.835195e-17, 
    2.915937e-17, 3.081571e-17, 3.20345e-17, 3.151684e-17, 3.118879e-17, 
    3.162733e-17, 3.210976e-17, 3.274404e-17, 3.388574e-17, 3.36038e-17, 
    3.268246e-17, 3.3102e-17, 3.392865e-17, 3.419855e-17, 3.612203e-17, 
    3.468164e-17, 3.436565e-17, 3.452245e-17, 3.397763e-17,
  7.165715e-17, 7.037917e-17, 6.645969e-17, 6.662802e-17, 6.64817e-17, 
    6.525509e-17, 6.625203e-17, 6.578296e-17, 6.857577e-17, 6.898922e-17, 
    6.839135e-17, 6.730585e-17, 6.755935e-17, 6.780705e-17, 6.450577e-17, 
    6.435216e-17, 6.418701e-17, 6.339181e-17, 6.408201e-17, 6.590877e-17, 
    6.839237e-17, 6.95192e-17, 7.059057e-17, 7.077082e-17, 7.223613e-17, 
    7.141246e-17, 7.249723e-17, 7.373002e-17, 7.37021e-17,
  1.124425e-16, 1.114116e-16, 1.152911e-16, 1.204139e-16, 1.224432e-16, 
    1.202093e-16, 1.17249e-16, 1.148774e-16, 1.111662e-16, 1.09014e-16, 
    1.088843e-16, 1.063054e-16, 1.039652e-16, 1.056993e-16, 1.01695e-16, 
    1.00501e-16, 1.030736e-16, 1.072217e-16, 1.08846e-16, 1.092401e-16, 
    1.116468e-16, 1.114391e-16, 1.128199e-16, 1.135062e-16, 1.112101e-16, 
    1.150295e-16, 1.146727e-16, 1.132895e-16, 1.118091e-16,
  1.676589e-16, 1.739366e-16, 1.866469e-16, 1.815216e-16, 1.886286e-16, 
    1.875146e-16, 1.868382e-16, 1.814179e-16, 1.987995e-16, 1.830764e-16, 
    1.801554e-16, 1.789939e-16, 1.781503e-16, 1.784478e-16, 1.695616e-16, 
    1.641607e-16, 1.728625e-16, 1.735046e-16, 1.596226e-16, 1.640641e-16, 
    1.659257e-16, 1.692865e-16, 1.747587e-16, 1.726167e-16, 1.723093e-16, 
    1.761571e-16, 1.737143e-16, 1.703615e-16, 1.705665e-16,
  2.56512e-16, 2.661117e-16, 2.628947e-16, 2.670689e-16, 2.701656e-16, 
    2.72974e-16, 2.77496e-16, 2.643248e-16, 2.611678e-16, 2.606825e-16, 
    2.531754e-16, 2.436036e-16, 2.295093e-16, 2.38817e-16, 2.214784e-16, 
    2.161636e-16, 2.127549e-16, 2.185745e-16, 2.247161e-16, 2.235008e-16, 
    2.228553e-16, 2.351843e-16, 2.415425e-16, 2.527427e-16, 2.515208e-16, 
    2.526907e-16, 2.491935e-16, 2.560796e-16, 2.639074e-16,
  2.961016e-16, 2.925044e-16, 2.779743e-16, 2.756996e-16, 2.722525e-16, 
    2.71046e-16, 2.667076e-16, 2.442615e-16, 2.35702e-16, 2.295207e-16, 
    2.302693e-16, 2.226042e-16, 2.062844e-16, 2.078262e-16, 2.114586e-16, 
    2.113109e-16, 2.120199e-16, 2.080604e-16, 2.174978e-16, 2.311295e-16, 
    2.450471e-16, 2.426363e-16, 2.389079e-16, 2.615756e-16, 2.606727e-16, 
    2.622719e-16, 2.726035e-16, 2.931522e-16, 3.08589e-16,
  2.664886e-16, 2.628072e-16, 2.621013e-16, 2.669651e-16, 2.666419e-16, 
    2.646928e-16, 2.529435e-16, 2.424186e-16, 2.338256e-16, 2.286057e-16, 
    2.205229e-16, 2.053865e-16, 1.994748e-16, 2.014716e-16, 2.020327e-16, 
    2.085713e-16, 2.161246e-16, 2.158581e-16, 2.215286e-16, 2.274456e-16, 
    2.322256e-16, 2.299961e-16, 2.317598e-16, 2.364071e-16, 2.246021e-16, 
    2.385106e-16, 2.501434e-16, 2.542209e-16, 2.600207e-16,
  2.018796e-16, 1.836969e-16, 1.808311e-16, 1.778647e-16, 1.822204e-16, 
    1.757158e-16, 1.786308e-16, 1.746654e-16, 1.800286e-16, 1.850251e-16, 
    1.871815e-16, 1.78256e-16, 1.680382e-16, 1.660473e-16, 1.687723e-16, 
    1.720524e-16, 1.643885e-16, 1.627149e-16, 1.61884e-16, 1.687316e-16, 
    1.739777e-16, 1.944978e-16, 1.936827e-16, 1.856658e-16, 1.762372e-16, 
    1.807263e-16, 1.915927e-16, 1.990098e-16, 1.980735e-16,
  1.17809e-16, 1.199605e-16, 1.192116e-16, 1.165059e-16, 1.092235e-16, 
    1.030513e-16, 9.993037e-17, 9.131381e-17, 8.497892e-17, 8.605351e-17, 
    8.508467e-17, 8.347328e-17, 8.820466e-17, 9.015688e-17, 8.924023e-17, 
    8.569841e-17, 9.100589e-17, 9.776665e-17, 9.714989e-17, 9.885807e-17, 
    1.007523e-16, 1.059095e-16, 1.163077e-16, 1.241008e-16, 1.25566e-16, 
    1.246511e-16, 1.240318e-16, 1.229528e-16, 1.200769e-16,
  7.95359e-17, 7.53846e-17, 7.51618e-17, 7.104201e-17, 6.667254e-17, 
    6.350997e-17, 6.215534e-17, 5.795849e-17, 5.298586e-17, 4.728739e-17, 
    4.620019e-17, 4.521274e-17, 4.308455e-17, 4.317583e-17, 4.1777e-17, 
    3.78217e-17, 3.688077e-17, 3.624524e-17, 3.692579e-17, 4.202935e-17, 
    4.787885e-17, 5.215456e-17, 5.568484e-17, 6.150812e-17, 6.546014e-17, 
    6.890868e-17, 7.453078e-17, 7.768626e-17, 7.85536e-17,
  3.789606e-17, 3.669976e-17, 3.928547e-17, 3.556165e-17, 3.231616e-17, 
    3.291956e-17, 3.619186e-17, 3.381148e-17, 3.31543e-17, 3.039143e-17, 
    2.687291e-17, 2.450798e-17, 2.208111e-17, 2.261259e-17, 2.021984e-17, 
    1.854772e-17, 1.715339e-17, 1.65847e-17, 1.524339e-17, 1.384286e-17, 
    1.352683e-17, 1.271694e-17, 1.241711e-17, 1.515112e-17, 2.3374e-17, 
    2.854035e-17, 3.325981e-17, 3.555191e-17, 3.668829e-17,
  7.377123e-18, 9.040106e-18, 1.120748e-17, 1.272003e-17, 1.46349e-17, 
    1.660446e-17, 2.015714e-17, 2.531048e-17, 2.659759e-17, 2.493653e-17, 
    2.286511e-17, 2.009993e-17, 1.713701e-17, 1.579538e-17, 1.451919e-17, 
    1.253337e-17, 1.144894e-17, 1.136122e-17, 8.96126e-18, 7.197902e-18, 
    5.961269e-18, 4.903587e-18, 4.309599e-18, 4.106762e-18, 4.173058e-18, 
    4.172901e-18, 4.860813e-18, 5.574401e-18, 6.457668e-18,
  2.940144e-18, 3.640027e-18, 4.932976e-18, 6.176662e-18, 7.096029e-18, 
    9.932484e-18, 1.217771e-17, 1.486681e-17, 1.780875e-17, 1.850241e-17, 
    1.875463e-17, 1.859685e-17, 1.735023e-17, 1.646515e-17, 1.481642e-17, 
    1.334479e-17, 1.206199e-17, 9.749803e-18, 7.477824e-18, 6.227391e-18, 
    4.753393e-18, 3.582653e-18, 3.36494e-18, 2.832212e-18, 2.266472e-18, 
    1.99366e-18, 1.910609e-18, 2.343849e-18, 2.832416e-18,
  2.497252e-18, 2.786942e-18, 3.288281e-18, 3.815723e-18, 4.61265e-18, 
    5.318598e-18, 6.070433e-18, 7.413504e-18, 8.712968e-18, 9.752924e-18, 
    1.039136e-17, 1.076927e-17, 1.081664e-17, 1.045702e-17, 9.719169e-18, 
    8.624976e-18, 7.333288e-18, 6.07042e-18, 5.446651e-18, 4.845043e-18, 
    4.012056e-18, 3.497684e-18, 3.284836e-18, 2.948488e-18, 2.705159e-18, 
    2.428389e-18, 2.288564e-18, 2.271353e-18, 2.378349e-18,
  2.335068e-19, 2.335068e-19, 2.335068e-19, 2.335068e-19, 2.335068e-19, 
    2.335068e-19, 2.335068e-19, 2.389021e-19, 2.389021e-19, 2.389021e-19, 
    2.389021e-19, 2.389021e-19, 2.389021e-19, 2.389021e-19, 2.410549e-19, 
    2.410549e-19, 2.410549e-19, 2.410549e-19, 2.410549e-19, 2.410549e-19, 
    2.410549e-19, 2.354581e-19, 2.354581e-19, 2.354581e-19, 2.354581e-19, 
    2.354581e-19, 2.354581e-19, 2.354581e-19, 2.335068e-19,
  4.396797e-19, 5.745231e-19, 6.913455e-19, 8.172092e-19, 1.007203e-18, 
    1.102303e-18, 1.136197e-18, 1.110544e-18, 9.686592e-19, 8.292545e-19, 
    7.620054e-19, 6.75499e-19, 5.716464e-19, 5.191885e-19, 4.772196e-19, 
    4.201365e-19, 3.614202e-19, 3.046351e-19, 2.652612e-19, 2.60987e-19, 
    2.828691e-19, 3.007027e-19, 3.056009e-19, 3.028018e-19, 2.835445e-19, 
    2.780156e-19, 2.994245e-19, 3.387148e-19, 3.969713e-19,
  4.279811e-18, 5.22291e-18, 5.480036e-18, 6.205282e-18, 6.85807e-18, 
    7.255761e-18, 7.508974e-18, 7.197593e-18, 7.173622e-18, 7.087698e-18, 
    6.921072e-18, 6.140906e-18, 5.42467e-18, 4.3577e-18, 3.24755e-18, 
    2.566933e-18, 2.314162e-18, 2.109469e-18, 1.659283e-18, 1.214128e-18, 
    8.230193e-19, 6.373858e-19, 6.751997e-19, 7.642937e-19, 7.953298e-19, 
    1.138093e-18, 2.255679e-18, 3.705268e-18, 3.979098e-18,
  2.341631e-17, 2.576996e-17, 2.575386e-17, 2.379277e-17, 2.32023e-17, 
    2.527585e-17, 2.681189e-17, 2.784341e-17, 2.802461e-17, 2.805042e-17, 
    2.77273e-17, 2.660993e-17, 2.599417e-17, 2.496126e-17, 2.232213e-17, 
    2.049858e-17, 1.890571e-17, 1.789113e-17, 1.784605e-17, 1.504488e-17, 
    1.454716e-17, 1.400686e-17, 1.297341e-17, 2.377292e-17, 3.122905e-17, 
    2.877274e-17, 1.721389e-17, 1.789456e-17, 1.998926e-17,
  1.067579e-16, 1.035442e-16, 9.786767e-17, 9.258308e-17, 9.464706e-17, 
    9.634311e-17, 9.378426e-17, 9.287373e-17, 9.552231e-17, 9.49405e-17, 
    9.869417e-17, 1.009295e-16, 9.983507e-17, 1.046625e-16, 1.042285e-16, 
    1.050662e-16, 1.077813e-16, 1.135305e-16, 1.176145e-16, 1.274556e-16, 
    1.306018e-16, 1.333518e-16, 1.347652e-16, 1.267263e-16, 1.274656e-16, 
    1.217086e-16, 1.200727e-16, 1.177597e-16, 1.114555e-16,
  2.680539e-16, 2.692678e-16, 2.594164e-16, 2.604455e-16, 2.568634e-16, 
    2.569912e-16, 2.551455e-16, 2.447808e-16, 2.497883e-16, 2.501823e-16, 
    2.356554e-16, 2.308922e-16, 2.281232e-16, 2.366644e-16, 2.336347e-16, 
    2.374987e-16, 2.354456e-16, 2.360899e-16, 2.494243e-16, 2.532708e-16, 
    2.672567e-16, 2.582616e-16, 2.59294e-16, 2.600205e-16, 2.592975e-16, 
    2.637387e-16, 2.69396e-16, 2.678164e-16, 2.731958e-16,
  4.425421e-16, 4.352795e-16, 4.448294e-16, 4.87146e-16, 4.829673e-16, 
    4.768413e-16, 4.917314e-16, 4.891677e-16, 4.681711e-16, 4.644354e-16, 
    4.530724e-16, 4.28984e-16, 4.299712e-16, 4.151016e-16, 3.935584e-16, 
    3.927808e-16, 3.796682e-16, 3.853449e-16, 4.058378e-16, 4.082596e-16, 
    4.122789e-16, 4.287886e-16, 4.427462e-16, 4.262842e-16, 4.116707e-16, 
    4.233166e-16, 4.360727e-16, 4.366612e-16, 4.365802e-16,
  8.159915e-16, 8.414362e-16, 8.734494e-16, 8.503762e-16, 8.38749e-16, 
    8.661025e-16, 8.417694e-16, 8.862944e-16, 9.053215e-16, 8.608762e-16, 
    8.526639e-16, 8.17425e-16, 7.900614e-16, 8.035625e-16, 7.990952e-16, 
    7.629073e-16, 7.509945e-16, 7.795861e-16, 7.890004e-16, 7.912354e-16, 
    7.852122e-16, 8.199144e-16, 8.142751e-16, 8.435106e-16, 8.342893e-16, 
    8.96109e-16, 8.788559e-16, 8.110053e-16, 7.959441e-16,
  1.243384e-15, 1.248319e-15, 1.280416e-15, 1.315563e-15, 1.292588e-15, 
    1.269097e-15, 1.246039e-15, 1.231218e-15, 1.255224e-15, 1.186175e-15, 
    1.107748e-15, 1.076941e-15, 1.069387e-15, 1.079702e-15, 1.074835e-15, 
    1.060815e-15, 1.069323e-15, 1.101849e-15, 1.107595e-15, 1.154503e-15, 
    1.170819e-15, 1.24906e-15, 1.268739e-15, 1.31958e-15, 1.307903e-15, 
    1.324602e-15, 1.274601e-15, 1.299945e-15, 1.282414e-15,
  1.396663e-15, 1.411299e-15, 1.391478e-15, 1.338858e-15, 1.354646e-15, 
    1.33696e-15, 1.277117e-15, 1.232253e-15, 1.229086e-15, 1.173576e-15, 
    1.150385e-15, 1.114943e-15, 1.074379e-15, 1.097641e-15, 1.054603e-15, 
    1.049788e-15, 1.058437e-15, 1.107762e-15, 1.124895e-15, 1.162151e-15, 
    1.243994e-15, 1.336985e-15, 1.354574e-15, 1.425712e-15, 1.39427e-15, 
    1.349359e-15, 1.378332e-15, 1.412687e-15, 1.405681e-15,
  1.177837e-15, 1.183015e-15, 1.196732e-15, 1.144875e-15, 1.193981e-15, 
    1.164782e-15, 1.177261e-15, 1.125919e-15, 1.084183e-15, 1.029891e-15, 
    9.770568e-16, 9.616387e-16, 9.676264e-16, 9.227652e-16, 9.388072e-16, 
    9.434761e-16, 9.613848e-16, 1.023498e-15, 1.066016e-15, 1.089022e-15, 
    1.141298e-15, 1.158524e-15, 1.194249e-15, 1.196432e-15, 1.194426e-15, 
    1.177216e-15, 1.140577e-15, 1.128847e-15, 1.139769e-15,
  7.976696e-16, 7.438908e-16, 7.332971e-16, 7.240816e-16, 7.353005e-16, 
    7.121352e-16, 6.78749e-16, 7.316325e-16, 7.560322e-16, 7.923576e-16, 
    7.588581e-16, 6.852285e-16, 6.571031e-16, 6.680201e-16, 6.891859e-16, 
    6.897871e-16, 6.895158e-16, 6.756509e-16, 6.786772e-16, 6.820244e-16, 
    7.397881e-16, 7.960585e-16, 8.047797e-16, 7.728573e-16, 7.544537e-16, 
    7.543642e-16, 7.961078e-16, 8.017373e-16, 8.160672e-16,
  3.919442e-16, 3.920635e-16, 3.948839e-16, 3.650768e-16, 3.559882e-16, 
    3.278077e-16, 3.181479e-16, 2.904532e-16, 2.820868e-16, 2.761911e-16, 
    2.624146e-16, 2.618695e-16, 2.799716e-16, 3.080787e-16, 3.05802e-16, 
    2.901128e-16, 3.106887e-16, 3.374783e-16, 3.241359e-16, 3.281263e-16, 
    3.356803e-16, 3.523198e-16, 3.880851e-16, 4.081502e-16, 4.215694e-16, 
    4.035548e-16, 4.031693e-16, 3.967603e-16, 3.96355e-16,
  2.212182e-16, 2.02893e-16, 2.030043e-16, 1.982809e-16, 1.949404e-16, 
    1.778165e-16, 1.648206e-16, 1.477486e-16, 1.389768e-16, 1.334983e-16, 
    1.272625e-16, 1.324282e-16, 1.370185e-16, 1.352115e-16, 1.346852e-16, 
    1.279315e-16, 1.324977e-16, 1.299361e-16, 1.356544e-16, 1.576054e-16, 
    1.733948e-16, 1.85032e-16, 2.006059e-16, 2.141428e-16, 2.000138e-16, 
    2.048435e-16, 2.163141e-16, 2.249202e-16, 2.303228e-16,
  1.004458e-16, 1.009754e-16, 1.008083e-16, 8.945005e-17, 8.338476e-17, 
    8.493621e-17, 8.443008e-17, 7.89096e-17, 7.944194e-17, 7.616285e-17, 
    7.271358e-17, 6.927762e-17, 6.937416e-17, 6.99129e-17, 6.193396e-17, 
    5.907037e-17, 5.853728e-17, 5.549668e-17, 5.191903e-17, 4.935326e-17, 
    4.873645e-17, 4.533732e-17, 4.522535e-17, 5.527138e-17, 7.725388e-17, 
    9.121147e-17, 9.618087e-17, 9.109359e-17, 9.074599e-17,
  1.635943e-17, 1.799083e-17, 2.504643e-17, 2.572588e-17, 3.337286e-17, 
    4.038382e-17, 4.65172e-17, 5.17831e-17, 5.38537e-17, 5.426689e-17, 
    5.172861e-17, 5.041679e-17, 4.532854e-17, 3.977343e-17, 3.770434e-17, 
    3.492991e-17, 3.321733e-17, 3.087589e-17, 2.719302e-17, 2.030788e-17, 
    1.71513e-17, 1.253845e-17, 1.013576e-17, 9.562291e-18, 9.382595e-18, 
    8.975842e-18, 1.041877e-17, 1.182191e-17, 1.519207e-17,
  6.292871e-18, 8.307251e-18, 9.466542e-18, 1.249014e-17, 1.32501e-17, 
    1.825446e-17, 2.502549e-17, 3.30578e-17, 3.88097e-17, 4.33717e-17, 
    4.332638e-17, 4.161617e-17, 3.765217e-17, 3.530735e-17, 3.353193e-17, 
    3.258803e-17, 3.113389e-17, 2.679301e-17, 1.990748e-17, 1.612549e-17, 
    1.222676e-17, 9.028441e-18, 7.416571e-18, 6.047376e-18, 4.985447e-18, 
    3.843186e-18, 3.625562e-18, 3.829954e-18, 4.999158e-18,
  4.705493e-18, 5.193153e-18, 6.187358e-18, 6.998874e-18, 8.244376e-18, 
    9.788204e-18, 1.257464e-17, 1.632954e-17, 1.962698e-17, 2.209064e-17, 
    2.407926e-17, 2.536451e-17, 2.550561e-17, 2.482328e-17, 2.328675e-17, 
    2.081385e-17, 1.823233e-17, 1.562959e-17, 1.41133e-17, 1.215658e-17, 
    9.532111e-18, 8.014392e-18, 7.023783e-18, 6.136113e-18, 4.6991e-18, 
    4.002696e-18, 3.993379e-18, 4.150758e-18, 4.429086e-18,
  7.670262e-19, 7.670262e-19, 7.670262e-19, 7.670262e-19, 7.670262e-19, 
    7.670262e-19, 7.670262e-19, 8.014739e-19, 8.014739e-19, 8.014739e-19, 
    8.014739e-19, 8.014739e-19, 8.014739e-19, 8.014739e-19, 8.446756e-19, 
    8.446756e-19, 8.446756e-19, 8.446756e-19, 8.446756e-19, 8.446756e-19, 
    8.446756e-19, 8.217599e-19, 8.217599e-19, 8.217599e-19, 8.217599e-19, 
    8.217599e-19, 8.217599e-19, 8.217599e-19, 7.670262e-19,
  8.44475e-19, 9.234996e-19, 1.130429e-18, 1.414845e-18, 1.889647e-18, 
    2.173232e-18, 2.284006e-18, 2.205619e-18, 2.010418e-18, 1.905944e-18, 
    1.83159e-18, 1.705106e-18, 1.58444e-18, 1.370553e-18, 1.181878e-18, 
    9.76602e-19, 8.239615e-19, 7.33699e-19, 6.603764e-19, 6.059334e-19, 
    6.041459e-19, 6.627752e-19, 8.271464e-19, 8.995825e-19, 9.320415e-19, 
    9.297337e-19, 7.730587e-19, 7.794052e-19, 8.193236e-19,
  6.632785e-18, 8.938266e-18, 1.114388e-17, 1.495444e-17, 1.874691e-17, 
    2.208152e-17, 2.295156e-17, 2.226172e-17, 1.96992e-17, 1.77646e-17, 
    1.685732e-17, 1.416945e-17, 1.189281e-17, 1.059994e-17, 8.541481e-18, 
    7.664504e-18, 7.388362e-18, 6.788336e-18, 5.709486e-18, 3.877528e-18, 
    2.031597e-18, 1.130512e-18, 1.323143e-18, 1.444564e-18, 1.47271e-18, 
    1.438658e-18, 1.762902e-18, 3.266643e-18, 5.195087e-18,
  6.353666e-17, 8.43087e-17, 8.316535e-17, 7.551666e-17, 7.897706e-17, 
    9.460628e-17, 9.204846e-17, 8.400775e-17, 7.552935e-17, 6.940425e-17, 
    6.936015e-17, 6.977877e-17, 6.634245e-17, 6.632689e-17, 6.870638e-17, 
    7.510794e-17, 7.618175e-17, 7.28688e-17, 7.269005e-17, 6.043392e-17, 
    4.301698e-17, 2.937455e-17, 2.044953e-17, 2.151583e-17, 3.86136e-17, 
    6.619737e-17, 4.987741e-17, 4.212393e-17, 4.964041e-17,
  2.38413e-16, 2.365768e-16, 2.149258e-16, 1.953167e-16, 1.640661e-16, 
    1.623396e-16, 1.584389e-16, 1.616385e-16, 1.661496e-16, 1.737618e-16, 
    1.791934e-16, 1.844385e-16, 1.869821e-16, 1.951451e-16, 2.092889e-16, 
    2.176442e-16, 2.164211e-16, 2.378906e-16, 2.556895e-16, 2.601746e-16, 
    2.951596e-16, 3.360057e-16, 3.75943e-16, 3.496112e-16, 3.350358e-16, 
    3.385703e-16, 2.913968e-16, 2.787913e-16, 2.703917e-16,
  8.576421e-16, 8.377082e-16, 8.439642e-16, 7.650124e-16, 7.342013e-16, 
    7.421794e-16, 7.288532e-16, 6.807521e-16, 6.649772e-16, 6.599712e-16, 
    6.242941e-16, 5.989526e-16, 5.969775e-16, 6.518427e-16, 6.806527e-16, 
    7.185107e-16, 7.389271e-16, 7.415904e-16, 7.559901e-16, 7.971532e-16, 
    8.583909e-16, 8.778801e-16, 8.333089e-16, 8.028656e-16, 7.988508e-16, 
    8.460077e-16, 8.582661e-16, 8.681575e-16, 8.8296e-16,
  1.636666e-15, 1.592595e-15, 1.566135e-15, 1.643685e-15, 1.647253e-15, 
    1.683378e-15, 1.644239e-15, 1.694609e-15, 1.677771e-15, 1.640281e-15, 
    1.660835e-15, 1.581196e-15, 1.560622e-15, 1.443251e-15, 1.460885e-15, 
    1.476566e-15, 1.436401e-15, 1.480034e-15, 1.490616e-15, 1.437093e-15, 
    1.460452e-15, 1.498049e-15, 1.469754e-15, 1.472323e-15, 1.432126e-15, 
    1.475945e-15, 1.521938e-15, 1.582343e-15, 1.626783e-15,
  3.515117e-15, 3.554146e-15, 3.55231e-15, 3.463045e-15, 3.495921e-15, 
    3.405194e-15, 3.513121e-15, 3.61426e-15, 3.545391e-15, 3.468316e-15, 
    3.351574e-15, 3.331949e-15, 3.195988e-15, 3.129567e-15, 3.230697e-15, 
    3.247257e-15, 3.277109e-15, 3.226109e-15, 3.353101e-15, 3.369677e-15, 
    3.417515e-15, 3.493835e-15, 3.609529e-15, 3.628192e-15, 3.600887e-15, 
    3.577862e-15, 3.666081e-15, 3.608504e-15, 3.58472e-15,
  5.746997e-15, 5.770759e-15, 5.664531e-15, 5.846544e-15, 5.82857e-15, 
    5.898612e-15, 5.696066e-15, 5.492152e-15, 5.461265e-15, 5.344424e-15, 
    5.01568e-15, 4.758948e-15, 4.656204e-15, 4.527216e-15, 4.555862e-15, 
    4.603294e-15, 4.622552e-15, 4.66277e-15, 4.983367e-15, 5.061627e-15, 
    5.107805e-15, 5.408236e-15, 5.752903e-15, 5.924205e-15, 5.966135e-15, 
    6.015398e-15, 6.006925e-15, 5.847371e-15, 5.723514e-15,
  5.464408e-15, 5.651675e-15, 5.570036e-15, 5.374245e-15, 5.399319e-15, 
    5.483378e-15, 5.542576e-15, 5.438699e-15, 5.313182e-15, 5.216136e-15, 
    5.025299e-15, 4.905075e-15, 4.596052e-15, 4.665696e-15, 4.689706e-15, 
    4.607448e-15, 4.475528e-15, 4.633202e-15, 4.669844e-15, 4.719712e-15, 
    4.902176e-15, 5.028769e-15, 5.125086e-15, 5.346781e-15, 5.455204e-15, 
    5.422888e-15, 5.191612e-15, 5.334118e-15, 5.41886e-15,
  3.802473e-15, 3.939032e-15, 4.050782e-15, 3.882274e-15, 3.8714e-15, 
    4.062369e-15, 4.015041e-15, 4.083019e-15, 4.034927e-15, 3.759931e-15, 
    3.598348e-15, 3.578088e-15, 3.469846e-15, 3.491726e-15, 3.449171e-15, 
    3.301824e-15, 3.232644e-15, 3.393232e-15, 3.616715e-15, 3.850785e-15, 
    3.882856e-15, 3.853729e-15, 3.905978e-15, 4.131501e-15, 4.213897e-15, 
    4.208235e-15, 4.094894e-15, 3.991083e-15, 3.867689e-15,
  2.555403e-15, 2.482492e-15, 2.561156e-15, 2.498715e-15, 2.414693e-15, 
    2.392282e-15, 2.382417e-15, 2.376025e-15, 2.494137e-15, 2.553298e-15, 
    2.327401e-15, 2.146655e-15, 2.177389e-15, 2.176368e-15, 2.199845e-15, 
    2.131653e-15, 2.060232e-15, 2.133421e-15, 2.282885e-15, 2.316552e-15, 
    2.410214e-15, 2.440826e-15, 2.492559e-15, 2.563358e-15, 2.653166e-15, 
    2.641249e-15, 2.612179e-15, 2.592196e-15, 2.695495e-15,
  1.129122e-15, 1.146288e-15, 1.139373e-15, 1.102928e-15, 1.087478e-15, 
    1.063484e-15, 1.043242e-15, 1.031017e-15, 9.758789e-16, 9.391443e-16, 
    8.877274e-16, 8.887397e-16, 8.82982e-16, 9.203918e-16, 9.127547e-16, 
    8.909711e-16, 9.419285e-16, 9.935119e-16, 9.976696e-16, 1.047897e-15, 
    1.085326e-15, 1.034971e-15, 1.047834e-15, 1.126753e-15, 1.263065e-15, 
    1.247372e-15, 1.250569e-15, 1.248401e-15, 1.153542e-15,
  5.853613e-16, 5.752449e-16, 5.668272e-16, 5.418769e-16, 5.723305e-16, 
    5.276566e-16, 4.66975e-16, 4.268718e-16, 4.407764e-16, 4.267582e-16, 
    4.294606e-16, 4.248508e-16, 4.278023e-16, 4.302192e-16, 4.173209e-16, 
    4.153222e-16, 4.616262e-16, 4.603606e-16, 4.613571e-16, 4.805943e-16, 
    4.914242e-16, 5.465544e-16, 5.305457e-16, 5.189016e-16, 5.261221e-16, 
    5.259724e-16, 5.543549e-16, 5.835653e-16, 5.997382e-16,
  2.030573e-16, 2.047122e-16, 2.041896e-16, 1.931857e-16, 1.939925e-16, 
    1.998536e-16, 2.002573e-16, 1.828885e-16, 1.989887e-16, 2.077214e-16, 
    1.911301e-16, 2.005699e-16, 1.917656e-16, 1.92328e-16, 1.78079e-16, 
    1.876039e-16, 1.883843e-16, 1.76367e-16, 1.651899e-16, 1.609081e-16, 
    1.643947e-16, 1.562179e-16, 1.49114e-16, 1.793944e-16, 1.942191e-16, 
    2.045784e-16, 2.05578e-16, 1.990503e-16, 1.944787e-16,
  2.703283e-17, 3.18638e-17, 4.620539e-17, 5.197194e-17, 6.742505e-17, 
    8.504253e-17, 1.06314e-16, 1.057996e-16, 1.162376e-16, 1.302546e-16, 
    1.239982e-16, 1.33176e-16, 1.419648e-16, 1.326072e-16, 1.289261e-16, 
    1.284567e-16, 1.155489e-16, 9.754946e-17, 8.242488e-17, 6.565506e-17, 
    4.977827e-17, 3.609896e-17, 2.870684e-17, 2.486103e-17, 2.134712e-17, 
    2.155363e-17, 2.413495e-17, 2.516516e-17, 2.601284e-17,
  9.190717e-18, 1.43732e-17, 1.811464e-17, 2.319429e-17, 2.504449e-17, 
    3.178349e-17, 4.753079e-17, 6.208184e-17, 7.844919e-17, 9.054216e-17, 
    9.446162e-17, 1.004311e-16, 9.627329e-17, 9.409752e-17, 9.26828e-17, 
    8.952568e-17, 7.703073e-17, 6.755589e-17, 5.633762e-17, 4.482383e-17, 
    3.424805e-17, 2.710416e-17, 2.075766e-17, 1.317766e-17, 9.407681e-18, 
    7.430578e-18, 7.002137e-18, 7.212046e-18, 7.686506e-18,
  7.970914e-18, 9.734601e-18, 1.168404e-17, 1.316588e-17, 1.63655e-17, 
    2.002944e-17, 2.307589e-17, 3.105201e-17, 4.050032e-17, 4.745707e-17, 
    5.204714e-17, 5.687141e-17, 5.95254e-17, 6.057866e-17, 5.875409e-17, 
    5.471106e-17, 4.907803e-17, 4.282681e-17, 3.811774e-17, 3.276096e-17, 
    2.595456e-17, 1.879961e-17, 1.437915e-17, 1.016442e-17, 7.397914e-18, 
    6.894311e-18, 6.537302e-18, 6.757348e-18, 7.375161e-18,
  3.003618e-18, 3.003618e-18, 3.003618e-18, 3.003618e-18, 3.003618e-18, 
    3.003618e-18, 3.003618e-18, 2.875658e-18, 2.875658e-18, 2.875658e-18, 
    2.875658e-18, 2.875658e-18, 2.875658e-18, 2.875658e-18, 2.728901e-18, 
    2.728901e-18, 2.728901e-18, 2.728901e-18, 2.728901e-18, 2.728901e-18, 
    2.728901e-18, 2.950492e-18, 2.950492e-18, 2.950492e-18, 2.950492e-18, 
    2.950492e-18, 2.950492e-18, 2.950492e-18, 3.003618e-18,
  2.536947e-18, 2.52326e-18, 2.679124e-18, 2.904627e-18, 3.59513e-18, 
    4.56193e-18, 5.436908e-18, 5.643946e-18, 5.73101e-18, 5.745638e-18, 
    5.691529e-18, 5.317043e-18, 5.054266e-18, 4.540417e-18, 3.744995e-18, 
    3.284421e-18, 3.047225e-18, 2.861767e-18, 2.49109e-18, 2.266563e-18, 
    2.007353e-18, 1.900554e-18, 2.337249e-18, 3.311246e-18, 3.428994e-18, 
    3.597148e-18, 3.325762e-18, 2.912662e-18, 2.617464e-18,
  1.208184e-17, 2.074201e-17, 2.818177e-17, 4.408647e-17, 5.676055e-17, 
    6.320341e-17, 7.003227e-17, 7.140824e-17, 7.355794e-17, 6.894122e-17, 
    6.396274e-17, 5.375949e-17, 4.412937e-17, 3.878892e-17, 2.973615e-17, 
    2.587847e-17, 2.222964e-17, 1.98255e-17, 1.666331e-17, 1.120455e-17, 
    5.793061e-18, 4.282769e-18, 5.252044e-18, 5.736711e-18, 6.312394e-18, 
    5.741675e-18, 4.631089e-18, 5.931974e-18, 9.171918e-18,
  2.764565e-16, 3.433845e-16, 3.580285e-16, 3.764547e-16, 4.069744e-16, 
    4.276034e-16, 3.824127e-16, 2.835018e-16, 2.269257e-16, 2.021829e-16, 
    2.094713e-16, 2.347765e-16, 2.512566e-16, 2.700979e-16, 2.718909e-16, 
    2.789007e-16, 2.741181e-16, 2.660747e-16, 2.609358e-16, 2.376021e-16, 
    1.657789e-16, 9.061644e-17, 3.871646e-17, 3.017515e-17, 4.26104e-17, 
    1.009792e-16, 1.264312e-16, 1.288295e-16, 1.812677e-16,
  6.761668e-16, 7.489805e-16, 6.628986e-16, 4.899101e-16, 3.349091e-16, 
    2.994283e-16, 2.962752e-16, 3.348548e-16, 3.480627e-16, 3.612635e-16, 
    3.732806e-16, 3.77935e-16, 3.739393e-16, 3.977822e-16, 4.353085e-16, 
    4.233393e-16, 4.091302e-16, 4.261722e-16, 4.142207e-16, 3.680185e-16, 
    4.567134e-16, 5.150711e-16, 6.750828e-16, 7.020569e-16, 8.420664e-16, 
    7.904819e-16, 7.727207e-16, 8.433647e-16, 7.53e-16,
  2.376646e-15, 2.208071e-15, 2.194052e-15, 1.982242e-15, 1.756918e-15, 
    1.688921e-15, 1.672358e-15, 1.683609e-15, 1.595708e-15, 1.427275e-15, 
    1.41308e-15, 1.338283e-15, 1.325404e-15, 1.451743e-15, 1.569179e-15, 
    1.630965e-15, 1.71282e-15, 1.809104e-15, 1.829315e-15, 2.039613e-15, 
    2.16006e-15, 2.476169e-15, 2.534352e-15, 2.317307e-15, 2.398421e-15, 
    2.660233e-15, 2.517564e-15, 2.663018e-15, 2.485924e-15,
  5.214645e-15, 5.326166e-15, 5.457358e-15, 5.577883e-15, 5.711609e-15, 
    5.515983e-15, 5.334892e-15, 5.324137e-15, 5.166048e-15, 5.104543e-15, 
    5.064759e-15, 4.888474e-15, 4.840156e-15, 5.010482e-15, 5.036255e-15, 
    4.977897e-15, 5.060409e-15, 5.209415e-15, 5.193076e-15, 5.150773e-15, 
    5.2837e-15, 5.359703e-15, 5.414546e-15, 5.304904e-15, 5.336699e-15, 
    5.33475e-15, 5.22459e-15, 5.480967e-15, 5.271088e-15,
  1.355664e-14, 1.303518e-14, 1.336635e-14, 1.294119e-14, 1.27768e-14, 
    1.243913e-14, 1.315956e-14, 1.384331e-14, 1.336183e-14, 1.292129e-14, 
    1.315004e-14, 1.285302e-14, 1.240486e-14, 1.245011e-14, 1.197898e-14, 
    1.191199e-14, 1.242702e-14, 1.264219e-14, 1.259228e-14, 1.293588e-14, 
    1.299867e-14, 1.360559e-14, 1.398021e-14, 1.422277e-14, 1.401917e-14, 
    1.419901e-14, 1.361068e-14, 1.333899e-14, 1.3662e-14,
  2.129468e-14, 2.185948e-14, 2.221619e-14, 2.257965e-14, 2.207272e-14, 
    2.190313e-14, 2.138597e-14, 2.180789e-14, 2.086355e-14, 2.019348e-14, 
    1.924083e-14, 1.798086e-14, 1.743315e-14, 1.754013e-14, 1.661234e-14, 
    1.640505e-14, 1.686531e-14, 1.684004e-14, 1.685929e-14, 1.754233e-14, 
    1.827877e-14, 1.855887e-14, 1.944795e-14, 1.986671e-14, 2.082404e-14, 
    2.162473e-14, 2.100023e-14, 2.188979e-14, 2.128882e-14,
  1.76382e-14, 1.674054e-14, 1.644602e-14, 1.660411e-14, 1.662991e-14, 
    1.764274e-14, 1.849025e-14, 1.832708e-14, 1.818013e-14, 1.769443e-14, 
    1.80852e-14, 1.758563e-14, 1.722739e-14, 1.747605e-14, 1.733917e-14, 
    1.684077e-14, 1.687277e-14, 1.670151e-14, 1.610361e-14, 1.608195e-14, 
    1.571928e-14, 1.555068e-14, 1.552753e-14, 1.661533e-14, 1.675003e-14, 
    1.65858e-14, 1.666192e-14, 1.647673e-14, 1.703754e-14,
  1.237115e-14, 1.22171e-14, 1.251531e-14, 1.21515e-14, 1.181016e-14, 
    1.17265e-14, 1.241713e-14, 1.273398e-14, 1.292524e-14, 1.255278e-14, 
    1.256102e-14, 1.246293e-14, 1.217752e-14, 1.225417e-14, 1.195467e-14, 
    1.130411e-14, 1.124843e-14, 1.119773e-14, 1.163212e-14, 1.199561e-14, 
    1.221443e-14, 1.217003e-14, 1.237315e-14, 1.280829e-14, 1.30009e-14, 
    1.316168e-14, 1.328011e-14, 1.311871e-14, 1.262733e-14,
  8.97803e-15, 8.917146e-15, 8.843161e-15, 8.793988e-15, 8.377156e-15, 
    8.050301e-15, 8.249594e-15, 7.939777e-15, 7.989411e-15, 8.060067e-15, 
    8.221092e-15, 7.891758e-15, 7.718391e-15, 7.681175e-15, 7.439659e-15, 
    7.574494e-15, 7.52166e-15, 7.329897e-15, 7.749687e-15, 7.727884e-15, 
    8.272223e-15, 8.603978e-15, 8.636541e-15, 8.807171e-15, 9.491552e-15, 
    9.31408e-15, 9.403438e-15, 9.592716e-15, 9.570406e-15,
  3.921993e-15, 3.943407e-15, 3.770898e-15, 3.701434e-15, 3.63796e-15, 
    3.70763e-15, 3.626248e-15, 3.48298e-15, 3.429476e-15, 3.580706e-15, 
    3.467716e-15, 3.287576e-15, 3.275576e-15, 3.401647e-15, 3.326874e-15, 
    3.484325e-15, 3.585982e-15, 3.651067e-15, 3.690516e-15, 3.725396e-15, 
    3.672535e-15, 3.881795e-15, 4.076403e-15, 4.150626e-15, 4.115737e-15, 
    4.156627e-15, 4.292682e-15, 4.063166e-15, 3.82945e-15,
  1.780318e-15, 1.842363e-15, 1.800419e-15, 1.829599e-15, 1.940817e-15, 
    1.939495e-15, 1.670934e-15, 1.55755e-15, 1.600762e-15, 1.542903e-15, 
    1.508376e-15, 1.453336e-15, 1.495482e-15, 1.522508e-15, 1.534817e-15, 
    1.624358e-15, 1.723811e-15, 1.67699e-15, 1.781297e-15, 1.635055e-15, 
    1.596835e-15, 1.477355e-15, 1.446778e-15, 1.544993e-15, 1.594689e-15, 
    1.621576e-15, 1.692826e-15, 1.740468e-15, 1.792613e-15,
  4.230788e-16, 4.358757e-16, 4.848929e-16, 5.153959e-16, 5.367594e-16, 
    5.87857e-16, 6.045089e-16, 6.166868e-16, 6.797091e-16, 6.790078e-16, 
    6.841207e-16, 6.530187e-16, 5.355358e-16, 5.202584e-16, 6.025331e-16, 
    6.156205e-16, 5.211555e-16, 4.873871e-16, 4.733827e-16, 4.922443e-16, 
    4.740726e-16, 4.932253e-16, 4.921419e-16, 5.129393e-16, 5.925503e-16, 
    6.014168e-16, 5.701033e-16, 5.136099e-16, 4.335843e-16,
  6.233884e-17, 7.444784e-17, 1.107426e-16, 1.353565e-16, 1.5621e-16, 
    2.362328e-16, 2.8366e-16, 2.947363e-16, 3.877034e-16, 4.208549e-16, 
    4.696255e-16, 4.896088e-16, 4.981409e-16, 5.043508e-16, 6.344493e-16, 
    6.241831e-16, 4.897128e-16, 3.922038e-16, 3.514014e-16, 2.480977e-16, 
    1.670121e-16, 1.311284e-16, 1.104503e-16, 7.500186e-17, 6.189196e-17, 
    6.41405e-17, 6.026111e-17, 6.550658e-17, 6.29058e-17,
  1.9038e-17, 2.638468e-17, 3.562998e-17, 4.975071e-17, 5.400541e-17, 
    6.80163e-17, 1.203462e-16, 1.616902e-16, 2.130365e-16, 2.652638e-16, 
    3.053332e-16, 3.424053e-16, 3.70072e-16, 3.825827e-16, 3.556054e-16, 
    3.306439e-16, 2.681593e-16, 2.521858e-16, 2.218105e-16, 1.926078e-16, 
    1.454861e-16, 1.163713e-16, 8.3733e-17, 4.33417e-17, 2.058229e-17, 
    1.492894e-17, 1.469294e-17, 1.543611e-17, 1.729803e-17,
  1.247012e-17, 1.682794e-17, 2.103061e-17, 2.292878e-17, 3.366398e-17, 
    4.620122e-17, 5.881645e-17, 8.081619e-17, 1.0732e-16, 1.346291e-16, 
    1.630661e-16, 1.749871e-16, 1.746523e-16, 1.69323e-16, 1.688682e-16, 
    1.641198e-16, 1.545916e-16, 1.385483e-16, 1.290342e-16, 1.166202e-16, 
    9.141332e-17, 6.278135e-17, 3.771707e-17, 2.310913e-17, 1.565975e-17, 
    1.163939e-17, 1.06648e-17, 1.031329e-17, 1.121224e-17,
  8.734008e-18, 8.734008e-18, 8.734008e-18, 8.734008e-18, 8.734008e-18, 
    8.734008e-18, 8.734008e-18, 8.250269e-18, 8.250269e-18, 8.250269e-18, 
    8.250269e-18, 8.250269e-18, 8.250269e-18, 8.250269e-18, 8.22487e-18, 
    8.22487e-18, 8.22487e-18, 8.22487e-18, 8.22487e-18, 8.22487e-18, 
    8.22487e-18, 8.65387e-18, 8.65387e-18, 8.65387e-18, 8.65387e-18, 
    8.65387e-18, 8.65387e-18, 8.65387e-18, 8.734008e-18,
  1.119383e-17, 1.005254e-17, 9.411438e-18, 9.245921e-18, 1.047868e-17, 
    1.305847e-17, 1.658797e-17, 1.892337e-17, 1.975829e-17, 1.969681e-17, 
    2.055594e-17, 1.840774e-17, 1.655163e-17, 1.452181e-17, 1.252356e-17, 
    1.168296e-17, 1.09159e-17, 1.004748e-17, 8.920244e-18, 8.277925e-18, 
    8.170921e-18, 8.110512e-18, 7.936524e-18, 9.433032e-18, 1.224387e-17, 
    1.291073e-17, 1.391962e-17, 1.381488e-17, 1.192452e-17,
  2.856497e-17, 4.527798e-17, 6.597526e-17, 1.093188e-16, 1.283164e-16, 
    1.404663e-16, 1.649964e-16, 1.854763e-16, 2.157414e-16, 2.087947e-16, 
    1.906992e-16, 1.687473e-16, 1.509245e-16, 1.360257e-16, 1.158327e-16, 
    1.122467e-16, 1.033982e-16, 6.886713e-17, 4.562074e-17, 2.764423e-17, 
    1.814145e-17, 1.672822e-17, 1.692721e-17, 2.282593e-17, 2.379854e-17, 
    2.775454e-17, 1.95375e-17, 1.73826e-17, 2.242318e-17,
  7.737218e-16, 9.209727e-16, 1.071927e-15, 1.302871e-15, 1.363315e-15, 
    1.37891e-15, 1.115547e-15, 8.08939e-16, 6.408109e-16, 5.681712e-16, 
    5.643951e-16, 6.550691e-16, 7.237847e-16, 7.417094e-16, 7.30375e-16, 
    7.122059e-16, 6.981414e-16, 7.094619e-16, 6.559506e-16, 5.915397e-16, 
    4.906288e-16, 3.064221e-16, 1.24436e-16, 8.953251e-17, 1.178198e-16, 
    1.654809e-16, 2.744906e-16, 3.743677e-16, 5.565663e-16,
  2.098232e-15, 2.198887e-15, 2.045122e-15, 1.326976e-15, 9.229739e-16, 
    8.202211e-16, 7.839056e-16, 8.471539e-16, 9.050489e-16, 9.44229e-16, 
    9.566744e-16, 9.660999e-16, 1.04577e-15, 1.113275e-15, 1.210971e-15, 
    1.145129e-15, 9.719991e-16, 9.027104e-16, 8.153484e-16, 7.400914e-16, 
    7.642448e-16, 9.508264e-16, 1.278511e-15, 1.345106e-15, 1.379161e-15, 
    1.563698e-15, 1.965718e-15, 2.334483e-15, 2.215802e-15,
  5.042064e-15, 4.344051e-15, 4.198157e-15, 4.040984e-15, 3.923949e-15, 
    3.68892e-15, 3.370668e-15, 3.495905e-15, 3.204308e-15, 2.771418e-15, 
    2.763652e-15, 2.752225e-15, 2.830799e-15, 3.052015e-15, 3.25077e-15, 
    3.325436e-15, 3.838365e-15, 4.46421e-15, 4.752401e-15, 5.245086e-15, 
    5.105344e-15, 5.83978e-15, 6.918e-15, 7.011631e-15, 6.273204e-15, 
    6.386594e-15, 5.533119e-15, 5.768776e-15, 5.202888e-15,
  1.682685e-14, 1.679181e-14, 1.679105e-14, 1.668354e-14, 1.626752e-14, 
    1.695766e-14, 1.683469e-14, 1.705952e-14, 1.709874e-14, 1.704233e-14, 
    1.583377e-14, 1.43291e-14, 1.483236e-14, 1.537243e-14, 1.502546e-14, 
    1.474341e-14, 1.524864e-14, 1.545926e-14, 1.607424e-14, 1.688134e-14, 
    1.728477e-14, 1.775016e-14, 1.831707e-14, 1.808967e-14, 1.788216e-14, 
    1.807024e-14, 1.806487e-14, 1.803172e-14, 1.747972e-14,
  4.850397e-14, 4.818309e-14, 4.749734e-14, 4.644341e-14, 4.76165e-14, 
    4.900307e-14, 4.82321e-14, 4.819645e-14, 4.749466e-14, 4.676038e-14, 
    4.539845e-14, 4.579097e-14, 4.547896e-14, 4.629029e-14, 4.71811e-14, 
    4.6721e-14, 4.618322e-14, 4.711497e-14, 4.877046e-14, 4.955947e-14, 
    5.158354e-14, 5.038568e-14, 5.249728e-14, 5.039683e-14, 5.096279e-14, 
    5.250879e-14, 5.130221e-14, 4.869142e-14, 4.743019e-14,
  7.386699e-14, 7.254275e-14, 7.564462e-14, 7.505777e-14, 7.723189e-14, 
    7.584327e-14, 7.583468e-14, 7.405479e-14, 7.466562e-14, 7.251698e-14, 
    7.058378e-14, 6.698255e-14, 6.308814e-14, 6.137488e-14, 5.944447e-14, 
    5.747524e-14, 5.807041e-14, 6.004083e-14, 6.030217e-14, 6.058386e-14, 
    5.948095e-14, 6.284922e-14, 6.531407e-14, 6.923634e-14, 6.848991e-14, 
    6.986729e-14, 7.211077e-14, 7.061701e-14, 7.27751e-14,
  5.257896e-14, 5.207723e-14, 5.132365e-14, 5.023228e-14, 5.097395e-14, 
    5.482493e-14, 5.662549e-14, 5.823876e-14, 5.766098e-14, 5.685269e-14, 
    5.913401e-14, 6.008174e-14, 6.11861e-14, 6.181786e-14, 6.104181e-14, 
    6.014978e-14, 5.912386e-14, 5.791598e-14, 5.748413e-14, 5.80489e-14, 
    5.656262e-14, 5.557152e-14, 5.668552e-14, 5.510302e-14, 5.196878e-14, 
    5.065716e-14, 5.071367e-14, 5.043525e-14, 5.082344e-14,
  4.394523e-14, 4.269025e-14, 4.265168e-14, 4.21068e-14, 4.204716e-14, 
    4.178435e-14, 4.410982e-14, 4.399076e-14, 4.376303e-14, 4.518524e-14, 
    4.658211e-14, 4.895846e-14, 4.793418e-14, 4.617921e-14, 4.573507e-14, 
    4.479953e-14, 4.356755e-14, 4.24399e-14, 4.287035e-14, 4.392602e-14, 
    4.370831e-14, 4.571709e-14, 4.740103e-14, 4.791437e-14, 4.68065e-14, 
    4.612603e-14, 4.723888e-14, 4.832394e-14, 4.65737e-14,
  3.796344e-14, 3.627628e-14, 3.540498e-14, 3.573298e-14, 3.544143e-14, 
    3.147618e-14, 3.150742e-14, 3.164812e-14, 3.187509e-14, 3.274039e-14, 
    3.183678e-14, 3.116144e-14, 3.14674e-14, 3.237815e-14, 3.022648e-14, 
    3.037549e-14, 2.934241e-14, 2.960312e-14, 3.103745e-14, 3.272574e-14, 
    3.262276e-14, 3.473678e-14, 3.561084e-14, 3.640776e-14, 3.775416e-14, 
    3.842071e-14, 3.922349e-14, 3.962299e-14, 3.839895e-14,
  1.53411e-14, 1.478194e-14, 1.499577e-14, 1.438672e-14, 1.410144e-14, 
    1.417851e-14, 1.411963e-14, 1.407129e-14, 1.39108e-14, 1.341646e-14, 
    1.278616e-14, 1.217721e-14, 1.245941e-14, 1.28095e-14, 1.304314e-14, 
    1.355744e-14, 1.414653e-14, 1.420515e-14, 1.446727e-14, 1.465103e-14, 
    1.480616e-14, 1.555184e-14, 1.680629e-14, 1.734467e-14, 1.766465e-14, 
    1.67425e-14, 1.640182e-14, 1.65543e-14, 1.556056e-14,
  7.089507e-15, 6.880067e-15, 6.302237e-15, 6.227132e-15, 6.04336e-15, 
    7.079252e-15, 7.071129e-15, 6.609357e-15, 5.328219e-15, 5.010725e-15, 
    5.00662e-15, 4.924362e-15, 5.270915e-15, 5.345741e-15, 5.457847e-15, 
    5.691454e-15, 6.141444e-15, 6.768329e-15, 6.251485e-15, 5.541569e-15, 
    5.120681e-15, 4.945681e-15, 5.266015e-15, 5.742211e-15, 6.053613e-15, 
    6.384102e-15, 6.510586e-15, 6.690532e-15, 7.33423e-15,
  8.403623e-16, 1.098398e-15, 1.359041e-15, 1.53147e-15, 1.756623e-15, 
    2.276375e-15, 2.766867e-15, 3.736069e-15, 3.938854e-15, 3.272766e-15, 
    3.156261e-15, 2.40376e-15, 1.846136e-15, 1.838424e-15, 2.216504e-15, 
    2.334814e-15, 1.78496e-15, 1.743638e-15, 1.780692e-15, 1.593913e-15, 
    1.326729e-15, 1.408547e-15, 1.417402e-15, 1.440721e-15, 1.59608e-15, 
    1.656104e-15, 1.550204e-15, 1.363288e-15, 1.005385e-15,
  1.848409e-16, 1.896889e-16, 2.712818e-16, 3.922719e-16, 4.773319e-16, 
    8.019902e-16, 1.143038e-15, 1.525826e-15, 1.63246e-15, 1.944391e-15, 
    2.425794e-15, 1.817547e-15, 1.666687e-15, 1.744048e-15, 2.300383e-15, 
    2.593002e-15, 2.439028e-15, 1.901924e-15, 1.578006e-15, 1.037315e-15, 
    8.612184e-16, 6.655044e-16, 6.621294e-16, 3.93483e-16, 2.079368e-16, 
    2.176117e-16, 1.927566e-16, 1.957126e-16, 1.965366e-16,
  5.189758e-17, 6.355377e-17, 8.815971e-17, 1.368304e-16, 1.536789e-16, 
    2.133759e-16, 3.838895e-16, 5.569987e-16, 8.987844e-16, 1.034229e-15, 
    1.243522e-15, 1.306538e-15, 1.440504e-15, 1.56792e-15, 1.583097e-15, 
    1.50662e-15, 1.136293e-15, 1.065655e-15, 9.43052e-16, 7.620213e-16, 
    8.426439e-16, 6.125081e-16, 3.798651e-16, 1.682224e-16, 6.357598e-17, 
    4.7287e-17, 4.595894e-17, 4.834403e-17, 5.268101e-17,
  2.76101e-17, 3.359918e-17, 4.084161e-17, 4.74853e-17, 8.344562e-17, 
    1.274191e-16, 1.977003e-16, 2.555351e-16, 3.43895e-16, 4.420307e-16, 
    5.803625e-16, 7.139062e-16, 7.642394e-16, 7.527896e-16, 7.514149e-16, 
    7.547122e-16, 7.434948e-16, 7.08042e-16, 6.740755e-16, 5.568949e-16, 
    4.172605e-16, 2.578331e-16, 1.319031e-16, 7.635234e-17, 4.661692e-17, 
    2.94983e-17, 2.645436e-17, 2.62431e-17, 2.6386e-17,
  2.687149e-17, 2.687149e-17, 2.687149e-17, 2.687149e-17, 2.687149e-17, 
    2.687149e-17, 2.687149e-17, 2.611712e-17, 2.611712e-17, 2.611712e-17, 
    2.611712e-17, 2.611712e-17, 2.611712e-17, 2.611712e-17, 2.413034e-17, 
    2.413034e-17, 2.413034e-17, 2.413034e-17, 2.413034e-17, 2.413034e-17, 
    2.413034e-17, 2.515423e-17, 2.515423e-17, 2.515423e-17, 2.515423e-17, 
    2.515423e-17, 2.515423e-17, 2.515423e-17, 2.687149e-17,
  5.017255e-17, 3.859873e-17, 3.409963e-17, 3.312649e-17, 3.567575e-17, 
    4.41543e-17, 6.068893e-17, 7.018471e-17, 6.955474e-17, 7.018625e-17, 
    7.619723e-17, 6.870437e-17, 6.354007e-17, 5.786471e-17, 4.790173e-17, 
    4.190792e-17, 3.914115e-17, 3.535817e-17, 3.201101e-17, 2.961831e-17, 
    2.666259e-17, 2.547436e-17, 2.576304e-17, 2.815803e-17, 3.682958e-17, 
    4.901115e-17, 5.829244e-17, 6.077426e-17, 5.568069e-17,
  8.800179e-17, 1.320592e-16, 1.765664e-16, 2.777932e-16, 3.087972e-16, 
    3.433749e-16, 3.859038e-16, 4.442549e-16, 4.972769e-16, 5.055924e-16, 
    4.843085e-16, 4.861941e-16, 4.737244e-16, 4.396924e-16, 4.063529e-16, 
    3.884819e-16, 4.019508e-16, 3.303117e-16, 1.914854e-16, 1.226366e-16, 
    8.787614e-17, 8.389844e-17, 7.607824e-17, 8.894539e-17, 1.066372e-16, 
    1.3439e-16, 9.362519e-17, 6.81256e-17, 6.679837e-17,
  1.484252e-15, 2.008759e-15, 2.217674e-15, 2.885049e-15, 3.095663e-15, 
    2.855084e-15, 2.428918e-15, 1.872598e-15, 1.505978e-15, 1.409212e-15, 
    1.444866e-15, 1.528458e-15, 1.608629e-15, 1.745386e-15, 1.823623e-15, 
    1.758921e-15, 1.62353e-15, 1.745972e-15, 1.867036e-15, 1.673797e-15, 
    1.324206e-15, 1.103804e-15, 4.864054e-16, 3.220907e-16, 4.003392e-16, 
    4.864004e-16, 6.423419e-16, 8.13704e-16, 1.113501e-15,
  5.090076e-15, 5.350379e-15, 4.680086e-15, 3.568623e-15, 2.92282e-15, 
    2.416518e-15, 2.167201e-15, 2.315833e-15, 2.394786e-15, 2.419362e-15, 
    2.397075e-15, 2.563824e-15, 2.827918e-15, 2.935704e-15, 3.333856e-15, 
    3.47412e-15, 3.281385e-15, 2.356225e-15, 1.958678e-15, 1.921842e-15, 
    1.796456e-15, 2.477648e-15, 3.400355e-15, 3.755005e-15, 3.203418e-15, 
    3.817429e-15, 4.766539e-15, 5.328569e-15, 4.874336e-15,
  9.475428e-15, 7.947951e-15, 7.377373e-15, 7.728377e-15, 8.101716e-15, 
    9.005032e-15, 8.556684e-15, 7.546062e-15, 6.676439e-15, 5.693852e-15, 
    5.31498e-15, 5.685647e-15, 6.161172e-15, 6.465603e-15, 6.50081e-15, 
    8.305437e-15, 9.985193e-15, 1.285945e-14, 1.441445e-14, 1.41697e-14, 
    1.461207e-14, 1.627435e-14, 1.887373e-14, 2.011325e-14, 1.634365e-14, 
    1.271054e-14, 1.058902e-14, 1.102712e-14, 1.035596e-14,
  5.081729e-14, 5.047598e-14, 4.639122e-14, 4.344996e-14, 4.197128e-14, 
    4.401689e-14, 4.641965e-14, 4.864645e-14, 5.415336e-14, 5.320037e-14, 
    5.211281e-14, 5.066484e-14, 5.040904e-14, 4.968439e-14, 4.842795e-14, 
    4.887862e-14, 4.806128e-14, 4.910995e-14, 4.890803e-14, 4.948845e-14, 
    5.296328e-14, 5.59058e-14, 5.656356e-14, 5.630107e-14, 5.476711e-14, 
    5.592133e-14, 5.603403e-14, 5.463951e-14, 5.216075e-14,
  1.799018e-13, 1.751258e-13, 1.761932e-13, 1.843758e-13, 1.84459e-13, 
    1.877795e-13, 1.835436e-13, 1.78339e-13, 1.811025e-13, 1.758112e-13, 
    1.749309e-13, 1.71334e-13, 1.696361e-13, 1.692202e-13, 1.705744e-13, 
    1.704524e-13, 1.741999e-13, 1.71321e-13, 1.786812e-13, 1.828673e-13, 
    1.899184e-13, 1.943562e-13, 1.970249e-13, 1.882836e-13, 1.889993e-13, 
    1.839395e-13, 1.83003e-13, 1.791939e-13, 1.745906e-13,
  2.478901e-13, 2.580736e-13, 2.54664e-13, 2.655779e-13, 2.612529e-13, 
    2.666026e-13, 2.695276e-13, 2.635146e-13, 2.631801e-13, 2.573969e-13, 
    2.5405e-13, 2.447145e-13, 2.322613e-13, 2.302243e-13, 2.250292e-13, 
    2.180078e-13, 2.107472e-13, 2.131977e-13, 2.236398e-13, 2.17066e-13, 
    2.242614e-13, 2.224752e-13, 2.377455e-13, 2.44768e-13, 2.430428e-13, 
    2.356711e-13, 2.339709e-13, 2.467133e-13, 2.416124e-13,
  1.750319e-13, 1.72849e-13, 1.714738e-13, 1.71427e-13, 1.664134e-13, 
    1.752092e-13, 1.829167e-13, 1.886622e-13, 1.86689e-13, 1.906077e-13, 
    1.930516e-13, 1.987161e-13, 2.074215e-13, 2.024745e-13, 2.027176e-13, 
    1.99904e-13, 1.957773e-13, 1.930866e-13, 1.931296e-13, 1.970001e-13, 
    1.977758e-13, 1.900722e-13, 1.874721e-13, 1.847602e-13, 1.819483e-13, 
    1.796344e-13, 1.734568e-13, 1.759591e-13, 1.763728e-13,
  1.696469e-13, 1.651874e-13, 1.657175e-13, 1.615574e-13, 1.676515e-13, 
    1.689789e-13, 1.703573e-13, 1.773609e-13, 1.736033e-13, 1.817526e-13, 
    1.873471e-13, 1.937405e-13, 1.893371e-13, 1.954105e-13, 1.880888e-13, 
    1.912646e-13, 1.826002e-13, 1.7684e-13, 1.788453e-13, 1.850088e-13, 
    1.922453e-13, 1.946933e-13, 1.911287e-13, 1.900505e-13, 1.881947e-13, 
    1.853298e-13, 1.876589e-13, 1.813415e-13, 1.757007e-13,
  1.505674e-13, 1.498298e-13, 1.508776e-13, 1.480709e-13, 1.431402e-13, 
    1.340817e-13, 1.286993e-13, 1.293693e-13, 1.386338e-13, 1.348408e-13, 
    1.362427e-13, 1.364283e-13, 1.332791e-13, 1.347899e-13, 1.346651e-13, 
    1.320565e-13, 1.286296e-13, 1.277137e-13, 1.320083e-13, 1.433558e-13, 
    1.610342e-13, 1.619993e-13, 1.621914e-13, 1.603385e-13, 1.604645e-13, 
    1.653965e-13, 1.701728e-13, 1.678377e-13, 1.59637e-13,
  6.682358e-14, 6.555709e-14, 6.187284e-14, 6.17591e-14, 6.201143e-14, 
    6.086854e-14, 5.673462e-14, 5.958079e-14, 5.404509e-14, 4.711778e-14, 
    4.693842e-14, 4.401822e-14, 4.343305e-14, 4.416607e-14, 4.692669e-14, 
    4.746289e-14, 4.89764e-14, 4.935189e-14, 5.570504e-14, 5.621872e-14, 
    6.322807e-14, 6.948601e-14, 7.577603e-14, 8.487226e-14, 8.193961e-14, 
    8.078586e-14, 7.638334e-14, 7.194645e-14, 6.967549e-14,
  2.93408e-14, 2.640468e-14, 2.205499e-14, 2.007191e-14, 2.097814e-14, 
    2.387727e-14, 2.673851e-14, 2.197151e-14, 1.647125e-14, 1.389968e-14, 
    1.456369e-14, 1.471772e-14, 1.583888e-14, 1.661856e-14, 1.681401e-14, 
    1.815116e-14, 1.847791e-14, 2.063707e-14, 1.897008e-14, 1.641118e-14, 
    1.537096e-14, 1.521893e-14, 1.629776e-14, 2.101098e-14, 2.599149e-14, 
    2.775643e-14, 2.695131e-14, 2.963219e-14, 3.262969e-14,
  2.94944e-15, 3.038688e-15, 3.995147e-15, 5.00636e-15, 6.359135e-15, 
    9.954069e-15, 1.383079e-14, 1.795585e-14, 1.844955e-14, 1.919721e-14, 
    1.453392e-14, 8.063401e-15, 6.487712e-15, 6.453888e-15, 7.292774e-15, 
    8.189375e-15, 6.938516e-15, 5.901228e-15, 6.066177e-15, 5.213456e-15, 
    3.811584e-15, 4.129742e-15, 3.877522e-15, 4.473366e-15, 3.449284e-15, 
    3.700266e-15, 5.723887e-15, 6.44466e-15, 4.603309e-15,
  5.41085e-16, 5.668676e-16, 8.479871e-16, 1.134389e-15, 1.782731e-15, 
    3.067204e-15, 5.65433e-15, 8.427393e-15, 9.491781e-15, 9.54484e-15, 
    8.073339e-15, 6.976666e-15, 6.780152e-15, 6.692877e-15, 7.18689e-15, 
    9.021799e-15, 8.911403e-15, 7.161373e-15, 5.689253e-15, 4.276502e-15, 
    3.970311e-15, 4.412729e-15, 3.601714e-15, 2.076729e-15, 9.026948e-16, 
    7.649561e-16, 6.35036e-16, 5.81842e-16, 5.718458e-16,
  1.730182e-16, 1.772975e-16, 2.220296e-16, 4.623206e-16, 5.172082e-16, 
    6.899495e-16, 1.350613e-15, 2.290332e-15, 3.48275e-15, 4.243105e-15, 
    4.448743e-15, 4.790698e-15, 5.360811e-15, 5.944451e-15, 6.391494e-15, 
    6.358319e-15, 5.14554e-15, 4.111077e-15, 3.403477e-15, 2.994206e-15, 
    3.652704e-15, 2.580503e-15, 1.844188e-15, 7.428763e-16, 2.017391e-16, 
    1.481493e-16, 1.424124e-16, 1.593154e-16, 1.914529e-16,
  8.907942e-17, 8.659936e-17, 9.690875e-17, 1.072808e-16, 2.176455e-16, 
    3.951072e-16, 5.916936e-16, 9.015333e-16, 1.485889e-15, 1.886938e-15, 
    2.317796e-15, 2.759971e-15, 3.048223e-15, 3.167589e-15, 3.309998e-15, 
    3.411878e-15, 3.472614e-15, 3.313405e-15, 3.006253e-15, 2.557117e-15, 
    1.883767e-15, 1.086777e-15, 6.105597e-16, 3.123846e-16, 1.643958e-16, 
    1.065265e-16, 1.000935e-16, 9.111465e-17, 9.147206e-17,
  7.383607e-17, 7.383607e-17, 7.383607e-17, 7.383607e-17, 7.383607e-17, 
    7.383607e-17, 7.383607e-17, 7.588738e-17, 7.588738e-17, 7.588738e-17, 
    7.588738e-17, 7.588738e-17, 7.588738e-17, 7.588738e-17, 7.320513e-17, 
    7.320513e-17, 7.320513e-17, 7.320513e-17, 7.320513e-17, 7.320513e-17, 
    7.320513e-17, 6.84138e-17, 6.84138e-17, 6.84138e-17, 6.84138e-17, 
    6.84138e-17, 6.84138e-17, 6.84138e-17, 7.383607e-17,
  2.501018e-16, 2.084324e-16, 1.742525e-16, 1.653075e-16, 1.725104e-16, 
    1.978337e-16, 2.146019e-16, 2.245512e-16, 2.217141e-16, 2.221126e-16, 
    2.319225e-16, 2.267844e-16, 2.308233e-16, 2.256854e-16, 1.950475e-16, 
    1.560523e-16, 1.367978e-16, 1.213721e-16, 1.050361e-16, 9.35256e-17, 
    8.164929e-17, 7.795302e-17, 8.14553e-17, 9.102194e-17, 1.018102e-16, 
    1.307054e-16, 1.747072e-16, 2.213811e-16, 2.573774e-16,
  2.989761e-16, 3.754976e-16, 4.792797e-16, 6.997171e-16, 8.274742e-16, 
    9.196405e-16, 9.500156e-16, 1.11873e-15, 1.344384e-15, 1.583092e-15, 
    1.553418e-15, 1.554637e-15, 1.370396e-15, 1.175779e-15, 1.116407e-15, 
    1.06094e-15, 1.033825e-15, 1.013289e-15, 7.237808e-16, 4.814708e-16, 
    3.824437e-16, 3.677953e-16, 3.174682e-16, 2.980608e-16, 4.16357e-16, 
    5.698923e-16, 4.931235e-16, 3.373518e-16, 3.046025e-16,
  3.987051e-15, 4.70506e-15, 4.853659e-15, 6.355605e-15, 6.675467e-15, 
    6.479253e-15, 5.980998e-15, 5.036464e-15, 3.909302e-15, 3.645242e-15, 
    3.929351e-15, 4.176608e-15, 4.594842e-15, 5.236908e-15, 5.678652e-15, 
    5.688317e-15, 5.353632e-15, 5.741407e-15, 7.028841e-15, 6.557136e-15, 
    4.561486e-15, 4.133197e-15, 2.182665e-15, 1.327928e-15, 1.427881e-15, 
    1.555667e-15, 1.704394e-15, 2.348289e-15, 3.231079e-15,
  1.236263e-14, 1.316262e-14, 1.149634e-14, 9.910228e-15, 8.699222e-15, 
    7.897612e-15, 6.776211e-15, 6.941289e-15, 6.903229e-15, 7.024486e-15, 
    7.707685e-15, 7.557875e-15, 8.331998e-15, 8.036516e-15, 9.232748e-15, 
    1.036489e-14, 1.026112e-14, 8.996301e-15, 7.00691e-15, 6.300115e-15, 
    6.742285e-15, 8.20348e-15, 7.95615e-15, 1.114219e-14, 9.308955e-15, 
    9.815479e-15, 1.064419e-14, 1.330644e-14, 1.247014e-14,
  2.577429e-14, 2.360577e-14, 2.098753e-14, 2.077284e-14, 1.973599e-14, 
    1.860701e-14, 2.294709e-14, 2.430131e-14, 2.044948e-14, 1.464956e-14, 
    1.234217e-14, 1.321995e-14, 1.363705e-14, 1.475548e-14, 1.383561e-14, 
    1.728637e-14, 2.069125e-14, 2.782386e-14, 3.932619e-14, 4.503695e-14, 
    4.971471e-14, 5.908124e-14, 6.299431e-14, 6.212372e-14, 5.307132e-14, 
    3.336949e-14, 2.793529e-14, 2.748666e-14, 2.683623e-14,
  1.477839e-13, 1.40324e-13, 1.371374e-13, 1.305816e-13, 1.363143e-13, 
    1.456641e-13, 1.585518e-13, 1.703306e-13, 1.68994e-13, 1.613662e-13, 
    1.568917e-13, 1.630667e-13, 1.627073e-13, 1.677581e-13, 1.678414e-13, 
    1.700282e-13, 1.782778e-13, 1.782997e-13, 1.789479e-13, 1.747848e-13, 
    1.913735e-13, 2.053036e-13, 1.957415e-13, 1.893126e-13, 1.839767e-13, 
    1.917227e-13, 1.736811e-13, 1.616812e-13, 1.519997e-13,
  6.65189e-13, 6.779523e-13, 6.890926e-13, 6.931121e-13, 6.944526e-13, 
    6.981915e-13, 6.939184e-13, 6.937533e-13, 7.016659e-13, 6.894226e-13, 
    6.714123e-13, 6.722708e-13, 6.527589e-13, 6.380022e-13, 6.456941e-13, 
    6.380116e-13, 6.437251e-13, 6.413891e-13, 6.690147e-13, 6.425792e-13, 
    6.724876e-13, 6.936525e-13, 6.878185e-13, 6.69987e-13, 6.539e-13, 
    6.625476e-13, 6.606087e-13, 6.586262e-13, 6.403109e-13,
  8.858567e-13, 9.244739e-13, 9.195089e-13, 9.353859e-13, 9.331222e-13, 
    9.318496e-13, 9.602513e-13, 9.84035e-13, 9.624169e-13, 9.331867e-13, 
    9.292964e-13, 9.061267e-13, 8.650404e-13, 8.537691e-13, 8.098744e-13, 
    8.227272e-13, 8.26195e-13, 8.150021e-13, 7.744012e-13, 7.787368e-13, 
    7.92843e-13, 8.563473e-13, 8.690981e-13, 8.69689e-13, 8.92751e-13, 
    8.975853e-13, 8.906833e-13, 9.171924e-13, 8.760116e-13,
  6.182424e-13, 6.199256e-13, 6.049398e-13, 6.027721e-13, 5.996894e-13, 
    6.240612e-13, 6.699328e-13, 6.834344e-13, 6.836104e-13, 7.082578e-13, 
    7.327451e-13, 7.446685e-13, 7.543834e-13, 7.517834e-13, 7.53837e-13, 
    7.225401e-13, 7.213557e-13, 7.114825e-13, 6.942197e-13, 6.999623e-13, 
    6.990895e-13, 6.844892e-13, 6.636687e-13, 6.423285e-13, 6.244333e-13, 
    6.117294e-13, 6.130742e-13, 5.995661e-13, 6.022365e-13,
  6.666926e-13, 6.866185e-13, 6.812681e-13, 6.78805e-13, 7.055355e-13, 
    6.853242e-13, 7.119106e-13, 7.124591e-13, 7.508633e-13, 7.722928e-13, 
    7.738644e-13, 7.971828e-13, 7.990468e-13, 7.798108e-13, 7.50265e-13, 
    7.378802e-13, 7.3577e-13, 7.323706e-13, 7.361384e-13, 7.832737e-13, 
    8.218035e-13, 8.052287e-13, 7.72088e-13, 7.547782e-13, 7.251725e-13, 
    7.264957e-13, 7.039448e-13, 6.652089e-13, 6.518792e-13,
  6.329076e-13, 6.479046e-13, 6.469948e-13, 6.285452e-13, 5.772873e-13, 
    5.796839e-13, 5.714863e-13, 6.121781e-13, 6.124267e-13, 5.717539e-13, 
    6.082341e-13, 6.211536e-13, 6.476057e-13, 6.4162e-13, 6.310768e-13, 
    6.122977e-13, 6.502494e-13, 6.96043e-13, 7.201533e-13, 7.017889e-13, 
    7.579999e-13, 7.248407e-13, 7.605533e-13, 7.353385e-13, 7.270535e-13, 
    7.059898e-13, 6.707415e-13, 6.364769e-13, 6.341525e-13,
  2.84468e-13, 2.782025e-13, 2.715471e-13, 2.419778e-13, 2.412963e-13, 
    2.389097e-13, 2.10148e-13, 2.274909e-13, 1.934148e-13, 1.646083e-13, 
    1.596907e-13, 1.623476e-13, 1.564161e-13, 1.688229e-13, 2.241577e-13, 
    2.05332e-13, 1.977972e-13, 1.974717e-13, 2.058135e-13, 2.483321e-13, 
    3.055664e-13, 3.457465e-13, 3.778221e-13, 3.822665e-13, 3.602815e-13, 
    3.57464e-13, 3.474317e-13, 3.224941e-13, 2.899746e-13,
  1.227025e-13, 1.083914e-13, 8.19397e-14, 7.260069e-14, 7.267576e-14, 
    8.640472e-14, 9.466298e-14, 7.509645e-14, 4.902842e-14, 4.18289e-14, 
    3.726237e-14, 4.132901e-14, 4.829377e-14, 4.470498e-14, 4.81292e-14, 
    4.775095e-14, 4.329699e-14, 4.593273e-14, 4.808128e-14, 4.464365e-14, 
    4.563986e-14, 5.239794e-14, 5.480632e-14, 1.0118e-13, 1.256601e-13, 
    1.407791e-13, 1.340648e-13, 1.407129e-13, 1.28448e-13,
  1.481996e-14, 1.199516e-14, 1.328604e-14, 1.8852e-14, 2.431976e-14, 
    3.759974e-14, 5.315307e-14, 6.599478e-14, 7.726485e-14, 7.064968e-14, 
    5.980225e-14, 4.235061e-14, 2.449972e-14, 2.036359e-14, 2.060556e-14, 
    2.345336e-14, 2.259152e-14, 1.965311e-14, 1.686608e-14, 1.877845e-14, 
    1.345469e-14, 1.316809e-14, 1.38328e-14, 1.366291e-14, 1.142628e-14, 
    1.669068e-14, 2.440881e-14, 3.001372e-14, 2.465187e-14,
  1.652194e-15, 1.593588e-15, 2.653303e-15, 4.797826e-15, 6.588349e-15, 
    1.14136e-14, 2.630939e-14, 3.923982e-14, 4.221602e-14, 4.225834e-14, 
    3.421603e-14, 2.916304e-14, 2.344394e-14, 2.176691e-14, 2.057343e-14, 
    2.569348e-14, 2.807195e-14, 2.188793e-14, 1.755446e-14, 1.624629e-14, 
    1.362709e-14, 1.64498e-14, 1.43265e-14, 6.81628e-15, 3.974741e-15, 
    2.451514e-15, 1.849074e-15, 1.805791e-15, 1.706181e-15,
  6.109428e-16, 5.782601e-16, 6.139181e-16, 1.575137e-15, 1.892902e-15, 
    2.196269e-15, 4.245322e-15, 8.961428e-15, 1.180176e-14, 1.789784e-14, 
    1.557862e-14, 1.531043e-14, 1.630063e-14, 1.838349e-14, 1.981983e-14, 
    1.956038e-14, 1.675889e-14, 1.339654e-14, 1.168442e-14, 1.162066e-14, 
    1.277312e-14, 9.276003e-15, 6.842952e-15, 3.082389e-15, 6.685897e-16, 
    5.351136e-16, 5.410137e-16, 5.664075e-16, 6.481799e-16,
  2.810055e-16, 2.38113e-16, 2.41286e-16, 2.830034e-16, 5.520364e-16, 
    1.144859e-15, 1.743434e-15, 3.495733e-15, 5.575969e-15, 6.723415e-15, 
    7.710395e-15, 9.306175e-15, 1.133034e-14, 1.211262e-14, 1.218543e-14, 
    1.211167e-14, 1.191106e-14, 1.117387e-14, 1.029541e-14, 9.093033e-15, 
    7.331919e-15, 4.576492e-15, 2.789987e-15, 1.27968e-15, 6.3639e-16, 
    4.490515e-16, 4.070042e-16, 3.517365e-16, 3.04301e-16,
  2.126669e-16, 2.126669e-16, 2.126669e-16, 2.126669e-16, 2.126669e-16, 
    2.126669e-16, 2.126669e-16, 2.243801e-16, 2.243801e-16, 2.243801e-16, 
    2.243801e-16, 2.243801e-16, 2.243801e-16, 2.243801e-16, 2.248969e-16, 
    2.248969e-16, 2.248969e-16, 2.248969e-16, 2.248969e-16, 2.248969e-16, 
    2.248969e-16, 2.111497e-16, 2.111497e-16, 2.111497e-16, 2.111497e-16, 
    2.111497e-16, 2.111497e-16, 2.111497e-16, 2.126669e-16,
  7.605858e-16, 7.466835e-16, 6.729833e-16, 6.358399e-16, 6.134617e-16, 
    6.309512e-16, 6.316342e-16, 6.221874e-16, 5.726888e-16, 5.225819e-16, 
    5.665097e-16, 5.739489e-16, 5.895007e-16, 5.846301e-16, 5.177976e-16, 
    4.420898e-16, 4.110245e-16, 4.004354e-16, 3.52682e-16, 3.193157e-16, 
    3.084224e-16, 2.987024e-16, 2.950234e-16, 2.941826e-16, 2.830987e-16, 
    3.028715e-16, 3.709463e-16, 5.798291e-16, 7.502217e-16,
  1.167597e-15, 1.426215e-15, 1.584836e-15, 1.851936e-15, 1.971143e-15, 
    1.952809e-15, 2.133073e-15, 2.608556e-15, 3.642657e-15, 4.641742e-15, 
    4.748086e-15, 4.589571e-15, 3.751285e-15, 3.283855e-15, 2.938364e-15, 
    2.796482e-15, 2.527908e-15, 2.435171e-15, 1.938723e-15, 1.37792e-15, 
    1.2272e-15, 1.194873e-15, 1.09691e-15, 9.703173e-16, 1.259125e-15, 
    2.091734e-15, 1.933411e-15, 1.246599e-15, 1.048386e-15,
  1.282097e-14, 1.371037e-14, 1.365825e-14, 1.703347e-14, 1.841186e-14, 
    1.852946e-14, 1.645967e-14, 1.413294e-14, 1.140182e-14, 1.00865e-14, 
    9.951981e-15, 1.143394e-14, 1.43483e-14, 1.807749e-14, 2.212762e-14, 
    2.591796e-14, 2.132227e-14, 2.151481e-14, 2.461676e-14, 2.350265e-14, 
    1.677412e-14, 1.440847e-14, 9.313796e-15, 5.196144e-15, 5.851567e-15, 
    5.62052e-15, 5.88956e-15, 8.181204e-15, 1.118074e-14,
  4.345227e-14, 3.95392e-14, 3.59904e-14, 3.068668e-14, 2.717662e-14, 
    2.575617e-14, 2.181836e-14, 2.156757e-14, 2.212783e-14, 2.320754e-14, 
    2.696611e-14, 2.749781e-14, 2.806032e-14, 2.593497e-14, 2.648319e-14, 
    3.041783e-14, 3.266176e-14, 4.661891e-14, 4.078196e-14, 2.658079e-14, 
    2.502848e-14, 3.32477e-14, 2.954999e-14, 3.397118e-14, 3.83359e-14, 
    3.527375e-14, 3.261673e-14, 3.839156e-14, 4.120496e-14,
  7.764124e-14, 7.903087e-14, 7.50917e-14, 7.411136e-14, 6.815122e-14, 
    5.455933e-14, 5.516119e-14, 7.429867e-14, 7.106971e-14, 4.315937e-14, 
    3.646019e-14, 4.062561e-14, 4.509593e-14, 4.643399e-14, 4.940244e-14, 
    4.848523e-14, 5.154604e-14, 6.420252e-14, 8.457049e-14, 1.179868e-13, 
    1.591215e-13, 2.013633e-13, 2.255488e-13, 2.284253e-13, 1.672139e-13, 
    1.119646e-13, 1.024266e-13, 9.299073e-14, 8.658038e-14,
  4.966774e-13, 4.786222e-13, 4.480871e-13, 4.709384e-13, 5.34652e-13, 
    5.284038e-13, 5.630728e-13, 5.623338e-13, 5.331731e-13, 5.234923e-13, 
    5.161293e-13, 4.929902e-13, 5.012058e-13, 5.093697e-13, 5.238225e-13, 
    5.798549e-13, 5.918877e-13, 5.914753e-13, 5.684461e-13, 6.062123e-13, 
    7.123695e-13, 6.621006e-13, 6.627242e-13, 6.741534e-13, 6.521358e-13, 
    6.063888e-13, 5.462562e-13, 5.374434e-13, 5.26217e-13,
  2.637334e-12, 2.637975e-12, 2.644188e-12, 2.543401e-12, 2.586847e-12, 
    2.634418e-12, 2.592343e-12, 2.61499e-12, 2.540438e-12, 2.580571e-12, 
    2.57786e-12, 2.479439e-12, 2.450931e-12, 2.424724e-12, 2.448541e-12, 
    2.466252e-12, 2.466813e-12, 2.506538e-12, 2.562448e-12, 2.571095e-12, 
    2.654498e-12, 2.686154e-12, 2.50158e-12, 2.45552e-12, 2.427911e-12, 
    2.390132e-12, 2.450411e-12, 2.45524e-12, 2.60804e-12,
  3.493049e-12, 3.617384e-12, 3.600898e-12, 3.582718e-12, 3.623084e-12, 
    3.544514e-12, 3.610686e-12, 3.607896e-12, 3.484956e-12, 3.514298e-12, 
    3.548039e-12, 3.577735e-12, 3.467259e-12, 3.344933e-12, 3.285618e-12, 
    3.233945e-12, 3.186245e-12, 3.093946e-12, 3.218793e-12, 3.172364e-12, 
    3.238224e-12, 3.37054e-12, 3.477039e-12, 3.489259e-12, 3.427903e-12, 
    3.352786e-12, 3.479893e-12, 3.385511e-12, 3.412669e-12,
  2.203521e-12, 2.214585e-12, 2.1199e-12, 2.297639e-12, 2.408937e-12, 
    2.389936e-12, 2.373058e-12, 2.417734e-12, 2.559269e-12, 2.622658e-12, 
    2.633771e-12, 2.728942e-12, 2.685244e-12, 2.624805e-12, 2.559267e-12, 
    2.442448e-12, 2.462582e-12, 2.366398e-12, 2.315521e-12, 2.371042e-12, 
    2.201259e-12, 2.206926e-12, 2.126623e-12, 2.074642e-12, 2.136813e-12, 
    2.143946e-12, 2.097945e-12, 2.04411e-12, 2.034929e-12,
  2.74193e-12, 2.824954e-12, 2.758088e-12, 2.910032e-12, 2.888307e-12, 
    2.864588e-12, 3.001575e-12, 3.113005e-12, 3.09829e-12, 3.23901e-12, 
    3.228402e-12, 3.262179e-12, 3.13408e-12, 3.016902e-12, 3.175739e-12, 
    3.177854e-12, 3.123167e-12, 3.001527e-12, 2.992286e-12, 3.078373e-12, 
    2.949921e-12, 2.878401e-12, 2.77232e-12, 2.707291e-12, 2.666093e-12, 
    2.695236e-12, 2.621124e-12, 2.646968e-12, 2.726068e-12,
  2.762807e-12, 2.795467e-12, 2.782711e-12, 2.725547e-12, 2.597411e-12, 
    2.573163e-12, 2.609261e-12, 2.585508e-12, 2.628245e-12, 2.602822e-12, 
    2.657365e-12, 2.784289e-12, 2.776184e-12, 2.888335e-12, 2.820802e-12, 
    2.755624e-12, 3.192191e-12, 3.378641e-12, 3.151804e-12, 3.024924e-12, 
    3.172899e-12, 3.298324e-12, 3.121246e-12, 2.981395e-12, 3.004748e-12, 
    2.846707e-12, 2.715339e-12, 2.692154e-12, 2.568397e-12,
  1.087746e-12, 1.024048e-12, 9.88129e-13, 8.469232e-13, 8.84722e-13, 
    8.861442e-13, 7.406136e-13, 7.629887e-13, 6.42556e-13, 5.826264e-13, 
    5.395482e-13, 5.989999e-13, 5.332126e-13, 6.636317e-13, 9.413924e-13, 
    9.729772e-13, 7.811036e-13, 8.020588e-13, 9.930741e-13, 1.209087e-12, 
    1.341784e-12, 1.529816e-12, 1.506919e-12, 1.47151e-12, 1.308133e-12, 
    1.388528e-12, 1.341886e-12, 1.232138e-12, 1.149628e-12,
  4.297259e-13, 4.202702e-13, 3.307923e-13, 2.792092e-13, 2.742376e-13, 
    3.648994e-13, 3.683204e-13, 2.846391e-13, 1.791006e-13, 1.542895e-13, 
    1.241857e-13, 1.329948e-13, 1.353611e-13, 1.130098e-13, 1.585447e-13, 
    1.467802e-13, 9.957361e-14, 9.842425e-14, 1.066585e-13, 1.05296e-13, 
    1.211599e-13, 1.700193e-13, 2.666646e-13, 5.881757e-13, 6.613219e-13, 
    6.365541e-13, 5.691745e-13, 4.678321e-13, 4.739282e-13,
  8.216365e-14, 4.187926e-14, 6.357837e-14, 7.3357e-14, 7.952687e-14, 
    1.240943e-13, 1.957253e-13, 1.951202e-13, 2.772577e-13, 2.250274e-13, 
    1.740345e-13, 1.580423e-13, 9.576763e-14, 6.505628e-14, 5.765086e-14, 
    6.574204e-14, 9.29072e-14, 7.489686e-14, 6.068459e-14, 6.455509e-14, 
    6.026767e-14, 4.635779e-14, 4.504615e-14, 4.032698e-14, 4.716329e-14, 
    9.26333e-14, 1.109451e-13, 1.280348e-13, 1.141627e-13,
  4.752543e-15, 4.254256e-15, 8.018483e-15, 1.48031e-14, 2.200128e-14, 
    3.596584e-14, 8.676546e-14, 1.354145e-13, 1.2778e-13, 1.347902e-13, 
    1.368074e-13, 1.163363e-13, 6.975951e-14, 6.195671e-14, 5.417759e-14, 
    6.915656e-14, 9.62534e-14, 8.074516e-14, 5.735823e-14, 6.0361e-14, 
    3.84787e-14, 4.054818e-14, 4.467919e-14, 2.007185e-14, 1.334157e-14, 
    8.69008e-15, 6.112402e-15, 5.181265e-15, 5.110852e-15,
  2.671211e-15, 2.216625e-15, 1.830755e-15, 5.652012e-15, 5.832492e-15, 
    7.979114e-15, 1.102604e-14, 3.42667e-14, 4.080466e-14, 5.761818e-14, 
    4.979668e-14, 4.713418e-14, 4.356165e-14, 5.039428e-14, 5.535388e-14, 
    6.290672e-14, 5.537125e-14, 4.579972e-14, 4.306664e-14, 3.842567e-14, 
    4.060365e-14, 2.906527e-14, 2.560993e-14, 1.250103e-14, 2.188226e-15, 
    1.680895e-15, 1.693863e-15, 1.873247e-15, 2.38036e-15,
  8.961511e-16, 7.12187e-16, 6.974944e-16, 6.64063e-16, 1.122245e-15, 
    3.332786e-15, 5.277067e-15, 1.092967e-14, 1.788988e-14, 1.983185e-14, 
    2.247748e-14, 2.951666e-14, 3.484096e-14, 3.579993e-14, 3.598674e-14, 
    3.557985e-14, 3.407367e-14, 3.213367e-14, 3.102893e-14, 3.174665e-14, 
    2.431945e-14, 1.680898e-14, 1.087817e-14, 5.040786e-15, 2.022024e-15, 
    1.50123e-15, 1.367475e-15, 1.169203e-15, 9.80995e-16,
  7.15242e-16, 7.15242e-16, 7.15242e-16, 7.15242e-16, 7.15242e-16, 
    7.15242e-16, 7.15242e-16, 7.307335e-16, 7.307335e-16, 7.307335e-16, 
    7.307335e-16, 7.307335e-16, 7.307335e-16, 7.307335e-16, 7.345109e-16, 
    7.345109e-16, 7.345109e-16, 7.345109e-16, 7.345109e-16, 7.345109e-16, 
    7.345109e-16, 7.2787e-16, 7.2787e-16, 7.2787e-16, 7.2787e-16, 7.2787e-16, 
    7.2787e-16, 7.2787e-16, 7.15242e-16,
  2.029833e-15, 2.382652e-15, 2.387313e-15, 2.182593e-15, 2.062252e-15, 
    1.970156e-15, 1.850174e-15, 1.702376e-15, 1.420806e-15, 1.36142e-15, 
    1.409594e-15, 1.451119e-15, 1.462043e-15, 1.446669e-15, 1.324731e-15, 
    1.215254e-15, 1.217635e-15, 1.265989e-15, 1.22396e-15, 1.159849e-15, 
    1.115986e-15, 1.025437e-15, 9.460654e-16, 8.879689e-16, 8.037537e-16, 
    7.466268e-16, 8.276008e-16, 1.086445e-15, 1.871303e-15,
  3.628464e-15, 4.523035e-15, 5.625334e-15, 6.120078e-15, 6.043067e-15, 
    5.550798e-15, 5.579388e-15, 6.089234e-15, 7.967162e-15, 9.720523e-15, 
    1.059216e-14, 1.105662e-14, 9.885105e-15, 8.622902e-15, 7.993408e-15, 
    7.708596e-15, 6.769428e-15, 5.841892e-15, 4.64494e-15, 3.494125e-15, 
    3.285346e-15, 3.066331e-15, 2.873816e-15, 2.755819e-15, 2.784559e-15, 
    5.992736e-15, 7.38252e-15, 5.337068e-15, 3.719275e-15,
  4.644193e-14, 5.32926e-14, 4.541672e-14, 4.741118e-14, 5.993346e-14, 
    6.710151e-14, 5.382127e-14, 4.2083e-14, 3.665094e-14, 3.586504e-14, 
    3.385629e-14, 3.963234e-14, 6.198763e-14, 8.323373e-14, 1.17373e-13, 
    1.510129e-13, 1.247349e-13, 8.232528e-14, 8.625218e-14, 8.879415e-14, 
    5.885326e-14, 4.801045e-14, 3.757206e-14, 1.854847e-14, 2.280856e-14, 
    2.076377e-14, 2.171258e-14, 3.228795e-14, 3.997152e-14,
  1.610682e-13, 1.624569e-13, 1.27851e-13, 9.903589e-14, 9.32064e-14, 
    8.963574e-14, 7.990506e-14, 7.460017e-14, 7.126703e-14, 7.665814e-14, 
    9.13069e-14, 1.060162e-13, 9.194265e-14, 8.56597e-14, 9.137166e-14, 
    1.076324e-13, 1.517751e-13, 1.938337e-13, 2.020582e-13, 1.412742e-13, 
    9.851099e-14, 1.365866e-13, 1.266334e-13, 1.355203e-13, 1.536416e-13, 
    1.227319e-13, 1.197321e-13, 1.379565e-13, 1.412052e-13,
  3.004467e-13, 3.076456e-13, 3.100136e-13, 2.810274e-13, 2.613976e-13, 
    2.116678e-13, 1.899651e-13, 1.906604e-13, 1.918169e-13, 1.40263e-13, 
    1.235e-13, 1.242385e-13, 1.441887e-13, 1.463261e-13, 1.512159e-13, 
    1.523577e-13, 1.713781e-13, 2.063493e-13, 2.451663e-13, 2.280582e-13, 
    3.144872e-13, 4.958327e-13, 6.638169e-13, 6.332881e-13, 5.178402e-13, 
    4.008479e-13, 3.603429e-13, 3.15526e-13, 3.351452e-13,
  1.692729e-12, 1.632824e-12, 1.55817e-12, 1.624438e-12, 1.682181e-12, 
    1.608675e-12, 1.656616e-12, 1.704127e-12, 1.718532e-12, 1.685943e-12, 
    1.728769e-12, 1.631856e-12, 1.615704e-12, 1.543622e-12, 1.630573e-12, 
    1.771786e-12, 1.894571e-12, 1.886588e-12, 1.837634e-12, 2.04257e-12, 
    2.296057e-12, 2.200383e-12, 2.195547e-12, 2.271794e-12, 2.243673e-12, 
    1.90828e-12, 1.780647e-12, 1.778175e-12, 1.716337e-12,
  1.00883e-11, 1.011932e-11, 9.840899e-12, 9.804511e-12, 9.505607e-12, 
    9.347603e-12, 9.297179e-12, 9.478654e-12, 9.49024e-12, 9.573767e-12, 
    9.424137e-12, 9.252749e-12, 9.153396e-12, 9.397267e-12, 9.003394e-12, 
    8.935387e-12, 8.839525e-12, 9.058995e-12, 9.18604e-12, 9.519874e-12, 
    9.625092e-12, 9.51232e-12, 9.636695e-12, 9.533902e-12, 9.554112e-12, 
    9.42408e-12, 9.335041e-12, 9.656437e-12, 9.909276e-12,
  1.425785e-11, 1.432e-11, 1.435299e-11, 1.421532e-11, 1.446157e-11, 
    1.473796e-11, 1.458042e-11, 1.442195e-11, 1.448378e-11, 1.436655e-11, 
    1.405549e-11, 1.397172e-11, 1.357579e-11, 1.304933e-11, 1.284688e-11, 
    1.293773e-11, 1.292538e-11, 1.300747e-11, 1.320557e-11, 1.364042e-11, 
    1.338437e-11, 1.388565e-11, 1.388078e-11, 1.441481e-11, 1.454771e-11, 
    1.416054e-11, 1.392191e-11, 1.393332e-11, 1.422198e-11,
  9.760914e-12, 9.826088e-12, 9.906386e-12, 1.003361e-11, 1.016497e-11, 
    1.059484e-11, 1.075605e-11, 1.099695e-11, 1.133933e-11, 1.158469e-11, 
    1.136809e-11, 1.119274e-11, 1.096595e-11, 1.101331e-11, 1.114373e-11, 
    1.084898e-11, 1.087447e-11, 1.060753e-11, 1.057381e-11, 1.038191e-11, 
    9.850069e-12, 9.429726e-12, 9.264013e-12, 9.330248e-12, 9.423548e-12, 
    9.549308e-12, 9.426162e-12, 9.81587e-12, 9.87556e-12,
  1.084991e-11, 1.074842e-11, 1.122188e-11, 1.132746e-11, 1.133347e-11, 
    1.170864e-11, 1.177823e-11, 1.190633e-11, 1.219115e-11, 1.243239e-11, 
    1.24182e-11, 1.260402e-11, 1.195612e-11, 1.193136e-11, 1.264212e-11, 
    1.308911e-11, 1.325799e-11, 1.300381e-11, 1.360226e-11, 1.311156e-11, 
    1.307169e-11, 1.238498e-11, 1.167969e-11, 1.074713e-11, 9.970949e-12, 
    9.982582e-12, 1.021991e-11, 1.034717e-11, 1.094375e-11,
  1.017219e-11, 1.035972e-11, 1.030476e-11, 1.018759e-11, 9.994962e-12, 
    9.997604e-12, 9.583396e-12, 9.017225e-12, 9.537516e-12, 9.142176e-12, 
    9.582367e-12, 1.013678e-11, 1.040485e-11, 1.086294e-11, 1.120588e-11, 
    1.147188e-11, 1.215861e-11, 1.208519e-11, 1.18529e-11, 1.141378e-11, 
    1.249973e-11, 1.241488e-11, 1.163602e-11, 1.108186e-11, 1.026569e-11, 
    1.001868e-11, 1.009754e-11, 1.008131e-11, 1.008176e-11,
  3.291912e-12, 3.237509e-12, 2.938656e-12, 2.601822e-12, 3.118129e-12, 
    3.070901e-12, 2.434993e-12, 2.20825e-12, 2.087366e-12, 1.937722e-12, 
    1.606643e-12, 1.913362e-12, 1.992414e-12, 2.50313e-12, 2.689947e-12, 
    3.080544e-12, 2.57609e-12, 2.563276e-12, 3.486147e-12, 3.743826e-12, 
    4.503533e-12, 5.455231e-12, 4.536627e-12, 4.529463e-12, 4.184007e-12, 
    4.258373e-12, 4.086125e-12, 3.442248e-12, 3.30319e-12,
  1.565462e-12, 1.426001e-12, 1.169268e-12, 8.894114e-13, 8.333362e-13, 
    1.180991e-12, 1.11042e-12, 7.603651e-13, 5.57646e-13, 4.764761e-13, 
    3.792368e-13, 3.755485e-13, 6.473789e-13, 3.356768e-13, 4.569132e-13, 
    6.26181e-13, 2.625772e-13, 2.276979e-13, 2.599073e-13, 2.857232e-13, 
    3.903407e-13, 5.609176e-13, 1.23133e-12, 2.068958e-12, 1.995188e-12, 
    1.933799e-12, 1.528084e-12, 1.295284e-12, 1.613713e-12,
  4.014238e-13, 1.596671e-13, 1.7121e-13, 2.724776e-13, 3.081021e-13, 
    3.697557e-13, 6.672193e-13, 5.213857e-13, 6.273257e-13, 6.184451e-13, 
    4.921475e-13, 4.040723e-13, 3.198036e-13, 2.394507e-13, 2.259596e-13, 
    2.676463e-13, 2.993572e-13, 2.899862e-13, 1.958656e-13, 1.916531e-13, 
    1.93964e-13, 1.514285e-13, 1.336546e-13, 1.183331e-13, 1.460836e-13, 
    4.590527e-13, 5.307487e-13, 5.943396e-13, 5.382826e-13,
  1.386431e-14, 1.278971e-14, 1.58387e-14, 4.146252e-14, 6.18536e-14, 
    1.247736e-13, 2.407199e-13, 3.858581e-13, 3.401782e-13, 3.466219e-13, 
    3.642221e-13, 3.656277e-13, 2.267156e-13, 1.612792e-13, 1.404728e-13, 
    2.051808e-13, 2.716368e-13, 2.543297e-13, 1.693129e-13, 1.853623e-13, 
    1.125678e-13, 8.652326e-14, 1.204725e-13, 6.965918e-14, 3.801771e-14, 
    2.830141e-14, 1.847222e-14, 1.451943e-14, 1.441044e-14,
  8.936573e-15, 8.176493e-15, 5.896837e-15, 1.255228e-14, 1.716404e-14, 
    1.734683e-14, 2.991673e-14, 9.565883e-14, 1.416359e-13, 1.57586e-13, 
    1.482827e-13, 1.506885e-13, 1.462365e-13, 1.652069e-13, 1.709052e-13, 
    1.900179e-13, 1.912674e-13, 1.541999e-13, 1.454476e-13, 1.071891e-13, 
    1.030169e-13, 8.642208e-14, 7.793915e-14, 4.669611e-14, 8.050501e-15, 
    5.577533e-15, 5.657008e-15, 6.298866e-15, 7.912668e-15,
  2.362214e-15, 2.046984e-15, 2.218673e-15, 2.247455e-15, 2.028843e-15, 
    4.936175e-15, 1.171158e-14, 1.955988e-14, 5.124062e-14, 5.481229e-14, 
    5.868176e-14, 8.464112e-14, 1.022559e-13, 1.109526e-13, 1.047502e-13, 
    9.449422e-14, 8.365879e-14, 7.605024e-14, 8.092819e-14, 9.408124e-14, 
    6.67985e-14, 5.543164e-14, 4.263755e-14, 2.125768e-14, 7.82408e-15, 
    4.534042e-15, 3.987787e-15, 3.344648e-15, 2.64711e-15,
  2.061948e-15, 2.061948e-15, 2.061948e-15, 2.061948e-15, 2.061948e-15, 
    2.061948e-15, 2.061948e-15, 2.148945e-15, 2.148945e-15, 2.148945e-15, 
    2.148945e-15, 2.148945e-15, 2.148945e-15, 2.148945e-15, 2.160922e-15, 
    2.160922e-15, 2.160922e-15, 2.160922e-15, 2.160922e-15, 2.160922e-15, 
    2.160922e-15, 2.084252e-15, 2.084252e-15, 2.084252e-15, 2.084252e-15, 
    2.084252e-15, 2.084252e-15, 2.084252e-15, 2.061948e-15,
  4.043051e-15, 5.290443e-15, 5.696812e-15, 5.452914e-15, 5.452771e-15, 
    5.057839e-15, 4.325547e-15, 3.54304e-15, 3.313606e-15, 3.387942e-15, 
    3.863072e-15, 4.065323e-15, 4.153821e-15, 4.077624e-15, 3.903722e-15, 
    3.589989e-15, 3.524243e-15, 3.632108e-15, 3.592124e-15, 3.446876e-15, 
    3.178926e-15, 2.843076e-15, 2.403498e-15, 2.186173e-15, 1.92722e-15, 
    1.655366e-15, 1.613228e-15, 1.979854e-15, 3.415586e-15,
  1.103167e-14, 1.368977e-14, 1.729191e-14, 1.80135e-14, 1.622836e-14, 
    1.661658e-14, 1.738463e-14, 1.721031e-14, 2.042907e-14, 2.465233e-14, 
    2.70454e-14, 2.658762e-14, 2.442715e-14, 2.297198e-14, 2.310986e-14, 
    2.283363e-14, 2.030934e-14, 1.662354e-14, 1.259467e-14, 9.68209e-15, 
    9.551288e-15, 9.311459e-15, 8.16662e-15, 7.740435e-15, 7.348919e-15, 
    1.29086e-14, 2.011442e-14, 1.754799e-14, 1.263319e-14,
  1.347713e-13, 1.530042e-13, 1.540702e-13, 1.8067e-13, 2.237103e-13, 
    2.304911e-13, 1.603869e-13, 1.332714e-13, 1.197309e-13, 1.229764e-13, 
    1.156064e-13, 1.618512e-13, 2.762969e-13, 3.630697e-13, 4.665899e-13, 
    6.239085e-13, 5.481847e-13, 3.22387e-13, 3.065037e-13, 2.983702e-13, 
    2.033459e-13, 1.363172e-13, 1.210982e-13, 6.389908e-14, 7.960591e-14, 
    7.925054e-14, 8.80373e-14, 1.120613e-13, 1.183367e-13,
  6.218026e-13, 6.5195e-13, 5.723678e-13, 3.634135e-13, 3.224704e-13, 
    3.12151e-13, 2.886219e-13, 2.408557e-13, 2.236087e-13, 2.834018e-13, 
    3.601972e-13, 3.711149e-13, 2.949631e-13, 2.82122e-13, 3.358404e-13, 
    4.243086e-13, 5.473518e-13, 5.994079e-13, 5.601121e-13, 5.354524e-13, 
    3.348126e-13, 4.164022e-13, 4.844104e-13, 5.239512e-13, 5.633e-13, 
    4.44301e-13, 4.233362e-13, 5.428701e-13, 5.297526e-13,
  1.159119e-12, 1.148241e-12, 1.320756e-12, 1.275796e-12, 1.09302e-12, 
    7.993238e-13, 6.854458e-13, 6.527994e-13, 6.237775e-13, 5.502325e-13, 
    4.318363e-13, 4.30996e-13, 5.225915e-13, 5.891159e-13, 5.656047e-13, 
    4.812747e-13, 5.366187e-13, 7.291564e-13, 6.842953e-13, 6.205514e-13, 
    7.249298e-13, 1.241167e-12, 1.448635e-12, 1.681991e-12, 1.629565e-12, 
    1.538717e-12, 1.361075e-12, 1.221115e-12, 1.452234e-12,
  5.043735e-12, 4.776623e-12, 4.870509e-12, 5.042814e-12, 5.599399e-12, 
    5.203986e-12, 5.449231e-12, 5.589004e-12, 5.315286e-12, 5.572564e-12, 
    5.628878e-12, 5.394048e-12, 4.978434e-12, 4.855884e-12, 5.253429e-12, 
    5.539038e-12, 5.872726e-12, 6.094674e-12, 6.365652e-12, 7.338873e-12, 
    7.922384e-12, 7.684914e-12, 7.422274e-12, 7.3422e-12, 6.710269e-12, 
    5.910769e-12, 5.71155e-12, 5.982425e-12, 5.476639e-12,
  3.613577e-11, 3.538739e-11, 3.471502e-11, 3.410483e-11, 3.395407e-11, 
    3.425689e-11, 3.434482e-11, 3.365309e-11, 3.474592e-11, 3.43834e-11, 
    3.316825e-11, 3.297179e-11, 3.228258e-11, 3.307984e-11, 3.200817e-11, 
    3.240339e-11, 3.271136e-11, 3.287887e-11, 3.318499e-11, 3.376502e-11, 
    3.524811e-11, 3.515525e-11, 3.420146e-11, 3.507095e-11, 3.396491e-11, 
    3.524797e-11, 3.476167e-11, 3.580734e-11, 3.698093e-11,
  5.853026e-11, 5.848286e-11, 5.815752e-11, 5.846525e-11, 5.800462e-11, 
    5.816609e-11, 5.905768e-11, 5.861234e-11, 5.784774e-11, 5.602841e-11, 
    5.497615e-11, 5.496494e-11, 5.423331e-11, 5.333071e-11, 5.308612e-11, 
    5.234703e-11, 5.319759e-11, 5.448751e-11, 5.594816e-11, 5.685188e-11, 
    5.716665e-11, 5.862109e-11, 6.062206e-11, 6.050142e-11, 6.076828e-11, 
    6.002106e-11, 5.999481e-11, 5.911784e-11, 5.870313e-11,
  4.944149e-11, 4.87748e-11, 4.926397e-11, 4.845173e-11, 4.90257e-11, 
    5.001528e-11, 5.300366e-11, 5.527178e-11, 5.674224e-11, 5.69117e-11, 
    5.712061e-11, 5.599491e-11, 5.497924e-11, 5.512283e-11, 5.504502e-11, 
    5.697894e-11, 5.806943e-11, 5.885162e-11, 5.880246e-11, 5.826064e-11, 
    5.904441e-11, 6.182268e-11, 6.08198e-11, 5.94625e-11, 5.632949e-11, 
    5.205041e-11, 5.029168e-11, 5.026696e-11, 4.928764e-11,
  3.661148e-11, 3.63528e-11, 3.538706e-11, 3.562216e-11, 3.650324e-11, 
    3.693771e-11, 3.824032e-11, 3.868563e-11, 3.930374e-11, 4.093095e-11, 
    4.22719e-11, 4.450861e-11, 4.53486e-11, 4.463936e-11, 4.550522e-11, 
    4.612532e-11, 4.735728e-11, 4.768791e-11, 4.849888e-11, 4.96723e-11, 
    4.744105e-11, 4.639589e-11, 4.437905e-11, 4.127193e-11, 3.690653e-11, 
    3.477073e-11, 3.24229e-11, 3.36806e-11, 3.512498e-11,
  3.115363e-11, 3.212695e-11, 3.225056e-11, 3.115661e-11, 2.961056e-11, 
    3.02052e-11, 2.893236e-11, 2.910282e-11, 3.025807e-11, 2.885739e-11, 
    3.149015e-11, 3.547009e-11, 3.69018e-11, 3.78845e-11, 3.938787e-11, 
    3.932471e-11, 3.888226e-11, 3.793752e-11, 3.77938e-11, 3.627745e-11, 
    3.721573e-11, 3.701392e-11, 3.597891e-11, 3.530118e-11, 3.37776e-11, 
    3.07823e-11, 3.141282e-11, 3.142645e-11, 3.224353e-11,
  8.577298e-12, 8.686288e-12, 7.769629e-12, 7.147827e-12, 8.245024e-12, 
    7.680349e-12, 7.551604e-12, 6.013206e-12, 5.643028e-12, 5.587053e-12, 
    4.368123e-12, 5.791601e-12, 6.233997e-12, 8.23718e-12, 7.881425e-12, 
    8.076425e-12, 7.646826e-12, 8.275278e-12, 9.217412e-12, 1.000454e-11, 
    1.241258e-11, 1.325619e-11, 1.158593e-11, 1.086163e-11, 9.973597e-12, 
    9.714465e-12, 9.840121e-12, 8.89575e-12, 8.549067e-12,
  3.618763e-12, 3.633759e-12, 2.895731e-12, 1.796232e-12, 1.755063e-12, 
    2.610262e-12, 2.436336e-12, 1.548993e-12, 1.468733e-12, 1.399782e-12, 
    1.059316e-12, 9.881588e-13, 1.694531e-12, 1.068275e-12, 8.940878e-13, 
    1.502307e-12, 6.647208e-13, 6.21236e-13, 6.833738e-13, 6.644909e-13, 
    1.108538e-12, 1.732203e-12, 3.565309e-12, 3.922268e-12, 3.99939e-12, 
    4.120863e-12, 3.261254e-12, 2.947854e-12, 3.675237e-12,
  1.064946e-12, 4.500088e-13, 3.674046e-13, 7.622647e-13, 9.155589e-13, 
    9.115257e-13, 1.522332e-12, 1.133683e-12, 1.043958e-12, 1.191976e-12, 
    1.212765e-12, 9.158809e-13, 7.180732e-13, 7.2167e-13, 7.352731e-13, 
    7.275685e-13, 7.405168e-13, 7.056631e-13, 4.654416e-13, 4.647102e-13, 
    4.105905e-13, 3.763344e-13, 2.946911e-13, 2.610845e-13, 4.739797e-13, 
    1.136926e-12, 1.273666e-12, 1.441627e-12, 1.345326e-12,
  4.73346e-14, 4.335932e-14, 3.80569e-14, 7.756254e-14, 1.336005e-13, 
    2.698449e-13, 6.290456e-13, 8.767769e-13, 7.807036e-13, 7.502517e-13, 
    7.586108e-13, 7.766927e-13, 6.287356e-13, 4.428933e-13, 3.836523e-13, 
    4.597759e-13, 5.35242e-13, 4.819292e-13, 3.765353e-13, 3.805055e-13, 
    3.006981e-13, 2.067506e-13, 2.836148e-13, 2.153096e-13, 1.152152e-13, 
    7.829914e-14, 6.274565e-14, 5.344098e-14, 4.808188e-14,
  2.460083e-14, 2.261564e-14, 1.586761e-14, 2.066116e-14, 3.563479e-14, 
    3.450787e-14, 6.009659e-14, 2.553486e-13, 3.844839e-13, 3.748075e-13, 
    3.589326e-13, 4.169974e-13, 4.153077e-13, 4.428558e-13, 4.30821e-13, 
    4.043151e-13, 4.027228e-13, 3.60009e-13, 3.481466e-13, 2.699839e-13, 
    2.318064e-13, 2.047814e-13, 1.873143e-13, 1.211004e-13, 3.071338e-14, 
    2.135956e-14, 2.193628e-14, 2.30955e-14, 2.406276e-14,
  6.761017e-15, 5.073286e-15, 4.650426e-15, 5.187209e-15, 5.350327e-15, 
    5.565649e-15, 1.257339e-14, 2.159465e-14, 6.904876e-14, 1.223677e-13, 
    1.282403e-13, 2.31897e-13, 2.835589e-13, 2.809293e-13, 2.45642e-13, 
    2.148432e-13, 1.857055e-13, 1.702389e-13, 1.954002e-13, 2.12688e-13, 
    1.559528e-13, 1.195423e-13, 1.023396e-13, 6.446308e-14, 2.630799e-14, 
    1.281969e-14, 1.076093e-14, 9.420277e-15, 7.647993e-15,
  6.156443e-15, 6.156443e-15, 6.156443e-15, 6.156443e-15, 6.156443e-15, 
    6.156443e-15, 6.156443e-15, 6.436592e-15, 6.436592e-15, 6.436592e-15, 
    6.436592e-15, 6.436592e-15, 6.436592e-15, 6.436592e-15, 6.426741e-15, 
    6.426741e-15, 6.426741e-15, 6.426741e-15, 6.426741e-15, 6.426741e-15, 
    6.426741e-15, 6.192577e-15, 6.192577e-15, 6.192577e-15, 6.192577e-15, 
    6.192577e-15, 6.192577e-15, 6.192577e-15, 6.156443e-15,
  6.723339e-15, 1.066336e-14, 1.299736e-14, 1.25997e-14, 1.271361e-14, 
    1.05089e-14, 8.852269e-15, 9.269352e-15, 1.036299e-14, 1.065708e-14, 
    1.091347e-14, 1.101901e-14, 1.10738e-14, 1.097423e-14, 1.067168e-14, 
    1.043349e-14, 1.09894e-14, 1.184808e-14, 1.108151e-14, 1.007077e-14, 
    9.397117e-15, 8.08476e-15, 7.108847e-15, 5.85795e-15, 4.598178e-15, 
    3.787385e-15, 3.619942e-15, 3.891297e-15, 5.417765e-15,
  3.461073e-14, 3.286738e-14, 4.669447e-14, 5.209478e-14, 4.765386e-14, 
    4.973191e-14, 4.931281e-14, 4.980318e-14, 5.564667e-14, 6.558313e-14, 
    7.149248e-14, 7.18284e-14, 7.07491e-14, 6.840599e-14, 7.032049e-14, 
    7.348352e-14, 6.677143e-14, 5.504247e-14, 3.993299e-14, 3.283123e-14, 
    3.196637e-14, 3.118877e-14, 2.871515e-14, 3.006533e-14, 2.277175e-14, 
    2.741126e-14, 6.235907e-14, 6.70572e-14, 4.204666e-14,
  4.073626e-13, 5.913078e-13, 5.921721e-13, 6.241221e-13, 7.975812e-13, 
    7.80051e-13, 5.679854e-13, 5.068537e-13, 4.171847e-13, 3.66957e-13, 
    3.354507e-13, 5.122302e-13, 7.97258e-13, 1.022229e-12, 1.151306e-12, 
    1.392817e-12, 1.3422e-12, 1.071875e-12, 1.005674e-12, 8.747883e-13, 
    6.064826e-13, 3.843266e-13, 3.336184e-13, 2.200351e-13, 2.685583e-13, 
    3.159483e-13, 3.388004e-13, 3.301792e-13, 3.347829e-13,
  2.479364e-12, 2.489297e-12, 2.070118e-12, 1.366382e-12, 9.9682e-13, 
    1.005172e-12, 9.921671e-13, 8.647701e-13, 7.846999e-13, 9.947491e-13, 
    1.329259e-12, 1.186112e-12, 9.750379e-13, 9.912443e-13, 1.123703e-12, 
    1.316171e-12, 1.476239e-12, 1.483868e-12, 1.116201e-12, 1.167436e-12, 
    9.653312e-13, 1.018793e-12, 1.322451e-12, 1.662295e-12, 2.410947e-12, 
    2.332627e-12, 2.128052e-12, 2.416644e-12, 2.292577e-12,
  4.27055e-12, 4.006413e-12, 4.698131e-12, 4.47459e-12, 3.643431e-12, 
    2.504243e-12, 2.178755e-12, 2.048628e-12, 2.220554e-12, 2.064337e-12, 
    1.630469e-12, 1.763449e-12, 2.03634e-12, 2.115646e-12, 2.026223e-12, 
    1.762486e-12, 1.91142e-12, 2.794933e-12, 2.218169e-12, 1.946642e-12, 
    2.582121e-12, 4.746078e-12, 4.652662e-12, 5.462025e-12, 4.913229e-12, 
    5.721337e-12, 4.990881e-12, 4.474185e-12, 5.030904e-12,
  1.553e-11, 1.488053e-11, 1.495395e-11, 1.576457e-11, 1.814782e-11, 
    1.849972e-11, 1.802753e-11, 1.725558e-11, 1.593973e-11, 1.636406e-11, 
    1.668039e-11, 1.535833e-11, 1.605318e-11, 1.487903e-11, 1.603227e-11, 
    1.753522e-11, 1.861796e-11, 1.954785e-11, 1.910011e-11, 2.322255e-11, 
    2.595206e-11, 2.363673e-11, 2.296388e-11, 2.257042e-11, 2.086869e-11, 
    1.823103e-11, 1.737313e-11, 1.768871e-11, 1.672245e-11,
  1.244854e-10, 1.24653e-10, 1.248351e-10, 1.209204e-10, 1.197058e-10, 
    1.17533e-10, 1.211353e-10, 1.202631e-10, 1.199133e-10, 1.175871e-10, 
    1.210023e-10, 1.195843e-10, 1.145178e-10, 1.115415e-10, 1.112953e-10, 
    1.095559e-10, 1.11426e-10, 1.129516e-10, 1.219833e-10, 1.249135e-10, 
    1.244367e-10, 1.27178e-10, 1.266493e-10, 1.235526e-10, 1.228848e-10, 
    1.254329e-10, 1.227352e-10, 1.224685e-10, 1.251103e-10,
  2.311508e-10, 2.243579e-10, 2.256657e-10, 2.2487e-10, 2.307753e-10, 
    2.328581e-10, 2.297315e-10, 2.258645e-10, 2.196986e-10, 2.149682e-10, 
    2.096434e-10, 2.085006e-10, 2.014735e-10, 2.02137e-10, 2.026228e-10, 
    2.084307e-10, 2.1096e-10, 2.169916e-10, 2.233597e-10, 2.280121e-10, 
    2.405093e-10, 2.43329e-10, 2.448323e-10, 2.477561e-10, 2.435322e-10, 
    2.315534e-10, 2.314271e-10, 2.302433e-10, 2.304039e-10,
  2.093363e-10, 1.977114e-10, 1.952783e-10, 1.951067e-10, 2.064101e-10, 
    2.100488e-10, 2.093894e-10, 2.16032e-10, 2.276232e-10, 2.280565e-10, 
    2.2773e-10, 2.273884e-10, 2.217667e-10, 2.113105e-10, 2.125402e-10, 
    2.104817e-10, 2.12275e-10, 2.159051e-10, 2.219264e-10, 2.203527e-10, 
    2.302518e-10, 2.260511e-10, 2.371906e-10, 2.340281e-10, 2.459298e-10, 
    2.513956e-10, 2.278592e-10, 2.220331e-10, 2.099297e-10,
  1.04896e-10, 1.049801e-10, 1.083489e-10, 1.111687e-10, 1.172233e-10, 
    1.141616e-10, 1.162811e-10, 1.212064e-10, 1.273025e-10, 1.298811e-10, 
    1.36364e-10, 1.398679e-10, 1.469292e-10, 1.468113e-10, 1.412603e-10, 
    1.411216e-10, 1.438941e-10, 1.423497e-10, 1.364123e-10, 1.398869e-10, 
    1.40109e-10, 1.350031e-10, 1.317932e-10, 1.236447e-10, 1.238498e-10, 
    1.172264e-10, 1.088257e-10, 1.078569e-10, 1.036689e-10,
  9.317296e-11, 9.56813e-11, 9.585885e-11, 9.408985e-11, 9.44746e-11, 
    9.269778e-11, 9.020858e-11, 9.126456e-11, 9.359861e-11, 1.019118e-10, 
    1.178967e-10, 1.294457e-10, 1.251176e-10, 1.194808e-10, 1.180269e-10, 
    1.145545e-10, 1.133192e-10, 1.128678e-10, 1.105894e-10, 1.11451e-10, 
    1.094425e-10, 1.054237e-10, 1.020413e-10, 9.709467e-11, 1.003661e-10, 
    1.00334e-10, 9.64382e-11, 9.535361e-11, 9.343316e-11,
  2.163217e-11, 2.058137e-11, 1.926219e-11, 1.800049e-11, 1.949799e-11, 
    1.887863e-11, 1.901816e-11, 1.665785e-11, 1.622684e-11, 1.545332e-11, 
    1.498379e-11, 2.02271e-11, 2.176816e-11, 2.468515e-11, 2.705816e-11, 
    2.631135e-11, 2.346019e-11, 2.438966e-11, 2.42668e-11, 2.507719e-11, 
    2.874899e-11, 2.794623e-11, 2.616794e-11, 2.287123e-11, 2.167095e-11, 
    2.222439e-11, 2.245904e-11, 2.188283e-11, 2.186603e-11,
  5.783095e-12, 6.528608e-12, 5.847005e-12, 3.738481e-12, 3.794103e-12, 
    4.533237e-12, 4.500738e-12, 3.074576e-12, 3.400747e-12, 4.085594e-12, 
    3.308556e-12, 2.935747e-12, 2.584525e-12, 2.109791e-12, 2.269788e-12, 
    2.576349e-12, 1.631028e-12, 1.850421e-12, 1.644856e-12, 1.573253e-12, 
    2.519483e-12, 3.670857e-12, 4.996341e-12, 5.753311e-12, 6.086076e-12, 
    6.955426e-12, 7.49836e-12, 5.446991e-12, 5.86069e-12,
  1.31097e-12, 4.8942e-13, 6.43092e-13, 1.388401e-12, 2.068262e-12, 
    1.841256e-12, 2.530933e-12, 1.869271e-12, 1.525091e-12, 1.865455e-12, 
    2.349511e-12, 2.154887e-12, 1.828984e-12, 1.474981e-12, 1.323408e-12, 
    1.107609e-12, 1.103445e-12, 1.165611e-12, 1.041294e-12, 1.102962e-12, 
    9.488619e-13, 8.489402e-13, 6.824279e-13, 5.026624e-13, 7.152129e-13, 
    1.525928e-12, 1.862529e-12, 1.938032e-12, 1.664831e-12,
  1.569542e-13, 1.487297e-13, 1.249705e-13, 1.603185e-13, 2.163663e-13, 
    4.173737e-13, 9.160448e-13, 1.512346e-12, 1.362874e-12, 1.321847e-12, 
    1.281026e-12, 1.423528e-12, 1.54761e-12, 1.311286e-12, 1.151666e-12, 
    1.013442e-12, 1.087112e-12, 9.910627e-13, 8.629931e-13, 8.539326e-13, 
    8.351938e-13, 6.304622e-13, 7.383242e-13, 7.056961e-13, 4.271653e-13, 
    2.476272e-13, 2.488836e-13, 2.230806e-13, 1.619103e-13,
  5.8682e-14, 4.996121e-14, 4.222932e-14, 4.466077e-14, 7.37856e-14, 
    4.96509e-14, 9.182015e-14, 3.746161e-13, 6.992158e-13, 6.205926e-13, 
    6.403915e-13, 7.491477e-13, 8.264177e-13, 8.220107e-13, 8.208352e-13, 
    7.775613e-13, 7.532249e-13, 6.972289e-13, 6.978451e-13, 6.14484e-13, 
    5.401518e-13, 4.176568e-13, 3.829096e-13, 2.935083e-13, 1.223202e-13, 
    5.824863e-14, 5.698903e-14, 6.247439e-14, 6.289212e-14,
  2.073703e-14, 1.463847e-14, 9.435258e-15, 9.025382e-15, 1.15098e-14, 
    1.305977e-14, 1.550072e-14, 2.464514e-14, 6.371522e-14, 2.033925e-13, 
    2.277823e-13, 3.985203e-13, 5.115737e-13, 5.31214e-13, 5.294445e-13, 
    4.734428e-13, 4.143205e-13, 4.011756e-13, 4.620845e-13, 4.062227e-13, 
    2.974372e-13, 2.384161e-13, 1.9881e-13, 1.615915e-13, 8.189231e-14, 
    3.652356e-14, 2.902165e-14, 2.725968e-14, 2.376913e-14,
  1.635776e-14, 1.635776e-14, 1.635776e-14, 1.635776e-14, 1.635776e-14, 
    1.635776e-14, 1.635776e-14, 1.682564e-14, 1.682564e-14, 1.682564e-14, 
    1.682564e-14, 1.682564e-14, 1.682564e-14, 1.682564e-14, 1.714907e-14, 
    1.714907e-14, 1.714907e-14, 1.714907e-14, 1.714907e-14, 1.714907e-14, 
    1.714907e-14, 1.67932e-14, 1.67932e-14, 1.67932e-14, 1.67932e-14, 
    1.67932e-14, 1.67932e-14, 1.67932e-14, 1.635776e-14,
  1.210668e-14, 1.835511e-14, 2.236926e-14, 2.135892e-14, 2.343876e-14, 
    1.965376e-14, 2.195872e-14, 2.708513e-14, 3.306985e-14, 3.285043e-14, 
    3.193229e-14, 3.190902e-14, 3.282258e-14, 3.371617e-14, 3.482579e-14, 
    3.720249e-14, 4.163756e-14, 4.526552e-14, 4.190765e-14, 3.500705e-14, 
    3.091131e-14, 2.546907e-14, 2.14135e-14, 1.578672e-14, 1.093746e-14, 
    1.000861e-14, 9.993407e-15, 1.023597e-14, 1.077206e-14,
  1.363382e-13, 1.110952e-13, 1.372406e-13, 1.499684e-13, 1.317515e-13, 
    1.38751e-13, 1.468619e-13, 1.651763e-13, 1.813882e-13, 1.847455e-13, 
    2.053799e-13, 2.147248e-13, 2.269608e-13, 2.225753e-13, 2.338293e-13, 
    2.622452e-13, 2.525654e-13, 2.16535e-13, 1.547041e-13, 1.211608e-13, 
    1.165052e-13, 9.911115e-14, 9.797032e-14, 1.025558e-13, 7.642414e-14, 
    8.122723e-14, 1.549003e-13, 2.334579e-13, 1.69661e-13,
  1.092716e-12, 1.575002e-12, 1.815147e-12, 1.935074e-12, 1.981058e-12, 
    1.676467e-12, 1.510485e-12, 1.384517e-12, 1.136165e-12, 9.835688e-13, 
    9.93186e-13, 1.284697e-12, 1.780009e-12, 2.223132e-12, 2.354225e-12, 
    2.626865e-12, 2.904338e-12, 2.988469e-12, 2.759346e-12, 2.526402e-12, 
    1.886225e-12, 1.149733e-12, 9.836438e-13, 8.427818e-13, 9.178003e-13, 
    1.064248e-12, 9.510432e-13, 8.984169e-13, 9.876428e-13,
  5.9893e-12, 5.592848e-12, 4.629444e-12, 4.387946e-12, 3.468619e-12, 
    3.752379e-12, 3.602591e-12, 3.252828e-12, 2.941949e-12, 3.091704e-12, 
    3.653187e-12, 3.551436e-12, 2.802881e-12, 2.769493e-12, 3.051551e-12, 
    3.407434e-12, 4.075289e-12, 3.428076e-12, 2.450766e-12, 2.419746e-12, 
    2.465355e-12, 2.553053e-12, 2.773431e-12, 3.681124e-12, 6.388925e-12, 
    8.210673e-12, 7.715532e-12, 7.731316e-12, 6.457709e-12,
  1.492365e-11, 1.323065e-11, 1.286055e-11, 1.116254e-11, 9.258781e-12, 
    7.088434e-12, 6.456633e-12, 5.683355e-12, 6.41297e-12, 5.937219e-12, 
    5.615814e-12, 5.678389e-12, 5.597869e-12, 6.094498e-12, 5.73483e-12, 
    5.761928e-12, 8.72837e-12, 1.308647e-11, 1.099981e-11, 7.640041e-12, 
    9.367948e-12, 1.35223e-11, 1.487225e-11, 1.468746e-11, 1.25407e-11, 
    1.637171e-11, 1.522646e-11, 1.33011e-11, 1.440043e-11,
  5.143665e-11, 4.956928e-11, 5.075044e-11, 5.382945e-11, 5.394345e-11, 
    5.800401e-11, 5.297567e-11, 4.952759e-11, 4.793345e-11, 4.511085e-11, 
    4.340281e-11, 4.381727e-11, 4.687076e-11, 4.684704e-11, 4.847367e-11, 
    5.881539e-11, 6.115442e-11, 5.88437e-11, 5.594339e-11, 6.066733e-11, 
    6.786795e-11, 6.650783e-11, 6.998535e-11, 6.783687e-11, 6.777237e-11, 
    6.008791e-11, 5.510802e-11, 5.453418e-11, 5.152875e-11,
  4.277172e-10, 4.196186e-10, 4.372976e-10, 4.332273e-10, 4.299395e-10, 
    4.325865e-10, 4.341957e-10, 4.164256e-10, 4.22558e-10, 4.160669e-10, 
    4.133267e-10, 4.010813e-10, 4.001334e-10, 4.031616e-10, 4.032753e-10, 
    3.936536e-10, 3.88121e-10, 3.859652e-10, 4.083514e-10, 4.146528e-10, 
    4.303831e-10, 4.406416e-10, 4.421693e-10, 4.452841e-10, 4.28933e-10, 
    4.26332e-10, 4.336863e-10, 4.427121e-10, 4.390427e-10,
  8.44184e-10, 8.306493e-10, 8.361745e-10, 8.399375e-10, 8.631401e-10, 
    8.907983e-10, 8.759557e-10, 8.372391e-10, 8.106669e-10, 7.838505e-10, 
    7.620813e-10, 7.365344e-10, 7.392489e-10, 7.195393e-10, 7.19566e-10, 
    7.345238e-10, 7.742146e-10, 7.95723e-10, 8.200153e-10, 8.40419e-10, 
    8.525258e-10, 8.794926e-10, 8.708976e-10, 8.922619e-10, 8.958096e-10, 
    9.08111e-10, 8.844523e-10, 8.776954e-10, 8.617841e-10,
  8.227403e-10, 7.817755e-10, 7.638509e-10, 7.4271e-10, 7.626645e-10, 
    7.878233e-10, 8.118954e-10, 7.954721e-10, 8.175796e-10, 8.245811e-10, 
    8.114673e-10, 8.334446e-10, 8.144539e-10, 8.208637e-10, 8.083203e-10, 
    8.010889e-10, 8.114848e-10, 8.379274e-10, 7.919834e-10, 8.093504e-10, 
    8.571128e-10, 8.69968e-10, 8.699812e-10, 8.407059e-10, 8.625303e-10, 
    9.13394e-10, 8.794848e-10, 8.898772e-10, 8.505563e-10,
  3.70834e-10, 3.70409e-10, 3.744093e-10, 3.844639e-10, 4.173748e-10, 
    4.106704e-10, 4.259348e-10, 4.691624e-10, 4.672615e-10, 4.627553e-10, 
    4.572706e-10, 4.530829e-10, 4.661472e-10, 4.84841e-10, 4.786124e-10, 
    4.724889e-10, 4.850525e-10, 4.778831e-10, 4.732935e-10, 4.776405e-10, 
    4.698946e-10, 4.804031e-10, 4.644142e-10, 4.777561e-10, 4.486318e-10, 
    4.201984e-10, 3.950051e-10, 3.888944e-10, 3.74535e-10,
  3.207905e-10, 3.146872e-10, 3.172045e-10, 3.250392e-10, 3.209591e-10, 
    3.149457e-10, 3.255569e-10, 3.219534e-10, 3.435033e-10, 3.676762e-10, 
    3.924953e-10, 3.755539e-10, 3.778362e-10, 3.690913e-10, 3.595114e-10, 
    3.617789e-10, 3.632324e-10, 3.694381e-10, 3.550767e-10, 3.518549e-10, 
    3.50686e-10, 3.452081e-10, 3.4443e-10, 3.406641e-10, 3.377421e-10, 
    3.227665e-10, 3.310615e-10, 3.350879e-10, 3.254974e-10,
  5.812742e-11, 5.621844e-11, 5.465369e-11, 5.24011e-11, 5.525044e-11, 
    5.635327e-11, 5.736463e-11, 5.280655e-11, 4.924248e-11, 5.155519e-11, 
    6.08778e-11, 7.187038e-11, 7.950254e-11, 7.291224e-11, 7.992274e-11, 
    7.949523e-11, 7.046273e-11, 7.200735e-11, 6.750348e-11, 6.786323e-11, 
    7.64105e-11, 6.826789e-11, 6.621791e-11, 6.093497e-11, 5.963178e-11, 
    5.87702e-11, 6.053728e-11, 5.865252e-11, 5.859762e-11,
  1.400487e-11, 1.284302e-11, 1.195821e-11, 9.766854e-12, 9.28987e-12, 
    9.895576e-12, 9.451333e-12, 7.390185e-12, 7.955238e-12, 1.227578e-11, 
    9.788571e-12, 1.806767e-11, 6.767148e-12, 6.007278e-12, 7.195877e-12, 
    6.102163e-12, 4.852069e-12, 5.407868e-12, 4.876159e-12, 5.166968e-12, 
    6.830882e-12, 8.586885e-12, 1.01107e-11, 9.887743e-12, 1.25643e-11, 
    1.553803e-11, 1.910915e-11, 1.412929e-11, 1.371242e-11,
  2.336665e-12, 9.844267e-13, 1.304696e-12, 2.557369e-12, 4.139916e-12, 
    3.799345e-12, 4.511713e-12, 3.565324e-12, 2.660673e-12, 3.525971e-12, 
    4.896668e-12, 6.117633e-12, 7.388009e-12, 4.364852e-12, 2.972254e-12, 
    2.265878e-12, 2.194299e-12, 2.702723e-12, 2.797009e-12, 3.13025e-12, 
    2.791663e-12, 2.358525e-12, 2.448855e-12, 1.521325e-12, 1.711789e-12, 
    2.163862e-12, 4.050002e-12, 4.379743e-12, 3.171725e-12,
  6.186857e-13, 6.145067e-13, 5.401454e-13, 4.913732e-13, 4.63488e-13, 
    7.076279e-13, 1.088368e-12, 2.382264e-12, 2.335672e-12, 2.128632e-12, 
    2.257714e-12, 3.075637e-12, 5.233828e-12, 4.855034e-12, 3.911101e-12, 
    2.843299e-12, 2.606044e-12, 2.750765e-12, 2.643023e-12, 2.521332e-12, 
    2.4465e-12, 2.255445e-12, 2.531616e-12, 2.332639e-12, 2.586207e-12, 
    9.000105e-13, 8.584484e-13, 8.717838e-13, 6.431488e-13,
  1.577411e-13, 1.374694e-13, 1.260857e-13, 1.284456e-13, 1.610564e-13, 
    1.227553e-13, 1.560085e-13, 3.554288e-13, 1.019115e-12, 8.870821e-13, 
    1.120028e-12, 1.409701e-12, 2.074805e-12, 1.950479e-12, 1.967925e-12, 
    1.711266e-12, 1.59628e-12, 1.583582e-12, 1.765783e-12, 1.78198e-12, 
    1.760351e-12, 1.305085e-12, 1.318949e-12, 1.861187e-12, 4.769933e-13, 
    1.533161e-13, 1.460592e-13, 1.549264e-13, 1.630936e-13,
  6.008956e-14, 4.914627e-14, 3.363447e-14, 2.385075e-14, 2.62202e-14, 
    3.270473e-14, 4.010957e-14, 4.986277e-14, 9.031912e-14, 3.082481e-13, 
    4.322561e-13, 6.129064e-13, 8.252733e-13, 1.002581e-12, 1.114572e-12, 
    1.104672e-12, 1.069093e-12, 1.112911e-12, 1.172511e-12, 1.04269e-12, 
    9.86254e-13, 1.197981e-12, 7.716786e-13, 3.931833e-13, 3.134075e-13, 
    1.164762e-13, 8.119547e-14, 7.624158e-14, 6.592052e-14,
  5.917032e-14, 5.917032e-14, 5.917032e-14, 5.917032e-14, 5.917032e-14, 
    5.917032e-14, 5.917032e-14, 6.156307e-14, 6.156307e-14, 6.156307e-14, 
    6.156307e-14, 6.156307e-14, 6.156307e-14, 6.156307e-14, 6.361631e-14, 
    6.361631e-14, 6.361631e-14, 6.361631e-14, 6.361631e-14, 6.361631e-14, 
    6.361631e-14, 6.03476e-14, 6.03476e-14, 6.03476e-14, 6.03476e-14, 
    6.03476e-14, 6.03476e-14, 6.03476e-14, 5.917032e-14,
  3.814151e-14, 4.551538e-14, 5.634894e-14, 6.101387e-14, 6.366232e-14, 
    6.036607e-14, 7.759127e-14, 1.013419e-13, 1.298459e-13, 1.356434e-13, 
    1.324395e-13, 1.295364e-13, 1.316302e-13, 1.383725e-13, 1.464572e-13, 
    1.581142e-13, 1.690836e-13, 1.733244e-13, 1.566534e-13, 1.333355e-13, 
    1.172657e-13, 1.004317e-13, 7.430721e-14, 4.948534e-14, 3.956068e-14, 
    3.537782e-14, 3.422939e-14, 3.49479e-14, 3.815046e-14,
  5.66103e-13, 4.418419e-13, 5.026049e-13, 5.402492e-13, 4.445987e-13, 
    4.442284e-13, 5.101269e-13, 5.820214e-13, 5.684553e-13, 5.932019e-13, 
    6.041948e-13, 6.392032e-13, 7.007884e-13, 7.634954e-13, 9.198713e-13, 
    1.102698e-12, 1.096608e-12, 9.020081e-13, 6.315775e-13, 4.824887e-13, 
    4.637068e-13, 3.413681e-13, 3.712048e-13, 4.470246e-13, 4.25581e-13, 
    4.319589e-13, 4.281906e-13, 8.902256e-13, 7.666075e-13,
  3.433863e-12, 4.053249e-12, 4.038847e-12, 4.24527e-12, 4.261059e-12, 
    4.458771e-12, 4.980855e-12, 4.28633e-12, 3.193163e-12, 2.599628e-12, 
    2.667496e-12, 3.350491e-12, 4.285814e-12, 5.317675e-12, 5.928745e-12, 
    6.62686e-12, 7.646406e-12, 7.973384e-12, 7.339381e-12, 6.53591e-12, 
    5.831481e-12, 3.714759e-12, 3.045975e-12, 2.946642e-12, 3.484878e-12, 
    4.105756e-12, 3.06931e-12, 3.060711e-12, 3.122994e-12,
  1.435672e-11, 1.345237e-11, 1.378219e-11, 1.505199e-11, 1.364435e-11, 
    1.478301e-11, 1.478688e-11, 1.290627e-11, 1.063311e-11, 9.207708e-12, 
    9.615931e-12, 9.666717e-12, 7.693452e-12, 7.699864e-12, 8.275491e-12, 
    8.700558e-12, 1.083885e-11, 9.264873e-12, 6.753479e-12, 6.454738e-12, 
    6.652914e-12, 7.07954e-12, 7.572249e-12, 9.93754e-12, 1.387524e-11, 
    1.730775e-11, 2.055477e-11, 1.808285e-11, 1.516165e-11,
  4.534605e-11, 4.411045e-11, 3.358758e-11, 2.968824e-11, 2.488344e-11, 
    2.04401e-11, 1.949848e-11, 1.572868e-11, 1.70711e-11, 1.827997e-11, 
    1.836646e-11, 1.705406e-11, 1.498999e-11, 1.523881e-11, 1.520281e-11, 
    1.578494e-11, 4.302031e-11, 4.553608e-11, 4.481704e-11, 3.078681e-11, 
    3.597517e-11, 4.06182e-11, 4.012903e-11, 3.737242e-11, 3.532625e-11, 
    4.733532e-11, 3.997375e-11, 3.935065e-11, 4.558205e-11,
  1.911878e-10, 1.924632e-10, 1.883094e-10, 1.82535e-10, 1.879299e-10, 
    1.854896e-10, 1.691067e-10, 1.593203e-10, 1.497509e-10, 1.433777e-10, 
    1.35215e-10, 1.377481e-10, 1.397227e-10, 1.473759e-10, 1.815041e-10, 
    2.015309e-10, 1.836871e-10, 1.764801e-10, 1.720101e-10, 1.758359e-10, 
    2.080546e-10, 2.27149e-10, 2.237919e-10, 2.534802e-10, 2.473353e-10, 
    2.194779e-10, 1.897414e-10, 1.864632e-10, 1.90584e-10,
  1.523878e-09, 1.495385e-09, 1.490332e-09, 1.448054e-09, 1.467145e-09, 
    1.490534e-09, 1.494686e-09, 1.491832e-09, 1.45993e-09, 1.47023e-09, 
    1.430792e-09, 1.409179e-09, 1.368584e-09, 1.388174e-09, 1.398347e-09, 
    1.371521e-09, 1.388004e-09, 1.407643e-09, 1.443369e-09, 1.503575e-09, 
    1.514488e-09, 1.511639e-09, 1.51484e-09, 1.504418e-09, 1.486716e-09, 
    1.467e-09, 1.463924e-09, 1.528118e-09, 1.546045e-09,
  3.062874e-09, 2.990804e-09, 2.94258e-09, 3.041842e-09, 3.210229e-09, 
    3.205345e-09, 3.213154e-09, 3.080094e-09, 2.96905e-09, 2.86963e-09, 
    2.856805e-09, 2.705958e-09, 2.56181e-09, 2.534245e-09, 2.523675e-09, 
    2.580794e-09, 2.59454e-09, 2.6945e-09, 2.816252e-09, 2.955579e-09, 
    3.150299e-09, 3.198973e-09, 3.153354e-09, 3.212205e-09, 3.216169e-09, 
    3.046518e-09, 3.130457e-09, 3.171561e-09, 3.197586e-09,
  3.022062e-09, 2.919079e-09, 2.864481e-09, 2.856236e-09, 2.836339e-09, 
    2.832878e-09, 2.884744e-09, 2.965425e-09, 2.942195e-09, 2.977645e-09, 
    3.018095e-09, 3.048879e-09, 3.101289e-09, 3.066163e-09, 3.088545e-09, 
    3.05771e-09, 3.06878e-09, 3.111705e-09, 3.159483e-09, 3.193355e-09, 
    3.212644e-09, 3.208278e-09, 3.185747e-09, 3.147409e-09, 3.140856e-09, 
    3.146138e-09, 3.255337e-09, 3.249926e-09, 3.123942e-09,
  1.425392e-09, 1.450131e-09, 1.440532e-09, 1.467541e-09, 1.494972e-09, 
    1.515983e-09, 1.606622e-09, 1.65148e-09, 1.665853e-09, 1.645191e-09, 
    1.663748e-09, 1.660765e-09, 1.649713e-09, 1.663378e-09, 1.726012e-09, 
    1.778947e-09, 1.748773e-09, 1.811888e-09, 1.836609e-09, 1.850346e-09, 
    1.855069e-09, 1.816834e-09, 1.788345e-09, 1.75506e-09, 1.683885e-09, 
    1.620965e-09, 1.546008e-09, 1.471382e-09, 1.469125e-09,
  1.160142e-09, 1.156625e-09, 1.170351e-09, 1.132495e-09, 1.151038e-09, 
    1.132651e-09, 1.12581e-09, 1.136129e-09, 1.19842e-09, 1.228788e-09, 
    1.227948e-09, 1.170396e-09, 1.12685e-09, 1.111786e-09, 1.118953e-09, 
    1.149239e-09, 1.218981e-09, 1.253657e-09, 1.218677e-09, 1.148678e-09, 
    1.158163e-09, 1.10995e-09, 1.152565e-09, 1.141785e-09, 1.18355e-09, 
    1.203479e-09, 1.164443e-09, 1.117263e-09, 1.13343e-09,
  1.92031e-10, 1.947327e-10, 1.886019e-10, 1.918316e-10, 1.858229e-10, 
    2.058889e-10, 2.041146e-10, 1.934185e-10, 1.649301e-10, 1.89057e-10, 
    2.166253e-10, 2.278635e-10, 2.798289e-10, 2.447292e-10, 2.323847e-10, 
    2.399734e-10, 2.149305e-10, 2.096786e-10, 2.052553e-10, 2.062009e-10, 
    2.265159e-10, 2.13069e-10, 2.01526e-10, 2.12015e-10, 2.129788e-10, 
    2.032063e-10, 1.860758e-10, 1.980676e-10, 1.885559e-10,
  4.637613e-11, 3.568417e-11, 3.27589e-11, 2.800986e-11, 3.019658e-11, 
    3.216546e-11, 3.336909e-11, 2.009356e-11, 2.053607e-11, 3.481861e-11, 
    2.795379e-11, 8.458322e-11, 4.286141e-11, 2.164164e-11, 2.112551e-11, 
    1.918479e-11, 1.513903e-11, 1.6692e-11, 1.681495e-11, 2.100217e-11, 
    2.395543e-11, 2.623318e-11, 2.99649e-11, 2.691362e-11, 3.961955e-11, 
    4.690641e-11, 6.139163e-11, 5.039751e-11, 4.497401e-11,
  6.948698e-12, 4.063618e-12, 4.431984e-12, 9.299837e-12, 1.363394e-11, 
    1.038529e-11, 1.156971e-11, 1.205218e-11, 6.860728e-12, 8.662946e-12, 
    1.435188e-11, 1.712722e-11, 2.765897e-11, 1.38864e-11, 9.917286e-12, 
    6.150162e-12, 6.444457e-12, 8.377758e-12, 9.200686e-12, 9.935809e-12, 
    9.257246e-12, 8.19156e-12, 1.086584e-11, 7.414546e-12, 8.319964e-12, 
    7.956502e-12, 1.05929e-11, 1.340897e-11, 1.095405e-11,
  2.769653e-12, 2.818994e-12, 2.598739e-12, 2.207119e-12, 1.840516e-12, 
    1.859449e-12, 2.120114e-12, 5.10134e-12, 6.317728e-12, 5.145367e-12, 
    4.567254e-12, 8.353508e-12, 1.724847e-11, 1.302805e-11, 1.172228e-11, 
    8.887681e-12, 7.625169e-12, 9.100071e-12, 8.712392e-12, 9.086345e-12, 
    8.285854e-12, 7.47423e-12, 1.018522e-11, 9.107002e-12, 1.200876e-11, 
    4.9897e-12, 3.873847e-12, 3.902573e-12, 2.950048e-12,
  5.794246e-13, 5.597889e-13, 4.889311e-13, 4.428782e-13, 4.890814e-13, 
    5.315506e-13, 5.672111e-13, 6.632854e-13, 2.026544e-12, 2.259109e-12, 
    3.242689e-12, 3.788792e-12, 6.698639e-12, 6.606054e-12, 5.798043e-12, 
    5.491764e-12, 5.212256e-12, 5.642191e-12, 5.171662e-12, 5.969357e-12, 
    6.172366e-12, 4.892059e-12, 6.83352e-12, 9.799723e-12, 4.845375e-12, 
    6.03918e-13, 5.615115e-13, 5.964178e-13, 5.906543e-13,
  1.880761e-13, 1.563828e-13, 1.285416e-13, 9.681144e-14, 8.491198e-14, 
    9.505081e-14, 1.173824e-13, 1.445242e-13, 2.000842e-13, 5.504557e-13, 
    9.775452e-13, 1.32786e-12, 2.348034e-12, 3.611925e-12, 5.850328e-12, 
    5.739258e-12, 4.498252e-12, 3.972339e-12, 4.083476e-12, 4.41758e-12, 
    6.059163e-12, 9.146287e-12, 8.633352e-12, 3.071275e-12, 1.116304e-12, 
    5.705139e-13, 2.863359e-13, 2.516379e-13, 2.138004e-13,
  1.942057e-13, 1.942057e-13, 1.942057e-13, 1.942057e-13, 1.942057e-13, 
    1.942057e-13, 1.942057e-13, 1.941546e-13, 1.941546e-13, 1.941546e-13, 
    1.941546e-13, 1.941546e-13, 1.941546e-13, 1.941546e-13, 2.01842e-13, 
    2.01842e-13, 2.01842e-13, 2.01842e-13, 2.01842e-13, 2.01842e-13, 
    2.01842e-13, 2.013964e-13, 2.013964e-13, 2.013964e-13, 2.013964e-13, 
    2.013964e-13, 2.013964e-13, 2.013964e-13, 1.942057e-13,
  1.758452e-13, 1.729065e-13, 2.092253e-13, 2.437131e-13, 2.048088e-13, 
    2.130095e-13, 2.067976e-13, 2.891046e-13, 4.498696e-13, 5.169106e-13, 
    5.350272e-13, 5.335848e-13, 5.466786e-13, 5.577978e-13, 5.864527e-13, 
    6.728371e-13, 7.139098e-13, 6.847649e-13, 6.157917e-13, 5.25302e-13, 
    4.72364e-13, 3.97614e-13, 2.99572e-13, 2.05647e-13, 1.798301e-13, 
    1.688476e-13, 1.620577e-13, 1.65835e-13, 1.721449e-13,
  2.4505e-12, 1.631787e-12, 1.460944e-12, 1.594266e-12, 1.402467e-12, 
    1.449987e-12, 1.894951e-12, 2.131466e-12, 2.157986e-12, 1.981215e-12, 
    1.807931e-12, 2.051778e-12, 2.38916e-12, 2.833003e-12, 3.775556e-12, 
    4.643361e-12, 4.755952e-12, 3.510091e-12, 2.509065e-12, 2.075233e-12, 
    1.944211e-12, 1.269464e-12, 1.712431e-12, 2.109597e-12, 1.991371e-12, 
    1.844548e-12, 1.724206e-12, 2.89612e-12, 3.140906e-12,
  1.350035e-11, 1.280941e-11, 1.253122e-11, 1.192722e-11, 1.368128e-11, 
    1.726879e-11, 1.819933e-11, 1.564983e-11, 1.200688e-11, 9.383988e-12, 
    8.964783e-12, 1.03955e-11, 1.268624e-11, 1.59985e-11, 1.852975e-11, 
    2.075532e-11, 2.467166e-11, 2.436898e-11, 2.281123e-11, 1.958025e-11, 
    1.687807e-11, 1.264216e-11, 1.063844e-11, 9.545147e-12, 1.161006e-11, 
    1.477367e-11, 1.178064e-11, 1.094009e-11, 1.074947e-11,
  5.893695e-11, 5.591169e-11, 4.750653e-11, 4.623419e-11, 5.18728e-11, 
    5.73042e-11, 5.243514e-11, 4.535829e-11, 3.794935e-11, 3.343568e-11, 
    3.344677e-11, 3.16078e-11, 2.691486e-11, 2.646908e-11, 3.110368e-11, 
    2.965856e-11, 2.973665e-11, 3.181994e-11, 2.388753e-11, 2.293422e-11, 
    2.392288e-11, 2.50505e-11, 2.685225e-11, 3.289721e-11, 4.529122e-11, 
    5.212553e-11, 5.726226e-11, 5.803496e-11, 6.261353e-11,
  1.56913e-10, 1.563044e-10, 1.078015e-10, 1.085894e-10, 9.331231e-11, 
    7.444247e-11, 6.825913e-11, 5.262185e-11, 5.587328e-11, 6.512831e-11, 
    6.402579e-11, 5.933304e-11, 5.212078e-11, 4.546458e-11, 4.444029e-11, 
    5.871165e-11, 1.563839e-10, 1.513616e-10, 1.375609e-10, 1.181054e-10, 
    1.320867e-10, 1.289429e-10, 1.332482e-10, 1.375312e-10, 1.436549e-10, 
    1.454047e-10, 1.2019e-10, 1.308346e-10, 1.426616e-10,
  7.349885e-10, 7.805959e-10, 7.648744e-10, 6.839531e-10, 6.613251e-10, 
    6.646307e-10, 6.399026e-10, 5.952192e-10, 5.673786e-10, 5.456868e-10, 
    5.165776e-10, 5.003492e-10, 5.30356e-10, 5.77522e-10, 7.512057e-10, 
    6.402386e-10, 6.621026e-10, 6.66274e-10, 6.907059e-10, 7.118073e-10, 
    7.838597e-10, 8.016767e-10, 8.701335e-10, 1.003193e-09, 9.556005e-10, 
    8.86792e-10, 7.215005e-10, 6.997992e-10, 7.126213e-10,
  5.438717e-09, 5.334039e-09, 5.344595e-09, 5.410794e-09, 5.600136e-09, 
    5.436978e-09, 5.326188e-09, 5.391166e-09, 5.474399e-09, 5.282393e-09, 
    5.244857e-09, 5.127125e-09, 5.106267e-09, 5.153558e-09, 4.936147e-09, 
    4.818796e-09, 4.867148e-09, 4.940804e-09, 5.163492e-09, 5.330989e-09, 
    5.511793e-09, 5.508233e-09, 5.411535e-09, 5.524947e-09, 5.470097e-09, 
    5.530722e-09, 5.48422e-09, 5.610376e-09, 5.654465e-09,
  1.143585e-08, 1.124245e-08, 1.101094e-08, 1.125869e-08, 1.148749e-08, 
    1.187436e-08, 1.198084e-08, 1.162941e-08, 1.08999e-08, 1.046894e-08, 
    1.009726e-08, 9.975428e-09, 9.661542e-09, 9.523068e-09, 9.419829e-09, 
    9.349085e-09, 9.670122e-09, 9.791361e-09, 1.024898e-08, 1.065293e-08, 
    1.162891e-08, 1.200246e-08, 1.196427e-08, 1.178798e-08, 1.18266e-08, 
    1.203914e-08, 1.208731e-08, 1.178679e-08, 1.152166e-08,
  1.195156e-08, 1.144574e-08, 1.128327e-08, 1.126694e-08, 1.128052e-08, 
    1.08837e-08, 1.114463e-08, 1.149255e-08, 1.132897e-08, 1.12654e-08, 
    1.133056e-08, 1.176076e-08, 1.17283e-08, 1.188077e-08, 1.196982e-08, 
    1.189318e-08, 1.191549e-08, 1.171045e-08, 1.19824e-08, 1.197487e-08, 
    1.189956e-08, 1.19244e-08, 1.191151e-08, 1.149047e-08, 1.128579e-08, 
    1.139302e-08, 1.15331e-08, 1.206645e-08, 1.213464e-08,
  6.018321e-09, 5.77981e-09, 5.766452e-09, 5.843991e-09, 5.830386e-09, 
    5.888493e-09, 5.880593e-09, 6.004774e-09, 6.083254e-09, 5.958135e-09, 
    5.990808e-09, 6.027335e-09, 6.195555e-09, 6.40669e-09, 6.633037e-09, 
    6.796074e-09, 6.85012e-09, 6.969821e-09, 7.120603e-09, 7.012405e-09, 
    6.890942e-09, 6.925562e-09, 6.912463e-09, 6.838748e-09, 6.495707e-09, 
    6.086332e-09, 5.921045e-09, 5.82893e-09, 5.820438e-09,
  4.084544e-09, 4.078966e-09, 4.077133e-09, 4.119382e-09, 4.013303e-09, 
    3.983537e-09, 3.926468e-09, 3.995753e-09, 4.250106e-09, 4.175909e-09, 
    4.290797e-09, 4.174828e-09, 4.1858e-09, 4.069642e-09, 4.153936e-09, 
    4.258947e-09, 4.367193e-09, 4.368394e-09, 4.24049e-09, 4.15768e-09, 
    4.19791e-09, 4.185586e-09, 4.177197e-09, 4.098077e-09, 4.000131e-09, 
    3.951543e-09, 4.086571e-09, 4.089959e-09, 4.052418e-09,
  7.194602e-10, 7.386405e-10, 6.71702e-10, 6.791301e-10, 6.410162e-10, 
    7.340951e-10, 6.725817e-10, 6.262021e-10, 6.254062e-10, 7.057169e-10, 
    7.619793e-10, 7.814202e-10, 9.473299e-10, 8.001666e-10, 7.398949e-10, 
    7.58163e-10, 7.072832e-10, 6.997887e-10, 7.457872e-10, 7.394566e-10, 
    7.556277e-10, 7.062169e-10, 7.055306e-10, 8.038444e-10, 7.788743e-10, 
    7.6544e-10, 6.97561e-10, 6.96665e-10, 6.926794e-10,
  1.53867e-10, 1.082906e-10, 1.110031e-10, 9.471677e-11, 1.098433e-10, 
    1.039061e-10, 1.34778e-10, 6.287498e-11, 6.361658e-11, 1.021358e-10, 
    1.067247e-10, 2.161636e-10, 2.182994e-10, 7.88376e-11, 6.608421e-11, 
    6.540154e-11, 5.576669e-11, 6.055392e-11, 6.44944e-11, 8.682018e-11, 
    9.07547e-11, 9.883008e-11, 1.077392e-10, 1.027457e-10, 1.119224e-10, 
    1.396882e-10, 2.002964e-10, 1.907572e-10, 1.569468e-10,
  2.884651e-11, 1.992286e-11, 2.077668e-11, 3.236469e-11, 5.007995e-11, 
    3.604607e-11, 3.373368e-11, 4.609303e-11, 2.132259e-11, 2.309874e-11, 
    4.723488e-11, 5.820591e-11, 1.146062e-10, 4.902995e-11, 3.4185e-11, 
    2.047238e-11, 2.257405e-11, 3.076483e-11, 3.918403e-11, 3.567038e-11, 
    4.012937e-11, 3.244284e-11, 5.421758e-11, 3.909657e-11, 3.422127e-11, 
    3.195439e-11, 2.957973e-11, 3.927436e-11, 3.781446e-11,
  1.359036e-11, 1.464976e-11, 1.1291e-11, 8.755343e-12, 7.646872e-12, 
    7.029379e-12, 6.659604e-12, 1.34666e-11, 2.003464e-11, 1.713321e-11, 
    1.093673e-11, 2.397983e-11, 6.705653e-11, 3.576635e-11, 3.188174e-11, 
    2.911358e-11, 2.813374e-11, 3.11335e-11, 3.53056e-11, 3.936231e-11, 
    4.15093e-11, 3.375177e-11, 3.639988e-11, 4.277539e-11, 3.25351e-11, 
    3.677553e-11, 2.021343e-11, 2.167003e-11, 1.499785e-11,
  2.982712e-12, 2.547947e-12, 2.478941e-12, 2.211692e-12, 2.205449e-12, 
    2.457652e-12, 2.307728e-12, 2.5279e-12, 5.322417e-12, 8.130472e-12, 
    1.06736e-11, 1.359084e-11, 3.941575e-11, 2.691942e-11, 1.998726e-11, 
    1.989931e-11, 2.062295e-11, 2.764142e-11, 2.471526e-11, 2.567945e-11, 
    2.338524e-11, 2.112958e-11, 2.810372e-11, 4.491926e-11, 2.679709e-11, 
    2.895909e-12, 2.758955e-12, 3.338208e-12, 3.181835e-12,
  8.037118e-13, 6.251417e-13, 4.731035e-13, 4.091975e-13, 3.417937e-13, 
    2.987959e-13, 3.631113e-13, 5.106366e-13, 6.899678e-13, 1.202892e-12, 
    2.393705e-12, 5.831803e-12, 2.072816e-11, 3.265328e-11, 3.671987e-11, 
    2.75699e-11, 1.871093e-11, 1.604129e-11, 1.571734e-11, 1.723445e-11, 
    2.573676e-11, 3.718223e-11, 4.608854e-11, 3.086944e-11, 7.009089e-12, 
    2.139135e-12, 1.079698e-12, 9.491605e-13, 8.544831e-13,
  8.420157e-13, 8.420157e-13, 8.420157e-13, 8.420157e-13, 8.420157e-13, 
    8.420157e-13, 8.420157e-13, 8.397193e-13, 8.397193e-13, 8.397193e-13, 
    8.397193e-13, 8.397193e-13, 8.397193e-13, 8.397193e-13, 8.755359e-13, 
    8.755359e-13, 8.755359e-13, 8.755359e-13, 8.755359e-13, 8.755359e-13, 
    8.755359e-13, 8.630618e-13, 8.630618e-13, 8.630618e-13, 8.630618e-13, 
    8.630618e-13, 8.630618e-13, 8.630618e-13, 8.420157e-13,
  6.553611e-13, 6.849211e-13, 7.20393e-13, 8.86194e-13, 1.029096e-12, 
    8.533131e-13, 7.944347e-13, 1.102182e-12, 1.587667e-12, 2.138287e-12, 
    2.182723e-12, 2.138647e-12, 2.173124e-12, 2.244074e-12, 2.419293e-12, 
    2.703694e-12, 2.753117e-12, 2.64128e-12, 2.380171e-12, 2.071123e-12, 
    1.966038e-12, 1.610701e-12, 1.246266e-12, 9.173375e-13, 7.562218e-13, 
    6.767285e-13, 6.579085e-13, 6.663975e-13, 6.645006e-13,
  1.628506e-11, 1.052249e-11, 7.883649e-12, 6.147528e-12, 6.532227e-12, 
    7.061571e-12, 8.826784e-12, 9.781909e-12, 8.160058e-12, 6.621865e-12, 
    5.803215e-12, 6.427449e-12, 8.164493e-12, 1.033566e-11, 1.398474e-11, 
    1.73429e-11, 1.880311e-11, 1.432897e-11, 9.960267e-12, 8.779463e-12, 
    7.81727e-12, 5.177673e-12, 6.643669e-12, 8.282808e-12, 7.669287e-12, 
    7.379245e-12, 6.199839e-12, 1.041374e-11, 1.863974e-11,
  4.6495e-11, 4.316801e-11, 4.222657e-11, 4.097693e-11, 5.04659e-11, 
    6.377057e-11, 6.295481e-11, 5.546157e-11, 4.573706e-11, 3.371423e-11, 
    3.102146e-11, 3.249101e-11, 4.046215e-11, 5.167703e-11, 6.460575e-11, 
    7.254618e-11, 8.280897e-11, 8.25934e-11, 7.321262e-11, 6.702638e-11, 
    5.274764e-11, 4.133711e-11, 3.829538e-11, 3.435231e-11, 3.93807e-11, 
    5.771211e-11, 4.388524e-11, 3.670293e-11, 3.562721e-11,
  2.026678e-10, 1.781058e-10, 1.361492e-10, 1.315283e-10, 1.635052e-10, 
    1.73001e-10, 1.696974e-10, 1.438162e-10, 1.246757e-10, 1.26004e-10, 
    1.281871e-10, 1.145395e-10, 1.020992e-10, 1.079186e-10, 1.238873e-10, 
    1.198916e-10, 1.175319e-10, 1.19085e-10, 9.700066e-11, 8.996809e-11, 
    8.823884e-11, 9.129731e-11, 1.035443e-10, 1.25291e-10, 1.691478e-10, 
    1.706297e-10, 1.7008e-10, 2.13272e-10, 2.366109e-10,
  5.055454e-10, 4.888654e-10, 4.094301e-10, 4.61868e-10, 3.638387e-10, 
    2.615712e-10, 2.271953e-10, 2.012564e-10, 2.147787e-10, 2.52969e-10, 
    2.621768e-10, 2.297114e-10, 1.943623e-10, 1.685634e-10, 1.490331e-10, 
    2.454295e-10, 4.308117e-10, 4.816537e-10, 4.421094e-10, 4.308777e-10, 
    4.492922e-10, 4.441829e-10, 5.581336e-10, 5.367188e-10, 6.194996e-10, 
    5.10496e-10, 4.574799e-10, 4.297038e-10, 4.57674e-10,
  3.316515e-09, 3.317021e-09, 2.700181e-09, 2.411369e-09, 2.434281e-09, 
    2.446371e-09, 2.388454e-09, 2.304232e-09, 2.230921e-09, 2.121636e-09, 
    2.011993e-09, 2.045018e-09, 2.104665e-09, 2.39905e-09, 2.702e-09, 
    2.58916e-09, 2.720884e-09, 2.79622e-09, 2.99696e-09, 2.955726e-09, 
    3.15125e-09, 3.119872e-09, 3.623184e-09, 3.550073e-09, 3.656961e-09, 
    3.26725e-09, 2.801947e-09, 2.775844e-09, 2.95623e-09,
  2.072793e-08, 2.043436e-08, 2.005042e-08, 1.969458e-08, 2.0101e-08, 
    1.99024e-08, 1.99453e-08, 2.00838e-08, 2.003499e-08, 1.899594e-08, 
    1.946108e-08, 1.877162e-08, 1.831425e-08, 1.82832e-08, 1.815809e-08, 
    1.817882e-08, 1.832464e-08, 1.919557e-08, 1.926064e-08, 1.941527e-08, 
    1.943825e-08, 2.039146e-08, 2.072248e-08, 2.055404e-08, 2.046252e-08, 
    2.037718e-08, 2.062167e-08, 2.176195e-08, 2.147124e-08,
  4.570375e-08, 4.298544e-08, 4.414905e-08, 4.602275e-08, 4.799733e-08, 
    4.590562e-08, 4.508401e-08, 4.539028e-08, 4.104866e-08, 4.014858e-08, 
    3.985729e-08, 3.710056e-08, 3.672871e-08, 3.682928e-08, 3.537219e-08, 
    3.590803e-08, 3.522921e-08, 3.654992e-08, 3.846055e-08, 4.163607e-08, 
    4.372486e-08, 4.42326e-08, 4.580223e-08, 4.377639e-08, 4.484816e-08, 
    4.580922e-08, 4.546414e-08, 4.709612e-08, 4.823076e-08,
  4.459493e-08, 4.327429e-08, 4.160919e-08, 4.241586e-08, 3.990411e-08, 
    3.99055e-08, 4.05699e-08, 4.264082e-08, 4.225734e-08, 4.291777e-08, 
    4.525107e-08, 4.516562e-08, 4.471246e-08, 4.493933e-08, 4.481395e-08, 
    4.31525e-08, 4.292168e-08, 4.326456e-08, 4.380571e-08, 4.329944e-08, 
    4.17431e-08, 4.32573e-08, 4.399441e-08, 4.226136e-08, 4.10821e-08, 
    4.02167e-08, 4.098463e-08, 4.140525e-08, 4.450808e-08,
  2.374594e-08, 2.327088e-08, 2.353866e-08, 2.410599e-08, 2.402814e-08, 
    2.307611e-08, 2.306533e-08, 2.27537e-08, 2.325563e-08, 2.319952e-08, 
    2.340398e-08, 2.3381e-08, 2.44068e-08, 2.514734e-08, 2.606759e-08, 
    2.692019e-08, 2.767657e-08, 2.810563e-08, 2.845358e-08, 2.830755e-08, 
    2.865112e-08, 2.737109e-08, 2.66828e-08, 2.574627e-08, 2.501483e-08, 
    2.432336e-08, 2.414346e-08, 2.318118e-08, 2.375348e-08,
  1.545614e-08, 1.525819e-08, 1.484251e-08, 1.465405e-08, 1.474466e-08, 
    1.506249e-08, 1.480666e-08, 1.511784e-08, 1.572275e-08, 1.582834e-08, 
    1.587406e-08, 1.601345e-08, 1.54761e-08, 1.577194e-08, 1.600014e-08, 
    1.635738e-08, 1.676981e-08, 1.617021e-08, 1.56398e-08, 1.51969e-08, 
    1.533633e-08, 1.531585e-08, 1.534888e-08, 1.539074e-08, 1.574579e-08, 
    1.551599e-08, 1.531531e-08, 1.486246e-08, 1.513119e-08,
  2.467839e-09, 2.564819e-09, 2.361858e-09, 2.365526e-09, 2.276178e-09, 
    2.577283e-09, 2.296257e-09, 2.389428e-09, 2.372902e-09, 2.686618e-09, 
    2.93817e-09, 3.004506e-09, 3.470839e-09, 3.036723e-09, 2.843995e-09, 
    3.098891e-09, 2.949227e-09, 2.915315e-09, 3.002165e-09, 2.954342e-09, 
    2.617976e-09, 2.457765e-09, 2.535766e-09, 3.04472e-09, 3.11184e-09, 
    2.964697e-09, 2.624876e-09, 2.668024e-09, 2.503954e-09,
  4.86213e-10, 3.436035e-10, 3.968929e-10, 3.257351e-10, 3.684678e-10, 
    3.44378e-10, 4.924957e-10, 2.262349e-10, 2.205205e-10, 3.251776e-10, 
    4.521111e-10, 6.687133e-10, 8.163377e-10, 4.006184e-10, 2.704251e-10, 
    2.237643e-10, 2.257057e-10, 2.553589e-10, 2.679287e-10, 3.531551e-10, 
    3.556092e-10, 3.790656e-10, 4.417746e-10, 4.237794e-10, 3.61533e-10, 
    4.882225e-10, 6.04717e-10, 6.207478e-10, 5.443656e-10,
  1.361019e-10, 9.931866e-11, 8.865723e-11, 1.064581e-10, 1.677109e-10, 
    1.547512e-10, 1.198345e-10, 1.813146e-10, 8.093465e-11, 6.580163e-11, 
    1.286725e-10, 2.680643e-10, 4.928583e-10, 2.06075e-10, 1.17061e-10, 
    7.618719e-11, 9.219921e-11, 1.13528e-10, 1.500928e-10, 1.258937e-10, 
    1.564527e-10, 1.322878e-10, 1.83533e-10, 1.594829e-10, 1.490535e-10, 
    1.411106e-10, 1.184397e-10, 1.357437e-10, 1.454259e-10,
  6.262858e-11, 5.670274e-11, 5.597818e-11, 4.438657e-11, 3.543338e-11, 
    3.318323e-11, 3.388639e-11, 4.389635e-11, 6.660113e-11, 6.885708e-11, 
    4.001335e-11, 7.710174e-11, 3.835593e-10, 1.366289e-10, 1.043555e-10, 
    9.70947e-11, 1.142528e-10, 1.069453e-10, 1.48119e-10, 1.794518e-10, 
    2.041515e-10, 1.599743e-10, 1.307774e-10, 1.462947e-10, 1.491234e-10, 
    1.095448e-10, 1.109535e-10, 9.412295e-11, 8.103427e-11,
  1.51403e-11, 1.257706e-11, 1.258149e-11, 1.13973e-11, 9.740546e-12, 
    9.319819e-12, 9.369177e-12, 9.911029e-12, 1.426448e-11, 2.662007e-11, 
    3.259561e-11, 5.111343e-11, 2.25398e-10, 1.389535e-10, 8.306032e-11, 
    8.0278e-11, 9.322561e-11, 1.54963e-10, 1.414991e-10, 1.433625e-10, 
    1.299167e-10, 9.743424e-11, 9.613991e-11, 1.572198e-10, 1.133716e-10, 
    2.408542e-11, 1.609107e-11, 1.865087e-11, 1.640495e-11,
  3.330078e-12, 2.584504e-12, 1.518241e-12, 1.466582e-12, 1.511332e-12, 
    1.178789e-12, 1.278014e-12, 1.663787e-12, 2.222941e-12, 3.083459e-12, 
    6.194783e-12, 3.567134e-11, 1.065048e-10, 1.498536e-10, 1.384498e-10, 
    1.126179e-10, 9.521945e-11, 8.5058e-11, 7.415642e-11, 6.488794e-11, 
    8.969963e-11, 1.170276e-10, 1.419496e-10, 1.42043e-10, 5.10872e-11, 
    6.203353e-12, 3.354552e-12, 3.371486e-12, 3.520438e-12,
  3.676693e-12, 3.676693e-12, 3.676693e-12, 3.676693e-12, 3.676693e-12, 
    3.676693e-12, 3.676693e-12, 3.746194e-12, 3.746194e-12, 3.746194e-12, 
    3.746194e-12, 3.746194e-12, 3.746194e-12, 3.746194e-12, 3.76394e-12, 
    3.76394e-12, 3.76394e-12, 3.76394e-12, 3.76394e-12, 3.76394e-12, 
    3.76394e-12, 3.631839e-12, 3.631839e-12, 3.631839e-12, 3.631839e-12, 
    3.631839e-12, 3.631839e-12, 3.631839e-12, 3.676693e-12,
  3.377821e-12, 3.22574e-12, 3.216524e-12, 3.122472e-12, 3.79542e-12, 
    4.286585e-12, 3.567903e-12, 3.214454e-12, 4.600643e-12, 7.099779e-12, 
    8.023826e-12, 8.375715e-12, 8.910624e-12, 9.26011e-12, 9.853724e-12, 
    1.082038e-11, 1.172114e-11, 1.146891e-11, 9.600736e-12, 8.002547e-12, 
    7.592419e-12, 6.91413e-12, 5.578319e-12, 4.303883e-12, 3.720069e-12, 
    3.48828e-12, 3.389959e-12, 3.406254e-12, 3.397672e-12,
  5.262788e-11, 4.092758e-11, 2.622542e-11, 2.33427e-11, 2.892694e-11, 
    3.192336e-11, 3.160079e-11, 3.391835e-11, 2.76873e-11, 2.024075e-11, 
    1.834468e-11, 2.149476e-11, 2.731022e-11, 3.561627e-11, 4.819212e-11, 
    5.935002e-11, 6.715163e-11, 5.967984e-11, 4.101723e-11, 3.620524e-11, 
    3.225951e-11, 2.220446e-11, 2.432748e-11, 3.126885e-11, 2.976955e-11, 
    2.997534e-11, 2.517428e-11, 2.752218e-11, 5.181211e-11,
  1.483365e-10, 1.412262e-10, 1.366332e-10, 1.453062e-10, 1.835706e-10, 
    2.284798e-10, 2.201775e-10, 1.903501e-10, 1.691794e-10, 1.229264e-10, 
    1.045137e-10, 1.078781e-10, 1.321531e-10, 1.694831e-10, 2.241078e-10, 
    2.530852e-10, 2.724267e-10, 2.739547e-10, 2.38885e-10, 2.208432e-10, 
    1.873308e-10, 1.476023e-10, 1.202369e-10, 1.274759e-10, 1.376358e-10, 
    1.980669e-10, 1.734133e-10, 1.350999e-10, 1.523909e-10,
  6.286491e-10, 5.38033e-10, 4.694997e-10, 4.431693e-10, 5.024046e-10, 
    5.045977e-10, 5.715618e-10, 5.042607e-10, 4.260122e-10, 4.232256e-10, 
    4.409463e-10, 4.081244e-10, 3.949613e-10, 5.026735e-10, 4.483833e-10, 
    4.329112e-10, 4.760164e-10, 4.98186e-10, 3.852848e-10, 3.165852e-10, 
    2.980903e-10, 3.204382e-10, 3.679641e-10, 4.775116e-10, 6.860936e-10, 
    5.90453e-10, 5.471458e-10, 6.506033e-10, 6.888078e-10,
  1.708894e-09, 1.536859e-09, 1.758344e-09, 1.741147e-09, 1.407312e-09, 
    9.352322e-10, 7.900327e-10, 7.535756e-10, 8.270161e-10, 1.018036e-09, 
    1.012913e-09, 9.371481e-10, 7.725171e-10, 6.86711e-10, 5.665701e-10, 
    7.811791e-10, 1.175976e-09, 1.431353e-09, 1.496239e-09, 1.583897e-09, 
    1.625465e-09, 1.69949e-09, 2.14685e-09, 2.20318e-09, 2.337174e-09, 
    1.752237e-09, 1.592316e-09, 1.510139e-09, 1.547266e-09,
  1.276888e-08, 1.140725e-08, 1.027366e-08, 9.040038e-09, 9.222997e-09, 
    9.023948e-09, 9.932624e-09, 9.930322e-09, 9.58865e-09, 8.993962e-09, 
    8.625478e-09, 8.724482e-09, 9.102357e-09, 1.084053e-08, 1.041905e-08, 
    1.009648e-08, 1.090123e-08, 1.124288e-08, 1.169854e-08, 1.196332e-08, 
    1.202324e-08, 1.305937e-08, 1.435387e-08, 1.317411e-08, 1.319692e-08, 
    1.207721e-08, 1.03514e-08, 1.11311e-08, 1.194689e-08,
  7.961338e-08, 7.705933e-08, 7.766547e-08, 7.80451e-08, 7.624872e-08, 
    7.526444e-08, 7.477374e-08, 7.379544e-08, 7.273159e-08, 7.2256e-08, 
    7.261127e-08, 7.031463e-08, 6.976247e-08, 6.858008e-08, 6.751471e-08, 
    6.665471e-08, 6.754853e-08, 6.918739e-08, 7.316763e-08, 7.592654e-08, 
    7.859754e-08, 7.977182e-08, 7.870553e-08, 7.823175e-08, 7.762231e-08, 
    7.675347e-08, 7.889007e-08, 8.054924e-08, 8.146272e-08,
  1.816839e-07, 1.817518e-07, 1.736884e-07, 1.730962e-07, 1.809221e-07, 
    1.869851e-07, 1.817918e-07, 1.794425e-07, 1.690099e-07, 1.569783e-07, 
    1.494193e-07, 1.468786e-07, 1.401546e-07, 1.36914e-07, 1.285911e-07, 
    1.309164e-07, 1.323925e-07, 1.404277e-07, 1.468749e-07, 1.553644e-07, 
    1.690069e-07, 1.789727e-07, 1.751373e-07, 1.78013e-07, 1.763237e-07, 
    1.817973e-07, 1.800545e-07, 1.837806e-07, 1.800513e-07,
  1.553324e-07, 1.534192e-07, 1.481962e-07, 1.42296e-07, 1.435917e-07, 
    1.362825e-07, 1.466706e-07, 1.52378e-07, 1.534458e-07, 1.605065e-07, 
    1.714725e-07, 1.698285e-07, 1.714561e-07, 1.709204e-07, 1.691454e-07, 
    1.612092e-07, 1.642792e-07, 1.663936e-07, 1.613349e-07, 1.557273e-07, 
    1.448056e-07, 1.519761e-07, 1.531514e-07, 1.523085e-07, 1.509581e-07, 
    1.499639e-07, 1.44893e-07, 1.489929e-07, 1.506237e-07,
  9.869061e-08, 9.51712e-08, 9.84518e-08, 1.032162e-07, 9.866022e-08, 
    9.585597e-08, 9.163242e-08, 9.02793e-08, 9.352014e-08, 9.353246e-08, 
    9.483365e-08, 9.723926e-08, 9.950266e-08, 1.022636e-07, 1.064418e-07, 
    1.042065e-07, 1.060606e-07, 1.08137e-07, 1.099074e-07, 1.08425e-07, 
    1.096763e-07, 1.055546e-07, 1.035882e-07, 1.030709e-07, 9.876479e-08, 
    9.42024e-08, 9.532474e-08, 9.791425e-08, 9.800382e-08,
  5.471589e-08, 5.625258e-08, 5.520476e-08, 5.822796e-08, 5.594546e-08, 
    5.691577e-08, 5.587282e-08, 5.682453e-08, 6.108422e-08, 6.366798e-08, 
    6.495914e-08, 6.457228e-08, 6.457405e-08, 6.530107e-08, 6.175807e-08, 
    6.049304e-08, 6.001884e-08, 5.897683e-08, 5.842151e-08, 5.861786e-08, 
    5.826803e-08, 5.947475e-08, 5.810876e-08, 5.724025e-08, 5.642964e-08, 
    5.591692e-08, 5.76292e-08, 5.783062e-08, 5.630101e-08,
  9.111134e-09, 9.420307e-09, 8.975838e-09, 8.719872e-09, 8.352171e-09, 
    9.459607e-09, 8.908291e-09, 9.497189e-09, 1.049358e-08, 1.125911e-08, 
    1.165142e-08, 1.324031e-08, 1.380238e-08, 1.267113e-08, 1.222529e-08, 
    1.314091e-08, 1.209697e-08, 1.240774e-08, 1.132577e-08, 1.096073e-08, 
    9.920655e-09, 9.706725e-09, 9.754403e-09, 1.12233e-08, 1.112298e-08, 
    1.066059e-08, 9.850744e-09, 9.818649e-09, 9.057888e-09,
  1.800085e-09, 1.391778e-09, 1.445249e-09, 1.16371e-09, 1.247793e-09, 
    1.16745e-09, 1.765569e-09, 8.377147e-10, 8.201496e-10, 1.06406e-09, 
    1.836239e-09, 2.449499e-09, 3.087838e-09, 1.677385e-09, 1.319136e-09, 
    8.73919e-10, 1.071262e-09, 1.105605e-09, 1.161662e-09, 1.281217e-09, 
    1.359837e-09, 1.520518e-09, 1.74921e-09, 1.768551e-09, 1.484568e-09, 
    1.903181e-09, 2.286894e-09, 2.314627e-09, 2.035882e-09,
  6.703084e-10, 4.469323e-10, 3.758803e-10, 4.251772e-10, 6.492026e-10, 
    5.847692e-10, 3.925388e-10, 6.091136e-10, 3.243844e-10, 2.046679e-10, 
    3.424559e-10, 9.74645e-10, 1.462001e-09, 7.473844e-10, 4.655491e-10, 
    3.207641e-10, 3.304677e-10, 4.055739e-10, 5.289962e-10, 4.065876e-10, 
    5.681681e-10, 5.341802e-10, 5.818289e-10, 5.144066e-10, 5.188776e-10, 
    6.511163e-10, 5.919628e-10, 6.269048e-10, 7.201404e-10,
  2.59103e-10, 2.694522e-10, 3.022927e-10, 2.443226e-10, 1.833533e-10, 
    1.60745e-10, 1.487228e-10, 1.707459e-10, 2.120875e-10, 2.282929e-10, 
    1.609906e-10, 2.723094e-10, 1.112342e-09, 5.285591e-10, 3.674957e-10, 
    3.675132e-10, 3.956472e-10, 3.677754e-10, 5.503708e-10, 7.140341e-10, 
    8.103843e-10, 6.286975e-10, 3.761569e-10, 3.785662e-10, 5.545259e-10, 
    4.042438e-10, 3.968211e-10, 3.944108e-10, 3.207003e-10,
  7.61731e-11, 6.699986e-11, 6.448232e-11, 5.323366e-11, 4.217847e-11, 
    3.520562e-11, 3.626855e-11, 3.962779e-11, 4.416589e-11, 8.733009e-11, 
    9.177143e-11, 2.274281e-10, 7.987364e-10, 5.40919e-10, 3.215614e-10, 
    3.236327e-10, 4.225426e-10, 7.128122e-10, 7.004197e-10, 6.310944e-10, 
    4.755497e-10, 3.40578e-10, 2.348211e-10, 4.156211e-10, 4.79196e-10, 
    2.080079e-10, 1.068149e-10, 1.053751e-10, 8.619635e-11,
  1.889591e-11, 1.881533e-11, 1.352321e-11, 7.119413e-12, 5.151481e-12, 
    5.194423e-12, 4.606104e-12, 5.503132e-12, 7.275751e-12, 9.690472e-12, 
    1.51929e-11, 1.664525e-10, 3.8003e-10, 4.960568e-10, 4.96864e-10, 
    4.534913e-10, 3.922243e-10, 3.422179e-10, 3.120144e-10, 2.733645e-10, 
    2.834328e-10, 3.303655e-10, 3.652482e-10, 4.197046e-10, 2.888315e-10, 
    3.623621e-11, 1.820749e-11, 1.998578e-11, 1.899129e-11,
  1.324723e-11, 1.324723e-11, 1.324723e-11, 1.324723e-11, 1.324723e-11, 
    1.324723e-11, 1.324723e-11, 1.374285e-11, 1.374285e-11, 1.374285e-11, 
    1.374285e-11, 1.374285e-11, 1.374285e-11, 1.374285e-11, 1.40417e-11, 
    1.40417e-11, 1.40417e-11, 1.40417e-11, 1.40417e-11, 1.40417e-11, 
    1.40417e-11, 1.323722e-11, 1.323722e-11, 1.323722e-11, 1.323722e-11, 
    1.323722e-11, 1.323722e-11, 1.323722e-11, 1.324723e-11,
  1.279997e-11, 1.367475e-11, 1.280501e-11, 1.329609e-11, 1.624156e-11, 
    1.478281e-11, 1.459576e-11, 1.589183e-11, 1.703747e-11, 2.263458e-11, 
    3.199734e-11, 3.311347e-11, 3.344642e-11, 3.440241e-11, 3.739285e-11, 
    4.158478e-11, 4.595575e-11, 4.464498e-11, 3.71155e-11, 3.253966e-11, 
    3.174826e-11, 2.926559e-11, 2.493191e-11, 2.051343e-11, 1.593569e-11, 
    1.429312e-11, 1.213169e-11, 1.203869e-11, 1.259534e-11,
  1.837668e-10, 1.646415e-10, 1.244651e-10, 1.052144e-10, 1.249327e-10, 
    1.383068e-10, 1.249681e-10, 1.136774e-10, 8.930785e-11, 6.638006e-11, 
    5.733447e-11, 6.623592e-11, 8.769981e-11, 1.189527e-10, 1.59696e-10, 
    1.9248e-10, 2.13949e-10, 2.146475e-10, 1.640735e-10, 1.471667e-10, 
    1.322727e-10, 9.616777e-11, 9.568404e-11, 1.185718e-10, 1.114113e-10, 
    1.057056e-10, 9.370286e-11, 9.521179e-11, 1.587718e-10,
  4.775433e-10, 4.737329e-10, 4.518098e-10, 5.158797e-10, 7.902419e-10, 
    8.762348e-10, 7.806858e-10, 6.561077e-10, 6.121315e-10, 4.344856e-10, 
    3.742509e-10, 3.73016e-10, 4.510534e-10, 5.849e-10, 7.832368e-10, 
    9.236604e-10, 9.573279e-10, 9.206756e-10, 8.525766e-10, 7.886551e-10, 
    6.658571e-10, 5.529042e-10, 4.175889e-10, 4.087862e-10, 4.354287e-10, 
    7.302648e-10, 5.86995e-10, 4.710614e-10, 5.293543e-10,
  2.164291e-09, 1.827773e-09, 1.554673e-09, 1.564875e-09, 1.67043e-09, 
    1.83886e-09, 1.956933e-09, 1.762205e-09, 1.468578e-09, 1.407148e-09, 
    1.457232e-09, 1.516731e-09, 1.561346e-09, 1.87003e-09, 1.520347e-09, 
    1.364805e-09, 1.460967e-09, 1.655788e-09, 1.53418e-09, 1.067909e-09, 
    9.855227e-10, 1.111327e-09, 1.306863e-09, 1.853239e-09, 2.606198e-09, 
    2.390495e-09, 1.904466e-09, 1.969894e-09, 2.229624e-09,
  5.534251e-09, 5.522676e-09, 6.603767e-09, 6.667318e-09, 6.464697e-09, 
    4.49144e-09, 3.321238e-09, 3.366337e-09, 3.506999e-09, 4.128839e-09, 
    4.142674e-09, 3.85583e-09, 3.193898e-09, 2.702592e-09, 2.282728e-09, 
    2.350332e-09, 2.881422e-09, 3.604059e-09, 4.516814e-09, 5.41092e-09, 
    5.494043e-09, 6.756459e-09, 8.429965e-09, 8.263699e-09, 9.191157e-09, 
    6.841507e-09, 6.319146e-09, 5.294225e-09, 4.610525e-09,
  4.455088e-08, 4.197866e-08, 4.289013e-08, 3.877317e-08, 3.846639e-08, 
    3.548353e-08, 3.719368e-08, 3.77936e-08, 3.837382e-08, 3.723565e-08, 
    3.765693e-08, 3.681395e-08, 3.919342e-08, 4.247797e-08, 4.130987e-08, 
    4.201651e-08, 4.279169e-08, 4.57436e-08, 4.526606e-08, 4.361706e-08, 
    4.693256e-08, 5.103601e-08, 5.235537e-08, 5.082961e-08, 4.916778e-08, 
    4.521979e-08, 4.053598e-08, 4.292029e-08, 4.515462e-08,
  3.160604e-07, 3.001348e-07, 2.958415e-07, 2.954098e-07, 2.946587e-07, 
    2.918555e-07, 2.937049e-07, 2.892983e-07, 2.794821e-07, 2.804956e-07, 
    2.751248e-07, 2.609632e-07, 2.606051e-07, 2.616769e-07, 2.664722e-07, 
    2.694397e-07, 2.772993e-07, 2.828126e-07, 2.937366e-07, 3.022028e-07, 
    3.037314e-07, 3.189252e-07, 3.195537e-07, 3.107731e-07, 3.14286e-07, 
    3.152243e-07, 3.216828e-07, 3.315843e-07, 3.278062e-07,
  7.691157e-07, 7.272314e-07, 7.350553e-07, 7.711274e-07, 7.402722e-07, 
    7.374882e-07, 7.394258e-07, 7.197755e-07, 6.83168e-07, 6.551327e-07, 
    6.180652e-07, 5.60528e-07, 5.246368e-07, 5.067884e-07, 4.958024e-07, 
    4.875431e-07, 4.947603e-07, 5.105933e-07, 5.53699e-07, 6.250455e-07, 
    6.693562e-07, 6.966467e-07, 7.212882e-07, 6.801471e-07, 6.70338e-07, 
    6.85178e-07, 7.163832e-07, 7.841746e-07, 7.780795e-07,
  5.696019e-07, 5.595261e-07, 5.361804e-07, 5.215161e-07, 5.149014e-07, 
    5.345823e-07, 5.836964e-07, 5.798377e-07, 5.8405e-07, 6.255764e-07, 
    6.623579e-07, 6.653392e-07, 6.532004e-07, 6.522204e-07, 6.468456e-07, 
    6.281654e-07, 6.247279e-07, 6.059993e-07, 5.744153e-07, 5.467805e-07, 
    5.422056e-07, 5.404632e-07, 5.549732e-07, 5.856602e-07, 5.742944e-07, 
    5.552004e-07, 5.538806e-07, 5.435032e-07, 5.566687e-07,
  3.942932e-07, 3.992241e-07, 4.220844e-07, 4.5096e-07, 4.369823e-07, 
    4.034264e-07, 3.904528e-07, 3.717018e-07, 3.795607e-07, 3.964601e-07, 
    4.039609e-07, 4.152372e-07, 4.098e-07, 4.10838e-07, 4.089699e-07, 
    4.050181e-07, 4.042115e-07, 4.262945e-07, 4.239152e-07, 4.341005e-07, 
    4.182203e-07, 3.969045e-07, 4.026748e-07, 3.946616e-07, 3.992442e-07, 
    4.076529e-07, 4.239765e-07, 4.073551e-07, 3.89544e-07,
  2.232776e-07, 2.212536e-07, 2.177144e-07, 2.184888e-07, 2.21795e-07, 
    2.190513e-07, 2.312807e-07, 2.251745e-07, 2.419911e-07, 2.568846e-07, 
    2.741967e-07, 2.718994e-07, 2.604661e-07, 2.540228e-07, 2.452657e-07, 
    2.365476e-07, 2.391342e-07, 2.283902e-07, 2.311248e-07, 2.338584e-07, 
    2.311497e-07, 2.288831e-07, 2.297374e-07, 2.302614e-07, 2.313564e-07, 
    2.238192e-07, 2.174971e-07, 2.175646e-07, 2.24886e-07,
  3.493678e-08, 3.619082e-08, 3.53947e-08, 3.530322e-08, 3.329839e-08, 
    3.658929e-08, 3.550468e-08, 3.781304e-08, 4.119403e-08, 4.418918e-08, 
    5.313703e-08, 5.933076e-08, 6.405787e-08, 5.537418e-08, 5.229231e-08, 
    4.851302e-08, 4.400672e-08, 4.453865e-08, 4.487818e-08, 4.27771e-08, 
    4.025614e-08, 4.121613e-08, 4.214672e-08, 4.386543e-08, 4.771857e-08, 
    4.326985e-08, 3.986102e-08, 3.888948e-08, 3.487724e-08,
  6.949661e-09, 6.29253e-09, 5.792078e-09, 5.199573e-09, 5.26247e-09, 
    4.526108e-09, 6.356424e-09, 3.573482e-09, 3.115123e-09, 4.330615e-09, 
    7.581459e-09, 9.213765e-09, 1.315657e-08, 8.937937e-09, 6.698775e-09, 
    4.314244e-09, 5.101976e-09, 5.031878e-09, 5.157428e-09, 5.299292e-09, 
    5.49197e-09, 6.464179e-09, 7.308243e-09, 7.414738e-09, 6.738254e-09, 
    6.846934e-09, 9.648643e-09, 1.022117e-08, 8.493268e-09,
  2.935085e-09, 1.970294e-09, 1.607341e-09, 1.723704e-09, 2.131652e-09, 
    1.97218e-09, 1.361919e-09, 2.130205e-09, 1.20173e-09, 7.615001e-10, 
    1.015048e-09, 3.240156e-09, 4.59402e-09, 3.036458e-09, 1.559254e-09, 
    1.482363e-09, 1.268163e-09, 1.557786e-09, 2.012393e-09, 1.676342e-09, 
    1.958067e-09, 2.774385e-09, 1.855192e-09, 1.698624e-09, 1.719132e-09, 
    2.339803e-09, 2.68168e-09, 2.879799e-09, 3.012118e-09,
  1.172638e-09, 1.38148e-09, 1.209935e-09, 1.021668e-09, 7.993425e-10, 
    7.039225e-10, 6.375195e-10, 6.132556e-10, 6.732043e-10, 7.804475e-10, 
    5.843572e-10, 9.545503e-10, 2.389894e-09, 2.178276e-09, 1.443896e-09, 
    1.227589e-09, 1.665152e-09, 1.270809e-09, 1.59216e-09, 2.081831e-09, 
    2.742738e-09, 2.152017e-09, 1.405103e-09, 9.905767e-10, 1.369018e-09, 
    1.648344e-09, 1.243409e-09, 1.567569e-09, 1.417403e-09,
  3.503583e-10, 3.056169e-10, 3.46717e-10, 2.662904e-10, 1.843755e-10, 
    1.392092e-10, 1.4161e-10, 1.507515e-10, 1.518995e-10, 2.451543e-10, 
    2.666958e-10, 9.47336e-10, 1.94187e-09, 1.53312e-09, 1.169098e-09, 
    1.142889e-09, 1.416091e-09, 2.074956e-09, 2.232368e-09, 2.055349e-09, 
    1.347746e-09, 9.159689e-10, 7.20553e-10, 1.016381e-09, 1.606647e-09, 
    1.171944e-09, 4.519651e-10, 4.732389e-10, 4.368466e-10,
  7.383747e-11, 8.023393e-11, 8.661303e-11, 5.268435e-11, 1.870813e-11, 
    1.877167e-11, 1.90595e-11, 1.941075e-11, 2.318278e-11, 3.002501e-11, 
    4.438264e-11, 7.246992e-10, 1.459475e-09, 1.580307e-09, 1.280996e-09, 
    9.774793e-10, 7.961721e-10, 6.682507e-10, 6.442158e-10, 7.384704e-10, 
    8.586855e-10, 9.164592e-10, 9.554757e-10, 1.040409e-09, 1.087058e-09, 
    4.089315e-10, 1.049863e-10, 9.059279e-11, 7.453991e-11,
  5.244899e-11, 5.244899e-11, 5.244899e-11, 5.244899e-11, 5.244899e-11, 
    5.244899e-11, 5.244899e-11, 5.369144e-11, 5.369144e-11, 5.369144e-11, 
    5.369144e-11, 5.369144e-11, 5.369144e-11, 5.369144e-11, 5.58296e-11, 
    5.58296e-11, 5.58296e-11, 5.58296e-11, 5.58296e-11, 5.58296e-11, 
    5.58296e-11, 5.330524e-11, 5.330524e-11, 5.330524e-11, 5.330524e-11, 
    5.330524e-11, 5.330524e-11, 5.330524e-11, 5.244899e-11,
  4.140589e-11, 4.331211e-11, 5.113443e-11, 6.258781e-11, 6.226193e-11, 
    6.318115e-11, 6.326607e-11, 5.846448e-11, 6.190243e-11, 8.410475e-11, 
    1.060693e-10, 1.123909e-10, 1.209901e-10, 1.307922e-10, 1.423054e-10, 
    1.492159e-10, 1.514597e-10, 1.433431e-10, 1.179793e-10, 1.208025e-10, 
    1.361774e-10, 1.269946e-10, 1.151132e-10, 9.976192e-11, 7.54141e-11, 
    5.583534e-11, 4.243301e-11, 4.025896e-11, 4.109338e-11,
  4.37375e-10, 4.449321e-10, 3.515405e-10, 3.699837e-10, 4.579273e-10, 
    4.616418e-10, 4.331114e-10, 3.644903e-10, 2.833551e-10, 2.290238e-10, 
    2.072341e-10, 2.359212e-10, 2.980625e-10, 4.106116e-10, 5.551829e-10, 
    6.538408e-10, 6.790355e-10, 7.347193e-10, 6.386323e-10, 5.582065e-10, 
    4.937685e-10, 3.650846e-10, 3.391886e-10, 3.822116e-10, 4.050797e-10, 
    3.748794e-10, 3.150324e-10, 2.851855e-10, 3.710255e-10,
  1.562617e-09, 1.522092e-09, 1.569437e-09, 2.009191e-09, 3.018443e-09, 
    3.099794e-09, 2.563985e-09, 2.216162e-09, 1.901526e-09, 1.435231e-09, 
    1.289724e-09, 1.310442e-09, 1.673924e-09, 2.210053e-09, 2.722194e-09, 
    3.244359e-09, 3.498907e-09, 3.209228e-09, 3.058249e-09, 2.900643e-09, 
    2.447577e-09, 2.152218e-09, 1.854203e-09, 1.409411e-09, 1.313609e-09, 
    2.144339e-09, 1.840765e-09, 1.599616e-09, 1.726512e-09,
  6.789359e-09, 6.233404e-09, 5.702014e-09, 5.655676e-09, 5.749855e-09, 
    6.154321e-09, 6.902968e-09, 6.185653e-09, 4.737585e-09, 4.773844e-09, 
    5.42285e-09, 5.752139e-09, 6.670938e-09, 7.104174e-09, 6.213513e-09, 
    5.280246e-09, 5.021208e-09, 5.029607e-09, 4.95925e-09, 3.843126e-09, 
    3.512742e-09, 4.059485e-09, 4.932672e-09, 6.76213e-09, 8.938849e-09, 
    9.377482e-09, 7.255359e-09, 6.315175e-09, 6.649816e-09,
  1.773266e-08, 2.071844e-08, 2.188928e-08, 2.464021e-08, 2.448922e-08, 
    1.76731e-08, 1.502427e-08, 1.503473e-08, 1.67028e-08, 1.806747e-08, 
    1.934768e-08, 1.611888e-08, 1.480314e-08, 1.247867e-08, 9.746345e-09, 
    8.623469e-09, 9.045003e-09, 1.175708e-08, 1.589204e-08, 1.9918e-08, 
    2.134589e-08, 2.782828e-08, 3.349369e-08, 3.471821e-08, 3.918224e-08, 
    3.206932e-08, 2.603093e-08, 2.058682e-08, 1.745526e-08,
  1.763573e-07, 1.714738e-07, 1.734014e-07, 1.6454e-07, 1.537447e-07, 
    1.460446e-07, 1.500457e-07, 1.476044e-07, 1.444784e-07, 1.372262e-07, 
    1.392954e-07, 1.480527e-07, 1.711945e-07, 1.726507e-07, 1.674535e-07, 
    1.780998e-07, 1.726517e-07, 1.675644e-07, 1.596552e-07, 1.614374e-07, 
    1.926995e-07, 2.159205e-07, 2.14371e-07, 1.953146e-07, 1.84107e-07, 
    1.827549e-07, 1.68437e-07, 1.626672e-07, 1.652794e-07,
  1.336835e-06, 1.272012e-06, 1.251172e-06, 1.237804e-06, 1.160355e-06, 
    1.13391e-06, 1.111117e-06, 1.070542e-06, 1.069485e-06, 1.039658e-06, 
    1.020289e-06, 1.02588e-06, 1.017566e-06, 1.019202e-06, 9.938941e-07, 
    1.017542e-06, 1.066527e-06, 1.13291e-06, 1.245069e-06, 1.324971e-06, 
    1.370035e-06, 1.327344e-06, 1.336664e-06, 1.304513e-06, 1.280277e-06, 
    1.240483e-06, 1.285757e-06, 1.341211e-06, 1.348801e-06,
  3.124788e-06, 3.041088e-06, 2.944334e-06, 2.988007e-06, 3.255929e-06, 
    3.18146e-06, 3.183814e-06, 3.113624e-06, 2.852081e-06, 2.764763e-06, 
    2.419913e-06, 2.207024e-06, 2.033436e-06, 2.007274e-06, 1.938095e-06, 
    1.968262e-06, 2.001807e-06, 2.080607e-06, 2.245668e-06, 2.452992e-06, 
    2.718261e-06, 2.806717e-06, 2.759249e-06, 2.733547e-06, 2.630365e-06, 
    2.685101e-06, 2.670197e-06, 2.907975e-06, 3.185064e-06,
  2.088071e-06, 2.05229e-06, 2.02179e-06, 1.958536e-06, 2.004934e-06, 
    2.096615e-06, 2.294262e-06, 2.309843e-06, 2.401981e-06, 2.480546e-06, 
    2.580656e-06, 2.680162e-06, 2.672765e-06, 2.624786e-06, 2.634169e-06, 
    2.49911e-06, 2.342744e-06, 2.306404e-06, 2.330001e-06, 2.209122e-06, 
    2.114611e-06, 2.174293e-06, 2.176983e-06, 2.146589e-06, 2.160425e-06, 
    2.140449e-06, 2.025552e-06, 2.017863e-06, 2.050097e-06,
  1.657461e-06, 1.651397e-06, 1.75067e-06, 1.779341e-06, 1.760179e-06, 
    1.647463e-06, 1.59535e-06, 1.494822e-06, 1.527274e-06, 1.630044e-06, 
    1.833996e-06, 1.737526e-06, 1.66991e-06, 1.667933e-06, 1.613529e-06, 
    1.584419e-06, 1.591296e-06, 1.648637e-06, 1.677494e-06, 1.618784e-06, 
    1.623668e-06, 1.671109e-06, 1.678828e-06, 1.744409e-06, 1.656121e-06, 
    1.64902e-06, 1.684161e-06, 1.726914e-06, 1.732283e-06,
  8.99956e-07, 8.550221e-07, 8.840532e-07, 8.865091e-07, 8.934677e-07, 
    8.729012e-07, 9.124449e-07, 9.842533e-07, 9.966519e-07, 1.121934e-06, 
    1.165357e-06, 1.12158e-06, 1.109598e-06, 1.029609e-06, 9.722578e-07, 
    9.479405e-07, 9.29824e-07, 9.330435e-07, 9.305342e-07, 9.536664e-07, 
    9.09228e-07, 9.300476e-07, 9.210056e-07, 9.049791e-07, 8.835888e-07, 
    9.037229e-07, 9.165783e-07, 9.092326e-07, 8.760837e-07,
  1.661902e-07, 1.611254e-07, 1.539318e-07, 1.440226e-07, 1.352036e-07, 
    1.517503e-07, 1.482326e-07, 1.55195e-07, 1.73629e-07, 1.882896e-07, 
    2.341251e-07, 2.751611e-07, 2.904553e-07, 2.444272e-07, 2.126134e-07, 
    2.091514e-07, 1.938208e-07, 1.92104e-07, 1.893113e-07, 1.893479e-07, 
    1.906419e-07, 1.87731e-07, 1.847551e-07, 1.924125e-07, 2.02897e-07, 
    1.882604e-07, 1.764275e-07, 1.749806e-07, 1.668647e-07,
  3.192675e-08, 3.062391e-08, 2.728744e-08, 2.476642e-08, 2.492172e-08, 
    2.107056e-08, 2.673683e-08, 1.760864e-08, 1.304322e-08, 1.591163e-08, 
    2.738117e-08, 3.944419e-08, 5.531634e-08, 4.770852e-08, 3.111484e-08, 
    2.297399e-08, 2.384466e-08, 2.282969e-08, 2.17789e-08, 2.33679e-08, 
    2.300184e-08, 2.718706e-08, 3.035033e-08, 3.236028e-08, 3.107715e-08, 
    3.066168e-08, 4.074964e-08, 4.433391e-08, 3.576337e-08,
  1.045593e-08, 8.93608e-09, 6.730947e-09, 5.883358e-09, 6.729794e-09, 
    7.070566e-09, 4.75961e-09, 6.53364e-09, 4.160505e-09, 2.783412e-09, 
    3.247139e-09, 1.124502e-08, 1.297211e-08, 1.418131e-08, 6.259382e-09, 
    5.637345e-09, 5.078543e-09, 5.207259e-09, 6.111024e-09, 6.377958e-09, 
    7.429109e-09, 1.099392e-08, 9.980393e-09, 6.160931e-09, 6.863269e-09, 
    8.275486e-09, 9.842926e-09, 9.807711e-09, 1.050989e-08,
  6.808033e-09, 5.16194e-09, 4.426107e-09, 3.697706e-09, 3.118647e-09, 
    2.913986e-09, 2.581547e-09, 2.143983e-09, 2.344391e-09, 2.368806e-09, 
    1.926056e-09, 3.083094e-09, 7.075351e-09, 7.397666e-09, 5.43104e-09, 
    4.176298e-09, 5.935144e-09, 4.469247e-09, 4.457049e-09, 6.5668e-09, 
    7.954494e-09, 7.250043e-09, 4.268011e-09, 3.161339e-09, 4.139166e-09, 
    4.885789e-09, 5.280772e-09, 6.113498e-09, 6.607348e-09,
  1.902502e-09, 1.660951e-09, 1.886605e-09, 1.464643e-09, 8.180874e-10, 
    5.107267e-10, 4.942908e-10, 4.910282e-10, 4.673136e-10, 5.102955e-10, 
    8.317595e-10, 2.662513e-09, 4.78596e-09, 4.767144e-09, 4.476306e-09, 
    4.193857e-09, 4.64428e-09, 5.654683e-09, 6.041687e-09, 5.742131e-09, 
    4.282156e-09, 2.38739e-09, 2.484031e-09, 3.084946e-09, 5.017641e-09, 
    4.950444e-09, 2.108376e-09, 1.932011e-09, 2.088817e-09,
  2.418147e-10, 2.222336e-10, 2.699969e-10, 2.376773e-10, 8.781467e-11, 
    6.434552e-11, 6.844529e-11, 7.33834e-11, 8.13801e-11, 9.816808e-11, 
    2.517389e-10, 2.640925e-09, 5.281692e-09, 4.069087e-09, 2.418171e-09, 
    2.071913e-09, 1.899401e-09, 1.716337e-09, 1.623613e-09, 1.692309e-09, 
    2.264643e-09, 2.583844e-09, 2.371729e-09, 2.847565e-09, 2.676651e-09, 
    1.942095e-09, 5.383615e-10, 3.328229e-10, 2.683598e-10,
  1.622715e-10, 1.622715e-10, 1.622715e-10, 1.622715e-10, 1.622715e-10, 
    1.622715e-10, 1.622715e-10, 1.839868e-10, 1.839868e-10, 1.839868e-10, 
    1.839868e-10, 1.839868e-10, 1.839868e-10, 1.839868e-10, 1.833026e-10, 
    1.833026e-10, 1.833026e-10, 1.833026e-10, 1.833026e-10, 1.833026e-10, 
    1.833026e-10, 1.657024e-10, 1.657024e-10, 1.657024e-10, 1.657024e-10, 
    1.657024e-10, 1.657024e-10, 1.657024e-10, 1.622715e-10,
  1.585583e-10, 1.691203e-10, 1.900374e-10, 2.239702e-10, 2.250211e-10, 
    2.541655e-10, 2.456832e-10, 2.215112e-10, 2.305658e-10, 2.648936e-10, 
    3.249016e-10, 3.661749e-10, 4.091454e-10, 4.500538e-10, 4.862798e-10, 
    5.039575e-10, 4.876353e-10, 4.567628e-10, 3.942612e-10, 4.313176e-10, 
    5.117261e-10, 4.974809e-10, 4.782202e-10, 4.311665e-10, 3.509549e-10, 
    2.611861e-10, 1.867177e-10, 1.617179e-10, 1.52809e-10,
  9.332589e-10, 1.044291e-09, 9.578669e-10, 1.104115e-09, 1.385187e-09, 
    1.42055e-09, 1.186185e-09, 1.025523e-09, 8.598623e-10, 8.305299e-10, 
    8.060949e-10, 8.560544e-10, 1.080608e-09, 1.51726e-09, 2.031922e-09, 
    2.685832e-09, 3.175914e-09, 2.994616e-09, 2.381613e-09, 2.102194e-09, 
    1.89696e-09, 1.442719e-09, 1.260141e-09, 1.306149e-09, 1.469938e-09, 
    1.416178e-09, 1.075421e-09, 9.17744e-10, 9.183546e-10,
  5.306374e-09, 5.102025e-09, 6.604921e-09, 7.422509e-09, 1.07122e-08, 
    1.108146e-08, 9.355228e-09, 7.916994e-09, 6.069858e-09, 5.144402e-09, 
    5.177312e-09, 5.405377e-09, 6.306492e-09, 8.467147e-09, 9.943124e-09, 
    1.174997e-08, 1.320635e-08, 1.205724e-08, 1.110529e-08, 1.078755e-08, 
    9.660906e-09, 8.679315e-09, 7.428013e-09, 6.519814e-09, 5.076433e-09, 
    6.568114e-09, 6.79057e-09, 5.716765e-09, 5.919939e-09,
  2.316408e-08, 2.361251e-08, 2.218329e-08, 2.233909e-08, 2.327497e-08, 
    2.009382e-08, 2.343926e-08, 2.203184e-08, 1.711785e-08, 1.657598e-08, 
    1.925906e-08, 2.363826e-08, 2.91994e-08, 3.278373e-08, 2.8506e-08, 
    2.35005e-08, 2.028295e-08, 1.734148e-08, 1.601081e-08, 1.50524e-08, 
    1.310074e-08, 1.608248e-08, 2.024134e-08, 2.818406e-08, 3.402686e-08, 
    3.483959e-08, 2.98436e-08, 2.449894e-08, 2.073894e-08,
  6.838152e-08, 7.679954e-08, 8.315831e-08, 9.519916e-08, 9.246574e-08, 
    6.761136e-08, 5.972333e-08, 7.240966e-08, 8.0002e-08, 8.827534e-08, 
    9.636526e-08, 7.561622e-08, 6.975861e-08, 6.90787e-08, 5.282456e-08, 
    3.919063e-08, 3.625249e-08, 4.771435e-08, 6.547525e-08, 7.604663e-08, 
    8.97237e-08, 1.015735e-07, 1.345346e-07, 1.568531e-07, 1.478089e-07, 
    1.358933e-07, 1.131433e-07, 8.885227e-08, 7.592572e-08,
  7.682044e-07, 7.390652e-07, 7.18534e-07, 6.954937e-07, 6.670508e-07, 
    6.918224e-07, 6.625446e-07, 6.99116e-07, 6.819175e-07, 5.877837e-07, 
    5.374523e-07, 5.360086e-07, 5.953642e-07, 6.388121e-07, 6.977842e-07, 
    7.022859e-07, 6.905183e-07, 6.427061e-07, 6.129753e-07, 6.500018e-07, 
    7.74332e-07, 8.61241e-07, 8.380715e-07, 8.001592e-07, 7.764282e-07, 
    7.477738e-07, 7.061457e-07, 7.189594e-07, 7.171897e-07,
  5.589536e-06, 5.463667e-06, 5.264319e-06, 5.296768e-06, 5.137537e-06, 
    4.877162e-06, 4.761608e-06, 4.522473e-06, 4.315926e-06, 4.217973e-06, 
    3.934439e-06, 3.80264e-06, 3.876421e-06, 4.063848e-06, 4.120173e-06, 
    4.3329e-06, 4.375021e-06, 4.481504e-06, 4.850085e-06, 4.992824e-06, 
    5.432761e-06, 6.01279e-06, 5.67604e-06, 5.541924e-06, 5.469371e-06, 
    5.565076e-06, 5.461333e-06, 5.566809e-06, 5.670974e-06,
  1.344018e-05, 1.313988e-05, 1.285153e-05, 1.342401e-05, 1.257417e-05, 
    1.307075e-05, 1.318154e-05, 1.317653e-05, 1.308817e-05, 1.210487e-05, 
    1.066395e-05, 9.415737e-06, 8.411877e-06, 7.668657e-06, 7.352041e-06, 
    7.291512e-06, 7.713614e-06, 7.970725e-06, 8.841411e-06, 9.765909e-06, 
    1.050934e-05, 1.150545e-05, 1.188279e-05, 1.115007e-05, 1.032585e-05, 
    1.040464e-05, 1.072679e-05, 1.183504e-05, 1.297929e-05,
  8.116502e-06, 8.261085e-06, 8.105574e-06, 8.036064e-06, 8.100833e-06, 
    8.761672e-06, 9.727156e-06, 9.383039e-06, 9.905858e-06, 1.045354e-05, 
    1.118874e-05, 1.135409e-05, 1.108745e-05, 1.096379e-05, 1.074961e-05, 
    1.102381e-05, 1.077107e-05, 1.023554e-05, 9.445995e-06, 8.969525e-06, 
    9.000944e-06, 8.523041e-06, 8.369605e-06, 8.151079e-06, 8.202073e-06, 
    8.131223e-06, 8.054409e-06, 7.965538e-06, 8.082175e-06,
  7.146969e-06, 7.131592e-06, 7.441524e-06, 7.195715e-06, 7.039195e-06, 
    7.100466e-06, 6.715929e-06, 6.648513e-06, 6.601826e-06, 6.64489e-06, 
    7.614957e-06, 7.276041e-06, 6.964783e-06, 6.589557e-06, 6.199732e-06, 
    5.943902e-06, 6.007194e-06, 6.683341e-06, 6.668914e-06, 6.659175e-06, 
    6.252618e-06, 6.344747e-06, 6.901159e-06, 6.90001e-06, 7.044302e-06, 
    7.191982e-06, 7.225687e-06, 6.983199e-06, 6.656243e-06,
  4.061072e-06, 3.913286e-06, 3.830904e-06, 3.77266e-06, 3.67993e-06, 
    3.817903e-06, 3.873626e-06, 3.959987e-06, 4.259522e-06, 4.605311e-06, 
    5.126461e-06, 4.996905e-06, 4.927612e-06, 4.348779e-06, 4.305974e-06, 
    4.166976e-06, 4.167054e-06, 4.149516e-06, 4.170062e-06, 4.21427e-06, 
    4.211389e-06, 4.022114e-06, 4.151418e-06, 4.069261e-06, 4.156898e-06, 
    4.060119e-06, 3.978017e-06, 3.989465e-06, 4.01804e-06,
  8.063567e-07, 8.071477e-07, 7.66125e-07, 7.253243e-07, 6.562699e-07, 
    6.601111e-07, 6.662564e-07, 6.332767e-07, 7.038608e-07, 8.440879e-07, 
    1.005609e-06, 1.193731e-06, 1.301834e-06, 1.040767e-06, 8.879441e-07, 
    8.637148e-07, 8.458375e-07, 7.918061e-07, 8.153522e-07, 8.612583e-07, 
    8.670227e-07, 9.202574e-07, 9.543044e-07, 9.705423e-07, 1.023179e-06, 
    9.721763e-07, 8.793232e-07, 8.840254e-07, 8.150092e-07,
  1.592991e-07, 1.691394e-07, 1.413934e-07, 1.366099e-07, 1.332661e-07, 
    1.226399e-07, 1.30194e-07, 9.413067e-08, 6.517659e-08, 6.139352e-08, 
    9.350769e-08, 1.512545e-07, 2.021083e-07, 2.330508e-07, 1.356102e-07, 
    1.222455e-07, 1.206177e-07, 9.926956e-08, 1.037108e-07, 1.039007e-07, 
    9.535385e-08, 1.077644e-07, 1.288175e-07, 1.431171e-07, 1.459871e-07, 
    1.344401e-07, 1.665106e-07, 1.748127e-07, 1.571222e-07,
  3.930822e-08, 3.495694e-08, 2.837766e-08, 2.266562e-08, 2.470491e-08, 
    2.697628e-08, 1.983157e-08, 2.308382e-08, 1.740231e-08, 1.08857e-08, 
    1.11555e-08, 3.744363e-08, 4.066368e-08, 7.246395e-08, 3.514583e-08, 
    2.152954e-08, 2.060719e-08, 1.975035e-08, 2.138276e-08, 2.318738e-08, 
    2.698763e-08, 3.11639e-08, 4.131489e-08, 2.876743e-08, 3.082953e-08, 
    3.804426e-08, 3.74354e-08, 3.991509e-08, 4.168255e-08,
  3.053588e-08, 2.185405e-08, 1.640272e-08, 1.167267e-08, 1.117358e-08, 
    1.139517e-08, 1.001051e-08, 7.903878e-09, 8.185562e-09, 7.585321e-09, 
    6.928133e-09, 8.997233e-09, 2.423045e-08, 2.313835e-08, 2.038272e-08, 
    1.604748e-08, 1.74711e-08, 1.548041e-08, 1.452885e-08, 2.252672e-08, 
    2.872023e-08, 2.466623e-08, 1.220257e-08, 9.799709e-09, 1.317659e-08, 
    1.584245e-08, 2.422792e-08, 2.986031e-08, 3.519302e-08,
  8.90819e-09, 8.994399e-09, 1.424264e-08, 1.093282e-08, 4.76829e-09, 
    2.335255e-09, 2.065539e-09, 1.87074e-09, 1.687323e-09, 1.467902e-09, 
    2.366981e-09, 6.989342e-09, 1.627122e-08, 1.658609e-08, 1.784105e-08, 
    1.568202e-08, 1.606683e-08, 1.752054e-08, 1.812629e-08, 1.597627e-08, 
    1.2253e-08, 7.641264e-09, 7.239632e-09, 8.221268e-09, 1.398941e-08, 
    1.746288e-08, 9.89379e-09, 6.731459e-09, 8.149394e-09,
  9.597005e-10, 7.635509e-10, 7.830676e-10, 8.104333e-10, 5.015431e-10, 
    2.556535e-10, 2.367174e-10, 2.404195e-10, 3.160388e-10, 5.055462e-10, 
    1.862832e-09, 6.446129e-09, 1.241406e-08, 8.638141e-09, 5.368755e-09, 
    4.99367e-09, 4.733913e-09, 4.526773e-09, 4.174431e-09, 4.060154e-09, 
    4.751166e-09, 5.614974e-09, 6.022522e-09, 7.368488e-09, 7.025156e-09, 
    6.98532e-09, 3.47854e-09, 1.429425e-09, 1.067422e-09,
  6.46474e-10, 6.46474e-10, 6.46474e-10, 6.46474e-10, 6.46474e-10, 
    6.46474e-10, 6.46474e-10, 6.785218e-10, 6.785218e-10, 6.785218e-10, 
    6.785218e-10, 6.785218e-10, 6.785218e-10, 6.785218e-10, 6.933575e-10, 
    6.933575e-10, 6.933575e-10, 6.933575e-10, 6.933575e-10, 6.933575e-10, 
    6.933575e-10, 6.835973e-10, 6.835973e-10, 6.835973e-10, 6.835973e-10, 
    6.835973e-10, 6.835973e-10, 6.835973e-10, 6.46474e-10,
  6.118613e-10, 5.785175e-10, 6.241016e-10, 8.131224e-10, 9.329554e-10, 
    9.176082e-10, 9.026159e-10, 8.589836e-10, 9.408242e-10, 9.441588e-10, 
    1.05206e-09, 1.166345e-09, 1.367207e-09, 1.68166e-09, 1.821084e-09, 
    1.767771e-09, 1.706907e-09, 1.63601e-09, 1.680587e-09, 1.947628e-09, 
    2.126457e-09, 2.128141e-09, 2.04871e-09, 1.923627e-09, 1.680893e-09, 
    1.358932e-09, 1.01653e-09, 7.586856e-10, 6.241506e-10,
  2.417557e-09, 2.186461e-09, 2.472341e-09, 3.046639e-09, 3.571e-09, 
    4.099298e-09, 3.524665e-09, 3.315833e-09, 3.067666e-09, 2.97787e-09, 
    2.999895e-09, 3.200602e-09, 4.542786e-09, 5.543621e-09, 8.2861e-09, 
    1.203994e-08, 1.355445e-08, 1.263486e-08, 1.104143e-08, 7.959776e-09, 
    7.369497e-09, 5.926116e-09, 5.032128e-09, 4.91932e-09, 5.419968e-09, 
    5.481442e-09, 4.298652e-09, 3.784864e-09, 2.910466e-09,
  2.149365e-08, 2.022445e-08, 2.305058e-08, 2.794061e-08, 3.701775e-08, 
    4.166406e-08, 3.421858e-08, 2.666016e-08, 2.071503e-08, 1.963744e-08, 
    2.117663e-08, 2.400109e-08, 2.68467e-08, 3.230166e-08, 3.782488e-08, 
    4.387971e-08, 5.106534e-08, 5.001051e-08, 4.328048e-08, 4.250378e-08, 
    4.046958e-08, 3.37136e-08, 2.627055e-08, 2.412913e-08, 2.263082e-08, 
    2.418503e-08, 2.317286e-08, 1.945673e-08, 2.141971e-08,
  8.429728e-08, 9.200811e-08, 8.919281e-08, 8.860584e-08, 9.404967e-08, 
    9.086035e-08, 8.848025e-08, 8.145302e-08, 6.865383e-08, 6.625467e-08, 
    7.976652e-08, 1.002885e-07, 1.278952e-07, 1.397158e-07, 1.284453e-07, 
    1.118392e-07, 8.778119e-08, 7.076418e-08, 6.089348e-08, 6.142998e-08, 
    5.160589e-08, 5.872617e-08, 1.035924e-07, 1.341319e-07, 1.464077e-07, 
    1.428956e-07, 1.177042e-07, 1.016733e-07, 8.351844e-08,
  3.053478e-07, 3.133003e-07, 3.466044e-07, 3.802129e-07, 3.727287e-07, 
    3.232142e-07, 2.669517e-07, 2.826973e-07, 3.713347e-07, 4.242995e-07, 
    4.937409e-07, 4.265054e-07, 4.108516e-07, 4.014772e-07, 3.04148e-07, 
    2.144024e-07, 1.684475e-07, 1.848036e-07, 2.532299e-07, 3.128739e-07, 
    3.891029e-07, 5.365858e-07, 5.857424e-07, 6.275419e-07, 5.878534e-07, 
    5.684769e-07, 5.495187e-07, 4.484835e-07, 3.420669e-07,
  3.285689e-06, 3.337527e-06, 3.32169e-06, 3.239278e-06, 3.228058e-06, 
    3.371318e-06, 3.586694e-06, 3.633249e-06, 3.274316e-06, 2.943892e-06, 
    2.625347e-06, 2.321632e-06, 2.138559e-06, 2.108093e-06, 2.256036e-06, 
    2.53232e-06, 2.61536e-06, 2.73059e-06, 2.652483e-06, 2.840658e-06, 
    3.170408e-06, 3.3358e-06, 3.374687e-06, 3.225543e-06, 3.199461e-06, 
    3.33852e-06, 3.142339e-06, 3.115322e-06, 3.284891e-06,
  2.559235e-05, 2.454828e-05, 2.474096e-05, 2.375653e-05, 2.310402e-05, 
    2.187643e-05, 2.108048e-05, 1.972546e-05, 1.890704e-05, 1.752905e-05, 
    1.680819e-05, 1.642836e-05, 1.630375e-05, 1.625433e-05, 1.63136e-05, 
    1.662863e-05, 1.806321e-05, 1.911994e-05, 2.062277e-05, 2.299271e-05, 
    2.38738e-05, 2.30619e-05, 2.447429e-05, 2.239786e-05, 2.313079e-05, 
    2.228755e-05, 2.412747e-05, 2.520458e-05, 2.550228e-05,
  5.655004e-05, 5.549475e-05, 5.508085e-05, 5.399436e-05, 5.633978e-05, 
    5.79419e-05, 5.954029e-05, 5.830745e-05, 5.650365e-05, 5.111366e-05, 
    4.285688e-05, 3.595049e-05, 3.376975e-05, 3.296857e-05, 3.275877e-05, 
    3.290465e-05, 3.396445e-05, 3.594537e-05, 3.720706e-05, 3.950438e-05, 
    4.162651e-05, 4.59066e-05, 4.863346e-05, 4.659381e-05, 4.541215e-05, 
    4.26093e-05, 4.345484e-05, 4.865551e-05, 5.290163e-05,
  3.28444e-05, 3.365815e-05, 3.39223e-05, 3.270019e-05, 3.395194e-05, 
    3.808575e-05, 4.120198e-05, 4.054995e-05, 4.303857e-05, 4.50655e-05, 
    4.819731e-05, 5.008452e-05, 5.07513e-05, 4.856371e-05, 4.89089e-05, 
    4.571059e-05, 4.294803e-05, 3.985473e-05, 3.826087e-05, 3.59114e-05, 
    3.369303e-05, 3.303291e-05, 3.30993e-05, 3.442529e-05, 3.491629e-05, 
    3.346404e-05, 3.149329e-05, 3.11551e-05, 3.165457e-05,
  3.077891e-05, 3.194812e-05, 3.332246e-05, 3.239668e-05, 3.026112e-05, 
    2.898937e-05, 2.865165e-05, 2.780123e-05, 2.855512e-05, 3.218418e-05, 
    3.525646e-05, 3.270089e-05, 3.102463e-05, 2.917675e-05, 2.80436e-05, 
    2.692233e-05, 2.697751e-05, 2.710573e-05, 2.691844e-05, 2.524663e-05, 
    2.626013e-05, 2.741217e-05, 2.820807e-05, 2.901594e-05, 2.824885e-05, 
    2.980213e-05, 3.149993e-05, 3.119525e-05, 3.081362e-05,
  1.938493e-05, 2.007581e-05, 1.816188e-05, 1.80809e-05, 1.707896e-05, 
    1.658163e-05, 1.650411e-05, 1.718051e-05, 1.839922e-05, 2.00732e-05, 
    2.129062e-05, 2.129916e-05, 2.040174e-05, 1.768904e-05, 1.796636e-05, 
    1.785498e-05, 1.7258e-05, 1.711586e-05, 1.814645e-05, 1.881525e-05, 
    1.900051e-05, 1.926894e-05, 1.949997e-05, 1.960706e-05, 1.953049e-05, 
    1.967126e-05, 1.995509e-05, 1.982443e-05, 1.950706e-05,
  5.225524e-06, 4.686692e-06, 4.27339e-06, 3.976557e-06, 3.529802e-06, 
    3.39167e-06, 3.019901e-06, 2.659875e-06, 2.748658e-06, 3.561707e-06, 
    4.923451e-06, 5.293288e-06, 6.021138e-06, 5.022111e-06, 4.295655e-06, 
    4.094344e-06, 3.927275e-06, 3.82022e-06, 3.776295e-06, 4.106487e-06, 
    4.273345e-06, 4.208618e-06, 4.332198e-06, 4.601595e-06, 4.762459e-06, 
    5.086115e-06, 5.01258e-06, 5.132019e-06, 5.157808e-06,
  8.331973e-07, 9.088626e-07, 7.901817e-07, 7.587134e-07, 7.625624e-07, 
    7.275262e-07, 6.770298e-07, 5.888936e-07, 4.159197e-07, 2.887022e-07, 
    3.52475e-07, 5.930833e-07, 7.862209e-07, 1.055115e-06, 6.816239e-07, 
    5.439935e-07, 5.421877e-07, 5.065983e-07, 5.141389e-07, 5.44338e-07, 
    4.369997e-07, 4.556723e-07, 5.417555e-07, 6.557678e-07, 6.863957e-07, 
    7.013592e-07, 8.663795e-07, 8.785532e-07, 8.02668e-07,
  1.701414e-07, 1.364094e-07, 1.242223e-07, 9.649514e-08, 9.523259e-08, 
    9.424958e-08, 8.337638e-08, 9.440458e-08, 8.749619e-08, 5.662403e-08, 
    4.648087e-08, 1.107251e-07, 1.390221e-07, 2.333095e-07, 2.169938e-07, 
    1.084871e-07, 1.026784e-07, 1.102803e-07, 1.218315e-07, 1.179292e-07, 
    1.08222e-07, 1.108589e-07, 1.302688e-07, 1.272302e-07, 1.328881e-07, 
    1.503523e-07, 1.582778e-07, 1.509898e-07, 1.75774e-07,
  1.132192e-07, 8.832136e-08, 6.004774e-08, 4.594892e-08, 3.903762e-08, 
    3.619778e-08, 3.925181e-08, 2.931277e-08, 2.676091e-08, 2.430223e-08, 
    2.248814e-08, 3.250652e-08, 6.510128e-08, 6.554749e-08, 9.04141e-08, 
    6.078037e-08, 6.183365e-08, 6.055279e-08, 5.538182e-08, 7.358705e-08, 
    1.223232e-07, 7.461262e-08, 3.841554e-08, 3.169643e-08, 3.467479e-08, 
    5.069944e-08, 8.423425e-08, 1.09336e-07, 1.439632e-07,
  3.242388e-08, 6.472403e-08, 7.294163e-08, 5.614135e-08, 2.786367e-08, 
    1.082809e-08, 7.984522e-09, 6.502737e-09, 6.01946e-09, 5.478976e-09, 
    6.359568e-09, 1.856238e-08, 4.430236e-08, 4.790034e-08, 6.056227e-08, 
    6.01857e-08, 6.661559e-08, 7.429473e-08, 6.80332e-08, 6.006431e-08, 
    3.436522e-08, 2.491155e-08, 1.790696e-08, 1.826207e-08, 3.036561e-08, 
    4.67871e-08, 4.029318e-08, 2.487721e-08, 2.608352e-08,
  5.124903e-09, 3.712481e-09, 2.648835e-09, 2.529924e-09, 2.130692e-09, 
    1.384257e-09, 1.027818e-09, 1.301187e-09, 2.211742e-09, 4.787329e-09, 
    1.074102e-08, 1.724071e-08, 2.484499e-08, 1.938999e-08, 1.388271e-08, 
    1.210194e-08, 1.143587e-08, 1.163438e-08, 1.070714e-08, 9.575355e-09, 
    9.250304e-09, 9.562821e-09, 1.10096e-08, 1.431449e-08, 2.067311e-08, 
    2.481011e-08, 1.843618e-08, 1.008969e-08, 6.271585e-09,
  3.054962e-09, 3.054962e-09, 3.054962e-09, 3.054962e-09, 3.054962e-09, 
    3.054962e-09, 3.054962e-09, 3.103097e-09, 3.103097e-09, 3.103097e-09, 
    3.103097e-09, 3.103097e-09, 3.103097e-09, 3.103097e-09, 3.222405e-09, 
    3.222405e-09, 3.222405e-09, 3.222405e-09, 3.222405e-09, 3.222405e-09, 
    3.222405e-09, 3.307464e-09, 3.307464e-09, 3.307464e-09, 3.307464e-09, 
    3.307464e-09, 3.307464e-09, 3.307464e-09, 3.054962e-09,
  3.581226e-09, 2.907362e-09, 2.298477e-09, 2.60409e-09, 3.212041e-09, 
    3.614548e-09, 3.533132e-09, 3.744092e-09, 3.899314e-09, 3.798711e-09, 
    4.131361e-09, 4.653924e-09, 5.115234e-09, 6.606071e-09, 9.169251e-09, 
    6.453729e-09, 6.395201e-09, 6.670883e-09, 7.521558e-09, 9.222489e-09, 
    9.539631e-09, 9.155902e-09, 8.750851e-09, 8.302822e-09, 7.592765e-09, 
    6.879036e-09, 5.718342e-09, 4.521633e-09, 3.741596e-09,
  1.308698e-08, 9.547453e-09, 8.754015e-09, 1.072183e-08, 1.145907e-08, 
    1.350164e-08, 1.474401e-08, 1.289629e-08, 1.188729e-08, 1.190035e-08, 
    1.161282e-08, 1.303321e-08, 1.948353e-08, 2.87164e-08, 3.48188e-08, 
    4.360319e-08, 4.387145e-08, 4.296537e-08, 4.502854e-08, 3.59853e-08, 
    3.089203e-08, 2.443598e-08, 2.040322e-08, 1.864943e-08, 1.966216e-08, 
    2.005436e-08, 1.821726e-08, 1.449146e-08, 1.340405e-08,
  9.554034e-08, 9.467323e-08, 8.680088e-08, 1.124974e-07, 1.339974e-07, 
    1.407278e-07, 1.246513e-07, 8.933541e-08, 7.632609e-08, 6.893689e-08, 
    6.999334e-08, 9.962342e-08, 1.114794e-07, 1.386022e-07, 1.559353e-07, 
    1.70533e-07, 1.982771e-07, 1.947577e-07, 1.703631e-07, 1.565603e-07, 
    1.471165e-07, 1.328193e-07, 1.028491e-07, 9.337997e-08, 1.00734e-07, 
    1.026087e-07, 9.037691e-08, 7.5975e-08, 7.818959e-08,
  3.579464e-07, 3.932971e-07, 3.615649e-07, 3.487501e-07, 3.822755e-07, 
    4.001098e-07, 3.783069e-07, 3.37443e-07, 2.905931e-07, 2.675705e-07, 
    3.373677e-07, 4.155857e-07, 5.536522e-07, 5.660298e-07, 5.612023e-07, 
    5.197976e-07, 3.744586e-07, 3.244982e-07, 2.755765e-07, 2.753762e-07, 
    2.237204e-07, 2.177866e-07, 4.183633e-07, 6.462227e-07, 6.181087e-07, 
    5.579793e-07, 4.499366e-07, 4.569479e-07, 3.866307e-07,
  1.417414e-06, 1.385026e-06, 1.560105e-06, 1.611075e-06, 1.702238e-06, 
    1.664747e-06, 1.541892e-06, 1.255568e-06, 1.576535e-06, 2.485092e-06, 
    2.987193e-06, 2.549044e-06, 2.119e-06, 2.855016e-06, 1.794087e-06, 
    1.093998e-06, 1.044553e-06, 8.111238e-07, 1.142266e-06, 1.326771e-06, 
    1.756124e-06, 3.114413e-06, 3.040393e-06, 2.282772e-06, 2.487054e-06, 
    2.607187e-06, 2.62027e-06, 2.450876e-06, 1.629262e-06,
  1.619237e-05, 1.558847e-05, 1.399656e-05, 1.52184e-05, 1.467499e-05, 
    1.587439e-05, 1.805876e-05, 1.94677e-05, 2.007907e-05, 1.785926e-05, 
    1.432161e-05, 1.190471e-05, 1.017779e-05, 8.116315e-06, 7.716275e-06, 
    8.056596e-06, 9.120643e-06, 1.008263e-05, 1.162976e-05, 1.215952e-05, 
    1.308777e-05, 1.379521e-05, 1.460606e-05, 1.518134e-05, 1.393756e-05, 
    1.280547e-05, 1.347095e-05, 1.371244e-05, 1.487497e-05,
  0.0001138842, 0.0001164106, 0.0001121129, 0.0001136466, 0.0001147988, 
    0.0001121901, 0.000108053, 0.0001016508, 8.525946e-05, 7.703801e-05, 
    6.727094e-05, 6.34753e-05, 6.460924e-05, 6.634217e-05, 6.83979e-05, 
    7.090419e-05, 6.962627e-05, 7.139769e-05, 7.768303e-05, 8.528531e-05, 
    9.212326e-05, 0.0001019959, 9.882567e-05, 0.0001028202, 9.857088e-05, 
    9.998229e-05, 0.0001001957, 0.0001067446, 0.0001126301,
  0.0002278669, 0.0002227437, 0.00022076, 0.0002198084, 0.0002301981, 
    0.0002553038, 0.000276833, 0.0002829647, 0.0002748319, 0.0002529485, 
    0.0002025485, 0.000169623, 0.0001395376, 0.0001289726, 0.0001282289, 
    0.0001320913, 0.0001383753, 0.000146682, 0.0001651538, 0.0001758628, 
    0.0001904954, 0.0001985763, 0.0002005598, 0.0001905644, 0.0001887683, 
    0.0001776558, 0.0001857921, 0.0002140258, 0.000226667,
  0.0001405185, 0.0001564331, 0.0001525466, 0.0001500761, 0.0001579384, 
    0.0001697839, 0.0001845804, 0.0001829047, 0.0001927694, 0.0002148414, 
    0.0002316182, 0.0002360069, 0.0002217366, 0.0002147875, 0.0001873444, 
    0.000187629, 0.0001754125, 0.0001695604, 0.0001513132, 0.0001464797, 
    0.0001382949, 0.0001351309, 0.0001392858, 0.0001420427, 0.0001496773, 
    0.000145932, 0.0001414977, 0.000139156, 0.0001360768,
  0.0001482726, 0.0001474636, 0.000148861, 0.0001470361, 0.0001472279, 
    0.0001421478, 0.0001432816, 0.0001312555, 0.0001386412, 0.0001504174, 
    0.0001523289, 0.0001465059, 0.0001287483, 0.0001201781, 0.0001155643, 
    0.0001053464, 0.0001056852, 0.0001062789, 0.0001114935, 0.0001096314, 
    0.0001053947, 0.0001157107, 0.0001214495, 0.0001260502, 0.0001275394, 
    0.0001331718, 0.0001297282, 0.0001362098, 0.0001476319,
  9.985224e-05, 9.818448e-05, 9.642545e-05, 8.842001e-05, 8.055176e-05, 
    7.600943e-05, 7.188954e-05, 6.962434e-05, 7.536724e-05, 8.817139e-05, 
    9.873931e-05, 9.372274e-05, 8.81611e-05, 8.011382e-05, 8.232534e-05, 
    7.951356e-05, 7.449454e-05, 7.559839e-05, 7.90405e-05, 8.380603e-05, 
    8.892811e-05, 8.775101e-05, 9.089857e-05, 9.257182e-05, 9.890284e-05, 
    9.984026e-05, 0.0001009929, 0.0001065726, 0.0001031663,
  2.940975e-05, 3.06821e-05, 2.924437e-05, 2.760597e-05, 2.381181e-05, 
    2.129335e-05, 1.79582e-05, 1.455696e-05, 1.246604e-05, 1.386442e-05, 
    1.919307e-05, 2.155402e-05, 2.686339e-05, 2.246577e-05, 1.975612e-05, 
    1.910273e-05, 1.827858e-05, 1.857958e-05, 1.773781e-05, 1.868666e-05, 
    2.008434e-05, 2.204074e-05, 2.322022e-05, 2.336581e-05, 2.429353e-05, 
    2.480501e-05, 2.459025e-05, 2.636431e-05, 2.782821e-05,
  4.657332e-06, 5.500008e-06, 4.644799e-06, 4.301738e-06, 4.29835e-06, 
    4.762327e-06, 4.431484e-06, 3.7659e-06, 2.956759e-06, 1.661766e-06, 
    1.551215e-06, 2.349619e-06, 3.599725e-06, 4.00672e-06, 3.576771e-06, 
    2.765312e-06, 2.800823e-06, 2.454486e-06, 2.705391e-06, 2.798859e-06, 
    2.179133e-06, 2.120781e-06, 2.161636e-06, 2.738104e-06, 3.472067e-06, 
    3.292845e-06, 4.064625e-06, 4.292532e-06, 4.240426e-06,
  8.713608e-07, 7.182032e-07, 7.003656e-07, 4.523389e-07, 3.808682e-07, 
    4.172144e-07, 4.022474e-07, 3.97518e-07, 4.758961e-07, 3.65848e-07, 
    2.501839e-07, 3.49001e-07, 5.327606e-07, 7.207331e-07, 9.973855e-07, 
    5.8072e-07, 6.667142e-07, 7.780121e-07, 7.48451e-07, 6.713821e-07, 
    5.979319e-07, 5.010478e-07, 4.495307e-07, 5.387317e-07, 5.736548e-07, 
    6.52559e-07, 6.990572e-07, 6.449443e-07, 7.718519e-07,
  3.812606e-07, 3.534955e-07, 2.58171e-07, 1.728989e-07, 1.468149e-07, 
    1.186587e-07, 1.334054e-07, 1.01957e-07, 9.632718e-08, 8.80321e-08, 
    8.457112e-08, 1.12514e-07, 1.961341e-07, 2.61244e-07, 3.762125e-07, 
    2.661305e-07, 2.30607e-07, 2.835963e-07, 3.066505e-07, 3.327446e-07, 
    5.300516e-07, 2.101594e-07, 1.233925e-07, 1.094499e-07, 1.228926e-07, 
    1.765743e-07, 2.652579e-07, 3.569533e-07, 4.416487e-07,
  1.399226e-07, 2.351021e-07, 2.183318e-07, 1.792664e-07, 1.094762e-07, 
    4.436249e-08, 2.684447e-08, 2.035171e-08, 1.942574e-08, 2.034669e-08, 
    2.445658e-08, 4.970251e-08, 1.096133e-07, 1.448873e-07, 1.83609e-07, 
    2.297223e-07, 2.432483e-07, 2.936701e-07, 2.667189e-07, 2.097594e-07, 
    1.114662e-07, 6.737277e-08, 4.940244e-08, 4.921847e-08, 8.042773e-08, 
    1.101497e-07, 1.180022e-07, 1.025635e-07, 9.488353e-08,
  2.968208e-08, 2.371813e-08, 1.559774e-08, 1.164079e-08, 1.040564e-08, 
    9.265791e-09, 8.869697e-09, 1.294054e-08, 1.973523e-08, 2.983754e-08, 
    3.918061e-08, 4.992997e-08, 6.573669e-08, 6.032472e-08, 4.568562e-08, 
    3.792593e-08, 3.394757e-08, 3.201162e-08, 3.017989e-08, 2.711279e-08, 
    2.448184e-08, 2.372164e-08, 2.847093e-08, 4.307459e-08, 6.263332e-08, 
    6.835497e-08, 5.593371e-08, 4.270297e-08, 3.325527e-08,
  1.791809e-08, 1.791809e-08, 1.791809e-08, 1.791809e-08, 1.791809e-08, 
    1.791809e-08, 1.791809e-08, 1.818239e-08, 1.818239e-08, 1.818239e-08, 
    1.818239e-08, 1.818239e-08, 1.818239e-08, 1.818239e-08, 1.926133e-08, 
    1.926133e-08, 1.926133e-08, 1.926133e-08, 1.926133e-08, 1.926133e-08, 
    1.926133e-08, 1.93107e-08, 1.93107e-08, 1.93107e-08, 1.93107e-08, 
    1.93107e-08, 1.93107e-08, 1.93107e-08, 1.791809e-08,
  2.71468e-08, 2.06764e-08, 1.588722e-08, 1.583925e-08, 1.636993e-08, 
    1.55509e-08, 1.543723e-08, 1.561616e-08, 1.709113e-08, 1.853268e-08, 
    2.084583e-08, 2.118746e-08, 2.214556e-08, 2.672878e-08, 5.273789e-08, 
    2.940147e-08, 2.908183e-08, 3.045029e-08, 3.081473e-08, 3.72896e-08, 
    4.286993e-08, 4.311036e-08, 4.001123e-08, 3.767905e-08, 3.424321e-08, 
    3.040942e-08, 2.559504e-08, 2.504835e-08, 2.705218e-08,
  6.412903e-08, 5.194434e-08, 4.545376e-08, 4.813239e-08, 5.360016e-08, 
    5.609579e-08, 6.031107e-08, 5.970351e-08, 5.088902e-08, 5.383848e-08, 
    5.572981e-08, 6.055124e-08, 1.090393e-07, 1.467877e-07, 1.941874e-07, 
    1.801971e-07, 1.913793e-07, 1.891713e-07, 1.601417e-07, 1.684422e-07, 
    1.354941e-07, 1.091857e-07, 9.149944e-08, 7.770522e-08, 7.578721e-08, 
    7.626685e-08, 7.758353e-08, 6.841617e-08, 5.634354e-08,
  3.82901e-07, 3.589969e-07, 3.263047e-07, 3.935411e-07, 4.912898e-07, 
    5.398541e-07, 4.739246e-07, 3.575797e-07, 2.859173e-07, 2.304546e-07, 
    2.294147e-07, 3.278062e-07, 4.364996e-07, 6.369309e-07, 7.078261e-07, 
    7.528109e-07, 7.90221e-07, 7.992745e-07, 6.701931e-07, 5.877399e-07, 
    5.25504e-07, 4.985325e-07, 4.384919e-07, 3.736747e-07, 4.700829e-07, 
    4.820592e-07, 4.05109e-07, 3.230183e-07, 3.661501e-07,
  1.732327e-06, 1.505687e-06, 1.565872e-06, 1.356308e-06, 1.442986e-06, 
    1.665509e-06, 1.581567e-06, 1.403382e-06, 1.206916e-06, 1.092674e-06, 
    1.173813e-06, 1.711668e-06, 2.241719e-06, 2.766398e-06, 2.819628e-06, 
    2.730269e-06, 1.912801e-06, 1.65234e-06, 1.588263e-06, 1.241192e-06, 
    1.001145e-06, 1.019268e-06, 1.59115e-06, 2.497012e-06, 2.71344e-06, 
    2.379472e-06, 1.907459e-06, 1.937359e-06, 1.71902e-06,
  6.857916e-06, 6.623152e-06, 7.046643e-06, 7.561587e-06, 8.523535e-06, 
    9.213892e-06, 9.145784e-06, 6.950218e-06, 6.972482e-06, 1.151969e-05, 
    1.903582e-05, 1.746378e-05, 1.239751e-05, 1.432153e-05, 1.367463e-05, 
    6.661901e-06, 5.843168e-06, 5.036706e-06, 5.717117e-06, 6.18176e-06, 
    6.742411e-06, 9.956975e-06, 1.593416e-05, 1.056281e-05, 1.172288e-05, 
    1.091463e-05, 1.12753e-05, 1.152976e-05, 8.087678e-06,
  7.103811e-05, 7.639545e-05, 6.941776e-05, 6.55863e-05, 7.07197e-05, 
    7.237397e-05, 7.593301e-05, 9.911447e-05, 0.0001149483, 0.0001222308, 
    0.0001089776, 8.430998e-05, 6.218026e-05, 4.870558e-05, 3.812617e-05, 
    3.202686e-05, 3.110211e-05, 3.454844e-05, 4.352513e-05, 5.355327e-05, 
    6.212266e-05, 6.323693e-05, 6.646346e-05, 6.853689e-05, 6.383812e-05, 
    5.991131e-05, 5.476456e-05, 5.528493e-05, 6.229966e-05,
  0.0005026255, 0.0005383856, 0.0005820679, 0.0005704137, 0.0005610148, 
    0.0005689244, 0.0005679756, 0.0005437363, 0.0005221288, 0.0004295447, 
    0.0003856705, 0.0003252951, 0.000272149, 0.0002586712, 0.0002678485, 
    0.0002761481, 0.0003029675, 0.0003036702, 0.0003183436, 0.0003460893, 
    0.0003542703, 0.0003641169, 0.0003803707, 0.0003802846, 0.0004071265, 
    0.0004322437, 0.0004603371, 0.0004787222, 0.0005012499,
  0.001071642, 0.00106212, 0.0009876871, 0.0009918702, 0.001064363, 
    0.001171776, 0.00125599, 0.001303133, 0.001282277, 0.00115828, 
    0.0009033677, 0.0008138836, 0.000749265, 0.0006991827, 0.00065105, 
    0.0006335598, 0.0006426464, 0.0006365438, 0.0006566491, 0.0006984479, 
    0.0007610882, 0.000832142, 0.0008558376, 0.0008330115, 0.0008013861, 
    0.0007774531, 0.0008378287, 0.0009353179, 0.00106509,
  0.0006047648, 0.0007455685, 0.0007247492, 0.0007058837, 0.0006994859, 
    0.0007444977, 0.0008282368, 0.0008764768, 0.001064545, 0.001093307, 
    0.001171024, 0.001128658, 0.001087982, 0.001067531, 0.0009490382, 
    0.0008556883, 0.0007478361, 0.000627317, 0.0005624818, 0.0005363121, 
    0.0005467079, 0.0006159827, 0.0006374991, 0.0006562482, 0.0006875644, 
    0.0006286713, 0.0006020621, 0.0005957494, 0.0005504105,
  0.0007526026, 0.0007280798, 0.0007090027, 0.0006703076, 0.0006267031, 
    0.0006839794, 0.0007078661, 0.0006807218, 0.0007370504, 0.0007786804, 
    0.0007827651, 0.0006932266, 0.0005779873, 0.0005164427, 0.0005006746, 
    0.0004733724, 0.0004696846, 0.0004554639, 0.0004644937, 0.0004779813, 
    0.0005187451, 0.0005391822, 0.0005579012, 0.0005303005, 0.0005226998, 
    0.0005442062, 0.0005865506, 0.0006476609, 0.0006974675,
  0.0005884529, 0.00058623, 0.0005917031, 0.000570021, 0.0005345077, 
    0.0004474689, 0.0003732447, 0.00033627, 0.0003260605, 0.0003536905, 
    0.0004658289, 0.0004274212, 0.0003710331, 0.0003394519, 0.0003504292, 
    0.0003489062, 0.0003250805, 0.0003097386, 0.0003272635, 0.0003589626, 
    0.0003807193, 0.0003803226, 0.0003867736, 0.0003964315, 0.0004266196, 
    0.0004598598, 0.0004855555, 0.0005397369, 0.0005826757,
  0.000183321, 0.0001779574, 0.0001736184, 0.0001680071, 0.0001597602, 
    0.0001567913, 0.0001302696, 9.941e-05, 8.10999e-05, 7.21846e-05, 
    7.560852e-05, 9.653856e-05, 0.0001130267, 9.730745e-05, 7.84834e-05, 
    7.634088e-05, 7.355274e-05, 7.123694e-05, 6.224653e-05, 6.450518e-05, 
    8.013757e-05, 7.83287e-05, 0.0001050197, 0.0001177911, 0.0001308745, 
    0.0001425841, 0.000146447, 0.0001570787, 0.0001695725,
  2.228268e-05, 2.965594e-05, 3.053874e-05, 2.864921e-05, 3.019737e-05, 
    2.677301e-05, 2.863411e-05, 2.60992e-05, 2.117658e-05, 1.262687e-05, 
    8.922665e-06, 1.073246e-05, 1.499926e-05, 1.607379e-05, 1.593766e-05, 
    1.322255e-05, 1.488649e-05, 1.265771e-05, 1.297617e-05, 1.599175e-05, 
    1.148205e-05, 8.786707e-06, 9.289798e-06, 1.063083e-05, 1.510112e-05, 
    1.520174e-05, 1.740568e-05, 2.024331e-05, 2.191513e-05,
  3.657796e-06, 3.619326e-06, 3.649004e-06, 2.619923e-06, 1.770385e-06, 
    1.77429e-06, 1.942504e-06, 2.280844e-06, 2.208107e-06, 2.393163e-06, 
    1.728832e-06, 1.499407e-06, 2.267973e-06, 2.728625e-06, 3.708777e-06, 
    3.462623e-06, 3.527794e-06, 4.38959e-06, 3.949958e-06, 3.406925e-06, 
    3.317997e-06, 2.200226e-06, 1.631638e-06, 2.064834e-06, 2.506105e-06, 
    2.695379e-06, 3.082878e-06, 3.131942e-06, 3.520087e-06,
  1.548222e-06, 1.361687e-06, 1.015827e-06, 7.285617e-07, 5.666636e-07, 
    4.345245e-07, 4.60977e-07, 3.992393e-07, 3.386461e-07, 4.285066e-07, 
    4.028844e-07, 4.391459e-07, 8.109528e-07, 9.381466e-07, 1.318083e-06, 
    1.213475e-06, 1.039992e-06, 1.352063e-06, 1.520501e-06, 1.642018e-06, 
    1.7372e-06, 9.846052e-07, 3.991157e-07, 4.011842e-07, 4.595964e-07, 
    7.182707e-07, 9.687486e-07, 1.31252e-06, 1.543847e-06,
  4.830134e-07, 5.667947e-07, 5.80221e-07, 4.917657e-07, 3.286951e-07, 
    1.811315e-07, 1.085573e-07, 7.484342e-08, 6.720605e-08, 7.023712e-08, 
    1.056242e-07, 1.597987e-07, 3.20429e-07, 4.752983e-07, 5.540907e-07, 
    6.237195e-07, 7.084175e-07, 8.503073e-07, 7.467443e-07, 5.964078e-07, 
    3.659842e-07, 1.861406e-07, 1.641133e-07, 1.762777e-07, 2.51009e-07, 
    3.081943e-07, 3.482979e-07, 3.948116e-07, 4.209622e-07,
  1.024337e-07, 1.022907e-07, 9.612882e-08, 7.25325e-08, 6.312586e-08, 
    5.973508e-08, 5.605207e-08, 6.391955e-08, 7.219843e-08, 7.569618e-08, 
    8.377786e-08, 1.037992e-07, 1.429335e-07, 1.741267e-07, 1.844704e-07, 
    1.511173e-07, 1.274789e-07, 1.131945e-07, 1.029519e-07, 9.810611e-08, 
    9.798986e-08, 1.009697e-07, 1.180808e-07, 1.447855e-07, 1.829271e-07, 
    1.755461e-07, 1.425079e-07, 1.227551e-07, 1.090297e-07,
  9.061949e-08, 9.061949e-08, 9.061949e-08, 9.061949e-08, 9.061949e-08, 
    9.061949e-08, 9.061949e-08, 9.504182e-08, 9.504182e-08, 9.504182e-08, 
    9.504182e-08, 9.504182e-08, 9.504182e-08, 9.504182e-08, 1.008396e-07, 
    1.008396e-07, 1.008396e-07, 1.008396e-07, 1.008396e-07, 1.008396e-07, 
    1.008396e-07, 9.794519e-08, 9.794519e-08, 9.794519e-08, 9.794519e-08, 
    9.794519e-08, 9.794519e-08, 9.794519e-08, 9.061949e-08,
  1.183366e-07, 1.092687e-07, 8.644223e-08, 9.670116e-08, 1.082746e-07, 
    1.026963e-07, 9.667684e-08, 8.022158e-08, 8.947291e-08, 9.383368e-08, 
    1.322908e-07, 1.327722e-07, 1.162118e-07, 1.247042e-07, 2.332239e-07, 
    1.853548e-07, 1.735948e-07, 1.829824e-07, 1.710654e-07, 1.665762e-07, 
    1.703526e-07, 1.744074e-07, 1.647739e-07, 1.555777e-07, 1.391508e-07, 
    1.217627e-07, 1.047012e-07, 9.912244e-08, 1.148166e-07,
  1.870818e-07, 1.943856e-07, 2.077866e-07, 1.959021e-07, 2.436256e-07, 
    2.936226e-07, 2.757191e-07, 2.48388e-07, 2.229938e-07, 2.240376e-07, 
    2.417164e-07, 3.098695e-07, 4.480865e-07, 5.556531e-07, 9.805083e-07, 
    9.829614e-07, 1.022348e-06, 1.045296e-06, 7.201036e-07, 7.688625e-07, 
    6.428862e-07, 4.897621e-07, 4.132352e-07, 3.491918e-07, 3.284463e-07, 
    3.301319e-07, 3.175439e-07, 2.685258e-07, 2.050658e-07,
  1.535192e-06, 1.400418e-06, 1.273354e-06, 1.434005e-06, 1.948109e-06, 
    2.228074e-06, 1.854644e-06, 1.577104e-06, 1.256233e-06, 9.634008e-07, 
    8.581546e-07, 1.010342e-06, 1.775504e-06, 2.79732e-06, 3.347656e-06, 
    3.50649e-06, 3.805822e-06, 3.575681e-06, 3.376903e-06, 2.406305e-06, 
    1.943782e-06, 1.636042e-06, 1.578325e-06, 1.506922e-06, 1.963673e-06, 
    2.081883e-06, 1.852666e-06, 1.572295e-06, 1.5099e-06,
  7.986347e-06, 6.507472e-06, 6.132796e-06, 5.871644e-06, 6.370186e-06, 
    6.983778e-06, 8.062311e-06, 6.445098e-06, 5.345873e-06, 4.347525e-06, 
    4.729688e-06, 6.727566e-06, 9.759612e-06, 1.173353e-05, 1.415931e-05, 
    1.382086e-05, 1.077748e-05, 8.241486e-06, 8.742946e-06, 6.489266e-06, 
    5.267496e-06, 4.94611e-06, 6.671981e-06, 1.008199e-05, 1.173044e-05, 
    1.078435e-05, 8.86925e-06, 8.378336e-06, 7.944509e-06,
  3.741634e-05, 3.791827e-05, 3.38436e-05, 3.390461e-05, 3.778507e-05, 
    4.952046e-05, 4.355112e-05, 3.264962e-05, 2.844092e-05, 4.520891e-05, 
    8.451742e-05, 9.483779e-05, 7.57174e-05, 6.649122e-05, 8.600955e-05, 
    3.835044e-05, 3.151619e-05, 3.04522e-05, 3.293849e-05, 2.933393e-05, 
    2.925619e-05, 3.861019e-05, 5.479786e-05, 6.9663e-05, 6.655179e-05, 
    5.197664e-05, 4.449458e-05, 4.712892e-05, 4.178297e-05,
  0.0002812668, 0.0002968236, 0.0002915395, 0.0003035218, 0.0003155148, 
    0.000320948, 0.0003376384, 0.0004148333, 0.0005753012, 0.0006213234, 
    0.0006693253, 0.000555969, 0.0003913532, 0.000297907, 0.0002745816, 
    0.0001832956, 0.0001436544, 0.0001432917, 0.0001606979, 0.0002043622, 
    0.0002629138, 0.0003165119, 0.0003115912, 0.000324391, 0.0002765596, 
    0.0002445896, 0.0002240731, 0.0002162061, 0.0002281069,
  0.002071399, 0.002154562, 0.00233518, 0.002522249, 0.002652827, 
    0.002715019, 0.003024712, 0.003130569, 0.002813086, 0.002351175, 
    0.002011224, 0.001767193, 0.001374527, 0.001099443, 0.0009950747, 
    0.0009153487, 0.000909667, 0.001088204, 0.001161366, 0.001303012, 
    0.00157965, 0.001729015, 0.001457861, 0.001359583, 0.001266419, 
    0.001271339, 0.001592037, 0.001800822, 0.002040705,
  0.004497685, 0.004729622, 0.00488846, 0.004848433, 0.005126763, 
    0.005760604, 0.006355843, 0.006443349, 0.006571122, 0.005858281, 
    0.004914318, 0.003664161, 0.003115234, 0.002726856, 0.002654261, 
    0.002421972, 0.002267489, 0.002483597, 0.00263953, 0.003175858, 
    0.003553526, 0.003769014, 0.003829744, 0.003462756, 0.003369475, 
    0.003559868, 0.003720439, 0.004276456, 0.004342408,
  0.002868561, 0.003381341, 0.003187185, 0.002918705, 0.003035189, 
    0.003248068, 0.003375265, 0.004118864, 0.005036579, 0.006403663, 
    0.006491314, 0.006276541, 0.005332251, 0.003793914, 0.003211306, 
    0.002733702, 0.002459809, 0.002291036, 0.002533001, 0.002637718, 
    0.002561903, 0.002922314, 0.003134214, 0.00314685, 0.003194603, 
    0.003010041, 0.003013289, 0.002835523, 0.002851326,
  0.003244642, 0.003594751, 0.003545063, 0.00332352, 0.003368918, 
    0.003573818, 0.00316511, 0.003235193, 0.003523904, 0.004310485, 
    0.003800378, 0.002903585, 0.002491385, 0.002097087, 0.002035358, 
    0.002015273, 0.002005291, 0.001924923, 0.002134632, 0.002149322, 
    0.002269077, 0.002306136, 0.002460561, 0.002584083, 0.002584049, 
    0.002357796, 0.002365405, 0.002823751, 0.003120565,
  0.002698024, 0.002790766, 0.003209459, 0.003314377, 0.003430093, 
    0.003107162, 0.002646887, 0.001970077, 0.001718503, 0.001707382, 
    0.002198266, 0.001943465, 0.001537134, 0.001361568, 0.001309345, 
    0.001292506, 0.001139148, 0.001057618, 0.001091168, 0.001287549, 
    0.001330885, 0.00147991, 0.001504803, 0.001605722, 0.001712159, 
    0.001710818, 0.001810459, 0.002056555, 0.002373994,
  0.0009371924, 0.001102091, 0.001164961, 0.001145079, 0.001085605, 
    0.001108943, 0.001127533, 0.000778069, 0.0006023013, 0.0004354126, 
    0.0003609943, 0.0004698857, 0.0005768019, 0.0004504048, 0.0003400808, 
    0.0002740051, 0.0002927695, 0.0002631601, 0.0002364141, 0.0002453063, 
    0.0002860482, 0.0002486167, 0.0003184114, 0.0004338168, 0.00047294, 
    0.0005158493, 0.0005969657, 0.0006773862, 0.0007824798,
  0.000131433, 0.0001586027, 0.0001765275, 0.0001704433, 0.0001935799, 
    0.0001903382, 0.0001895641, 0.0001958452, 0.0001420017, 9.637146e-05, 
    5.616056e-05, 5.789784e-05, 6.877448e-05, 6.7075e-05, 6.069476e-05, 
    5.297246e-05, 5.644279e-05, 5.470807e-05, 5.666544e-05, 7.524589e-05, 
    6.272626e-05, 4.428726e-05, 3.5793e-05, 4.390581e-05, 5.36355e-05, 
    6.186822e-05, 8.305036e-05, 9.672964e-05, 0.0001197078,
  1.539331e-05, 1.667773e-05, 1.942214e-05, 1.892974e-05, 1.062616e-05, 
    6.999628e-06, 9.249211e-06, 1.184091e-05, 1.33681e-05, 1.419267e-05, 
    1.260847e-05, 8.214353e-06, 1.104361e-05, 1.297116e-05, 1.32141e-05, 
    1.331933e-05, 1.307987e-05, 1.620233e-05, 1.646364e-05, 1.619506e-05, 
    1.519044e-05, 9.952602e-06, 6.302261e-06, 6.538516e-06, 9.907004e-06, 
    1.039408e-05, 1.203376e-05, 1.454319e-05, 1.630504e-05,
  7.135474e-06, 5.528878e-06, 3.838366e-06, 2.837922e-06, 2.376901e-06, 
    1.800359e-06, 1.722979e-06, 1.792648e-06, 1.652616e-06, 2.052357e-06, 
    2.343533e-06, 2.734769e-06, 3.246596e-06, 3.369252e-06, 4.520386e-06, 
    4.188271e-06, 4.497398e-06, 5.389119e-06, 6.467757e-06, 6.560084e-06, 
    5.362871e-06, 3.416598e-06, 1.669052e-06, 1.617858e-06, 1.898325e-06, 
    2.945603e-06, 4.452419e-06, 5.174924e-06, 5.564161e-06,
  1.695786e-06, 2.192612e-06, 2.592085e-06, 1.669902e-06, 8.529676e-07, 
    5.668206e-07, 4.294734e-07, 3.699758e-07, 3.765234e-07, 4.68659e-07, 
    6.515388e-07, 7.302112e-07, 1.027027e-06, 1.491808e-06, 1.488333e-06, 
    1.79731e-06, 1.869135e-06, 2.169892e-06, 2.178339e-06, 1.98081e-06, 
    1.322376e-06, 6.755853e-07, 6.739481e-07, 7.298665e-07, 8.371218e-07, 
    1.012181e-06, 1.297219e-06, 1.604642e-06, 1.612607e-06,
  3.971998e-07, 3.840788e-07, 3.948661e-07, 3.48236e-07, 2.818892e-07, 
    2.661642e-07, 2.263666e-07, 2.17107e-07, 1.922862e-07, 1.98382e-07, 
    2.274467e-07, 2.683327e-07, 3.516147e-07, 4.376369e-07, 4.76174e-07, 
    4.692602e-07, 4.332043e-07, 3.911677e-07, 3.702059e-07, 3.778342e-07, 
    3.781343e-07, 3.758464e-07, 3.769659e-07, 4.088743e-07, 4.625193e-07, 
    4.42733e-07, 3.993491e-07, 3.922073e-07, 3.969847e-07,
  3.910738e-07, 3.910738e-07, 3.910738e-07, 3.910738e-07, 3.910738e-07, 
    3.910738e-07, 3.910738e-07, 4.346903e-07, 4.346903e-07, 4.346903e-07, 
    4.346903e-07, 4.346903e-07, 4.346903e-07, 4.346903e-07, 4.632075e-07, 
    4.632075e-07, 4.632075e-07, 4.632075e-07, 4.632075e-07, 4.632075e-07, 
    4.632075e-07, 4.265738e-07, 4.265738e-07, 4.265738e-07, 4.265738e-07, 
    4.265738e-07, 4.265738e-07, 4.265738e-07, 3.910738e-07,
  4.410547e-07, 4.059652e-07, 3.454443e-07, 3.707498e-07, 4.535263e-07, 
    5.569883e-07, 5.969354e-07, 5.366724e-07, 4.468295e-07, 4.404915e-07, 
    4.687868e-07, 5.444889e-07, 7.663212e-07, 1.013941e-06, 1.288082e-06, 
    1.372039e-06, 1.251338e-06, 1.191726e-06, 1.089913e-06, 9.411962e-07, 
    8.410308e-07, 8.108173e-07, 7.925929e-07, 7.254269e-07, 6.105645e-07, 
    5.390531e-07, 4.749809e-07, 4.308712e-07, 4.226821e-07,
  6.564947e-07, 5.314922e-07, 6.239518e-07, 7.81848e-07, 1.035939e-06, 
    1.281981e-06, 1.211109e-06, 1.028227e-06, 8.164123e-07, 7.535356e-07, 
    8.072277e-07, 9.428992e-07, 1.27212e-06, 2.778307e-06, 3.79419e-06, 
    5.39071e-06, 5.668851e-06, 4.683456e-06, 3.446616e-06, 2.805966e-06, 
    2.351554e-06, 2.108586e-06, 2.099371e-06, 1.83811e-06, 1.981497e-06, 
    1.833074e-06, 1.631059e-06, 1.212869e-06, 8.763192e-07,
  6.018156e-06, 6.378437e-06, 6.040689e-06, 5.850732e-06, 6.670659e-06, 
    7.165407e-06, 6.364396e-06, 5.516777e-06, 4.715578e-06, 3.859479e-06, 
    3.337339e-06, 3.940345e-06, 6.515131e-06, 1.119058e-05, 1.7661e-05, 
    1.813035e-05, 2.026597e-05, 2.031539e-05, 1.662898e-05, 1.073954e-05, 
    8.184882e-06, 6.669129e-06, 5.974003e-06, 6.043207e-06, 7.841105e-06, 
    8.248429e-06, 8.418458e-06, 7.514509e-06, 6.360896e-06,
  3.432363e-05, 2.821878e-05, 2.587908e-05, 2.520565e-05, 2.711136e-05, 
    2.787074e-05, 3.402031e-05, 3.059135e-05, 2.542516e-05, 1.957701e-05, 
    2.1059e-05, 2.908908e-05, 4.625833e-05, 5.300336e-05, 7.620621e-05, 
    6.853922e-05, 4.550812e-05, 4.640307e-05, 4.385228e-05, 3.037128e-05, 
    2.646901e-05, 2.319317e-05, 2.595895e-05, 4.356681e-05, 4.855556e-05, 
    4.756626e-05, 4.401184e-05, 3.870526e-05, 3.605364e-05,
  0.0001716195, 0.0001544989, 0.0001434452, 0.0001480508, 0.0001709666, 
    0.0001872034, 0.0001967104, 0.000146761, 0.000137919, 0.0002027993, 
    0.0003198586, 0.0003999034, 0.000388052, 0.0003341132, 0.000540648, 
    0.0002270332, 0.0001686041, 0.0001547117, 0.0001387703, 0.0001245034, 
    0.0001313816, 0.0001730224, 0.0001949101, 0.0003464979, 0.0003653903, 
    0.0002624048, 0.0001921074, 0.0001956831, 0.0001832964,
  0.001118709, 0.001272899, 0.001227609, 0.00128652, 0.001607117, 
    0.001290808, 0.001588521, 0.002215034, 0.002697919, 0.003440364, 
    0.004673822, 0.004852229, 0.002895876, 0.001957626, 0.001367881, 
    0.001168232, 0.0007514696, 0.0005899513, 0.0006536777, 0.000857694, 
    0.001126852, 0.001312064, 0.001626181, 0.001765268, 0.001594834, 
    0.001029622, 0.0009818558, 0.0008410643, 0.0008671722,
  0.007452739, 0.007185334, 0.007255337, 0.007966638, 0.009564025, 
    0.01102051, 0.01415402, 0.01759347, 0.02027783, 0.01725335, 0.01446331, 
    0.01341225, 0.01027388, 0.008289333, 0.005738638, 0.005053023, 
    0.003840068, 0.003073005, 0.003585742, 0.003997945, 0.005245731, 
    0.007592754, 0.008416506, 0.006877793, 0.00605247, 0.00414311, 
    0.004422022, 0.005792944, 0.006932247,
  0.01949148, 0.01942202, 0.01879972, 0.01931803, 0.02056898, 0.02282324, 
    0.02779266, 0.03279817, 0.03740406, 0.03501067, 0.02806137, 0.02366241, 
    0.02009042, 0.01771023, 0.01470585, 0.01308398, 0.01090956, 0.008988741, 
    0.009025245, 0.01249249, 0.01692722, 0.0203417, 0.02102949, 0.01825234, 
    0.01431263, 0.01354813, 0.01475771, 0.01759778, 0.01968597,
  0.01883477, 0.01788144, 0.01510716, 0.01473064, 0.01403649, 0.01595392, 
    0.01686907, 0.02022485, 0.02544972, 0.03186211, 0.03182641, 0.03069232, 
    0.02319022, 0.01779361, 0.01542486, 0.01405365, 0.0120863, 0.01133122, 
    0.01137725, 0.0145683, 0.01790944, 0.01689817, 0.01739926, 0.01635698, 
    0.01540127, 0.01461672, 0.01567126, 0.01615849, 0.01898404,
  0.01562633, 0.01683931, 0.0184469, 0.01833703, 0.01968504, 0.020882, 
    0.01911842, 0.01998535, 0.01992125, 0.02353803, 0.02041527, 0.01671008, 
    0.01556379, 0.01347362, 0.01234358, 0.01103908, 0.01015956, 0.009072511, 
    0.009446359, 0.01033969, 0.01200114, 0.01129426, 0.01050755, 0.01076099, 
    0.01146, 0.01204741, 0.01271583, 0.01370907, 0.01431638,
  0.01021313, 0.01301803, 0.01490443, 0.0162467, 0.01720472, 0.01885353, 
    0.01647976, 0.01323888, 0.01028658, 0.009590394, 0.0109035, 0.009083379, 
    0.007991472, 0.007261583, 0.006036533, 0.005257403, 0.004842893, 
    0.003905069, 0.003514645, 0.003896781, 0.004550443, 0.005473833, 
    0.005732589, 0.006468038, 0.006888149, 0.006929707, 0.007377981, 
    0.007389418, 0.008315637,
  0.00317433, 0.00424039, 0.005828946, 0.005999609, 0.007327912, 0.007179089, 
    0.007489548, 0.006688286, 0.004373177, 0.003385531, 0.002410407, 
    0.002471105, 0.002871429, 0.002232208, 0.00154132, 0.001189842, 
    0.001226444, 0.001113727, 0.001026412, 0.001056627, 0.001200857, 
    0.001051757, 0.001033433, 0.001308283, 0.001539912, 0.00167278, 
    0.001948298, 0.002059228, 0.002656515,
  0.0005518539, 0.0007674319, 0.0009016304, 0.0008303613, 0.001033843, 
    0.001098663, 0.001227856, 0.001287221, 0.0009601003, 0.0006499632, 
    0.0004737366, 0.0003026572, 0.0003572621, 0.0003407757, 0.0002597884, 
    0.0002040338, 0.0001998108, 0.0002136656, 0.0002505227, 0.0003110338, 
    0.0003317869, 0.0002590406, 0.0001706229, 0.0001639861, 0.0001921534, 
    0.0002001163, 0.0002640757, 0.0003823443, 0.0004659991,
  6.226839e-05, 7.84029e-05, 9.750402e-05, 9.573129e-05, 6.901319e-05, 
    3.774286e-05, 4.322815e-05, 5.532237e-05, 8.421734e-05, 6.662794e-05, 
    8.407434e-05, 5.780928e-05, 4.773463e-05, 6.957959e-05, 6.671669e-05, 
    5.625657e-05, 5.122814e-05, 6.244919e-05, 6.065466e-05, 7.200114e-05, 
    7.351435e-05, 5.572894e-05, 2.779416e-05, 2.781808e-05, 3.791445e-05, 
    3.989022e-05, 4.06105e-05, 5.721488e-05, 6.425974e-05,
  2.500319e-05, 2.724267e-05, 1.510465e-05, 1.233129e-05, 9.113277e-06, 
    9.459781e-06, 7.473139e-06, 6.804735e-06, 7.903566e-06, 8.8795e-06, 
    1.110754e-05, 1.652362e-05, 1.652752e-05, 1.666535e-05, 1.539392e-05, 
    1.522676e-05, 1.816694e-05, 1.989695e-05, 2.457782e-05, 2.346965e-05, 
    1.790096e-05, 1.001501e-05, 6.665911e-06, 6.620216e-06, 8.158062e-06, 
    1.232738e-05, 2.21782e-05, 2.628829e-05, 2.288353e-05,
  6.439181e-06, 8.988295e-06, 9.919502e-06, 6.22791e-06, 3.213823e-06, 
    2.104068e-06, 1.740643e-06, 1.579474e-06, 1.80591e-06, 1.895879e-06, 
    3.047129e-06, 3.363233e-06, 4.183748e-06, 5.126863e-06, 4.884214e-06, 
    5.626297e-06, 5.375781e-06, 6.884164e-06, 6.497512e-06, 5.455167e-06, 
    4.289705e-06, 3.080861e-06, 3.073024e-06, 3.350719e-06, 3.640816e-06, 
    4.179469e-06, 5.615425e-06, 6.021293e-06, 5.803793e-06,
  1.63077e-06, 1.55808e-06, 1.447771e-06, 1.394828e-06, 1.315658e-06, 
    1.208028e-06, 1.070629e-06, 8.991969e-07, 7.342558e-07, 7.753026e-07, 
    8.380801e-07, 9.493882e-07, 1.176211e-06, 1.316424e-06, 1.362318e-06, 
    1.427366e-06, 1.499602e-06, 1.483195e-06, 1.385069e-06, 1.333658e-06, 
    1.298451e-06, 1.332123e-06, 1.334408e-06, 1.322082e-06, 1.209641e-06, 
    1.172352e-06, 1.210525e-06, 1.329408e-06, 1.556482e-06,
  1.3234e-06, 1.3234e-06, 1.3234e-06, 1.3234e-06, 1.3234e-06, 1.3234e-06, 
    1.3234e-06, 1.366308e-06, 1.366308e-06, 1.366308e-06, 1.366308e-06, 
    1.366308e-06, 1.366308e-06, 1.366308e-06, 1.513811e-06, 1.513811e-06, 
    1.513811e-06, 1.513811e-06, 1.513811e-06, 1.513811e-06, 1.513811e-06, 
    1.467425e-06, 1.467425e-06, 1.467425e-06, 1.467425e-06, 1.467425e-06, 
    1.467425e-06, 1.467425e-06, 1.3234e-06,
  1.73945e-06, 1.61254e-06, 1.46913e-06, 1.730807e-06, 1.964488e-06, 
    2.177181e-06, 2.538739e-06, 2.670899e-06, 2.31698e-06, 2.199701e-06, 
    2.350039e-06, 2.599399e-06, 2.865291e-06, 3.424765e-06, 4.304818e-06, 
    5.048229e-06, 4.841793e-06, 4.27177e-06, 3.9777e-06, 3.757532e-06, 
    3.800109e-06, 3.911997e-06, 3.826141e-06, 3.434695e-06, 2.845934e-06, 
    2.438788e-06, 2.097874e-06, 1.770059e-06, 1.697566e-06,
  3.287275e-06, 2.378988e-06, 2.378023e-06, 2.878243e-06, 3.815531e-06, 
    5.362547e-06, 5.388747e-06, 4.706076e-06, 3.562273e-06, 3.113219e-06, 
    3.266542e-06, 3.61013e-06, 4.425086e-06, 8.3503e-06, 1.46787e-05, 
    2.345562e-05, 2.565633e-05, 2.16652e-05, 1.734747e-05, 1.332399e-05, 
    1.163178e-05, 1.032391e-05, 9.512472e-06, 8.584278e-06, 1.056051e-05, 
    9.124326e-06, 8.168905e-06, 5.629962e-06, 3.957565e-06,
  2.090809e-05, 2.240924e-05, 2.052563e-05, 2.143625e-05, 2.110561e-05, 
    2.238731e-05, 2.099206e-05, 1.848991e-05, 1.754392e-05, 1.400186e-05, 
    1.211663e-05, 1.383097e-05, 2.150254e-05, 3.591165e-05, 6.551049e-05, 
    8.338291e-05, 8.591395e-05, 8.552925e-05, 7.318983e-05, 5.108154e-05, 
    3.717578e-05, 2.90078e-05, 2.376136e-05, 2.625363e-05, 3.021772e-05, 
    3.086755e-05, 3.087871e-05, 2.845208e-05, 2.485613e-05,
  0.000123171, 0.0001154735, 0.0001034988, 0.000100648, 0.0001157453, 
    0.0001069807, 0.0001423976, 0.0001380726, 0.0001302426, 0.0001093178, 
    0.0001005933, 0.0001387939, 0.0002010928, 0.0002454243, 0.0003020799, 
    0.0002892675, 0.0001940102, 0.0002144406, 0.0001779244, 0.0001580891, 
    0.0001338528, 0.0001063197, 9.83225e-05, 0.0001439203, 0.000173724, 
    0.0001916313, 0.0001690238, 0.0001527818, 0.0001288559,
  0.0006285995, 0.0005967958, 0.0006349491, 0.0006961833, 0.0006845467, 
    0.0008061209, 0.0007367617, 0.0007283798, 0.0005980674, 0.0008332891, 
    0.001533378, 0.001832879, 0.00211175, 0.001634158, 0.002085424, 
    0.001120913, 0.000726097, 0.0007422671, 0.0005599044, 0.0005682221, 
    0.0005358777, 0.000627319, 0.0007599611, 0.001224598, 0.001425326, 
    0.001008129, 0.0008468765, 0.0006668367, 0.0006738735,
  0.004124932, 0.005404924, 0.005846321, 0.005020593, 0.009866067, 
    0.00761139, 0.00619548, 0.009660126, 0.01291215, 0.02138877, 0.03486179, 
    0.03442677, 0.02145248, 0.01155157, 0.00844209, 0.005824681, 0.004163191, 
    0.002999574, 0.002587633, 0.003240239, 0.004173159, 0.004216204, 
    0.006772719, 0.007720848, 0.008215923, 0.004494862, 0.003742609, 
    0.003188898, 0.00346851,
  0.02954921, 0.03007048, 0.02874692, 0.03045371, 0.03567606, 0.04204634, 
    0.05392737, 0.0825033, 0.1158382, 0.1422217, 0.1415511, 0.1288542, 
    0.09839997, 0.07114491, 0.05067324, 0.04425953, 0.0323385, 0.01735658, 
    0.0131019, 0.01378914, 0.01866686, 0.02604187, 0.03191096, 0.03731759, 
    0.03031764, 0.02249082, 0.01455873, 0.01761421, 0.02535304,
  0.08344446, 0.08918867, 0.07647, 0.06558863, 0.07446221, 0.07746589, 
    0.1070147, 0.1397832, 0.1912298, 0.1917906, 0.1772437, 0.1740642, 
    0.1674481, 0.1503732, 0.1203922, 0.09395126, 0.0834659, 0.05517508, 
    0.04103266, 0.03743289, 0.05665835, 0.07568156, 0.09006109, 0.1046428, 
    0.08383802, 0.06213288, 0.04976743, 0.05689393, 0.07387655,
  0.09771463, 0.08595162, 0.07767142, 0.0637164, 0.06465667, 0.06834033, 
    0.07931276, 0.1026997, 0.1260133, 0.1516786, 0.149469, 0.1268075, 
    0.1080788, 0.1143854, 0.1009645, 0.08859338, 0.06962825, 0.05814754, 
    0.04804625, 0.05217496, 0.07042608, 0.09095672, 0.08786, 0.07548781, 
    0.06407022, 0.06044358, 0.05565878, 0.06473558, 0.08075333,
  0.08105019, 0.08955313, 0.09600978, 0.1175539, 0.1107196, 0.1061723, 
    0.1088132, 0.1198286, 0.1275552, 0.1385208, 0.1197676, 0.101732, 
    0.09987725, 0.1023896, 0.08434328, 0.0687878, 0.06262485, 0.0545673, 
    0.04784694, 0.04772657, 0.05598434, 0.05480087, 0.04382125, 0.04107906, 
    0.03891033, 0.0391788, 0.04691132, 0.05769989, 0.07044402,
  0.04996426, 0.07346113, 0.09182876, 0.1332652, 0.1518865, 0.1455325, 
    0.134312, 0.1172746, 0.1003414, 0.07344613, 0.06344508, 0.05689697, 
    0.04943045, 0.04365898, 0.03240657, 0.02655828, 0.02558435, 0.02111807, 
    0.01809187, 0.01858248, 0.01921338, 0.02113384, 0.01978041, 0.02074282, 
    0.02083634, 0.0206275, 0.02398067, 0.03093991, 0.03910503,
  0.01517344, 0.01934489, 0.03282657, 0.03965298, 0.04470644, 0.05103618, 
    0.0651328, 0.05514346, 0.04131472, 0.02256236, 0.01594264, 0.01455472, 
    0.01496147, 0.01147989, 0.00695509, 0.004982351, 0.005141952, 
    0.004762025, 0.005317635, 0.006725546, 0.006559984, 0.006124514, 
    0.004508431, 0.004094, 0.004184844, 0.005186001, 0.005626538, 
    0.006319284, 0.008882782,
  0.001874969, 0.002907493, 0.00362826, 0.003767324, 0.004477799, 
    0.004401552, 0.005472181, 0.006458018, 0.005599887, 0.003823362, 
    0.00301129, 0.001927105, 0.001735026, 0.001618658, 0.00130872, 
    0.0008241594, 0.0007035352, 0.000840188, 0.00102026, 0.001506633, 
    0.00173375, 0.001589658, 0.000949108, 0.0006637887, 0.0006383574, 
    0.000585922, 0.0006643576, 0.001228459, 0.001545837,
  0.0002396338, 0.0002465136, 0.0003116334, 0.0003613248, 0.0004275852, 
    0.0001795877, 0.0002033644, 0.0002557764, 0.0003749822, 0.0003922429, 
    0.0004625626, 0.000424381, 0.0002794083, 0.0003092937, 0.0002841264, 
    0.0002759667, 0.0002315426, 0.0002580775, 0.0002436767, 0.0002884789, 
    0.0003039551, 0.0002520822, 0.0001363594, 0.0001138526, 0.0001448213, 
    0.0001625672, 0.0001689453, 0.0001775228, 0.0002442508,
  8.080937e-05, 8.451218e-05, 6.807793e-05, 5.012442e-05, 3.997398e-05, 
    5.001961e-05, 3.859799e-05, 2.805607e-05, 2.761326e-05, 5.07486e-05, 
    4.441156e-05, 6.845007e-05, 8.535261e-05, 8.29379e-05, 5.45402e-05, 
    5.674642e-05, 7.61559e-05, 7.787342e-05, 8.680955e-05, 7.166424e-05, 
    5.746049e-05, 3.657447e-05, 2.69047e-05, 2.573869e-05, 3.403872e-05, 
    4.719462e-05, 7.948512e-05, 9.640151e-05, 7.466049e-05,
  2.30036e-05, 2.869851e-05, 2.842404e-05, 2.219352e-05, 1.604142e-05, 
    1.227224e-05, 9.397685e-06, 8.004704e-06, 1.48857e-05, 1.190742e-05, 
    1.084451e-05, 1.620168e-05, 2.099505e-05, 1.937552e-05, 1.941819e-05, 
    1.800821e-05, 1.924095e-05, 2.127068e-05, 2.041138e-05, 1.798158e-05, 
    1.495376e-05, 1.325863e-05, 1.182677e-05, 1.396973e-05, 1.551746e-05, 
    1.86572e-05, 2.431577e-05, 2.688413e-05, 2.128355e-05,
  5.123246e-06, 5.314817e-06, 4.751331e-06, 4.490432e-06, 4.790541e-06, 
    4.772239e-06, 4.613094e-06, 4.06555e-06, 3.492023e-06, 3.406995e-06, 
    3.428612e-06, 3.756245e-06, 4.216111e-06, 4.564802e-06, 4.947768e-06, 
    5.943522e-06, 6.318757e-06, 6.492091e-06, 6.469404e-06, 5.991557e-06, 
    5.639042e-06, 5.685768e-06, 5.864757e-06, 5.754404e-06, 5.116541e-06, 
    4.661605e-06, 4.106047e-06, 4.402501e-06, 4.943079e-06,
  4.982602e-06, 4.982602e-06, 4.982602e-06, 4.982602e-06, 4.982602e-06, 
    4.982602e-06, 4.982602e-06, 5.526211e-06, 5.526211e-06, 5.526211e-06, 
    5.526211e-06, 5.526211e-06, 5.526211e-06, 5.526211e-06, 6.526013e-06, 
    6.526013e-06, 6.526013e-06, 6.526013e-06, 6.526013e-06, 6.526013e-06, 
    6.526013e-06, 6.171131e-06, 6.171131e-06, 6.171131e-06, 6.171131e-06, 
    6.171131e-06, 6.171131e-06, 6.171131e-06, 4.982602e-06,
  7.986441e-06, 6.262919e-06, 5.278067e-06, 6.065005e-06, 6.644432e-06, 
    6.996243e-06, 8.209572e-06, 9.007616e-06, 9.699518e-06, 9.547504e-06, 
    9.963617e-06, 1.009874e-05, 1.059738e-05, 1.144293e-05, 1.542506e-05, 
    1.836236e-05, 1.784009e-05, 1.603312e-05, 1.352798e-05, 1.208636e-05, 
    1.205889e-05, 1.376547e-05, 1.388367e-05, 1.286958e-05, 1.074097e-05, 
    9.673255e-06, 8.916053e-06, 8.634237e-06, 8.115997e-06,
  1.292433e-05, 1.076493e-05, 1.021004e-05, 1.205192e-05, 1.556489e-05, 
    2.430903e-05, 2.183874e-05, 1.983854e-05, 1.565074e-05, 1.3567e-05, 
    1.363481e-05, 1.500293e-05, 1.831669e-05, 3.569146e-05, 4.862679e-05, 
    5.662816e-05, 7.004857e-05, 6.649803e-05, 5.438888e-05, 4.46983e-05, 
    4.953741e-05, 3.813317e-05, 3.362947e-05, 3.490644e-05, 3.900802e-05, 
    3.75838e-05, 3.507712e-05, 2.648793e-05, 1.527348e-05,
  6.217645e-05, 6.676521e-05, 7.042397e-05, 7.014372e-05, 6.845426e-05, 
    6.993265e-05, 7.195863e-05, 6.665519e-05, 5.894127e-05, 4.872152e-05, 
    4.424337e-05, 4.532744e-05, 7.123894e-05, 0.0001073991, 0.0001631713, 
    0.0002810297, 0.0002821016, 0.0002570099, 0.0002342247, 0.000159807, 
    0.0001324531, 9.795801e-05, 8.84148e-05, 9.048112e-05, 9.789285e-05, 
    9.575279e-05, 9.810804e-05, 8.948157e-05, 7.738759e-05,
  0.0003874861, 0.0003544746, 0.0003245987, 0.0003611074, 0.000418408, 
    0.0004051533, 0.0005096535, 0.0005122, 0.0004382827, 0.0003886229, 
    0.0003302566, 0.000418621, 0.0005706433, 0.0007387822, 0.0009585271, 
    0.001155509, 0.0009405469, 0.0008464204, 0.0006609228, 0.0006367156, 
    0.0005170662, 0.0003796352, 0.0003090315, 0.0004172086, 0.0005256479, 
    0.0005295657, 0.0005084414, 0.0004772597, 0.0004119786,
  0.00220815, 0.002267671, 0.002782476, 0.003211862, 0.002790258, 
    0.002780349, 0.002733568, 0.002642947, 0.00252833, 0.002861251, 
    0.005916861, 0.008949547, 0.008243847, 0.008542441, 0.007396252, 
    0.005467146, 0.003721029, 0.003101959, 0.00272916, 0.002550633, 
    0.002039147, 0.00196759, 0.002549741, 0.003024823, 0.003811212, 
    0.003325668, 0.003052611, 0.002195719, 0.002131804,
  0.01477234, 0.02110229, 0.03051009, 0.02382245, 0.02947551, 0.05254068, 
    0.03068686, 0.02998789, 0.0546329, 0.1015257, 0.1302961, 0.1409537, 
    0.08977944, 0.04193787, 0.04158982, 0.03075907, 0.02077079, 0.01599269, 
    0.01393036, 0.009287789, 0.01199311, 0.01400131, 0.01915342, 0.02367249, 
    0.02433057, 0.01543672, 0.01254773, 0.01139886, 0.0119583,
  0.121314, 0.1770098, 0.1682612, 0.1977144, 0.1984849, 0.1634095, 0.1899083, 
    0.2749911, 0.4275504, 0.5765548, 0.5848227, 0.6509278, 0.4266742, 
    0.2973732, 0.2488638, 0.2149411, 0.1503729, 0.09725434, 0.05262775, 
    0.04162002, 0.0470254, 0.06292883, 0.1064055, 0.1394726, 0.1471806, 
    0.1413174, 0.09767798, 0.0598942, 0.07946666,
  0.3260903, 0.4215398, 0.3418452, 0.2578601, 0.243899, 0.2591084, 0.3219357, 
    0.4718196, 0.7183074, 0.8196427, 0.8903558, 0.8168785, 0.5960495, 
    0.5033721, 0.4016334, 0.3347943, 0.2905739, 0.2142758, 0.148114, 
    0.1203684, 0.1245415, 0.1883744, 0.2536057, 0.3984669, 0.472297, 
    0.3193674, 0.1900213, 0.1883404, 0.2387342,
  0.3222488, 0.345912, 0.2976267, 0.2458962, 0.2178338, 0.2384866, 0.2896935, 
    0.4014648, 0.5082588, 0.6678485, 0.626653, 0.4431909, 0.3431145, 
    0.3353717, 0.292775, 0.256635, 0.2233084, 0.1938208, 0.1589072, 
    0.1375979, 0.1654879, 0.2426108, 0.2894401, 0.2345383, 0.2163168, 
    0.1867461, 0.1771226, 0.2026465, 0.2353837,
  0.2701201, 0.3212734, 0.3743362, 0.4396182, 0.4265669, 0.4722129, 
    0.6212417, 0.5691191, 0.6720929, 0.6303249, 0.4733044, 0.3963095, 
    0.3559827, 0.3321672, 0.2735825, 0.2419196, 0.2064789, 0.2028503, 
    0.1831731, 0.1881274, 0.2014102, 0.2092718, 0.1716177, 0.139804, 
    0.1180175, 0.1021157, 0.1227645, 0.173571, 0.2382364,
  0.1937866, 0.2685547, 0.4027433, 0.5412939, 0.6815836, 0.7408749, 
    0.9800639, 0.918053, 0.6992592, 0.4755604, 0.3235988, 0.2829891, 
    0.240864, 0.1803958, 0.133057, 0.1095789, 0.09784525, 0.103508, 
    0.09368137, 0.1122347, 0.1286625, 0.09165227, 0.06646831, 0.05574027, 
    0.04851574, 0.04710087, 0.05310863, 0.08261327, 0.1450417,
  0.04831269, 0.1080308, 0.1566802, 0.2080197, 0.2122028, 0.2724968, 
    0.3830541, 0.4253675, 0.3513045, 0.1331801, 0.0919389, 0.07022505, 
    0.07368075, 0.05187338, 0.03083534, 0.02058462, 0.02177364, 0.02441585, 
    0.02767953, 0.04280759, 0.03999362, 0.03348469, 0.02199235, 0.01621201, 
    0.01372097, 0.01113143, 0.009676412, 0.01174074, 0.02615422,
  0.006077854, 0.009277286, 0.01439481, 0.01546822, 0.01462059, 0.01661167, 
    0.02418915, 0.03011855, 0.02712764, 0.01889674, 0.01303844, 0.009869716, 
    0.008030677, 0.006743796, 0.005703347, 0.003379527, 0.002427531, 
    0.002831416, 0.004108842, 0.005648913, 0.01081542, 0.008603291, 
    0.003993669, 0.002712632, 0.002370878, 0.002020251, 0.001971992, 
    0.0024787, 0.004487696,
  0.0007761811, 0.000820259, 0.001101986, 0.001105134, 0.001867692, 
    0.0007366454, 0.0005985544, 0.0009590388, 0.001541065, 0.002218737, 
    0.001983512, 0.002341806, 0.00161853, 0.00166225, 0.001080694, 
    0.0009932842, 0.0009554274, 0.0008152666, 0.0009041089, 0.001000188, 
    0.00114827, 0.0009805437, 0.000549344, 0.0003539261, 0.0004702717, 
    0.0006216479, 0.0005908455, 0.0005217953, 0.0006486828,
  0.0002231253, 0.0003352022, 0.0002809554, 0.0001976461, 0.0001749455, 
    0.0001947488, 0.000191995, 0.0001594264, 0.0001240362, 0.0002077378, 
    0.0002219236, 0.0002142512, 0.0003748079, 0.0003496521, 0.0002282856, 
    0.0001969096, 0.0002488384, 0.0002896595, 0.0002763809, 0.0002172849, 
    0.0001755991, 0.0001388126, 9.828565e-05, 0.0001063892, 0.0001204163, 
    0.0001482882, 0.0002302778, 0.0002214757, 0.0001853802,
  0.0001083043, 0.0001021379, 9.135695e-05, 7.339274e-05, 6.822259e-05, 
    5.85765e-05, 3.696285e-05, 3.649786e-05, 7.011426e-05, 9.18286e-05, 
    6.690211e-05, 6.553826e-05, 7.832828e-05, 6.973179e-05, 6.258869e-05, 
    5.976632e-05, 6.176009e-05, 7.103374e-05, 7.851738e-05, 7.924785e-05, 
    6.297453e-05, 6.103553e-05, 5.570574e-05, 6.198908e-05, 6.5057e-05, 
    6.157376e-05, 8.265243e-05, 0.0001175811, 0.0001269821,
  1.635153e-05, 1.631225e-05, 1.351051e-05, 1.264726e-05, 1.390967e-05, 
    1.568156e-05, 1.634693e-05, 1.604595e-05, 1.842041e-05, 1.992387e-05, 
    2.021192e-05, 2.131304e-05, 2.396156e-05, 2.663866e-05, 2.469077e-05, 
    2.808955e-05, 2.798109e-05, 2.798072e-05, 2.859461e-05, 2.676823e-05, 
    2.563894e-05, 2.588125e-05, 2.665907e-05, 2.553076e-05, 2.284092e-05, 
    2.244675e-05, 1.688392e-05, 1.546625e-05, 1.555852e-05,
  2.935227e-05, 2.935227e-05, 2.935227e-05, 2.935227e-05, 2.935227e-05, 
    2.935227e-05, 2.935227e-05, 3.334714e-05, 3.334714e-05, 3.334714e-05, 
    3.334714e-05, 3.334714e-05, 3.334714e-05, 3.334714e-05, 3.53019e-05, 
    3.53019e-05, 3.53019e-05, 3.53019e-05, 3.53019e-05, 3.53019e-05, 
    3.53019e-05, 3.179367e-05, 3.179367e-05, 3.179367e-05, 3.179367e-05, 
    3.179367e-05, 3.179367e-05, 3.179367e-05, 2.935227e-05,
  3.047991e-05, 2.411587e-05, 2.047352e-05, 2.339991e-05, 2.551687e-05, 
    2.672872e-05, 2.725869e-05, 3.122108e-05, 3.439101e-05, 3.398027e-05, 
    2.981207e-05, 3.225447e-05, 3.517936e-05, 4.586507e-05, 5.978618e-05, 
    6.303831e-05, 6.10985e-05, 5.80309e-05, 5.083224e-05, 4.529075e-05, 
    4.424357e-05, 4.7279e-05, 4.811815e-05, 4.705337e-05, 4.784316e-05, 
    4.078125e-05, 3.624224e-05, 3.567553e-05, 3.187944e-05,
  5.406208e-05, 4.444905e-05, 3.536118e-05, 4.067398e-05, 6.056978e-05, 
    8.01169e-05, 7.9195e-05, 6.6878e-05, 5.868575e-05, 5.088164e-05, 
    4.832811e-05, 4.725313e-05, 7.230965e-05, 0.0001490234, 0.0001727734, 
    0.000195732, 0.0002237097, 0.0002040199, 0.0001652233, 0.000129708, 
    0.0001342402, 0.0001215685, 0.0001166253, 0.000119636, 0.0001332663, 
    0.0001259151, 0.0001132526, 9.282662e-05, 6.179068e-05,
  0.0001848384, 0.0002145793, 0.0002132142, 0.0001919166, 0.0001837403, 
    0.0002028012, 0.0002242102, 0.0001974887, 0.0001618832, 0.0001330413, 
    0.0001295049, 0.0001298199, 0.0002481896, 0.0002753414, 0.0004689964, 
    0.0007502983, 0.0008128975, 0.0007410048, 0.0006791193, 0.000425958, 
    0.0003727461, 0.0003061611, 0.00027668, 0.0002423538, 0.0002568654, 
    0.0002489276, 0.0002695061, 0.0002515719, 0.0002381991,
  0.0009748826, 0.0008799213, 0.0009389571, 0.001106936, 0.001405389, 
    0.00136006, 0.001346195, 0.001521082, 0.001253271, 0.001050578, 
    0.00095615, 0.0009175416, 0.001306638, 0.002109928, 0.003032705, 
    0.003627947, 0.003420908, 0.002876621, 0.001996734, 0.001998314, 
    0.001689687, 0.001220646, 0.001126595, 0.001254472, 0.001284942, 
    0.001377078, 0.001258138, 0.001160446, 0.0009984417,
  0.006418148, 0.006583762, 0.007935216, 0.01094883, 0.01127657, 0.01039606, 
    0.008497961, 0.01062004, 0.009227043, 0.009382683, 0.01647542, 
    0.03007039, 0.03231633, 0.02812529, 0.02150681, 0.02110357, 0.01568026, 
    0.009994403, 0.008573784, 0.008220362, 0.006369435, 0.005423788, 
    0.006188662, 0.007825295, 0.00955802, 0.009026857, 0.009182122, 
    0.007261837, 0.006523652,
  0.04664625, 0.07812366, 0.1341806, 0.1502497, 0.1232589, 0.1620332, 
    0.1338082, 0.1089575, 0.1535336, 0.2989458, 0.3441401, 0.351092, 
    0.2261425, 0.1167757, 0.110188, 0.1126332, 0.07387798, 0.05993442, 
    0.04903524, 0.0275834, 0.02644951, 0.03642258, 0.04529636, 0.05586151, 
    0.05690354, 0.04173727, 0.04275412, 0.05454192, 0.03930861,
  0.4555076, 0.8712304, 1.017288, 0.8094289, 0.7509468, 0.5017159, 0.4343675, 
    0.6417668, 1.076709, 1.405842, 1.349956, 1.293417, 0.9290713, 0.6371328, 
    0.5684965, 0.50477, 0.38744, 0.2674194, 0.1590987, 0.1064232, 0.1005721, 
    0.128378, 0.2156807, 0.4824941, 0.9331773, 0.7671235, 0.4683741, 
    0.2415526, 0.2571344,
  1.036237, 1.696504, 1.278671, 0.7870897, 0.6400939, 0.653, 0.7162932, 
    1.113547, 1.719945, 2.007167, 2.046761, 1.860532, 1.069884, 0.8002956, 
    0.6687541, 0.5916716, 0.5240971, 0.4379974, 0.3170877, 0.2558515, 
    0.2331527, 0.3194841, 0.529961, 1.085259, 1.907877, 1.503564, 0.7322393, 
    0.5088012, 0.6698413,
  0.9046398, 1.256732, 1.021531, 0.6968352, 0.5943331, 0.6520702, 0.8443553, 
    1.134753, 1.666828, 1.963314, 1.58299, 1.086507, 0.626411, 0.5289338, 
    0.4675404, 0.3961743, 0.3727735, 0.3594162, 0.3216689, 0.2682104, 
    0.3299706, 0.4386631, 0.6801477, 0.716096, 0.6620712, 0.567152, 0.486546, 
    0.5614217, 0.6248659,
  0.8007393, 0.901966, 0.9271196, 0.9451062, 1.072286, 1.397636, 1.919398, 
    1.877093, 2.111483, 1.656696, 1.118699, 0.8138177, 0.6445256, 0.5594528, 
    0.4884135, 0.4527167, 0.3948968, 0.3873593, 0.4046301, 0.4195677, 
    0.5114963, 0.6505358, 0.5977207, 0.4821747, 0.4126762, 0.3334203, 
    0.3614953, 0.4871599, 0.6292731,
  0.4689272, 0.6661001, 0.8719653, 1.088675, 1.554346, 1.930576, 2.805089, 
    2.904836, 2.340496, 1.722188, 1.034127, 0.7636473, 0.6819696, 0.4949741, 
    0.3773965, 0.3020655, 0.2541015, 0.2691118, 0.2574847, 0.3331728, 
    0.4784313, 0.4146811, 0.2120228, 0.1676763, 0.1199537, 0.1119173, 
    0.145728, 0.2268116, 0.377267,
  0.09269791, 0.2604438, 0.3951948, 0.476306, 0.6563831, 0.7766813, 1.249866, 
    1.607244, 1.164699, 0.5631208, 0.3605298, 0.2814887, 0.272652, 0.1771292, 
    0.1129903, 0.07936489, 0.06966168, 0.07584458, 0.09432267, 0.1323042, 
    0.171746, 0.1254861, 0.07591234, 0.05912538, 0.04687207, 0.03179147, 
    0.02403786, 0.02256774, 0.06001075,
  0.01402991, 0.02603762, 0.04403608, 0.04405783, 0.04485161, 0.05236808, 
    0.080226, 0.1101779, 0.1006021, 0.07047875, 0.0491229, 0.04527427, 
    0.03400081, 0.02696835, 0.02293304, 0.01563989, 0.009869672, 0.0103542, 
    0.01594803, 0.02128975, 0.04131662, 0.03398672, 0.01472445, 0.01057518, 
    0.008280241, 0.007589854, 0.00677408, 0.005988553, 0.009092282,
  0.002007801, 0.002570332, 0.002949648, 0.00306251, 0.004611332, 
    0.001828623, 0.001828964, 0.002853838, 0.005077061, 0.008074441, 
    0.007254592, 0.01020782, 0.008217363, 0.009787684, 0.005558036, 
    0.003666007, 0.002848074, 0.002747883, 0.003053892, 0.003228725, 
    0.004012752, 0.003304123, 0.001775998, 0.001214818, 0.001330842, 
    0.001705936, 0.001801478, 0.001543509, 0.001653608,
  0.0004743918, 0.0009487085, 0.0009447235, 0.0007526722, 0.0006861138, 
    0.000645501, 0.0006440052, 0.000608496, 0.0005138862, 0.0006593751, 
    0.0009318946, 0.0008476169, 0.001327663, 0.001388891, 0.0009507688, 
    0.000702676, 0.0006880193, 0.0009082353, 0.0008044338, 0.0006603841, 
    0.0005699511, 0.0004721925, 0.0004205999, 0.0003884146, 0.00043575, 
    0.0004947036, 0.0006474954, 0.0006147663, 0.0004700288,
  0.0004648232, 0.0003591554, 0.0003257682, 0.0002396143, 0.0002100804, 
    0.0001881918, 0.0001236791, 0.0001462948, 0.0001629119, 0.0002904097, 
    0.0002054191, 0.0001828381, 0.0002230616, 0.0002845008, 0.0002564088, 
    0.0001728128, 0.000165535, 0.000223142, 0.0002933956, 0.0003522536, 
    0.0002742168, 0.0002602799, 0.0002290425, 0.0002278543, 0.000244105, 
    0.0001809917, 0.0002131664, 0.0003155439, 0.0004636266,
  5.427276e-05, 5.615482e-05, 5.155138e-05, 5.048201e-05, 5.120334e-05, 
    5.241163e-05, 4.988893e-05, 5.236441e-05, 8.069186e-05, 9.439173e-05, 
    9.677431e-05, 0.0001111769, 0.0001184305, 0.0001268358, 0.0001150742, 
    9.782699e-05, 9.806317e-05, 0.0001156989, 0.0001165539, 0.0001025236, 
    9.611568e-05, 9.653138e-05, 9.471318e-05, 0.0001014128, 0.000100757, 
    9.018627e-05, 7.908783e-05, 5.956752e-05, 5.386362e-05,
  0.0001150029, 0.0001150029, 0.0001150029, 0.0001150029, 0.0001150029, 
    0.0001150029, 0.0001150029, 0.000113149, 0.000113149, 0.000113149, 
    0.000113149, 0.000113149, 0.000113149, 0.000113149, 0.0001353594, 
    0.0001353594, 0.0001353594, 0.0001353594, 0.0001353594, 0.0001353594, 
    0.0001353594, 0.0001275914, 0.0001275914, 0.0001275914, 0.0001275914, 
    0.0001275914, 0.0001275914, 0.0001275914, 0.0001150029,
  0.0001219315, 8.384464e-05, 6.776017e-05, 7.259792e-05, 7.82757e-05, 
    8.33143e-05, 9.158899e-05, 9.61891e-05, 9.977754e-05, 9.664273e-05, 
    8.312333e-05, 8.44224e-05, 0.0001044413, 0.0001718162, 0.0002387789, 
    0.0001951671, 0.0001903077, 0.0001800757, 0.0001509312, 0.0001350045, 
    0.0001355158, 0.0001293227, 0.0001550057, 0.0001913333, 0.0001856738, 
    0.0001734642, 0.0001516213, 0.0001394416, 0.0001196334,
  0.0001665085, 0.0001531541, 0.0001195574, 0.0001307752, 0.0001616008, 
    0.0001962319, 0.0002232654, 0.0001864748, 0.0001536254, 0.0001459481, 
    0.0001312605, 0.0001178782, 0.0002505403, 0.0004073786, 0.0004916808, 
    0.00059793, 0.0006274773, 0.0005860259, 0.0004739988, 0.0003836472, 
    0.0003363072, 0.0003622061, 0.0003446964, 0.0003366039, 0.0003450996, 
    0.0003386227, 0.0003031741, 0.0002524118, 0.0001944624,
  0.0005754139, 0.0005673803, 0.0004564365, 0.0003794883, 0.0004408821, 
    0.0005047971, 0.0005545735, 0.0005598257, 0.0004167088, 0.0003195624, 
    0.0002989345, 0.0003719511, 0.0006394009, 0.000710686, 0.0009497795, 
    0.001661805, 0.002035279, 0.001865142, 0.001602775, 0.001170592, 
    0.0009659554, 0.0007892511, 0.0007830528, 0.0007732486, 0.0008054275, 
    0.0007486285, 0.0006794439, 0.0006920312, 0.0006440434,
  0.002532065, 0.00270646, 0.002847697, 0.003036924, 0.003651455, 
    0.003406806, 0.003069331, 0.003773004, 0.00315228, 0.002663254, 
    0.00243743, 0.002096478, 0.003307952, 0.005752977, 0.007901028, 
    0.009373361, 0.00890078, 0.007162376, 0.004661494, 0.005178688, 
    0.005454328, 0.004068214, 0.003801491, 0.003338796, 0.002853718, 
    0.003179696, 0.003006051, 0.002758889, 0.002579623,
  0.01905699, 0.01835746, 0.02014994, 0.03096063, 0.04287278, 0.04032161, 
    0.03182432, 0.03213884, 0.02575159, 0.03034987, 0.04166999, 0.07093152, 
    0.07592306, 0.06657612, 0.05315321, 0.05361023, 0.04031906, 0.02587311, 
    0.02519749, 0.02294764, 0.01754518, 0.01385519, 0.0136373, 0.0167367, 
    0.02068214, 0.02073647, 0.03116787, 0.0255454, 0.0226441,
  0.1418884, 0.2535851, 0.5066687, 0.6107607, 0.5127795, 0.352557, 0.2903349, 
    0.2659598, 0.3361427, 0.6090474, 0.6955134, 0.6035402, 0.4480371, 
    0.2480368, 0.215465, 0.234081, 0.1790749, 0.1483521, 0.1099801, 
    0.07524139, 0.05868022, 0.06609374, 0.08775257, 0.1007543, 0.129711, 
    0.09854319, 0.1752163, 0.2295502, 0.1484366,
  1.177276, 2.652151, 3.031745, 2.087207, 1.70086, 1.060266, 0.8343976, 
    1.120385, 1.756211, 2.384391, 2.242843, 1.884305, 1.465307, 1.032867, 
    0.9244298, 0.8339514, 0.6778408, 0.5091593, 0.3251129, 0.220867, 
    0.1966661, 0.2546344, 0.4078533, 1.368959, 2.906799, 2.351337, 1.282383, 
    0.6992236, 0.7381107,
  2.145927, 4.271271, 3.640004, 1.899289, 1.271254, 1.241527, 1.327047, 
    1.922836, 2.820471, 3.076268, 2.959101, 2.891632, 1.472164, 0.9966911, 
    0.8002306, 0.7309625, 0.6957909, 0.6221963, 0.4822226, 0.4051234, 
    0.3809438, 0.4671724, 0.8953834, 2.487567, 5.103821, 4.041335, 1.936956, 
    1.062786, 1.414388,
  1.980835, 3.511164, 2.789576, 1.425198, 1.252771, 1.315839, 1.653938, 
    2.234958, 3.464939, 4.090401, 2.48449, 1.708954, 0.8311047, 0.6143361, 
    0.5454822, 0.4755023, 0.4531328, 0.4485264, 0.4408815, 0.4111092, 
    0.5272612, 0.7210018, 1.293937, 1.940026, 1.800631, 1.623482, 1.350393, 
    1.311661, 1.4357,
  2.207705, 2.460757, 2.051984, 1.752708, 2.098118, 2.607553, 3.309859, 
    3.466844, 3.786687, 2.79731, 1.782972, 1.096718, 0.8529496, 0.670893, 
    0.6111083, 0.575659, 0.5380238, 0.542555, 0.6185738, 0.6835339, 
    0.9983572, 1.392662, 1.634057, 1.526163, 1.284225, 1.028927, 1.009387, 
    1.25613, 1.646746,
  1.070203, 1.33432, 1.494691, 1.759715, 2.523604, 3.389715, 4.496558, 
    4.431119, 4.32593, 3.220327, 2.008953, 1.292392, 1.089583, 0.8405684, 
    0.7183388, 0.5991089, 0.520301, 0.4596872, 0.4670761, 0.6340275, 
    1.088144, 0.986698, 0.5400342, 0.4484653, 0.305274, 0.2710098, 0.4286085, 
    0.706214, 0.9163578,
  0.1545267, 0.4554891, 0.6786671, 0.7947892, 1.167211, 1.447904, 2.324744, 
    2.84179, 2.062198, 1.334079, 0.9651392, 0.8364146, 0.7415418, 0.4889532, 
    0.3176191, 0.234552, 0.1762349, 0.1588047, 0.2145283, 0.2660937, 
    0.3086475, 0.3187583, 0.1987167, 0.1662644, 0.129846, 0.1146338, 
    0.0708166, 0.07160568, 0.09114972,
  0.02763772, 0.05551404, 0.08825795, 0.1008011, 0.1113399, 0.1201299, 
    0.1738537, 0.2556672, 0.2869275, 0.2044669, 0.1436618, 0.1564301, 
    0.1149479, 0.08426274, 0.07857973, 0.05839581, 0.0364445, 0.03561674, 
    0.04661055, 0.05403572, 0.09170254, 0.08737092, 0.04223328, 0.03217904, 
    0.02816475, 0.02802155, 0.0234027, 0.02124523, 0.01918881,
  0.005375721, 0.005510323, 0.007476003, 0.007193087, 0.009507135, 
    0.003387264, 0.004052122, 0.006224926, 0.01262643, 0.01955758, 
    0.01901948, 0.03442308, 0.02975851, 0.02548715, 0.02127149, 0.0127646, 
    0.01027613, 0.01130815, 0.009645113, 0.007678063, 0.0104576, 0.008560043, 
    0.006111179, 0.004502436, 0.004344718, 0.00479358, 0.005903027, 
    0.004967837, 0.005089973,
  0.001230654, 0.001437897, 0.002339808, 0.002235241, 0.001767431, 
    0.001234512, 0.001162248, 0.001266588, 0.001381749, 0.001311625, 
    0.002185629, 0.002034387, 0.003523752, 0.006519084, 0.003701159, 
    0.002188318, 0.001996799, 0.002454909, 0.002494008, 0.001934247, 
    0.001595247, 0.001414893, 0.001538312, 0.001275228, 0.001376764, 
    0.00169051, 0.00186477, 0.001751935, 0.001382693,
  0.0008587951, 0.0006977961, 0.0006908674, 0.0007476669, 0.0006969412, 
    0.0005626276, 0.000497193, 0.0005107956, 0.000489669, 0.0005287396, 
    0.0004770544, 0.000489955, 0.0006158678, 0.0008266997, 0.001127714, 
    0.0006613613, 0.0006667296, 0.0007170973, 0.0008243272, 0.001072987, 
    0.00103103, 0.001036491, 0.0008064064, 0.0007412686, 0.0006653566, 
    0.0005650251, 0.0005249251, 0.0008394592, 0.0009162041,
  0.0002124791, 0.0002082748, 0.000194651, 0.0001793109, 0.0001635365, 
    0.0001512928, 0.0001419957, 0.0001427794, 0.0002128393, 0.0002389187, 
    0.0002482597, 0.0002783116, 0.0003225864, 0.0003607353, 0.0003385181, 
    0.0003236332, 0.0003236396, 0.0004051807, 0.0004156118, 0.0003969272, 
    0.0003786236, 0.0003835284, 0.0003951322, 0.0004124613, 0.0003936607, 
    0.0003112199, 0.000278153, 0.0002541703, 0.0002174985,
  0.001580484, 0.001580484, 0.001580484, 0.001580484, 0.001580484, 
    0.001580484, 0.001580484, 0.001493644, 0.001493644, 0.001493644, 
    0.001493644, 0.001493644, 0.001493644, 0.001493644, 0.001840477, 
    0.001840477, 0.001840477, 0.001840477, 0.001840477, 0.001840477, 
    0.001840477, 0.001658431, 0.001658431, 0.001658431, 0.001658431, 
    0.001658431, 0.001658431, 0.001658431, 0.001580484,
  0.0005094475, 0.0003166444, 0.0002399866, 0.000232933, 0.0002351684, 
    0.0002453342, 0.0002642254, 0.000279362, 0.0002831479, 0.0002654165, 
    0.0002585209, 0.0002747364, 0.0004658028, 0.001207772, 0.000922161, 
    0.0005919959, 0.0005776747, 0.0004864129, 0.0004130391, 0.0004041005, 
    0.0004231986, 0.000429955, 0.0004824032, 0.0007978925, 0.0009300404, 
    0.0007476318, 0.0006548059, 0.0005292806, 0.0005203041,
  0.0006054715, 0.0004887122, 0.0004587613, 0.0004451837, 0.000428638, 
    0.0005072936, 0.0005525953, 0.000450355, 0.0003824894, 0.0003562069, 
    0.0003123943, 0.000299488, 0.0005719723, 0.000956103, 0.001173509, 
    0.001327511, 0.001288156, 0.001349939, 0.001256919, 0.001089154, 
    0.0009957647, 0.001040808, 0.001014544, 0.0009376235, 0.001072527, 
    0.001082905, 0.0008878937, 0.0008140437, 0.0006773545,
  0.001295175, 0.001186509, 0.0009185589, 0.0008178464, 0.001036572, 
    0.001214648, 0.001340871, 0.001373149, 0.001030726, 0.0007648026, 
    0.0007446239, 0.0007963044, 0.001579102, 0.00176904, 0.00207793, 
    0.003910816, 0.004801326, 0.004180556, 0.003771002, 0.002640771, 
    0.002240035, 0.002337083, 0.002253378, 0.002103422, 0.001960097, 
    0.001843648, 0.001827786, 0.001694385, 0.001415854,
  0.006961389, 0.006289882, 0.006636178, 0.007956707, 0.01144392, 0.01083854, 
    0.007573372, 0.009185911, 0.007385067, 0.00568483, 0.004293622, 
    0.00461515, 0.009712781, 0.01608883, 0.01983575, 0.01876065, 0.01866458, 
    0.01422826, 0.01048927, 0.01179639, 0.01189154, 0.01117277, 0.009908752, 
    0.007677461, 0.007603322, 0.007665419, 0.01121002, 0.009961697, 
    0.008411449,
  0.07535709, 0.05560476, 0.06350586, 0.1032577, 0.1265818, 0.1364115, 
    0.1072714, 0.0847914, 0.06952918, 0.08015566, 0.116415, 0.1346577, 
    0.1294144, 0.1214164, 0.1092899, 0.1072823, 0.0832921, 0.05489032, 
    0.06289847, 0.05790957, 0.04285448, 0.03305787, 0.02803599, 0.03165111, 
    0.04929824, 0.0606252, 0.09596177, 0.0953524, 0.078535,
  0.3944621, 0.6993607, 1.426851, 1.411543, 1.127284, 0.7326498, 0.563819, 
    0.5300629, 0.6199071, 0.9986335, 1.083316, 0.9284907, 0.7422689, 
    0.4580857, 0.3866082, 0.4099921, 0.3288087, 0.2775288, 0.2156224, 
    0.1622581, 0.1235491, 0.1160565, 0.1397562, 0.1749916, 0.3425147, 
    0.2781511, 0.5361204, 0.6452662, 0.4442227,
  2.150586, 4.973696, 5.810345, 3.626312, 2.691199, 1.759424, 1.318869, 
    1.544982, 2.28852, 3.067115, 3.02232, 2.43122, 1.971802, 1.406171, 
    1.245571, 1.11806, 0.9505062, 0.755119, 0.5179077, 0.3703791, 0.3314427, 
    0.4003606, 0.7199643, 2.952328, 5.695574, 4.538196, 2.671431, 1.542595, 
    1.411821,
  3.630293, 7.754515, 6.92725, 3.373362, 2.065215, 1.721906, 1.833915, 
    2.605708, 3.750361, 3.852066, 3.547425, 3.698649, 1.845379, 1.070945, 
    0.8545272, 0.7813402, 0.7881691, 0.7545725, 0.6050852, 0.5612222, 
    0.5431006, 0.6595535, 1.507852, 4.83143, 8.343967, 6.897871, 3.425492, 
    1.926538, 2.3394,
  3.556195, 6.790874, 5.699396, 2.350365, 2.011144, 1.947465, 2.285791, 
    3.15218, 4.998835, 6.384584, 2.922505, 2.008731, 0.9340983, 0.6380356, 
    0.5672219, 0.5167897, 0.4932446, 0.507417, 0.5264923, 0.5457768, 
    0.7263605, 1.172394, 2.200186, 4.22486, 3.938222, 3.374203, 2.923099, 
    2.566793, 2.635635,
  4.592996, 5.458025, 4.097816, 2.713217, 2.939263, 3.459235, 4.25457, 
    4.556525, 5.062462, 3.681779, 2.244201, 1.298302, 0.9328591, 0.7124712, 
    0.6609232, 0.6355134, 0.6204843, 0.6510146, 0.8212858, 0.9632015, 
    1.46293, 2.169981, 3.103409, 3.394793, 2.774088, 2.298118, 2.283682, 
    2.732953, 3.726723,
  1.973805, 2.22693, 2.40899, 2.566699, 3.375231, 4.477416, 5.640049, 
    5.759037, 5.738905, 4.411582, 2.801348, 1.781302, 1.388843, 1.144179, 
    1.042778, 0.9515355, 0.8226511, 0.6774509, 0.7164302, 0.9920224, 
    1.842137, 1.66472, 1.097936, 0.9216244, 0.7537667, 0.6593578, 1.01922, 
    1.792734, 1.876346,
  0.2630745, 0.684691, 0.9579034, 1.109262, 1.574347, 2.018528, 3.126827, 
    3.785121, 3.059104, 2.436967, 1.901743, 1.615308, 1.491327, 1.089826, 
    0.8296589, 0.5868082, 0.4155922, 0.3328947, 0.4008181, 0.4558316, 
    0.546069, 0.607638, 0.5307879, 0.5046313, 0.3996671, 0.3874219, 
    0.2144794, 0.1876213, 0.1938992,
  0.06067614, 0.09686025, 0.1452944, 0.1822353, 0.1993875, 0.21504, 
    0.2916742, 0.4763438, 0.5585863, 0.4356972, 0.3617471, 0.3847968, 
    0.3160199, 0.2249951, 0.2360832, 0.2080248, 0.1398498, 0.1039801, 
    0.1090673, 0.1146012, 0.1657911, 0.1802924, 0.1157401, 0.1037936, 
    0.1126847, 0.1080077, 0.1039451, 0.0854777, 0.05886786,
  0.01563546, 0.01223122, 0.01663202, 0.01461217, 0.01449284, 0.007044686, 
    0.006309222, 0.008364682, 0.02075057, 0.03366857, 0.03641582, 0.06508306, 
    0.06876563, 0.04914443, 0.05149369, 0.03422356, 0.03123657, 0.03627523, 
    0.0263409, 0.01808429, 0.02168995, 0.01922062, 0.01652811, 0.01235473, 
    0.01237745, 0.01532743, 0.01866636, 0.01522932, 0.01623837,
  0.003521952, 0.003158769, 0.004397222, 0.005208588, 0.003850227, 
    0.002716466, 0.002393847, 0.002200984, 0.001938004, 0.002071428, 
    0.003125905, 0.00338961, 0.009770365, 0.0207173, 0.009989598, 
    0.006314492, 0.005033693, 0.00561452, 0.006517424, 0.004905741, 
    0.00392035, 0.003938107, 0.00517847, 0.003872161, 0.004637908, 
    0.004651139, 0.005024297, 0.004406419, 0.003666075,
  0.001655085, 0.001346814, 0.001411114, 0.001722981, 0.001807779, 
    0.001408679, 0.001169646, 0.001057755, 0.001150102, 0.00091368, 
    0.001073651, 0.001185906, 0.001452094, 0.002641903, 0.00423435, 
    0.003218938, 0.002588127, 0.002925567, 0.002595128, 0.003259078, 
    0.003606794, 0.004043495, 0.003032903, 0.002763523, 0.002273812, 
    0.001559676, 0.001204234, 0.001986171, 0.001974489,
  0.0006877149, 0.0006874856, 0.0006466993, 0.0006179176, 0.0005806275, 
    0.0005284218, 0.0005221575, 0.0005363685, 0.0007755139, 0.0009282209, 
    0.001050148, 0.001103685, 0.000988615, 0.0009663245, 0.001030817, 
    0.001085114, 0.001147009, 0.001191355, 0.001289765, 0.001329818, 
    0.001307529, 0.001319311, 0.001413617, 0.001259618, 0.001156294, 
    0.0008222061, 0.0007148289, 0.000811205, 0.0007128643,
  0.006951712, 0.006951712, 0.006951712, 0.006951712, 0.006951712, 
    0.006951712, 0.006951712, 0.007636101, 0.007636101, 0.007636101, 
    0.007636101, 0.007636101, 0.007636101, 0.007636101, 0.01035031, 
    0.01035031, 0.01035031, 0.01035031, 0.01035031, 0.01035031, 0.01035031, 
    0.009275301, 0.009275301, 0.009275301, 0.009275301, 0.009275301, 
    0.009275301, 0.009275301, 0.006951712,
  0.001530386, 0.001031392, 0.000740075, 0.0007743145, 0.000667775, 
    0.0006535344, 0.0007233199, 0.000761823, 0.000729389, 0.0009396534, 
    0.00162787, 0.002665729, 0.003540572, 0.004279959, 0.003266488, 
    0.002488517, 0.002067192, 0.001526234, 0.001182669, 0.001299605, 
    0.001333298, 0.001459709, 0.00185952, 0.005240523, 0.006243953, 
    0.003983255, 0.002560997, 0.001903596, 0.001621531,
  0.002539031, 0.001914461, 0.001815103, 0.001733809, 0.001213313, 
    0.002057662, 0.002445892, 0.001017587, 0.0008879863, 0.0009217087, 
    0.0008383189, 0.0008045982, 0.001276709, 0.004172576, 0.007410894, 
    0.004793511, 0.0039892, 0.0043452, 0.003969897, 0.003487166, 0.003107211, 
    0.003103396, 0.002920989, 0.002971565, 0.00381688, 0.003578199, 
    0.002912198, 0.002699116, 0.003021501,
  0.002552466, 0.002174972, 0.001944421, 0.002158242, 0.002681151, 
    0.005537366, 0.005797823, 0.003970243, 0.002652339, 0.002201961, 
    0.001829988, 0.002982463, 0.007598225, 0.008276242, 0.00828844, 
    0.01270764, 0.0133588, 0.01136842, 0.01050217, 0.007105785, 0.005422061, 
    0.00724825, 0.007362254, 0.007193909, 0.006206431, 0.005392282, 
    0.008210535, 0.006201585, 0.003382562,
  0.02110928, 0.01881344, 0.01690788, 0.02480322, 0.04960823, 0.05232393, 
    0.03180238, 0.02940149, 0.02501366, 0.01447402, 0.009771085, 0.01212685, 
    0.02736207, 0.04182205, 0.05800786, 0.05106352, 0.03927739, 0.03208551, 
    0.03287132, 0.03046931, 0.03413464, 0.03241305, 0.02963417, 0.02276364, 
    0.02354573, 0.03356856, 0.06558359, 0.05059149, 0.03703017,
  0.2371364, 0.1831234, 0.1853961, 0.3246022, 0.3171057, 0.3759529, 
    0.3207823, 0.2233586, 0.1772228, 0.1780204, 0.2419719, 0.2496135, 
    0.231393, 0.2165736, 0.2281473, 0.2229831, 0.170752, 0.1218651, 
    0.1414367, 0.1356613, 0.1019615, 0.07645024, 0.06560864, 0.06021721, 
    0.1296164, 0.1808429, 0.3069121, 0.341568, 0.2671729,
  0.8531952, 1.40258, 2.725296, 2.475757, 1.876039, 1.277073, 0.9961599, 
    0.9300961, 0.9426039, 1.371761, 1.452451, 1.286746, 1.113205, 0.7467928, 
    0.6297265, 0.6612925, 0.5386244, 0.4789113, 0.3961928, 0.2908125, 
    0.2367287, 0.236556, 0.2651593, 0.428133, 0.8280236, 0.8743529, 1.193951, 
    1.329282, 0.9873758,
  3.23155, 7.326175, 8.099332, 4.953174, 3.622484, 2.396501, 1.733916, 
    1.919463, 2.66672, 3.459682, 3.60738, 2.89754, 2.37423, 1.746637, 
    1.455135, 1.305109, 1.136763, 0.960829, 0.7203938, 0.5587338, 0.4989164, 
    0.6253682, 1.292734, 5.013988, 7.830761, 6.567622, 4.279104, 2.734871, 
    2.218114,
  5.324015, 10.96564, 10.26986, 4.979702, 2.718161, 2.066092, 2.112337, 
    2.958978, 4.319996, 4.336878, 3.826365, 4.130176, 2.085821, 1.092664, 
    0.8475223, 0.7705789, 0.8179833, 0.8094718, 0.6975412, 0.6772824, 
    0.6683985, 0.8991938, 2.587984, 7.761147, 10.89518, 9.043403, 4.849286, 
    2.942418, 3.305575,
  5.679382, 10.59163, 9.25357, 3.378987, 2.706485, 2.400444, 2.664974, 
    3.439434, 6.090319, 8.156769, 3.069418, 2.14365, 0.9900059, 0.6411309, 
    0.5626385, 0.5315582, 0.5247582, 0.5642806, 0.6137373, 0.6875257, 
    0.9612522, 1.651265, 3.372937, 7.405557, 6.845757, 5.546163, 4.29983, 
    3.857741, 4.076531,
  7.232336, 9.087193, 6.960203, 3.717959, 3.742234, 3.902857, 4.713958, 
    5.113469, 5.795646, 4.236352, 2.533003, 1.445528, 0.9675586, 0.7351783, 
    0.6601478, 0.664639, 0.6625165, 0.7369902, 0.9287018, 1.198516, 1.783847, 
    2.687475, 4.377697, 5.555742, 4.511688, 3.699784, 4.048571, 4.939763, 
    6.635523,
  3.371907, 3.505473, 3.738691, 3.730545, 4.204821, 5.245625, 6.454237, 
    6.656936, 6.814035, 5.352244, 3.458818, 2.178901, 1.67685, 1.455926, 
    1.343213, 1.307253, 1.103516, 0.8955855, 0.9634458, 1.315263, 2.482009, 
    2.354138, 1.75424, 1.57909, 1.513795, 1.269844, 1.750568, 3.02697, 3.27692,
  0.5537164, 0.9738026, 1.26221, 1.412438, 1.850091, 2.413077, 3.582556, 
    4.442333, 3.949749, 3.59392, 3.077612, 2.608621, 2.516404, 2.068125, 
    1.779993, 1.287437, 0.9909655, 0.7562012, 0.7247404, 0.7620569, 
    0.9499828, 1.140528, 1.239736, 1.320704, 1.12036, 1.010108, 0.587431, 
    0.4715466, 0.4728314,
  0.1795035, 0.1894846, 0.2253042, 0.2555197, 0.2955032, 0.3335621, 
    0.4168984, 0.7368968, 0.8414015, 0.6591178, 0.7502964, 0.7842473, 
    0.7805684, 0.6342809, 0.7009932, 0.6767127, 0.5461736, 0.2889315, 
    0.2645402, 0.2500238, 0.2969857, 0.3658043, 0.4384147, 0.4636684, 
    0.5927147, 0.5511773, 0.4494694, 0.3404827, 0.2268965,
  0.0605882, 0.03773217, 0.03830818, 0.03608865, 0.0250191, 0.0195291, 
    0.01344806, 0.01268281, 0.03005841, 0.06492101, 0.09839439, 0.1478704, 
    0.1395275, 0.1005924, 0.1146165, 0.1111365, 0.1235818, 0.09186696, 
    0.07022019, 0.04290187, 0.05339237, 0.04892998, 0.04916945, 0.03110737, 
    0.04310425, 0.0608206, 0.08086527, 0.0697535, 0.06719052,
  0.01337002, 0.01086179, 0.01159219, 0.01346997, 0.01131754, 0.008139445, 
    0.006834511, 0.005354655, 0.00449373, 0.003885701, 0.00524183, 
    0.006891586, 0.02188932, 0.04040675, 0.02161255, 0.01373581, 0.0127255, 
    0.01551913, 0.01389591, 0.01167279, 0.0105549, 0.01185565, 0.0149102, 
    0.01132028, 0.01199381, 0.01330256, 0.01772988, 0.01714473, 0.01608658,
  0.004608718, 0.004963528, 0.00450792, 0.004839703, 0.005003836, 0.00434257, 
    0.003270304, 0.002381538, 0.002440563, 0.002274888, 0.002389997, 
    0.002587142, 0.00353222, 0.00654855, 0.01154401, 0.01236207, 0.007839254, 
    0.008656752, 0.008077242, 0.009350578, 0.009896703, 0.01148634, 
    0.01009756, 0.008202768, 0.006825745, 0.003862006, 0.002960089, 
    0.00600607, 0.005438817,
  0.002131521, 0.002157472, 0.001865509, 0.001752339, 0.001543059, 
    0.001479139, 0.001520037, 0.001611106, 0.002232866, 0.002463132, 
    0.00284106, 0.002860113, 0.002698356, 0.002607078, 0.002727808, 
    0.003070136, 0.003222935, 0.003275344, 0.003512267, 0.003799892, 
    0.003640714, 0.003524503, 0.003281673, 0.002821096, 0.00253357, 
    0.001901922, 0.001797295, 0.002180933, 0.002274455,
  0.01511111, 0.01511111, 0.01511111, 0.01511111, 0.01511111, 0.01511111, 
    0.01511111, 0.01532842, 0.01532842, 0.01532842, 0.01532842, 0.01532842, 
    0.01532842, 0.01532842, 0.01724832, 0.01724832, 0.01724832, 0.01724832, 
    0.01724832, 0.01724832, 0.01724832, 0.01702866, 0.01702866, 0.01702866, 
    0.01702866, 0.01702866, 0.01702866, 0.01702866, 0.01511111,
  0.005332128, 0.003749793, 0.002545513, 0.002938672, 0.00261324, 
    0.002235064, 0.002148724, 0.002166856, 0.002301289, 0.006398683, 
    0.009015989, 0.01178379, 0.01167777, 0.01527302, 0.01431668, 0.009887318, 
    0.007921777, 0.006023682, 0.004519053, 0.005368875, 0.006221745, 
    0.006785155, 0.01094038, 0.02583887, 0.0255541, 0.01728187, 0.01212632, 
    0.007325314, 0.005387528,
  0.008719712, 0.009821682, 0.01068908, 0.007641638, 0.004515855, 0.01208546, 
    0.01447073, 0.003161901, 0.002492201, 0.002936727, 0.002628392, 
    0.002740293, 0.00572158, 0.0264503, 0.03743208, 0.03354632, 0.01859061, 
    0.01604202, 0.01288449, 0.01100855, 0.01128451, 0.01086023, 0.0112468, 
    0.0124742, 0.01645541, 0.01469853, 0.01299971, 0.009921526, 0.008981682,
  0.008537212, 0.00650635, 0.006313365, 0.007414198, 0.01571261, 0.05233074, 
    0.04727796, 0.02348154, 0.01039855, 0.009853831, 0.006856558, 0.0161502, 
    0.02760033, 0.03185696, 0.03254415, 0.05928922, 0.06931079, 0.05720442, 
    0.04464773, 0.0309605, 0.02219535, 0.02159614, 0.02330087, 0.02366593, 
    0.02198995, 0.02410638, 0.03642888, 0.03289399, 0.01828178,
  0.1036178, 0.07059926, 0.06318419, 0.08857111, 0.1602776, 0.16979, 
    0.1442328, 0.1339012, 0.1019012, 0.05475314, 0.03858202, 0.05243208, 
    0.09798074, 0.1321438, 0.1675998, 0.1660781, 0.1180607, 0.1027401, 
    0.1210356, 0.1039265, 0.09716034, 0.08821299, 0.08550934, 0.06958503, 
    0.07743493, 0.1836627, 0.2838956, 0.2519748, 0.1703553,
  0.6277775, 0.4917445, 0.5154516, 0.7128973, 0.7447922, 0.874487, 0.7529864, 
    0.5429895, 0.4395549, 0.3751937, 0.4170209, 0.4469697, 0.4751739, 
    0.4546996, 0.4706634, 0.465358, 0.3773624, 0.2917335, 0.3061161, 
    0.3069096, 0.2413042, 0.1918984, 0.1651334, 0.131769, 0.2736953, 
    0.5832796, 0.8707004, 0.9174927, 0.8036583,
  1.592656, 2.182764, 3.929897, 3.64083, 2.80754, 1.981381, 1.589153, 
    1.458947, 1.346988, 1.731598, 1.852311, 1.6607, 1.52137, 1.145583, 
    0.9454076, 0.9723351, 0.8115549, 0.7077252, 0.6127631, 0.476232, 
    0.411156, 0.4581954, 0.5215827, 0.9326669, 1.592372, 1.886303, 2.301134, 
    2.247076, 1.888644,
  4.328771, 9.10191, 9.913984, 6.256444, 4.584117, 2.887891, 2.119515, 
    2.186603, 2.921224, 3.644874, 4.075247, 3.252454, 2.708067, 2.05036, 
    1.603024, 1.399006, 1.210954, 1.082679, 0.8692253, 0.7415267, 0.6561793, 
    0.9160462, 2.180344, 6.598634, 8.995624, 8.215826, 5.735483, 3.878997, 
    3.304462,
  6.791904, 13.90766, 13.4828, 6.639337, 3.349489, 2.275988, 2.157084, 
    2.976036, 4.602953, 4.585913, 3.992972, 4.339365, 2.223799, 1.062055, 
    0.8115653, 0.7443889, 0.8099909, 0.8261886, 0.7685893, 0.7592465, 
    0.773482, 1.162905, 3.797468, 10.78402, 12.58004, 10.42242, 6.033156, 
    3.879925, 4.284447,
  7.728687, 14.66736, 12.89356, 4.382424, 3.298981, 2.540939, 2.784657, 
    3.413242, 6.666172, 9.132317, 3.137887, 2.205638, 0.9995427, 0.6389977, 
    0.542868, 0.5254204, 0.5260392, 0.6054584, 0.667917, 0.8086473, 1.150521, 
    2.051379, 4.74472, 10.63109, 9.955057, 7.656169, 5.329571, 4.843908, 
    5.514168,
  9.893394, 12.06967, 10.07566, 4.732163, 4.500092, 4.040002, 4.762089, 
    5.178194, 6.089296, 4.576267, 2.696867, 1.532762, 0.9862981, 0.7496182, 
    0.6525042, 0.6793457, 0.7005761, 0.7893482, 0.9954547, 1.339441, 
    1.973162, 2.926935, 5.291141, 7.618023, 5.983488, 5.141035, 5.59586, 
    6.991391, 9.155485,
  4.722902, 5.168579, 5.396625, 5.114639, 5.302925, 5.936427, 7.049647, 
    7.189176, 7.586354, 5.895446, 4.048012, 2.506141, 1.947498, 1.760124, 
    1.642784, 1.612244, 1.336815, 1.105912, 1.171275, 1.598471, 2.865263, 
    2.986379, 2.343704, 2.163507, 2.265174, 2.081805, 2.587168, 4.060379, 
    4.842722,
  1.097959, 1.373605, 1.569541, 1.766557, 2.147713, 2.759139, 3.981376, 
    4.93033, 4.764506, 4.957766, 4.473251, 3.914511, 3.57866, 3.14167, 
    2.708625, 2.076839, 1.866637, 1.445539, 1.262802, 1.207472, 1.502797, 
    1.974808, 2.191031, 2.388562, 2.106984, 1.960495, 1.317439, 1.015823, 
    0.9657719,
  0.5431685, 0.507104, 0.4349629, 0.3568382, 0.5337634, 0.508694, 0.5477465, 
    1.033354, 1.096844, 0.9535319, 1.284278, 1.364323, 1.472617, 1.457678, 
    1.593458, 1.38738, 1.342641, 0.891848, 0.7299761, 0.5945635, 0.5353203, 
    0.8353323, 1.29098, 1.391222, 1.663778, 1.589531, 1.150371, 0.9160087, 
    0.6809665,
  0.2949945, 0.1681855, 0.184229, 0.1557972, 0.1452218, 0.1308788, 
    0.08261947, 0.04117641, 0.07828725, 0.2124044, 0.4313813, 0.4871961, 
    0.3915293, 0.3174828, 0.3714372, 0.4120969, 0.4476052, 0.3136238, 
    0.250396, 0.1497739, 0.1639251, 0.2000411, 0.2160901, 0.1364142, 
    0.185017, 0.2959647, 0.4168842, 0.3709425, 0.3269577,
  0.07401027, 0.04081625, 0.04241714, 0.05173058, 0.05331051, 0.04715138, 
    0.04087564, 0.03480924, 0.02597727, 0.0189082, 0.04481453, 0.04786512, 
    0.06785966, 0.08534419, 0.05890085, 0.05420921, 0.06571453, 0.06973681, 
    0.0412532, 0.05512821, 0.04064011, 0.04731156, 0.03892661, 0.03038224, 
    0.04103636, 0.07246731, 0.1069301, 0.09306551, 0.08609842,
  0.02216307, 0.02313466, 0.01976598, 0.02100315, 0.01996052, 0.01721523, 
    0.01320974, 0.01020971, 0.008856913, 0.02168541, 0.01277862, 0.01052848, 
    0.01358885, 0.02132009, 0.03415563, 0.03808559, 0.02814955, 0.02237181, 
    0.02354093, 0.02576366, 0.02484129, 0.02703611, 0.0238114, 0.02144214, 
    0.02377668, 0.010956, 0.008161938, 0.02862352, 0.02458872,
  0.007838026, 0.00796607, 0.007405359, 0.00730161, 0.006248452, 0.005771136, 
    0.005425583, 0.006962125, 0.01163417, 0.01694024, 0.01851421, 0.0173109, 
    0.01661338, 0.01355972, 0.01108314, 0.009571579, 0.009295111, 0.00824871, 
    0.008760868, 0.009532074, 0.01002717, 0.009395463, 0.008133234, 
    0.007051887, 0.006041236, 0.004392935, 0.004649817, 0.006522326, 
    0.007858324,
  0.02353415, 0.02353415, 0.02353415, 0.02353415, 0.02353415, 0.02353415, 
    0.02353415, 0.02269775, 0.02269775, 0.02269775, 0.02269775, 0.02269775, 
    0.02269775, 0.02269775, 0.0237714, 0.0237714, 0.0237714, 0.0237714, 
    0.0237714, 0.0237714, 0.0237714, 0.02511728, 0.02511728, 0.02511728, 
    0.02511728, 0.02511728, 0.02511728, 0.02511728, 0.02353415,
  0.01732665, 0.01451974, 0.01092764, 0.01141971, 0.01181054, 0.00911276, 
    0.007056473, 0.007091687, 0.009478845, 0.02025359, 0.02268932, 
    0.02666511, 0.02767241, 0.04419655, 0.05206429, 0.04176861, 0.03092688, 
    0.02296774, 0.0189069, 0.02212146, 0.02525388, 0.02647608, 0.04125503, 
    0.07634577, 0.07429758, 0.05712794, 0.04717719, 0.02875038, 0.01777375,
  0.03086604, 0.03627167, 0.0439208, 0.03887248, 0.02139945, 0.04966191, 
    0.060543, 0.01158498, 0.008035151, 0.0100975, 0.009856207, 0.01108332, 
    0.03624746, 0.09364606, 0.118249, 0.1180785, 0.07802685, 0.06653651, 
    0.05022051, 0.04020758, 0.04059121, 0.0384105, 0.04144266, 0.04873322, 
    0.06202899, 0.05743853, 0.05204935, 0.036892, 0.02800821,
  0.04385491, 0.0242077, 0.0244079, 0.0278333, 0.09145793, 0.2239785, 
    0.1887943, 0.1021499, 0.05255225, 0.04125241, 0.03109243, 0.05408435, 
    0.07076947, 0.1061487, 0.1274169, 0.2384775, 0.2776386, 0.223709, 
    0.1673012, 0.1194129, 0.08050494, 0.07193178, 0.06933281, 0.06853474, 
    0.07520705, 0.08830132, 0.1175309, 0.1262743, 0.08156952,
  0.3464734, 0.2243935, 0.1918407, 0.3035091, 0.4342381, 0.4981282, 
    0.5028173, 0.4316328, 0.2947577, 0.1756258, 0.165499, 0.209155, 
    0.2686572, 0.3473314, 0.4355422, 0.4449213, 0.3579618, 0.3087586, 
    0.3265221, 0.2883023, 0.2429672, 0.2119224, 0.2055686, 0.1767337, 
    0.2540092, 0.5075297, 0.7873107, 0.730244, 0.5276727,
  1.357823, 1.072331, 1.133348, 1.304299, 1.471144, 1.637677, 1.42277, 
    1.089821, 0.9239173, 0.7548452, 0.7568793, 0.8760127, 0.9365661, 
    1.002264, 0.8586157, 0.87931, 0.7304225, 0.6242987, 0.5757294, 0.5652615, 
    0.4559702, 0.4079597, 0.3672821, 0.2691979, 0.5847154, 1.449871, 
    1.831565, 1.836206, 1.653175,
  2.49289, 2.948062, 4.825466, 4.708982, 3.927885, 2.844235, 2.382258, 
    2.076773, 1.844008, 2.085083, 2.274374, 2.110822, 1.960709, 1.696643, 
    1.392047, 1.298038, 1.066514, 0.917613, 0.8174531, 0.6748152, 0.6288309, 
    0.6922973, 0.823892, 1.4953, 2.460922, 2.893613, 3.536166, 3.279494, 
    2.911586,
  5.382041, 10.27356, 11.26737, 7.65631, 5.593888, 3.31673, 2.424376, 
    2.344084, 3.023547, 3.711735, 4.4416, 3.543851, 2.926231, 2.266169, 
    1.737862, 1.45945, 1.235734, 1.126632, 0.9316456, 0.8470345, 0.7613146, 
    1.16213, 2.92222, 7.795585, 9.940176, 9.374944, 6.981789, 4.995313, 
    4.357917,
  8.073236, 16.3179, 15.86753, 8.183512, 3.922119, 2.391325, 2.108436, 
    2.814749, 4.667784, 4.696301, 4.042511, 4.371235, 2.317522, 1.034923, 
    0.7767179, 0.6977077, 0.7859499, 0.8230098, 0.7896282, 0.8097321, 
    0.8511522, 1.378672, 4.959991, 13.33864, 14.03979, 11.45049, 6.846908, 
    4.719218, 5.343144,
  9.275721, 17.63164, 15.75067, 5.553607, 3.798602, 2.54494, 2.731149, 
    3.262219, 7.056797, 9.726856, 3.1983, 2.188617, 0.9722338, 0.6148274, 
    0.5229236, 0.5139025, 0.5214535, 0.6151793, 0.7191636, 0.8827033, 
    1.265162, 2.331841, 6.073141, 13.62188, 12.47156, 9.151601, 6.107343, 
    5.733632, 6.598494,
  11.95797, 14.07066, 12.31996, 5.638963, 4.95838, 4.158165, 4.718024, 
    5.024546, 6.106493, 4.778955, 2.782161, 1.564873, 1.003134, 0.7630253, 
    0.6624467, 0.6839465, 0.7192651, 0.8170183, 1.04773, 1.427479, 2.081678, 
    3.086492, 6.075787, 9.236147, 7.252852, 6.282995, 6.727562, 8.22445, 
    11.21778,
  5.917679, 6.604487, 6.847071, 6.22732, 6.335303, 6.500968, 7.451329, 
    7.582521, 8.176217, 6.118811, 4.404107, 2.814383, 2.172489, 2.045825, 
    1.922672, 1.854195, 1.526494, 1.313978, 1.347567, 1.744885, 3.087026, 
    3.482632, 2.869658, 2.792555, 2.972546, 2.817377, 3.269418, 4.67794, 
    5.819546,
  1.609989, 1.859082, 1.917618, 2.257214, 2.625863, 3.186395, 4.396323, 
    5.320103, 5.533826, 6.568771, 5.872885, 5.198679, 4.463385, 3.988151, 
    3.429787, 2.715944, 2.678827, 2.161972, 1.805571, 1.683338, 2.156854, 
    2.771981, 3.103975, 3.303118, 2.909374, 2.85497, 2.169696, 1.74626, 
    1.588758,
  1.207652, 1.109382, 0.9553972, 0.5911633, 1.136937, 0.9219319, 0.7398592, 
    1.594353, 1.735268, 1.909252, 2.335205, 2.268797, 2.473677, 2.570107, 
    2.520659, 2.165592, 2.253219, 1.958469, 1.588018, 1.185207, 0.9567534, 
    1.682182, 2.315158, 2.574555, 2.857894, 2.702002, 2.061957, 1.737384, 
    1.368861,
  0.8877245, 0.5885301, 0.829977, 0.7074152, 0.869801, 0.6568743, 0.4950542, 
    0.205629, 0.4095557, 0.7689078, 1.104524, 1.161177, 1.026803, 0.9090542, 
    1.016558, 1.071, 1.13841, 0.8734968, 0.7498857, 0.4815964, 0.5301259, 
    0.7599933, 0.7280856, 0.523899, 0.6467641, 0.9341257, 1.132827, 1.039921, 
    0.9675555,
  0.2846027, 0.1664294, 0.2137938, 0.274426, 0.4094867, 0.3246445, 0.3006563, 
    0.2830704, 0.2617615, 0.2597193, 0.4341015, 0.3423256, 0.2634684, 
    0.3129709, 0.2667873, 0.3187004, 0.3056303, 0.259735, 0.1929989, 
    0.2526238, 0.2011062, 0.2168678, 0.1726306, 0.1687563, 0.2309225, 
    0.3434718, 0.4252971, 0.3694174, 0.3239535,
  0.103009, 0.101548, 0.08231499, 0.1049403, 0.1097331, 0.1315244, 0.1082484, 
    0.07945175, 0.06031414, 0.132409, 0.09998416, 0.08479741, 0.09563052, 
    0.125535, 0.1478921, 0.198015, 0.1467859, 0.102829, 0.1031347, 0.1166163, 
    0.09191502, 0.07968823, 0.07198068, 0.08229491, 0.1466346, 0.03998694, 
    0.02909199, 0.1347142, 0.1095761,
  0.03146236, 0.03225944, 0.03141638, 0.03085317, 0.03015892, 0.02807507, 
    0.0309916, 0.04569735, 0.07028128, 0.08788168, 0.09228004, 0.09687269, 
    0.09187279, 0.08031096, 0.0637767, 0.05126228, 0.0407432, 0.03287085, 
    0.0305048, 0.02949098, 0.02880926, 0.02774078, 0.02290078, 0.02396039, 
    0.02114848, 0.01316691, 0.01362019, 0.02334497, 0.03161585,
  0.04405832, 0.04405832, 0.04405832, 0.04405832, 0.04405832, 0.04405832, 
    0.04405832, 0.04054525, 0.04054525, 0.04054525, 0.04054525, 0.04054525, 
    0.04054525, 0.04054525, 0.0421253, 0.0421253, 0.0421253, 0.0421253, 
    0.0421253, 0.0421253, 0.0421253, 0.04619896, 0.04619896, 0.04619896, 
    0.04619896, 0.04619896, 0.04619896, 0.04619896, 0.04405832,
  0.04354375, 0.04125238, 0.03371315, 0.03129054, 0.03302769, 0.02843528, 
    0.02274302, 0.02432151, 0.03334702, 0.04319768, 0.04439432, 0.05031502, 
    0.05598873, 0.1088015, 0.1332852, 0.1219441, 0.09759084, 0.07311891, 
    0.06291329, 0.06230459, 0.06892236, 0.07151324, 0.09981437, 0.1713689, 
    0.1715105, 0.1404876, 0.1299333, 0.08583588, 0.04716579,
  0.08906865, 0.09643564, 0.1223603, 0.1273369, 0.07584698, 0.1260467, 
    0.1711024, 0.03944312, 0.02837037, 0.03598017, 0.03207678, 0.03715119, 
    0.14382, 0.2630139, 0.2940575, 0.2718403, 0.2258462, 0.2112851, 
    0.1551027, 0.1231678, 0.1159514, 0.1095004, 0.11243, 0.1311308, 0.171018, 
    0.1710875, 0.1533624, 0.1206662, 0.09279136,
  0.1371151, 0.08742693, 0.08047059, 0.09560757, 0.3053607, 0.4991068, 
    0.4287576, 0.2797031, 0.1643686, 0.1107, 0.1012867, 0.1417125, 0.2177124, 
    0.2888936, 0.3794164, 0.609482, 0.6572626, 0.5583572, 0.4313727, 
    0.3196446, 0.2161155, 0.1827245, 0.1696934, 0.1665646, 0.1901999, 
    0.2482662, 0.2813094, 0.2974462, 0.2064343,
  0.7769977, 0.5156301, 0.4241433, 0.6999621, 0.9232925, 1.062439, 1.065139, 
    0.901554, 0.5964005, 0.3994897, 0.3928484, 0.4807948, 0.5728465, 
    0.7709185, 0.9218338, 0.8957195, 0.8486324, 0.7291287, 0.6455215, 
    0.5871676, 0.4833588, 0.4196111, 0.3963672, 0.3528573, 0.5359851, 
    0.9445261, 1.433889, 1.397432, 1.062778,
  2.222106, 1.810468, 1.890722, 2.027647, 2.383504, 2.523572, 2.192064, 
    1.75064, 1.552252, 1.295742, 1.28257, 1.526071, 1.631054, 1.705752, 
    1.384468, 1.379801, 1.178272, 1.043079, 0.9136682, 0.8354012, 0.7060967, 
    0.6803238, 0.6114859, 0.4475697, 1.122218, 2.471177, 2.81274, 2.811507, 
    2.592448,
  3.278234, 3.610768, 5.545362, 5.539493, 4.917222, 3.727191, 3.16547, 
    2.677311, 2.287205, 2.354483, 2.584666, 2.567172, 2.449052, 2.27028, 
    1.915615, 1.624068, 1.324127, 1.130123, 0.9775351, 0.8421964, 0.778285, 
    0.8717252, 0.9781035, 1.761487, 2.967824, 3.864663, 4.670659, 4.317426, 
    3.782533,
  6.171607, 10.91545, 12.1925, 8.608304, 6.447398, 3.88148, 2.670992, 
    2.363581, 2.986024, 3.674123, 4.675293, 3.742503, 3.119538, 2.442461, 
    1.882425, 1.522181, 1.245315, 1.126841, 0.9569975, 0.8616595, 0.8033313, 
    1.344553, 3.165342, 8.124192, 10.61954, 10.22292, 7.786186, 5.794362, 
    5.155262,
  8.93085, 17.76401, 17.5106, 9.392919, 4.430055, 2.474141, 2.078725, 
    2.639961, 4.534021, 4.697206, 4.03776, 4.303308, 2.377828, 1.02412, 
    0.7494127, 0.6565402, 0.7489455, 0.8076556, 0.7570271, 0.7992892, 
    0.8855243, 1.470309, 5.750131, 15.02132, 15.21846, 12.13938, 7.371402, 
    5.389951, 6.193922,
  10.3419, 19.16615, 17.89554, 6.662904, 4.293016, 2.560222, 2.643575, 
    3.063097, 7.241293, 10.11052, 3.254551, 2.130368, 0.9302088, 0.5871961, 
    0.5023369, 0.50088, 0.5211457, 0.6111079, 0.7681209, 0.9273576, 1.291909, 
    2.515827, 7.045166, 15.85042, 14.1832, 9.857533, 6.577755, 6.495783, 
    7.472366,
  13.21543, 15.18117, 13.65226, 6.543843, 5.286088, 4.227055, 4.673527, 
    4.789721, 6.048709, 4.851265, 2.856988, 1.577836, 1.014968, 0.7656331, 
    0.6771786, 0.6851314, 0.7263031, 0.8229092, 1.074892, 1.468902, 2.12192, 
    3.152216, 6.786563, 10.37175, 8.23901, 7.03859, 7.372891, 8.812462, 
    12.4539,
  6.679238, 7.426672, 7.647952, 6.76588, 6.895083, 6.945659, 7.725692, 
    7.813612, 8.58879, 6.214727, 4.635169, 3.027474, 2.327358, 2.283427, 
    2.187071, 2.047568, 1.703882, 1.503039, 1.494019, 1.831733, 3.159446, 
    3.927698, 3.325815, 3.493592, 3.604414, 3.36302, 3.611125, 4.909204, 
    6.19916,
  2.032926, 2.305776, 2.317295, 2.926093, 3.20625, 3.660646, 4.84265, 
    5.660988, 6.27764, 8.35466, 7.275843, 6.226427, 5.278645, 4.734296, 
    3.95655, 3.261398, 3.27357, 2.702201, 2.210197, 2.08471, 2.778485, 
    3.380878, 4.024663, 3.995594, 3.365432, 3.434513, 2.866241, 2.432961, 
    2.224321,
  2.052665, 1.890823, 1.800772, 1.152723, 2.234412, 1.708895, 1.185657, 
    2.951475, 3.119673, 3.526094, 3.793704, 3.510403, 3.719295, 3.736811, 
    3.369959, 3.008449, 3.023537, 2.892155, 2.487192, 1.895316, 1.555815, 
    2.67172, 3.433439, 3.744849, 3.884118, 3.723169, 3.013107, 2.525849, 
    2.088498,
  1.703862, 1.482619, 1.964736, 2.023182, 2.426438, 2.057677, 1.51926, 
    0.913854, 1.440187, 1.912711, 2.207915, 2.134978, 2.122267, 1.92648, 
    1.993473, 2.056013, 1.987964, 1.577511, 1.504524, 1.032845, 1.292171, 
    1.687367, 1.656524, 1.186235, 1.446595, 1.762724, 1.95386, 1.983808, 
    1.817585,
  0.7746012, 0.587563, 0.8737028, 1.224193, 1.642957, 1.261504, 1.275329, 
    1.222695, 1.20638, 1.268003, 1.634604, 1.110498, 0.7737719, 0.9452256, 
    0.9508983, 0.9293041, 0.8136943, 0.7227362, 0.62331, 0.7153679, 
    0.6860409, 0.664832, 0.6916028, 0.6452168, 0.814597, 0.9399637, 1.024866, 
    0.9357134, 0.8377474,
  0.3710128, 0.3629012, 0.3381096, 0.5007275, 0.5429282, 0.587647, 0.5245665, 
    0.4123293, 0.32147, 0.4417665, 0.414926, 0.4071014, 0.4407092, 0.5125028, 
    0.5895595, 0.7003198, 0.5730571, 0.4230781, 0.426061, 0.4409941, 
    0.3316864, 0.2762543, 0.2875388, 0.3235202, 0.6024521, 0.1796778, 
    0.1019948, 0.4472797, 0.3871508,
  0.1200015, 0.1217746, 0.1227149, 0.1274106, 0.1304948, 0.129671, 0.1470409, 
    0.1700297, 0.2122687, 0.249078, 0.2636687, 0.261593, 0.2703258, 
    0.2752587, 0.2375327, 0.2011584, 0.1798808, 0.1639959, 0.1439373, 
    0.1231496, 0.1165135, 0.1137229, 0.09753983, 0.1141647, 0.1055171, 
    0.04751956, 0.0488555, 0.09495354, 0.1225981,
  0.08071082, 0.08071082, 0.08071082, 0.08071082, 0.08071082, 0.08071082, 
    0.08071082, 0.07622877, 0.07622877, 0.07622877, 0.07622877, 0.07622877, 
    0.07622877, 0.07622877, 0.07787628, 0.07787628, 0.07787628, 0.07787628, 
    0.07787628, 0.07787628, 0.07787628, 0.08297741, 0.08297741, 0.08297741, 
    0.08297741, 0.08297741, 0.08297741, 0.08297741, 0.08071082,
  0.09177209, 0.08587226, 0.0763882, 0.0673634, 0.07087537, 0.06532107, 
    0.05628275, 0.06440875, 0.07564017, 0.08069164, 0.08512881, 0.09966984, 
    0.1088848, 0.2138387, 0.2593633, 0.2472876, 0.2177646, 0.1768466, 
    0.1520493, 0.1410581, 0.1486063, 0.1473601, 0.1900543, 0.296037, 
    0.3014785, 0.2644227, 0.252014, 0.1774445, 0.1007247,
  0.1990761, 0.2112598, 0.2618232, 0.2701442, 0.180685, 0.2486603, 0.3250742, 
    0.1186253, 0.0969736, 0.1142467, 0.07381049, 0.09559183, 0.3233508, 
    0.5691997, 0.6031502, 0.5363937, 0.496557, 0.4560255, 0.3338142, 
    0.2742659, 0.2575813, 0.2421103, 0.2461818, 0.2707858, 0.3488727, 
    0.3612334, 0.3207927, 0.2850892, 0.222442,
  0.2929258, 0.2102416, 0.1916393, 0.2578033, 0.592626, 0.7989929, 0.724048, 
    0.5316787, 0.3470942, 0.2559559, 0.2698637, 0.34828, 0.5038077, 0.626334, 
    0.8180032, 1.115857, 1.174616, 1.033374, 0.816838, 0.6189668, 0.441486, 
    0.3474948, 0.3185686, 0.3262998, 0.3529034, 0.4516902, 0.4968972, 
    0.51771, 0.3961072,
  1.211326, 0.848639, 0.707123, 1.186771, 1.473964, 1.63599, 1.60319, 
    1.392597, 0.9841228, 0.6878771, 0.6833595, 0.800423, 0.9574479, 1.284583, 
    1.515357, 1.435699, 1.442528, 1.197292, 1.022906, 0.9221973, 0.7534289, 
    0.6735324, 0.6081228, 0.5554314, 0.7759966, 1.306079, 1.889402, 1.906487, 
    1.545048,
  2.877755, 2.425665, 2.595966, 2.750236, 3.242963, 3.28719, 2.833904, 
    2.393451, 2.17668, 1.855114, 1.839347, 2.167505, 2.349552, 2.45286, 
    2.036804, 1.908278, 1.674262, 1.430418, 1.216842, 1.084693, 0.9239119, 
    0.9029429, 0.8094769, 0.6293678, 1.637232, 3.222525, 3.50694, 3.615607, 
    3.319327,
  3.923971, 4.060248, 5.95982, 6.257867, 5.538871, 4.395675, 3.802013, 
    3.215719, 2.608429, 2.545143, 2.849895, 3.069555, 2.998919, 2.788551, 
    2.389709, 1.969493, 1.590984, 1.330783, 1.102806, 0.9591168, 0.8579391, 
    0.9439815, 1.028324, 1.756871, 3.192478, 4.620824, 5.408517, 5.137064, 
    4.424211,
  6.549183, 10.99764, 12.70147, 9.071527, 7.038162, 4.437501, 2.965088, 
    2.389318, 2.871005, 3.545969, 4.849615, 3.900488, 3.276691, 2.59408, 
    2.010925, 1.585225, 1.245234, 1.117103, 0.9704633, 0.84388, 0.8026852, 
    1.363225, 2.997618, 7.818314, 10.94515, 10.70442, 8.144175, 6.167489, 
    5.61585,
  9.189305, 17.91838, 18.51675, 10.15611, 4.939802, 2.634798, 2.107072, 
    2.539794, 4.254849, 4.595731, 3.988465, 4.115536, 2.447207, 1.02215, 
    0.728763, 0.6299145, 0.7149287, 0.7867177, 0.7178532, 0.773934, 
    0.8459571, 1.56195, 6.096308, 16.13019, 16.01598, 12.63363, 7.579506, 
    5.75605, 6.686267,
  10.91703, 20.2082, 19.10379, 7.311253, 4.791693, 2.682266, 2.576332, 
    2.903803, 7.378207, 10.25965, 3.285668, 2.064154, 0.903645, 0.558856, 
    0.4747156, 0.4884982, 0.5141832, 0.6012161, 0.7708431, 0.9427376, 
    1.248225, 2.616604, 7.601067, 17.0926, 15.17185, 10.03189, 6.747217, 
    6.821091, 8.097964,
  13.82625, 15.80731, 14.26532, 7.465805, 5.574113, 4.238484, 4.634077, 
    4.55997, 5.951771, 4.75701, 2.933461, 1.600044, 1.025609, 0.775983, 
    0.6913134, 0.6922045, 0.7268102, 0.8147818, 1.065004, 1.479301, 2.089037, 
    3.128736, 7.144079, 11.00892, 8.820794, 7.39422, 7.618247, 8.957538, 
    13.13255,
  6.906364, 7.66588, 7.787841, 6.86305, 7.106474, 7.219933, 7.758297, 
    7.937933, 8.81791, 6.23325, 4.813989, 3.192454, 2.455939, 2.475833, 
    2.368194, 2.173678, 1.83721, 1.650301, 1.607277, 1.876496, 3.109636, 
    4.26865, 3.522266, 3.830844, 3.914768, 3.563865, 3.636352, 4.852513, 
    6.112382,
  2.571446, 2.67318, 2.678671, 3.51612, 3.781162, 4.122192, 5.267681, 
    5.946747, 7.135581, 9.860818, 8.446424, 7.002515, 5.949853, 5.239192, 
    4.404627, 3.779557, 3.696739, 3.068014, 2.495443, 2.412719, 3.293378, 
    3.97145, 4.682057, 4.404889, 3.655493, 3.819284, 3.293746, 2.893315, 
    2.849962,
  2.844232, 2.764533, 2.981534, 2.211098, 3.729357, 2.858449, 2.106281, 
    4.861905, 4.952366, 5.347178, 5.53228, 4.871505, 4.900459, 4.781469, 
    4.211824, 3.773423, 3.603543, 3.517261, 3.109274, 2.509728, 2.173017, 
    3.640026, 4.418283, 4.777261, 4.691918, 4.50599, 3.770501, 3.193157, 
    2.780944,
  2.509405, 2.64339, 3.30407, 3.564104, 4.113014, 3.729035, 3.007977, 
    2.255697, 2.942712, 3.464773, 3.640634, 3.502054, 3.511987, 3.192944, 
    3.122575, 3.04387, 2.787568, 2.277079, 2.319682, 1.820633, 2.310623, 
    2.809855, 2.704653, 2.047027, 2.420127, 2.676208, 2.758184, 2.862318, 
    2.662495,
  1.562109, 1.427013, 2.182531, 2.672388, 3.094432, 2.818684, 2.832934, 
    2.668563, 2.447912, 2.777264, 3.168879, 2.259399, 1.650932, 2.002541, 
    2.076979, 1.78723, 1.495462, 1.425949, 1.24912, 1.36147, 1.484659, 
    1.380543, 1.567808, 1.41232, 1.799279, 1.838225, 1.843831, 1.729378, 
    1.579232,
  0.950395, 0.9237912, 1.012719, 1.395963, 1.421884, 1.387407, 1.284948, 
    1.104195, 0.911388, 1.111135, 0.9830497, 1.037938, 1.114591, 1.211123, 
    1.35051, 1.425741, 1.206574, 1.021391, 1.082467, 1.042918, 0.8027951, 
    0.7179716, 0.8012362, 0.8403285, 1.286327, 0.5529941, 0.3224928, 
    1.009932, 0.9688846,
  0.3753633, 0.3757688, 0.388393, 0.4103114, 0.4193218, 0.4210998, 0.4455628, 
    0.4827083, 0.530543, 0.565793, 0.5788566, 0.5827208, 0.6117056, 
    0.6273996, 0.5827948, 0.5417993, 0.5365022, 0.5108492, 0.4702306, 
    0.4322841, 0.4114461, 0.3995463, 0.3375311, 0.3611318, 0.3512372, 
    0.1838593, 0.1817371, 0.3196405, 0.3927347,
  0.1330787, 0.1330787, 0.1330787, 0.1330787, 0.1330787, 0.1330787, 
    0.1330787, 0.1283427, 0.1283427, 0.1283427, 0.1283427, 0.1283427, 
    0.1283427, 0.1283427, 0.1306274, 0.1306274, 0.1306274, 0.1306274, 
    0.1306274, 0.1306274, 0.1306274, 0.1362982, 0.1362982, 0.1362982, 
    0.1362982, 0.1362982, 0.1362982, 0.1362982, 0.1330787,
  0.1716765, 0.1484769, 0.1362556, 0.1249054, 0.1314096, 0.1232645, 
    0.1137184, 0.1212273, 0.1331175, 0.1340479, 0.1484156, 0.1724424, 
    0.1882564, 0.3380137, 0.4077721, 0.3982851, 0.3753088, 0.3234501, 
    0.2845097, 0.2635525, 0.268375, 0.2568586, 0.3067993, 0.4219744, 
    0.4342735, 0.4013499, 0.3822705, 0.2914293, 0.1838874,
  0.3498477, 0.3837142, 0.4324802, 0.4362815, 0.3162405, 0.3998937, 
    0.4904324, 0.2517542, 0.2167154, 0.2289109, 0.1489635, 0.1988777, 
    0.5341578, 0.9029784, 0.9554787, 0.8607975, 0.8173537, 0.7467905, 
    0.5667945, 0.4835503, 0.4523869, 0.4149168, 0.4205684, 0.4464623, 
    0.5692171, 0.5659886, 0.5355951, 0.4813122, 0.3887414,
  0.5268769, 0.3904783, 0.3524249, 0.4684101, 0.8635717, 1.057422, 0.9855074, 
    0.8141714, 0.5766236, 0.457911, 0.4944508, 0.6429992, 0.8770316, 
    1.049025, 1.339931, 1.607355, 1.647469, 1.495802, 1.246016, 0.9505928, 
    0.7016488, 0.5455236, 0.4988361, 0.5238608, 0.5624983, 0.67509, 
    0.7279848, 0.7927722, 0.6537728,
  1.536375, 1.129096, 0.992658, 1.5766, 1.875158, 2.015714, 1.974171, 
    1.73094, 1.301406, 0.9634368, 0.9415329, 1.092215, 1.320338, 1.782555, 
    2.037096, 2.004452, 1.913743, 1.605836, 1.402153, 1.212179, 0.9874421, 
    0.9033754, 0.7970868, 0.727111, 0.9708233, 1.51114, 2.159404, 2.159594, 
    1.896826,
  3.236833, 2.819775, 3.200279, 3.362239, 3.829865, 3.812462, 3.269907, 
    2.818087, 2.628976, 2.30798, 2.26498, 2.595264, 2.790681, 3.048232, 
    2.626348, 2.370205, 2.080429, 1.744679, 1.484264, 1.29706, 1.084828, 
    1.025897, 0.9217736, 0.795652, 2.01109, 3.633531, 3.767505, 3.952764, 
    3.667928,
  4.324335, 4.307743, 6.146826, 6.623487, 5.807827, 4.79972, 4.234104, 
    3.613942, 2.88036, 2.691244, 3.106373, 3.623516, 3.56126, 3.162463, 
    2.759979, 2.297647, 1.853252, 1.519913, 1.192801, 1.024145, 0.8967326, 
    0.9689401, 1.025089, 1.596571, 3.423965, 5.114696, 5.753984, 5.582607, 
    4.822219,
  6.444798, 10.35223, 12.58512, 9.080102, 7.324626, 4.837164, 3.248397, 
    2.485011, 2.748553, 3.392682, 4.970663, 4.026296, 3.40787, 2.749757, 
    2.124216, 1.640413, 1.26549, 1.110105, 0.9714741, 0.8200095, 0.7849033, 
    1.306426, 2.64868, 7.17881, 10.95783, 10.77759, 8.236727, 6.282749, 
    5.785271,
  9.006404, 17.13972, 18.84077, 10.40384, 5.27314, 2.853097, 2.180155, 
    2.482378, 3.908297, 4.414589, 3.862666, 3.872593, 2.497425, 1.03097, 
    0.7136157, 0.6110714, 0.6925162, 0.7495727, 0.6834853, 0.7420033, 
    0.7755857, 1.583856, 5.981533, 16.74541, 16.55175, 12.92523, 7.639911, 
    5.786067, 7.000722,
  11.11963, 20.68262, 19.48422, 7.482239, 5.195488, 2.877542, 2.556285, 
    2.791583, 7.370695, 10.14904, 3.309488, 1.988543, 0.896367, 0.5328207, 
    0.4590046, 0.4736237, 0.4983452, 0.5810398, 0.729308, 0.9292967, 
    1.213988, 2.621178, 7.542295, 17.69524, 15.37934, 9.718254, 6.723905, 
    6.958571, 8.25676,
  13.97083, 15.91008, 14.21786, 8.270159, 5.79038, 4.30502, 4.566159, 
    4.316864, 5.715101, 4.55466, 2.987031, 1.618902, 1.048573, 0.805638, 
    0.7129495, 0.7022437, 0.7192921, 0.8088117, 1.055708, 1.476609, 2.05375, 
    3.063584, 6.954849, 11.00173, 8.760146, 7.484859, 7.587631, 8.889332, 
    13.45108,
  6.703546, 7.400798, 7.618818, 6.489532, 7.028275, 7.246546, 7.685129, 
    8.047466, 8.943175, 6.232702, 4.959711, 3.380258, 2.608416, 2.629034, 
    2.471565, 2.266971, 1.946067, 1.778664, 1.675445, 1.883523, 3.012681, 
    4.468259, 3.517088, 3.72618, 3.745214, 3.469895, 3.541278, 4.616012, 
    5.763069,
  3.128495, 3.017413, 2.981841, 3.926428, 4.257659, 4.647546, 5.6175, 
    6.204237, 8.058701, 11.04338, 9.382921, 7.582377, 6.415586, 5.635734, 
    4.858216, 4.266398, 3.974862, 3.305888, 2.668948, 2.638109, 3.721826, 
    4.487069, 5.091783, 4.683568, 3.84395, 4.061883, 3.562732, 3.186822, 
    3.370731,
  3.580743, 3.551572, 4.173249, 3.537841, 5.424381, 4.295325, 3.522562, 
    6.81228, 7.107326, 7.394794, 7.259262, 6.288662, 6.082569, 5.776351, 
    5.023536, 4.35502, 4.09826, 3.893274, 3.451724, 2.926486, 2.731803, 
    4.665808, 5.234943, 5.557966, 5.30991, 5.083409, 4.321669, 3.692224, 
    3.391231,
  3.286343, 3.889346, 4.668254, 4.883482, 5.498586, 5.23183, 4.480425, 
    3.706926, 4.421587, 4.913239, 5.187113, 4.927904, 4.745597, 4.38127, 
    4.129901, 3.920918, 3.473779, 2.957074, 3.025636, 2.657884, 3.224154, 
    3.875843, 3.743662, 3.062897, 3.427432, 3.518641, 3.437896, 3.562225, 
    3.359967,
  2.361205, 2.39505, 3.41655, 3.887796, 4.376749, 4.379688, 4.389987, 
    4.151645, 3.828143, 4.320919, 4.566692, 3.458353, 2.86252, 3.156305, 
    3.117701, 2.685751, 2.244161, 2.155805, 1.920004, 2.1368, 2.350863, 
    2.18766, 2.393856, 2.313141, 2.815332, 2.799692, 2.691456, 2.57783, 
    2.402508,
  1.746856, 1.805592, 1.965909, 2.326404, 2.322961, 2.253111, 2.145404, 
    1.997015, 1.773356, 1.920561, 1.696966, 1.847973, 2.026001, 2.097253, 
    2.193568, 2.163557, 1.928939, 1.784625, 1.83882, 1.754875, 1.447198, 
    1.352459, 1.494917, 1.598848, 2.043369, 1.135627, 0.7260664, 1.744562, 
    1.798544,
  0.9181513, 0.9215679, 0.9586348, 0.9944266, 0.975172, 0.9546111, 0.9542877, 
    1.002681, 1.060242, 1.098237, 1.12171, 1.133821, 1.191036, 1.192435, 
    1.169778, 1.172066, 1.174936, 1.095523, 1.021406, 0.9633055, 0.9190491, 
    0.8971979, 0.7617536, 0.7874866, 0.7920572, 0.4930344, 0.5140378, 
    0.8066629, 0.95183,
  0.1946154, 0.1946154, 0.1946154, 0.1946154, 0.1946154, 0.1946154, 
    0.1946154, 0.1892021, 0.1892021, 0.1892021, 0.1892021, 0.1892021, 
    0.1892021, 0.1892021, 0.1965302, 0.1965302, 0.1965302, 0.1965302, 
    0.1965302, 0.1965302, 0.1965302, 0.202504, 0.202504, 0.202504, 0.202504, 
    0.202504, 0.202504, 0.202504, 0.1946154,
  0.272545, 0.2262737, 0.2057744, 0.1953246, 0.2088844, 0.1963222, 0.185475, 
    0.1894417, 0.2045034, 0.2059805, 0.2282314, 0.2600901, 0.2833823, 
    0.4597501, 0.5493384, 0.5505245, 0.5330765, 0.4788549, 0.4343566, 
    0.3974189, 0.3978107, 0.3771752, 0.416535, 0.5249157, 0.534869, 
    0.5064081, 0.481064, 0.3971444, 0.2927504,
  0.4984062, 0.5445061, 0.5866772, 0.5860522, 0.4668801, 0.5466439, 
    0.6230033, 0.3977668, 0.3521993, 0.3609512, 0.2797538, 0.3558944, 
    0.7715436, 1.169693, 1.237201, 1.160229, 1.130533, 1.041254, 0.8175888, 
    0.7048485, 0.6388047, 0.5629801, 0.5700341, 0.6084127, 0.7540456, 
    0.7239363, 0.733219, 0.6612487, 0.5396796,
  0.7351401, 0.5811215, 0.5360919, 0.6768522, 1.055496, 1.22464, 1.147056, 
    1.008473, 0.7672443, 0.6486959, 0.6948997, 0.913233, 1.267488, 1.470633, 
    1.89496, 2.023918, 1.999897, 1.809596, 1.578495, 1.238959, 0.9447227, 
    0.7374361, 0.6800733, 0.6995643, 0.778767, 0.8749229, 0.9262716, 
    1.001483, 0.8810419,
  1.733048, 1.329947, 1.218126, 1.800283, 2.092357, 2.210692, 2.190459, 
    1.88713, 1.497453, 1.163352, 1.135878, 1.28142, 1.659368, 2.262371, 
    2.556278, 2.505216, 2.23162, 1.936322, 1.689705, 1.433347, 1.173712, 
    1.079316, 0.9351228, 0.8585086, 1.130272, 1.609319, 2.269248, 2.307743, 
    2.071851,
  3.363508, 2.994412, 3.450411, 3.715993, 4.103307, 4.048148, 3.443135, 
    3.00747, 2.825602, 2.584506, 2.4719, 2.814361, 3.040449, 3.460483, 
    3.061959, 2.767344, 2.399308, 1.987735, 1.710574, 1.456706, 1.193736, 
    1.08847, 0.9860264, 0.9522752, 2.294541, 3.753757, 3.706577, 3.901232, 
    3.769786,
  4.513144, 4.382123, 6.16298, 6.692126, 5.787651, 4.95313, 4.391266, 
    3.87595, 3.138061, 2.793692, 3.397831, 4.006884, 4.028124, 3.392362, 
    3.033064, 2.565056, 2.102125, 1.686019, 1.270248, 1.057361, 0.9067522, 
    0.9601415, 0.9938592, 1.374483, 3.712596, 5.286367, 5.704573, 5.592571, 
    4.924725,
  6.121963, 9.282945, 11.84007, 8.631808, 7.341736, 5.090025, 3.577145, 
    2.581866, 2.68963, 3.318009, 5.011747, 4.102841, 3.568501, 2.913578, 
    2.24392, 1.704403, 1.287316, 1.100426, 0.9481202, 0.7965229, 0.7592892, 
    1.181451, 2.219078, 6.151409, 10.70534, 10.7439, 8.033927, 6.20491, 
    5.666893,
  8.621758, 15.96184, 18.61125, 10.16164, 5.442359, 3.070614, 2.286038, 
    2.432428, 3.559619, 4.124143, 3.647476, 3.638314, 2.49384, 1.085607, 
    0.698507, 0.5998842, 0.6779622, 0.7106737, 0.6544743, 0.7025661, 
    0.7078719, 1.466804, 5.585078, 16.6683, 16.8115, 12.93024, 7.575573, 
    5.689758, 6.979741,
  11.04755, 20.60197, 19.22957, 7.456471, 5.409341, 3.066556, 2.600021, 
    2.734727, 7.177102, 9.916286, 3.296832, 1.907164, 0.872951, 0.5152211, 
    0.4509457, 0.4547398, 0.4863935, 0.5594638, 0.685777, 0.891609, 1.158019, 
    2.477587, 6.810991, 17.31853, 14.60355, 9.105037, 6.551595, 6.954893, 
    8.154229,
  13.85165, 15.56899, 13.6649, 8.625851, 5.915653, 4.361215, 4.495153, 
    4.102986, 5.409892, 4.308475, 2.932981, 1.650393, 1.082649, 0.8532158, 
    0.7331027, 0.7169331, 0.7152905, 0.8087488, 1.053902, 1.464347, 2.016042, 
    3.006087, 6.514231, 10.45226, 8.102962, 7.304583, 7.321364, 8.664417, 
    13.49643,
  6.326561, 7.006079, 7.215897, 5.87921, 6.687404, 6.989439, 7.604631, 
    8.105766, 9.023234, 6.242763, 5.029125, 3.488681, 2.745351, 2.782414, 
    2.53342, 2.362065, 2.042073, 1.88948, 1.735194, 1.882132, 2.902127, 
    4.464179, 3.447152, 3.335023, 3.394376, 3.19518, 3.372147, 4.344656, 
    5.387192,
  3.613359, 3.311632, 3.251084, 4.290275, 4.654094, 5.124593, 5.968435, 
    6.47677, 9.054654, 11.95719, 10.01728, 7.906077, 6.662151, 5.931773, 
    5.265461, 4.619717, 4.147499, 3.430361, 2.733058, 2.746309, 4.021603, 
    4.845934, 5.337714, 4.855401, 3.958276, 4.192286, 3.790278, 3.340251, 
    3.757916,
  4.243879, 4.276568, 5.193917, 4.823467, 7.00869, 5.984853, 5.204048, 
    8.732668, 9.188703, 9.215751, 8.858329, 7.670772, 7.134367, 6.557612, 
    5.752995, 4.838466, 4.566204, 4.160093, 3.615338, 3.179881, 3.259906, 
    5.617774, 5.876964, 6.107175, 5.765235, 5.490509, 4.63633, 4.057524, 
    3.930264,
  3.905981, 4.916885, 5.704734, 6.09054, 6.568939, 6.404267, 5.675853, 
    5.084295, 5.723423, 6.228168, 6.707339, 6.119291, 5.825634, 5.387978, 
    4.953563, 4.65652, 4.082726, 3.523051, 3.610178, 3.493638, 3.961993, 
    4.913135, 4.718489, 4.037408, 4.311907, 4.222349, 3.999574, 4.086833, 
    3.910178,
  3.055896, 3.326744, 4.319734, 4.777446, 5.522528, 5.68697, 5.657909, 
    5.413011, 5.086527, 5.411013, 5.564834, 4.545703, 3.978623, 4.147812, 
    4.005154, 3.459238, 2.941521, 2.850663, 2.592618, 2.948951, 3.189868, 
    3.104215, 3.169784, 3.234386, 3.682366, 3.64001, 3.399117, 3.325437, 
    3.106395,
  2.596626, 2.741985, 2.879433, 3.148323, 3.171368, 3.086612, 3.080328, 
    3.019871, 2.769635, 2.732255, 2.484832, 2.744772, 3.029801, 2.990298, 
    3.006209, 2.808715, 2.612517, 2.537535, 2.527585, 2.376497, 2.065622, 
    1.99671, 2.186944, 2.390718, 2.75788, 1.825322, 1.271731, 2.486714, 
    2.622416,
  1.572363, 1.607865, 1.732246, 1.774177, 1.719716, 1.691543, 1.680005, 
    1.709298, 1.752451, 1.797269, 1.831884, 1.890454, 1.981797, 1.971193, 
    1.903803, 1.881563, 1.850433, 1.737492, 1.649884, 1.577185, 1.533002, 
    1.516898, 1.321111, 1.367812, 1.390356, 0.9998843, 1.06357, 1.448582, 
    1.602322,
  0.2565826, 0.2565826, 0.2565826, 0.2565826, 0.2565826, 0.2565826, 
    0.2565826, 0.2532023, 0.2532023, 0.2532023, 0.2532023, 0.2532023, 
    0.2532023, 0.2532023, 0.265802, 0.265802, 0.265802, 0.265802, 0.265802, 
    0.265802, 0.265802, 0.2714462, 0.2714462, 0.2714462, 0.2714462, 
    0.2714462, 0.2714462, 0.2714462, 0.2565826,
  0.3724229, 0.3113475, 0.2902049, 0.2764471, 0.2867877, 0.2739436, 
    0.2584454, 0.2647559, 0.2818916, 0.2885511, 0.3108221, 0.3499271, 
    0.3867388, 0.5556834, 0.6531422, 0.6675998, 0.6441711, 0.5939983, 
    0.5570177, 0.512965, 0.4976947, 0.4785304, 0.5084869, 0.5855984, 
    0.5832546, 0.5600885, 0.5394996, 0.4726706, 0.3994634,
  0.6183556, 0.6557678, 0.7015169, 0.6919683, 0.6075004, 0.6687728, 0.701507, 
    0.5285804, 0.4771799, 0.480458, 0.4440107, 0.5469179, 0.9455163, 
    1.301955, 1.398797, 1.341554, 1.327046, 1.234873, 0.9920167, 0.8558739, 
    0.764025, 0.66474, 0.6735297, 0.7162709, 0.8385455, 0.83434, 0.8968916, 
    0.8014784, 0.6560931,
  0.9161394, 0.749453, 0.697919, 0.8358834, 1.180656, 1.315931, 1.229416, 
    1.101279, 0.877135, 0.776937, 0.8250837, 1.105486, 1.558687, 1.83374, 
    2.262007, 2.287512, 2.19277, 1.978903, 1.763692, 1.406718, 1.102993, 
    0.8985882, 0.8133149, 0.8060481, 0.9419376, 1.03551, 1.099828, 1.143047, 
    1.056567,
  1.82421, 1.465989, 1.354007, 1.895628, 2.148026, 2.223038, 2.230709, 
    1.941462, 1.603423, 1.293819, 1.261695, 1.409982, 1.940847, 2.562914, 
    2.96179, 2.846814, 2.417059, 2.155337, 1.874679, 1.571276, 1.308264, 
    1.179286, 1.00872, 0.9617597, 1.23041, 1.678599, 2.335489, 2.417779, 
    2.146594,
  3.318294, 3.047669, 3.461979, 3.826959, 4.083542, 4.026097, 3.421729, 
    3.050916, 2.826159, 2.657658, 2.526943, 2.86861, 3.139304, 3.654318, 
    3.407893, 3.044446, 2.594993, 2.133091, 1.872898, 1.553947, 1.267372, 
    1.125232, 1.027523, 1.07108, 2.442934, 3.665151, 3.564583, 3.695397, 
    3.71213,
  4.480204, 4.372833, 6.109309, 6.607831, 5.648417, 4.916, 4.366673, 
    4.024415, 3.334454, 2.873489, 3.597715, 4.248627, 4.324492, 3.532603, 
    3.175902, 2.769902, 2.290696, 1.801182, 1.338707, 1.079304, 0.9218863, 
    0.9359596, 0.9372056, 1.154868, 3.844416, 5.168778, 5.465443, 5.366489, 
    4.781178,
  5.768852, 8.259574, 11.00966, 8.129182, 7.038859, 5.046632, 3.795972, 
    2.745662, 2.708864, 3.227034, 4.966936, 4.11199, 3.676101, 3.089081, 
    2.35495, 1.780756, 1.297139, 1.093068, 0.9197174, 0.775461, 0.7200921, 
    1.007856, 1.840884, 5.209528, 10.18896, 10.67389, 7.600768, 5.971227, 
    5.435805,
  8.132775, 14.48193, 17.94423, 9.559702, 5.519503, 3.259834, 2.410026, 
    2.39886, 3.259262, 3.736218, 3.416825, 3.432456, 2.423253, 1.148949, 
    0.7041299, 0.5905707, 0.6676944, 0.6809753, 0.6226659, 0.6598065, 
    0.6423874, 1.326353, 4.863555, 15.85105, 16.6685, 12.50877, 7.245654, 
    5.45911, 6.725656,
  10.50207, 19.85955, 18.04313, 7.328711, 5.450818, 3.27703, 2.683214, 
    2.687079, 6.758778, 9.490664, 3.208385, 1.826843, 0.8405729, 0.512862, 
    0.4465941, 0.4359003, 0.4737628, 0.5370029, 0.6470811, 0.8450962, 
    1.05771, 2.182846, 5.837395, 16.15635, 12.98738, 8.340603, 6.321928, 
    6.692098, 7.825662,
  13.51359, 14.86368, 12.95168, 8.799242, 5.864622, 4.406782, 4.431239, 
    3.983941, 5.137119, 4.062613, 2.845981, 1.680119, 1.121072, 0.9067357, 
    0.7625715, 0.7435375, 0.7177796, 0.8058957, 1.043772, 1.455185, 1.984097, 
    2.878126, 5.928409, 9.501247, 7.170805, 6.78935, 6.832322, 8.317949, 
    13.15473,
  6.015293, 6.575436, 6.593215, 5.210269, 6.276824, 6.515306, 7.409455, 
    7.994467, 8.96734, 6.198538, 4.967204, 3.503812, 2.81653, 2.900292, 
    2.590416, 2.463408, 2.122506, 1.970576, 1.77015, 1.870235, 2.74102, 
    4.338591, 3.313283, 2.992287, 2.93525, 2.849755, 3.155668, 4.066975, 
    5.040906,
  3.970571, 3.476727, 3.443116, 4.650577, 5.041082, 5.462388, 6.283245, 
    6.749118, 10.1817, 12.83167, 10.38406, 8.002528, 6.787604, 6.157584, 
    5.628221, 4.844558, 4.205315, 3.471622, 2.745767, 2.809139, 4.213446, 
    5.053631, 5.471472, 4.929437, 4.012293, 4.21577, 3.9447, 3.416323, 
    4.007053,
  4.793109, 4.891361, 6.082687, 6.007003, 8.269315, 7.486024, 6.91762, 
    10.55734, 10.97053, 10.89647, 10.36254, 8.815634, 7.973355, 7.165779, 
    6.343559, 5.234424, 4.897531, 4.353772, 3.699919, 3.35219, 3.809011, 
    6.170402, 6.285843, 6.449538, 6.068291, 5.751578, 4.848901, 4.321446, 
    4.366555,
  4.428134, 5.596155, 6.479706, 7.066633, 7.420906, 7.282653, 6.626321, 
    6.308638, 6.916953, 7.518704, 7.939589, 7.040371, 6.654356, 6.215273, 
    5.717312, 5.229169, 4.595657, 3.959339, 4.033051, 4.148101, 4.585637, 
    5.71571, 5.555292, 4.883295, 5.030816, 4.76985, 4.460426, 4.416492, 
    4.287646,
  3.577497, 4.012982, 4.951605, 5.515929, 6.390654, 6.660339, 6.661291, 
    6.464778, 6.123216, 6.224639, 6.45621, 5.44006, 4.94378, 4.875726, 
    4.70874, 4.090816, 3.525523, 3.423189, 3.208667, 3.621523, 3.771693, 
    3.796283, 3.786585, 3.944026, 4.34562, 4.347627, 3.944562, 3.886662, 
    3.589219,
  3.293842, 3.553718, 3.696906, 3.889072, 3.884048, 3.758919, 3.837691, 
    3.852591, 3.62765, 3.425493, 3.205763, 3.574082, 3.880061, 3.73308, 
    3.685625, 3.327829, 3.144995, 3.116229, 3.009947, 2.854655, 2.524876, 
    2.532498, 2.797795, 3.056955, 3.342407, 2.504572, 1.894223, 3.072246, 
    3.29179,
  2.205934, 2.257762, 2.419031, 2.446373, 2.409798, 2.441947, 2.490519, 
    2.504847, 2.517676, 2.559411, 2.602747, 2.700211, 2.778389, 2.723808, 
    2.619226, 2.540196, 2.455549, 2.304893, 2.22406, 2.157554, 2.129929, 
    2.11997, 1.890536, 1.946104, 2.005802, 1.602302, 1.671064, 2.062695, 
    2.222348,
  0.3135954, 0.3135954, 0.3135954, 0.3135954, 0.3135954, 0.3135954, 
    0.3135954, 0.3108048, 0.3108048, 0.3108048, 0.3108048, 0.3108048, 
    0.3108048, 0.3108048, 0.3277778, 0.3277778, 0.3277778, 0.3277778, 
    0.3277778, 0.3277778, 0.3277778, 0.3328542, 0.3328542, 0.3328542, 
    0.3328542, 0.3328542, 0.3328542, 0.3328542, 0.3135954,
  0.4482261, 0.3872498, 0.3714812, 0.3548845, 0.3603036, 0.3493512, 
    0.3272249, 0.3342814, 0.3533554, 0.368635, 0.3847704, 0.4264539, 
    0.4752624, 0.605049, 0.6946531, 0.7218022, 0.6924464, 0.6532481, 
    0.6276722, 0.5949988, 0.5656834, 0.5514166, 0.5736781, 0.6067263, 
    0.5886863, 0.5725276, 0.5657346, 0.5230679, 0.4743844,
  0.6981878, 0.7329848, 0.7703708, 0.7585392, 0.7173105, 0.7548752, 0.730512, 
    0.6255565, 0.5822493, 0.5734644, 0.5840588, 0.7081172, 1.008406, 
    1.315907, 1.439779, 1.403022, 1.402887, 1.314477, 1.073724, 0.9166301, 
    0.8190982, 0.7163976, 0.7185576, 0.7715449, 0.8640987, 0.8914078, 
    0.9997185, 0.8740836, 0.7266143,
  1.060854, 0.8842164, 0.8209924, 0.9288934, 1.242126, 1.337536, 1.244412, 
    1.13272, 0.9249645, 0.8328809, 0.8635679, 1.205536, 1.743833, 2.026335, 
    2.36134, 2.38381, 2.274622, 2.031579, 1.827118, 1.482579, 1.179253, 
    0.9936608, 0.8860659, 0.8627888, 1.054778, 1.129013, 1.23025, 1.254939, 
    1.175955,
  1.853321, 1.542892, 1.40504, 1.899572, 2.092299, 2.140604, 2.184746, 
    1.939323, 1.626812, 1.346028, 1.322294, 1.483177, 2.127397, 2.7331, 
    3.108907, 2.972083, 2.497937, 2.242482, 1.958752, 1.633833, 1.370071, 
    1.22677, 1.046118, 1.033837, 1.284226, 1.741557, 2.335955, 2.43716, 
    2.144946,
  3.12665, 2.967407, 3.342142, 3.732579, 3.92277, 3.854321, 3.27282, 
    2.993399, 2.733818, 2.606363, 2.488995, 2.829504, 3.138994, 3.725425, 
    3.620449, 3.16793, 2.698161, 2.217097, 1.969093, 1.597692, 1.305411, 
    1.140863, 1.046567, 1.137099, 2.509726, 3.475044, 3.383125, 3.385558, 
    3.499769,
  4.327167, 4.24766, 6.078471, 6.396536, 5.446119, 4.753006, 4.184693, 
    4.00842, 3.400142, 2.884688, 3.715088, 4.321806, 4.486976, 3.562486, 
    3.262067, 2.927943, 2.408981, 1.877165, 1.38598, 1.097834, 0.938483, 
    0.8926911, 0.8771327, 0.9676806, 3.825854, 4.977568, 5.080911, 4.943985, 
    4.511994,
  5.289886, 7.321214, 10.35581, 7.679375, 6.47566, 4.803793, 3.824533, 
    2.870813, 2.715877, 3.122276, 4.791545, 4.069474, 3.719916, 3.275766, 
    2.483381, 1.846403, 1.309446, 1.092008, 0.9090036, 0.7521217, 0.6732791, 
    0.8847029, 1.580411, 4.496429, 9.399604, 10.4039, 7.052663, 5.587336, 
    5.238038,
  7.568786, 12.95183, 16.85013, 8.701469, 5.343126, 3.405305, 2.50029, 
    2.344702, 2.944143, 3.318301, 3.221517, 3.220014, 2.282271, 1.18777, 
    0.7318332, 0.5971454, 0.65175, 0.6556804, 0.5915162, 0.6042992, 
    0.5999938, 1.201357, 3.987904, 14.34782, 16.01467, 11.82666, 6.681821, 
    5.241634, 6.33075,
  9.816138, 18.49056, 16.03991, 6.90653, 5.279884, 3.429034, 2.762042, 
    2.617266, 6.186564, 8.742911, 3.020597, 1.735363, 0.8171138, 0.5319191, 
    0.4458879, 0.4174635, 0.4491245, 0.5189599, 0.6151484, 0.7968667, 
    0.9244711, 1.825661, 4.802149, 14.15445, 11.00603, 7.400893, 6.115987, 
    6.323929, 7.324847,
  12.97645, 13.90906, 12.10898, 8.732548, 5.568367, 4.381463, 4.423173, 
    3.919677, 4.98812, 3.855026, 2.768252, 1.728221, 1.163408, 0.9554741, 
    0.798678, 0.7709298, 0.7200374, 0.8024533, 1.044604, 1.411007, 1.896282, 
    2.758566, 5.32181, 8.365319, 5.892754, 5.982018, 6.126791, 7.813483, 
    12.57136,
  5.68439, 6.087795, 5.884087, 4.628305, 5.875701, 5.975309, 7.06895, 
    7.665643, 8.790406, 6.105726, 4.826569, 3.45066, 2.8146, 2.974036, 
    2.686397, 2.585214, 2.184242, 2.060169, 1.79159, 1.837027, 2.60525, 
    4.112287, 3.111362, 2.784894, 2.504128, 2.587975, 2.982194, 3.808144, 
    4.624606,
  4.219858, 3.613202, 3.584191, 4.909483, 5.376372, 5.705929, 6.613315, 
    7.075901, 11.26971, 13.77246, 10.64717, 8.036753, 6.81761, 6.210262, 
    5.916296, 4.964904, 4.215569, 3.441391, 2.732642, 2.856247, 4.35845, 
    5.118994, 5.467711, 4.872158, 3.991363, 4.164944, 4.020387, 3.473786, 
    4.160182,
  5.163042, 5.331562, 6.780991, 6.995649, 9.084055, 8.590014, 8.502094, 
    12.14038, 12.4144, 12.32705, 11.63509, 9.792661, 8.676993, 7.622891, 
    6.810771, 5.550751, 5.126992, 4.478838, 3.762435, 3.506381, 4.138699, 
    6.455429, 6.484136, 6.667694, 6.245692, 5.861362, 4.933199, 4.494602, 
    4.63179,
  4.785144, 6.00626, 6.956026, 7.77942, 7.985301, 7.865797, 7.342469, 
    7.268659, 7.975486, 8.643974, 8.895267, 7.776951, 7.274741, 6.82941, 
    6.3626, 5.682857, 4.993686, 4.27755, 4.302801, 4.594637, 5.0822, 
    6.251255, 6.173875, 5.663871, 5.655987, 5.167533, 4.884112, 4.611746, 
    4.52724,
  3.98556, 4.55322, 5.439306, 6.037467, 6.976496, 7.428882, 7.372576, 
    7.192951, 6.921767, 6.892465, 7.191539, 6.200619, 5.687935, 5.42804, 
    5.192234, 4.607743, 3.990722, 3.857163, 3.714495, 4.053179, 4.193727, 
    4.243231, 4.336538, 4.579047, 4.820053, 4.89698, 4.396884, 4.305136, 
    3.971967,
  3.804318, 4.19997, 4.346646, 4.485344, 4.456432, 4.295829, 4.365797, 
    4.462391, 4.308909, 4.055781, 3.901777, 4.248356, 4.496099, 4.305739, 
    4.214332, 3.788826, 3.56288, 3.523534, 3.354793, 3.229579, 2.918486, 
    3.024291, 3.352449, 3.649258, 3.817241, 3.094713, 2.487627, 3.537621, 
    3.739271,
  2.80309, 2.868154, 3.021649, 3.070961, 3.035016, 3.114333, 3.242248, 
    3.227906, 3.223745, 3.244781, 3.322304, 3.440982, 3.462878, 3.340102, 
    3.213448, 3.076225, 2.96642, 2.802351, 2.744565, 2.688841, 2.675162, 
    2.632344, 2.414261, 2.470184, 2.561609, 2.170251, 2.238696, 2.623428, 
    2.805807,
  0.3573337, 0.3573337, 0.3573337, 0.3573337, 0.3573337, 0.3573337, 
    0.3573337, 0.3556668, 0.3556668, 0.3556668, 0.3556668, 0.3556668, 
    0.3556668, 0.3556668, 0.3765854, 0.3765854, 0.3765854, 0.3765854, 
    0.3765854, 0.3765854, 0.3765854, 0.3787483, 0.3787483, 0.3787483, 
    0.3787483, 0.3787483, 0.3787483, 0.3787483, 0.3573337,
  0.4966939, 0.4465986, 0.4357855, 0.4192985, 0.4241995, 0.4119187, 
    0.3838156, 0.3863123, 0.4080009, 0.4301301, 0.4391995, 0.4761153, 
    0.5307866, 0.6147001, 0.6817013, 0.7191311, 0.685828, 0.6672466, 
    0.6502914, 0.6318341, 0.6070783, 0.5946576, 0.6073497, 0.6025509, 
    0.584483, 0.5744196, 0.5799314, 0.5590674, 0.5221928,
  0.7479411, 0.7835767, 0.8045135, 0.7879732, 0.7875793, 0.7978412, 
    0.7261668, 0.6780594, 0.6447131, 0.6271645, 0.6649419, 0.7969289, 
    0.9951046, 1.262988, 1.396849, 1.38858, 1.401786, 1.306941, 1.064328, 
    0.908949, 0.8186511, 0.7285089, 0.7211126, 0.7872667, 0.8678579, 
    0.9074077, 1.011474, 0.893271, 0.7615919,
  1.169876, 0.9793001, 0.9051501, 0.9809896, 1.269539, 1.32041, 1.226954, 
    1.117363, 0.9210603, 0.8268226, 0.8410191, 1.197674, 1.789663, 2.086632, 
    2.295301, 2.351767, 2.255622, 2.019817, 1.795603, 1.495333, 1.194299, 
    1.018849, 0.8994786, 0.8710552, 1.115058, 1.193987, 1.33535, 1.321075, 
    1.232525,
  1.818099, 1.548232, 1.417926, 1.845296, 1.988779, 2.020202, 2.084154, 
    1.871261, 1.579873, 1.337659, 1.302416, 1.481068, 2.217654, 2.782648, 
    3.083961, 2.947424, 2.477314, 2.256196, 1.975357, 1.652725, 1.382992, 
    1.247497, 1.061148, 1.072792, 1.309454, 1.748937, 2.279864, 2.387301, 
    2.105837,
  2.928763, 2.807588, 3.146899, 3.540569, 3.698281, 3.599181, 3.044802, 
    2.838959, 2.599709, 2.499646, 2.389521, 2.743593, 3.082389, 3.707786, 
    3.698881, 3.168198, 2.716555, 2.255448, 2.027843, 1.598001, 1.323212, 
    1.143965, 1.048347, 1.164914, 2.518199, 3.314013, 3.191361, 3.090276, 
    3.210315,
  4.052326, 3.990871, 5.998713, 6.073409, 5.113338, 4.502188, 3.925563, 
    3.86121, 3.328056, 2.894797, 3.778588, 4.327656, 4.614592, 3.51504, 
    3.299289, 3.036062, 2.490311, 1.939376, 1.42567, 1.115831, 0.9481839, 
    0.8444828, 0.8340923, 0.8525819, 3.702116, 4.738176, 4.651279, 4.461081, 
    4.173814,
  4.856117, 6.544385, 9.875952, 7.170984, 5.950486, 4.445217, 3.728394, 
    2.840153, 2.673446, 3.016721, 4.63826, 4.087117, 3.707891, 3.359965, 
    2.577431, 1.887761, 1.330791, 1.093362, 0.9077008, 0.730046, 0.6316785, 
    0.7812184, 1.433621, 4.001374, 8.404162, 9.957454, 6.454655, 5.080522, 
    4.96924,
  6.803502, 11.54596, 15.16854, 7.655223, 4.9407, 3.439445, 2.502987, 
    2.254209, 2.640043, 2.994251, 3.023566, 2.99554, 2.096252, 1.16775, 
    0.7564597, 0.6013617, 0.6390882, 0.6295488, 0.5646639, 0.5541577, 
    0.5735253, 1.091198, 3.212409, 12.5389, 14.95101, 10.76776, 6.060796, 
    5.020254, 5.84602,
  9.156878, 16.86634, 13.75648, 6.429744, 4.939841, 3.404379, 2.77842, 
    2.589176, 5.467485, 7.921823, 2.820666, 1.71441, 0.8232948, 0.54184, 
    0.4502821, 0.4127717, 0.430758, 0.4903363, 0.5941761, 0.7163484, 
    0.8274844, 1.578841, 3.888193, 11.79472, 9.086185, 6.549367, 5.950558, 
    5.801906, 6.716882,
  12.46283, 12.94996, 11.25832, 8.418286, 5.170526, 4.175165, 4.459523, 
    3.925479, 4.864653, 3.70558, 2.676366, 1.765064, 1.194937, 1.003298, 
    0.8298463, 0.7978874, 0.7227326, 0.801281, 1.062826, 1.345798, 1.79927, 
    2.586556, 4.723338, 7.182444, 4.621014, 4.973638, 5.256808, 7.034984, 
    11.96995,
  5.177364, 5.662543, 5.183534, 4.23885, 5.446165, 5.481324, 6.741979, 
    7.290734, 8.587609, 5.91549, 4.645438, 3.342572, 2.780719, 3.053709, 
    2.814243, 2.715456, 2.227308, 2.139093, 1.80761, 1.826635, 2.505653, 
    3.900331, 2.900846, 2.641744, 2.272551, 2.463306, 2.876355, 3.572218, 
    4.229902,
  4.337062, 3.737019, 3.707244, 5.046673, 5.66501, 5.877451, 6.895313, 
    7.540392, 12.27483, 14.69695, 11.03805, 8.077131, 6.797976, 6.189944, 
    6.090915, 4.999241, 4.199789, 3.339666, 2.711379, 2.875732, 4.424964, 
    5.057068, 5.368913, 4.714163, 3.860003, 4.078603, 4.032753, 3.498918, 
    4.289751,
  5.365037, 5.592, 7.062568, 7.710495, 9.495026, 9.339396, 9.862405, 
    13.39428, 13.4796, 13.42531, 12.44807, 10.59621, 9.20472, 7.921189, 
    7.122692, 5.874124, 5.288649, 4.548816, 3.840523, 3.609383, 4.349987, 
    6.478112, 6.522534, 6.763171, 6.315531, 5.893634, 4.963551, 4.600412, 
    4.703093,
  5.004467, 6.310549, 7.25266, 8.142699, 8.342069, 8.284328, 7.854484, 
    7.986398, 8.881369, 9.42127, 9.524576, 8.494581, 7.744004, 7.168912, 
    6.765103, 5.987155, 5.263685, 4.440163, 4.440909, 4.848826, 5.437529, 
    6.600386, 6.565437, 6.301468, 6.197861, 5.459651, 5.180083, 4.734071, 
    4.615479,
  4.287146, 5.044636, 5.831223, 6.307312, 7.269538, 7.830215, 7.775174, 
    7.652949, 7.434062, 7.399539, 7.784902, 6.899799, 6.267261, 5.82459, 
    5.508509, 4.984733, 4.371324, 4.165915, 4.103254, 4.370166, 4.52359, 
    4.593207, 4.816099, 5.076902, 5.202541, 5.237221, 4.715032, 4.604174, 
    4.286886,
  4.153604, 4.588571, 4.849789, 4.915098, 4.860763, 4.727742, 4.794865, 
    4.957104, 4.92976, 4.717266, 4.654062, 4.924364, 5.0368, 4.796237, 
    4.64889, 4.198212, 3.921258, 3.854892, 3.646775, 3.522208, 3.253438, 
    3.418221, 3.823421, 4.130424, 4.192187, 3.582489, 3.009163, 3.873641, 
    4.033209,
  3.305804, 3.405578, 3.522728, 3.618836, 3.581192, 3.691701, 3.84938, 
    3.82249, 3.817555, 3.832755, 3.949963, 4.001007, 3.984398, 3.79981, 
    3.616568, 3.441191, 3.332619, 3.184796, 3.146609, 3.133665, 3.113272, 
    3.032887, 2.840009, 2.924325, 3.050075, 2.670644, 2.733836, 3.112308, 
    3.297194,
  0.3869947, 0.3869947, 0.3869947, 0.3869947, 0.3869947, 0.3869947, 
    0.3869947, 0.3861099, 0.3861099, 0.3861099, 0.3861099, 0.3861099, 
    0.3861099, 0.3861099, 0.4111116, 0.4111116, 0.4111116, 0.4111116, 
    0.4111116, 0.4111116, 0.4111116, 0.4098827, 0.4098827, 0.4098827, 
    0.4098827, 0.4098827, 0.4098827, 0.4098827, 0.3869947,
  0.5298803, 0.4908582, 0.4824181, 0.4653676, 0.4677014, 0.4528335, 
    0.4217181, 0.4193134, 0.4409229, 0.4617556, 0.4714307, 0.5016017, 
    0.5544473, 0.5912176, 0.6375644, 0.6753682, 0.6463356, 0.6466264, 
    0.6424264, 0.6340764, 0.6206135, 0.6096416, 0.6150358, 0.5818717, 
    0.5722456, 0.5762467, 0.5778863, 0.575899, 0.5565966,
  0.7682658, 0.8146847, 0.8161669, 0.7874765, 0.824182, 0.8115762, 0.7037604, 
    0.6950471, 0.6634052, 0.6415672, 0.6913599, 0.8183981, 0.9459172, 
    1.179748, 1.318041, 1.328203, 1.356968, 1.248023, 1.009683, 0.8762906, 
    0.7817258, 0.7141703, 0.6999786, 0.7738594, 0.8581585, 0.8989006, 
    0.9864667, 0.8840486, 0.7664448,
  1.237415, 1.029386, 0.95744, 1.017064, 1.270307, 1.280857, 1.179031, 
    1.073352, 0.8827737, 0.7887963, 0.787199, 1.116861, 1.724457, 2.01176, 
    2.153632, 2.250335, 2.163659, 1.958963, 1.713566, 1.455543, 1.159659, 
    0.9958478, 0.8745121, 0.8458973, 1.144531, 1.232874, 1.414838, 1.338003, 
    1.262708,
  1.758067, 1.51905, 1.409137, 1.760944, 1.874087, 1.898305, 1.948707, 
    1.760033, 1.506743, 1.288156, 1.240126, 1.435891, 2.194835, 2.748342, 
    2.978096, 2.834891, 2.381193, 2.224735, 1.953959, 1.637099, 1.367662, 
    1.24447, 1.057406, 1.073133, 1.325513, 1.736888, 2.181589, 2.294904, 
    2.01693,
  2.686187, 2.594962, 2.928937, 3.330089, 3.423534, 3.32258, 2.786524, 
    2.615919, 2.442151, 2.333045, 2.24732, 2.623107, 3.023158, 3.632329, 
    3.655555, 3.099509, 2.695899, 2.27843, 2.037899, 1.585482, 1.331547, 
    1.135172, 1.043901, 1.160522, 2.556102, 3.228199, 2.972814, 2.83776, 
    2.852815,
  3.756247, 3.680622, 5.870982, 5.721836, 4.766205, 4.175004, 3.652046, 
    3.619567, 3.193089, 2.866503, 3.845312, 4.302583, 4.596668, 3.455065, 
    3.229337, 3.064225, 2.530757, 2.007245, 1.453882, 1.133422, 0.9390707, 
    0.8258932, 0.7900772, 0.7868236, 3.663954, 4.533243, 4.243052, 4.050946, 
    3.771077,
  4.486189, 5.888312, 9.449544, 6.708745, 5.507944, 4.04037, 3.571831, 
    2.697358, 2.632085, 2.965649, 4.607267, 4.1226, 3.650454, 3.332875, 
    2.578905, 1.916052, 1.345147, 1.086637, 0.8973498, 0.6933653, 0.5875197, 
    0.7134641, 1.325686, 3.673361, 7.581203, 9.454205, 5.849279, 4.518951, 
    4.58415,
  6.206816, 10.42351, 13.42107, 6.666501, 4.477684, 3.286622, 2.399739, 
    2.174821, 2.417953, 2.841516, 2.858135, 2.894328, 2.006349, 1.154753, 
    0.7574437, 0.6015152, 0.6346709, 0.6060986, 0.5566756, 0.5122759, 
    0.5345792, 1.016376, 2.756848, 11.09385, 13.48511, 9.701226, 5.398929, 
    4.592051, 5.249519,
  8.639805, 15.1499, 12.15027, 5.901193, 4.371635, 3.221744, 2.695246, 
    2.575712, 4.918881, 7.371655, 2.701485, 1.752275, 0.8403745, 0.5351837, 
    0.4485206, 0.4229886, 0.4194395, 0.4745101, 0.583541, 0.6226185, 
    0.7535422, 1.364486, 3.233515, 9.62023, 7.810512, 5.88513, 5.506221, 
    5.3087, 6.127137,
  11.90191, 12.21576, 10.5165, 7.894486, 4.749619, 3.859342, 4.452585, 
    3.843468, 4.769235, 3.609087, 2.556039, 1.778349, 1.262493, 1.079204, 
    0.8704317, 0.8227703, 0.7322033, 0.8095463, 1.072487, 1.28951, 1.716879, 
    2.405239, 4.162897, 5.976659, 3.556567, 3.792105, 4.389462, 6.278717, 
    11.34247,
  4.771717, 5.218265, 4.573177, 3.955907, 5.119189, 5.230917, 6.519526, 
    6.953476, 8.294789, 5.697195, 4.428502, 3.212939, 2.725125, 3.086008, 
    2.876768, 2.840403, 2.255703, 2.157211, 1.808406, 1.85248, 2.420407, 
    3.744048, 2.722566, 2.491094, 2.153713, 2.367397, 2.808394, 3.420478, 
    3.966695,
  4.315838, 3.856175, 3.883156, 5.11483, 5.796987, 5.974132, 7.296989, 
    8.021047, 13.2106, 15.6597, 11.57093, 8.200194, 6.810119, 6.263166, 
    6.143094, 4.993193, 4.155776, 3.250299, 2.706781, 2.882009, 4.452586, 
    4.97849, 5.21539, 4.575049, 3.674065, 3.939368, 4.021144, 3.468545, 
    4.416263,
  5.483541, 5.724778, 7.152261, 8.083926, 9.660718, 9.742321, 11.03411, 
    14.3269, 14.1905, 14.17335, 12.90532, 11.11127, 9.537696, 8.091498, 
    7.258263, 6.087171, 5.422754, 4.556314, 3.883261, 3.667985, 4.530966, 
    6.467101, 6.508395, 6.784287, 6.404195, 5.923799, 4.981075, 4.655776, 
    4.671028,
  5.079101, 6.526263, 7.376982, 8.288281, 8.577842, 8.564452, 8.204212, 
    8.545364, 9.576447, 10.06996, 9.973728, 9.104105, 8.061205, 7.388882, 
    6.996598, 6.173189, 5.414089, 4.492687, 4.465283, 5.031491, 5.617768, 
    6.794438, 6.768955, 6.726278, 6.593637, 5.688128, 5.365894, 4.800898, 
    4.632135,
  4.462418, 5.414168, 6.155716, 6.535315, 7.451972, 8.047132, 8.091137, 
    7.956834, 7.777227, 7.807625, 8.285458, 7.55951, 6.727246, 6.160452, 
    5.744408, 5.230662, 4.68093, 4.395526, 4.356795, 4.615839, 4.842644, 
    4.883539, 5.13351, 5.486991, 5.585831, 5.470335, 4.951872, 4.807225, 
    4.47371,
  4.354774, 4.825869, 5.23085, 5.277304, 5.181819, 5.170692, 5.163972, 
    5.406967, 5.477799, 5.271403, 5.388093, 5.532262, 5.496423, 5.22952, 
    4.983691, 4.492716, 4.246394, 4.136923, 3.879686, 3.73116, 3.547204, 
    3.709803, 4.225697, 4.473199, 4.514786, 3.974554, 3.460964, 4.103034, 
    4.219481,
  3.682318, 3.81264, 3.938066, 4.052794, 4.051117, 4.117302, 4.287611, 
    4.26434, 4.24892, 4.305099, 4.407976, 4.45115, 4.398614, 4.190026, 
    3.969725, 3.76012, 3.639538, 3.47401, 3.4538, 3.490579, 3.464564, 
    3.333645, 3.186054, 3.314633, 3.491102, 3.135189, 3.170302, 3.520767, 
    3.675109,
  0.4063181, 0.4063181, 0.4063181, 0.4063181, 0.4063181, 0.4063181, 
    0.4063181, 0.4040863, 0.4040863, 0.4040863, 0.4040863, 0.4040863, 
    0.4040863, 0.4040863, 0.4330112, 0.4330112, 0.4330112, 0.4330112, 
    0.4330112, 0.4330112, 0.4330112, 0.4288161, 0.4288161, 0.4288161, 
    0.4288161, 0.4288161, 0.4288161, 0.4288161, 0.4063181,
  0.5524696, 0.516091, 0.5118719, 0.4953892, 0.4918867, 0.4720733, 0.4423701, 
    0.4372175, 0.4552123, 0.467464, 0.4842609, 0.5132982, 0.5583866, 
    0.5478745, 0.5723098, 0.6088678, 0.5911608, 0.6044787, 0.6130842, 
    0.6163658, 0.6119344, 0.6037437, 0.6063064, 0.552394, 0.5498299, 
    0.5607187, 0.5480241, 0.5712622, 0.5794358,
  0.7661672, 0.8164724, 0.8022296, 0.7687166, 0.828186, 0.8016014, 0.6676368, 
    0.6868777, 0.6539001, 0.6284357, 0.6816244, 0.7968997, 0.8892964, 
    1.081494, 1.22083, 1.249335, 1.273616, 1.171976, 0.9394592, 0.8181344, 
    0.7279369, 0.6775626, 0.6688615, 0.7456438, 0.8398799, 0.8727035, 
    0.936149, 0.8655689, 0.7639921,
  1.238918, 1.049627, 0.991456, 1.030395, 1.24812, 1.223404, 1.103085, 
    0.9966347, 0.8247172, 0.7274491, 0.7157559, 1.034997, 1.619938, 1.855293, 
    1.991028, 2.121408, 2.038362, 1.864869, 1.609475, 1.382445, 1.090269, 
    0.9441381, 0.8269373, 0.8001188, 1.160366, 1.251414, 1.466529, 1.343798, 
    1.271382,
  1.694623, 1.498016, 1.393188, 1.68583, 1.76202, 1.787514, 1.803523, 
    1.617931, 1.401588, 1.202363, 1.160517, 1.386469, 2.107254, 2.662128, 
    2.847751, 2.685365, 2.25217, 2.137208, 1.893412, 1.596708, 1.319596, 
    1.2158, 1.0444, 1.068898, 1.355935, 1.722067, 2.091944, 2.180856, 1.925887,
  2.413938, 2.353007, 2.708023, 3.152912, 3.155982, 3.007453, 2.545084, 
    2.39564, 2.261774, 2.127362, 2.072153, 2.491061, 2.966723, 3.480811, 
    3.545509, 2.976553, 2.609488, 2.259633, 1.98259, 1.569358, 1.329953, 
    1.116678, 1.031685, 1.124801, 2.664644, 3.149871, 2.707997, 2.605538, 
    2.502271,
  3.456517, 3.406567, 5.649008, 5.393715, 4.396222, 3.796417, 3.360025, 
    3.339635, 3.024961, 2.829676, 3.916727, 4.229856, 4.4614, 3.324037, 
    3.081544, 3.022609, 2.535949, 2.049407, 1.477084, 1.149989, 0.9277107, 
    0.8220723, 0.7452133, 0.7720719, 3.871741, 4.482104, 3.933373, 3.655013, 
    3.403889,
  4.096213, 5.46403, 9.024598, 6.180953, 5.072929, 3.635224, 3.33302, 
    2.539063, 2.59058, 2.870574, 4.686362, 4.177386, 3.649209, 3.254015, 
    2.511967, 1.942152, 1.361836, 1.081696, 0.8710083, 0.6426176, 0.5525271, 
    0.655349, 1.241569, 3.62393, 7.159085, 8.873251, 5.297437, 4.064016, 
    4.14676,
  5.720152, 9.753551, 11.83149, 5.785546, 3.938973, 3.018088, 2.209941, 
    2.068081, 2.328314, 2.787741, 2.778755, 2.905431, 2.014496, 1.146907, 
    0.7377005, 0.5972059, 0.6283028, 0.5930281, 0.5453409, 0.4766205, 
    0.4833081, 0.9821277, 2.633884, 10.17442, 12.21254, 8.925158, 4.679235, 
    3.989501, 4.55701,
  8.501921, 14.44274, 11.34628, 5.283751, 3.762039, 2.897996, 2.545104, 
    2.512191, 4.670762, 7.202798, 2.737453, 1.789891, 0.8638417, 0.5132426, 
    0.4337663, 0.42867, 0.4188074, 0.4789074, 0.5366921, 0.5739125, 
    0.6891719, 1.268999, 2.91082, 8.383323, 6.967878, 5.223785, 4.900808, 
    4.889149, 5.743676,
  11.80409, 11.70704, 9.97698, 7.359332, 4.423971, 3.627415, 4.340983, 
    3.794458, 4.669354, 3.520859, 2.426004, 1.813765, 1.317272, 1.133461, 
    0.9111944, 0.8460882, 0.7503468, 0.8589858, 1.086404, 1.252889, 1.624292, 
    2.268563, 3.716672, 5.152362, 2.784009, 3.034022, 3.763962, 5.819803, 
    11.01693,
  4.590545, 4.735527, 4.030645, 3.874843, 4.941304, 5.103782, 6.365418, 
    6.646311, 8.097039, 5.496777, 4.24774, 3.115155, 2.597831, 3.04992, 
    2.916536, 2.901668, 2.236368, 2.116992, 1.790118, 1.918148, 2.380051, 
    3.670782, 2.567922, 2.320536, 2.050668, 2.247459, 2.797374, 3.410963, 
    3.959697,
  4.318511, 4.023155, 4.130367, 5.134792, 5.889093, 6.086896, 7.785466, 
    8.440567, 14.12498, 16.74212, 12.19511, 8.398262, 6.866493, 6.346439, 
    6.133502, 4.992715, 4.1049, 3.172148, 2.716354, 2.918039, 4.442252, 
    4.888945, 5.080661, 4.432007, 3.438271, 3.775716, 3.93092, 3.426186, 
    4.484098,
  5.566497, 5.819813, 7.170215, 8.260795, 9.887776, 9.906002, 12.12307, 
    15.01411, 14.68762, 14.54252, 13.13158, 11.27365, 9.753181, 8.223851, 
    7.324569, 6.140965, 5.438665, 4.533123, 3.847369, 3.674269, 4.751924, 
    6.566624, 6.56952, 6.862216, 6.509682, 5.918052, 4.973302, 4.61712, 
    4.613155,
  5.077196, 6.73621, 7.375668, 8.18505, 8.780475, 8.745148, 8.397516, 
    8.934763, 10.03448, 10.58964, 10.42795, 9.505828, 8.327016, 7.486432, 
    7.093688, 6.253238, 5.464373, 4.512815, 4.416532, 5.095654, 5.724261, 
    6.958296, 6.94119, 7.115185, 6.984364, 5.865982, 5.493218, 4.814849, 
    4.593289,
  4.54708, 5.651777, 6.360433, 6.713666, 7.594659, 8.12616, 8.227796, 
    8.23875, 8.066879, 8.083734, 8.661042, 8.159006, 7.122173, 6.415854, 
    5.886059, 5.359709, 4.880732, 4.547071, 4.521997, 4.790252, 5.139929, 
    5.095964, 5.406665, 5.913767, 5.992633, 5.669036, 5.105142, 4.912621, 
    4.551921,
  4.482094, 5.010765, 5.493181, 5.632749, 5.542455, 5.584506, 5.511464, 
    5.805049, 5.904006, 5.702992, 6.007554, 6.013688, 5.874261, 5.539203, 
    5.176702, 4.68289, 4.487626, 4.338, 4.017893, 3.878643, 3.76283, 
    3.934382, 4.533186, 4.747231, 4.849538, 4.294651, 3.849456, 4.281031, 
    4.336045,
  3.97246, 4.11107, 4.259092, 4.412035, 4.434087, 4.453714, 4.603029, 4.6229, 
    4.60968, 4.714213, 4.817772, 4.836647, 4.757578, 4.524086, 4.271511, 
    4.044106, 3.913383, 3.702066, 3.694321, 3.76583, 3.725792, 3.615386, 
    3.495905, 3.662619, 3.882273, 3.552845, 3.559628, 3.8769, 3.992469,
  0.4189714, 0.4189714, 0.4189714, 0.4189714, 0.4189714, 0.4189714, 
    0.4189714, 0.414577, 0.414577, 0.414577, 0.414577, 0.414577, 0.414577, 
    0.414577, 0.4439672, 0.4439672, 0.4439672, 0.4439672, 0.4439672, 
    0.4439672, 0.4439672, 0.4375601, 0.4375601, 0.4375601, 0.4375601, 
    0.4375601, 0.4375601, 0.4375601, 0.4189714,
  0.5645616, 0.5260128, 0.5243974, 0.5082309, 0.4973058, 0.4723863, 0.447087, 
    0.4417417, 0.4542978, 0.4610513, 0.481159, 0.5125373, 0.5491251, 
    0.4942518, 0.4986415, 0.5324157, 0.5300849, 0.553212, 0.572929, 
    0.5856354, 0.5893241, 0.5850277, 0.5898454, 0.5283872, 0.5255132, 
    0.5338787, 0.5116067, 0.5517764, 0.5865842,
  0.7380154, 0.7861576, 0.7549483, 0.7341855, 0.8049628, 0.7697922, 
    0.6230972, 0.6649268, 0.628378, 0.6015803, 0.6534766, 0.7571615, 
    0.832913, 0.9766308, 1.113954, 1.161709, 1.162315, 1.083507, 0.8574058, 
    0.7505478, 0.6751445, 0.6422474, 0.6343662, 0.7171928, 0.8152735, 
    0.828687, 0.8964415, 0.8393486, 0.7555624,
  1.221521, 1.054209, 1.010157, 1.034018, 1.209514, 1.164486, 1.014281, 
    0.9042752, 0.7566153, 0.6563653, 0.6447473, 0.9516696, 1.512771, 
    1.684693, 1.837588, 1.968649, 1.885063, 1.742288, 1.492059, 1.284944, 
    1.001212, 0.8698477, 0.7662802, 0.7497495, 1.151477, 1.251433, 1.473988, 
    1.338635, 1.269263,
  1.649117, 1.489553, 1.384134, 1.615018, 1.657857, 1.670336, 1.654742, 
    1.470696, 1.283813, 1.100869, 1.069865, 1.326012, 2.014877, 2.565664, 
    2.673553, 2.531023, 2.120284, 2.012413, 1.799237, 1.517755, 1.26018, 
    1.174982, 1.011646, 1.047067, 1.380884, 1.738431, 2.011643, 2.080518, 
    1.849258,
  2.169664, 2.100346, 2.468229, 3.014914, 2.964663, 2.705606, 2.339561, 
    2.179971, 2.05003, 1.924952, 1.936936, 2.376239, 2.935885, 3.344393, 
    3.403379, 2.824575, 2.472211, 2.194083, 1.886362, 1.551056, 1.316581, 
    1.09008, 1.018114, 1.075243, 2.83568, 3.110444, 2.492966, 2.380564, 
    2.219688,
  3.109211, 3.160636, 5.483951, 5.290086, 4.021005, 3.453861, 3.0686, 
    3.080411, 2.835106, 2.800454, 3.958155, 4.232453, 4.371654, 3.18367, 
    2.910623, 2.930822, 2.510939, 2.032288, 1.480249, 1.158819, 0.9260142, 
    0.8051961, 0.7172971, 0.7970785, 4.473354, 4.586646, 3.722708, 3.283839, 
    3.078386,
  3.684158, 5.198661, 8.53481, 5.677136, 4.649188, 3.333247, 3.054308, 
    2.413353, 2.468755, 2.791112, 4.850606, 4.25465, 3.626009, 3.134149, 
    2.40412, 1.950008, 1.375801, 1.074417, 0.850394, 0.5954027, 0.5279132, 
    0.6013285, 1.198652, 3.699059, 7.282222, 8.271256, 4.77885, 3.710834, 
    3.717316,
  5.312043, 9.475636, 10.82062, 5.11491, 3.320616, 2.643835, 2.007238, 
    1.923968, 2.288188, 2.728958, 2.760875, 2.950648, 2.065229, 1.146996, 
    0.7162102, 0.5812763, 0.60359, 0.6002639, 0.5145606, 0.4512104, 
    0.4481377, 0.9640786, 2.714129, 10.20134, 11.37393, 8.386744, 3.950933, 
    3.377161, 3.99606,
  8.527891, 14.99853, 11.66886, 4.699756, 3.10208, 2.564714, 2.366687, 
    2.447421, 4.570858, 7.179401, 2.84375, 1.881077, 0.9060504, 0.4957482, 
    0.4119708, 0.4282327, 0.4250457, 0.4774615, 0.4911481, 0.5239237, 
    0.6709889, 1.300578, 2.962172, 8.407125, 6.642097, 4.860209, 4.394851, 
    4.498269, 5.582204,
  11.75752, 11.24902, 9.78978, 7.064486, 4.060159, 3.475826, 4.247898, 
    3.833164, 4.554053, 3.404072, 2.34178, 1.808406, 1.332976, 1.166193, 
    0.9214911, 0.8562815, 0.7686721, 0.914707, 1.08744, 1.238012, 1.594324, 
    2.170597, 3.481795, 4.790011, 2.346492, 2.620655, 3.555267, 5.619354, 
    11.20199,
  4.717316, 4.38677, 3.634278, 4.512675, 4.875973, 5.017183, 6.183745, 
    6.558915, 8.073638, 5.35818, 4.105919, 3.034636, 2.50035, 2.997408, 
    2.990018, 2.858171, 2.175008, 2.072541, 1.729105, 1.994588, 2.468733, 
    3.710301, 2.41853, 2.206231, 1.955973, 2.128954, 2.850697, 3.565183, 
    3.943911,
  4.398194, 4.261843, 4.466027, 5.226916, 6.060942, 6.305599, 8.553997, 
    8.97215, 15.14095, 18.0791, 12.97165, 8.760055, 7.032343, 6.415177, 
    6.200095, 5.049675, 4.040676, 3.07304, 2.694942, 2.981169, 4.486248, 
    4.899037, 5.026689, 4.319716, 3.218386, 3.597265, 3.805244, 3.382799, 
    4.702067,
  5.648211, 5.956864, 7.228202, 8.34698, 10.54998, 9.90854, 13.09242, 
    15.60901, 15.03603, 14.74528, 13.14677, 11.28483, 9.858543, 8.306419, 
    7.318143, 6.158341, 5.376708, 4.492085, 3.771413, 3.663769, 5.038512, 
    6.979496, 6.733927, 7.059786, 6.597561, 5.916109, 4.958306, 4.533891, 
    4.555377,
  5.090158, 6.905801, 7.328772, 8.020853, 9.001419, 8.855893, 8.546726, 
    9.239623, 10.33795, 11.06772, 10.95222, 9.980587, 8.609932, 7.571168, 
    7.118881, 6.26592, 5.419189, 4.498924, 4.35695, 5.068099, 5.815678, 
    7.18252, 7.22538, 7.591391, 7.481158, 5.983212, 5.569838, 4.81092, 
    4.556739,
  4.626311, 5.818754, 6.487061, 6.911988, 7.708619, 8.172148, 8.326512, 
    8.550749, 8.421659, 8.283244, 8.943885, 8.631275, 7.513484, 6.62217, 
    6.018332, 5.44996, 5.014791, 4.61739, 4.603454, 4.967507, 5.421058, 
    5.273451, 5.627664, 6.391903, 6.372619, 5.884762, 5.266056, 4.961861, 
    4.597216,
  4.611732, 5.172875, 5.65324, 5.998533, 5.875644, 5.942114, 5.889435, 
    6.165349, 6.193293, 6.02073, 6.53455, 6.466816, 6.215995, 5.73764, 
    5.324524, 4.799613, 4.672955, 4.492386, 4.140398, 3.995318, 3.96208, 
    4.220781, 4.746592, 5.023157, 5.190392, 4.55424, 4.164184, 4.46261, 
    4.464085,
  4.237833, 4.331197, 4.500961, 4.667979, 4.740453, 4.781846, 4.900989, 
    4.963908, 4.972466, 5.043707, 5.165343, 5.20401, 5.065022, 4.784535, 
    4.519473, 4.254891, 4.116239, 3.898517, 3.877839, 3.994943, 3.951903, 
    3.887653, 3.803921, 3.997542, 4.233637, 3.919108, 3.900451, 4.200957, 
    4.279215,
  0.425905, 0.425905, 0.425905, 0.425905, 0.425905, 0.425905, 0.425905, 
    0.4204995, 0.4204995, 0.4204995, 0.4204995, 0.4204995, 0.4204995, 
    0.4204995, 0.4467578, 0.4467578, 0.4467578, 0.4467578, 0.4467578, 
    0.4467578, 0.4467578, 0.4412242, 0.4412242, 0.4412242, 0.4412242, 
    0.4412242, 0.4412242, 0.4412242, 0.425905,
  0.564113, 0.530057, 0.5207566, 0.5050433, 0.4895195, 0.4624095, 0.4390124, 
    0.4338467, 0.4457589, 0.4530063, 0.4715842, 0.5044572, 0.5301836, 
    0.435087, 0.4315464, 0.4568202, 0.4685179, 0.500075, 0.5332416, 
    0.5527042, 0.5622931, 0.5597524, 0.5697527, 0.5089925, 0.5074323, 
    0.5053075, 0.4769928, 0.5235497, 0.5824617,
  0.6968728, 0.7372223, 0.6887696, 0.6863735, 0.7678621, 0.7272348, 
    0.5729074, 0.6315904, 0.5913292, 0.5612689, 0.6182272, 0.716569, 
    0.7741952, 0.878575, 1.00176, 1.079951, 1.056295, 0.9830385, 0.7725695, 
    0.6740468, 0.6218671, 0.6032844, 0.589219, 0.6846068, 0.7768254, 
    0.7757388, 0.8536984, 0.7979854, 0.7333153,
  1.198323, 1.051487, 1.006807, 1.032399, 1.156888, 1.098877, 0.9304851, 
    0.8156568, 0.685551, 0.5931445, 0.583994, 0.8714206, 1.409759, 1.557649, 
    1.69743, 1.810812, 1.731518, 1.618789, 1.365942, 1.18069, 0.9021493, 
    0.7892787, 0.7074906, 0.6959172, 1.114139, 1.248065, 1.470227, 1.326603, 
    1.257337,
  1.602401, 1.477784, 1.361436, 1.558523, 1.572717, 1.547301, 1.51284, 
    1.351424, 1.176175, 1.007224, 0.9811634, 1.257425, 1.954159, 2.453782, 
    2.507766, 2.359463, 1.993098, 1.881529, 1.690372, 1.425732, 1.199255, 
    1.115584, 0.9514676, 1.01924, 1.423604, 1.825426, 1.968176, 2.000143, 
    1.776928,
  1.957772, 1.85043, 2.19986, 2.940006, 2.860483, 2.503988, 2.177927, 
    1.973268, 1.842325, 1.739801, 1.838894, 2.320849, 2.932701, 3.251102, 
    3.213044, 2.652465, 2.317207, 2.098555, 1.781582, 1.491808, 1.297563, 
    1.063904, 0.9981801, 1.048983, 3.095766, 3.104795, 2.38999, 2.169295, 
    2.023532,
  2.760639, 2.949222, 5.503967, 5.312818, 3.69347, 3.155059, 2.787307, 
    2.816704, 2.624278, 2.728609, 4.10479, 4.435109, 4.416655, 3.100906, 
    2.785531, 2.812015, 2.449831, 1.969434, 1.464041, 1.156446, 0.9094204, 
    0.7810311, 0.7164965, 0.8453742, 5.445313, 4.787642, 3.590131, 2.949051, 
    2.762701,
  3.328213, 5.212458, 8.190663, 5.357174, 4.314324, 3.036119, 2.777689, 
    2.30536, 2.387911, 2.846202, 5.213918, 4.43908, 3.53791, 2.965867, 
    2.28923, 1.907862, 1.396311, 1.06445, 0.8331872, 0.5494332, 0.5046294, 
    0.5600894, 1.134206, 3.879444, 7.96808, 8.033537, 4.327168, 3.413702, 
    3.316184,
  4.976802, 9.774418, 10.11805, 4.96143, 2.793584, 2.281511, 1.842749, 
    1.790372, 2.264145, 2.678396, 2.725084, 2.984105, 2.114902, 1.159418, 
    0.7004098, 0.5380459, 0.5638273, 0.5794426, 0.4692259, 0.416178, 
    0.4463568, 1.003797, 3.185881, 10.83391, 10.91998, 8.019435, 3.286693, 
    2.973057, 3.652158,
  8.917571, 16.35399, 13.31098, 4.35854, 2.527346, 2.243621, 2.217202, 
    2.376215, 4.528516, 7.226473, 2.952044, 1.995818, 0.9656045, 0.4763672, 
    0.3919517, 0.4089408, 0.4239146, 0.4488552, 0.477747, 0.5034344, 
    0.7132643, 1.402056, 3.603505, 9.319353, 6.976336, 4.655815, 4.000398, 
    4.360735, 5.652401,
  11.83887, 10.96019, 9.981089, 7.254521, 3.937701, 3.337748, 4.321471, 
    3.956298, 4.497078, 3.290153, 2.307412, 1.781537, 1.321729, 1.153187, 
    0.8978322, 0.8533965, 0.7838681, 0.9637737, 1.094309, 1.255885, 1.611446, 
    2.144249, 3.439447, 4.656389, 2.135916, 2.512383, 3.519044, 5.796574, 
    11.52212,
  5.140694, 4.42563, 3.769322, 6.388581, 5.251503, 5.055125, 6.066626, 
    6.764594, 8.118363, 5.334785, 3.955445, 2.945068, 2.469239, 2.920655, 
    3.019509, 2.782628, 2.116132, 2.010154, 1.692511, 2.090916, 2.692352, 
    3.896195, 2.320188, 2.111695, 1.869761, 2.093259, 2.937865, 3.839659, 
    4.109233,
  4.701634, 4.644013, 4.800799, 5.490771, 6.504069, 6.811087, 9.737899, 
    9.59928, 16.28182, 19.50857, 13.6448, 9.381577, 7.383317, 6.540801, 
    6.233361, 5.161321, 3.968796, 3.003493, 2.690041, 3.106493, 4.716054, 
    5.147799, 5.122666, 4.299078, 3.04197, 3.357384, 3.745087, 3.466544, 
    5.201064,
  5.756841, 6.189521, 7.390791, 8.448756, 11.67509, 10.05101, 13.97928, 
    16.27182, 15.4587, 14.8564, 13.11095, 11.16926, 9.943859, 8.337862, 
    7.243612, 6.127251, 5.277791, 4.393085, 3.672121, 3.651997, 5.523285, 
    7.728263, 7.075026, 7.359825, 6.727585, 5.964988, 4.936149, 4.42577, 
    4.504972,
  5.197781, 7.1201, 7.317105, 7.970186, 9.272752, 9.051613, 8.68698, 
    9.449202, 10.65856, 11.52797, 11.49865, 10.48792, 8.963649, 7.718555, 
    7.09719, 6.253563, 5.341897, 4.474742, 4.293031, 5.038638, 6.029236, 
    7.567317, 7.589986, 8.204593, 8.090577, 6.114257, 5.648145, 4.79637, 
    4.521056,
  4.789189, 5.896593, 6.6146, 7.075071, 7.795819, 8.326873, 8.462237, 
    8.822946, 8.818628, 8.501199, 9.298094, 9.054947, 7.91118, 6.841478, 
    6.136436, 5.539635, 5.091698, 4.667686, 4.67193, 5.175913, 5.719337, 
    5.522986, 5.851164, 6.900108, 6.853678, 6.136084, 5.379181, 4.98087, 
    4.629347,
  4.792985, 5.364197, 5.767018, 6.319202, 6.213699, 6.32759, 6.356545, 
    6.511981, 6.449015, 6.370043, 7.028474, 6.872108, 6.422733, 5.860026, 
    5.439732, 4.86702, 4.884414, 4.611999, 4.263527, 4.129794, 4.194018, 
    4.51295, 5.005539, 5.335119, 5.481787, 4.776377, 4.425834, 4.637132, 
    4.569559,
  4.490253, 4.53273, 4.688076, 4.852588, 4.991216, 5.111407, 5.176473, 
    5.27133, 5.316943, 5.343281, 5.423104, 5.456057, 5.27659, 4.979962, 
    4.699605, 4.396465, 4.245219, 4.081581, 4.054819, 4.170108, 4.148232, 
    4.140636, 4.120323, 4.349818, 4.594123, 4.234713, 4.190642, 4.513084, 
    4.553108,
  0.4269015, 0.4269015, 0.4269015, 0.4269015, 0.4269015, 0.4269015, 
    0.4269015, 0.4208236, 0.4208236, 0.4208236, 0.4208236, 0.4208236, 
    0.4208236, 0.4208236, 0.443893, 0.443893, 0.443893, 0.443893, 0.443893, 
    0.443893, 0.443893, 0.442735, 0.442735, 0.442735, 0.442735, 0.442735, 
    0.442735, 0.442735, 0.4269015,
  0.5555304, 0.5293595, 0.5098624, 0.4888435, 0.4760394, 0.4501513, 
    0.4260468, 0.4235296, 0.4387484, 0.4457198, 0.4648426, 0.4933297, 
    0.5055276, 0.3778798, 0.3764961, 0.3948286, 0.4108503, 0.4501859, 
    0.4951703, 0.518007, 0.5344962, 0.532171, 0.5439293, 0.4900929, 
    0.4900643, 0.4757888, 0.446551, 0.4948997, 0.5673892,
  0.6589624, 0.67634, 0.6229459, 0.6310374, 0.7299908, 0.6806448, 0.520874, 
    0.5895184, 0.5464784, 0.5136406, 0.5736611, 0.674392, 0.7070565, 
    0.7866451, 0.8920172, 0.9870722, 0.9588225, 0.879346, 0.6928622, 
    0.6010391, 0.5662948, 0.5596555, 0.5403095, 0.6499117, 0.7317795, 
    0.73264, 0.7942693, 0.7610003, 0.7045888,
  1.169679, 1.037623, 0.9947408, 1.018576, 1.09592, 1.033252, 0.8606576, 
    0.7451351, 0.6222381, 0.5381275, 0.5306345, 0.7947119, 1.329575, 
    1.454076, 1.578301, 1.658399, 1.579413, 1.473892, 1.232782, 1.059401, 
    0.8080426, 0.7094167, 0.6519777, 0.642719, 1.070729, 1.258382, 1.47163, 
    1.32456, 1.236239,
  1.566159, 1.45286, 1.337795, 1.498722, 1.520665, 1.454413, 1.388476, 
    1.2443, 1.068367, 0.9230072, 0.9030143, 1.188345, 1.918871, 2.350124, 
    2.354999, 2.167145, 1.848119, 1.754098, 1.575292, 1.326094, 1.136871, 
    1.043, 0.8880897, 0.9924706, 1.488462, 1.942583, 1.971484, 1.936923, 
    1.746385,
  1.81192, 1.665563, 1.975539, 2.92328, 2.832319, 2.370101, 2.007054, 
    1.782846, 1.650231, 1.560129, 1.777212, 2.329927, 3.052078, 3.204997, 
    3.015132, 2.460882, 2.15129, 1.985708, 1.692412, 1.416167, 1.243226, 
    1.02675, 0.9671146, 1.021677, 3.57546, 3.211066, 2.36849, 2.046668, 
    1.895583,
  2.465483, 2.807289, 5.786424, 5.545609, 3.4479, 2.908359, 2.557348, 
    2.537732, 2.428154, 2.609013, 4.542434, 4.906236, 4.676952, 3.171898, 
    2.721242, 2.681448, 2.347071, 1.878068, 1.414547, 1.140674, 0.8741688, 
    0.7571033, 0.7196311, 0.9359157, 6.690842, 5.088043, 3.508191, 2.72937, 
    2.503336,
  3.060947, 5.826855, 8.091804, 5.248998, 4.101255, 2.755693, 2.56073, 
    2.195998, 2.362829, 2.981421, 5.824724, 4.708407, 3.496197, 2.728604, 
    2.126799, 1.800239, 1.39707, 1.043489, 0.7960482, 0.5378286, 0.5031544, 
    0.5501498, 1.057133, 4.079216, 9.166537, 7.969213, 4.004428, 3.107512, 
    3.014899,
  4.869037, 10.33123, 10.05473, 5.151015, 2.491477, 1.972059, 1.701457, 
    1.701596, 2.20068, 2.675002, 2.763067, 3.0507, 2.160253, 1.172605, 
    0.6733555, 0.4904421, 0.5384364, 0.5385569, 0.4301637, 0.3885939, 
    0.5344524, 1.228795, 4.2483, 11.71032, 10.75997, 8.032099, 2.759496, 
    2.591142, 3.33441,
  9.923697, 18.23907, 16.00036, 4.292064, 2.183867, 1.941485, 2.069979, 
    2.341054, 4.585671, 7.209995, 3.027524, 2.069993, 1.027926, 0.4638813, 
    0.3694859, 0.3842845, 0.410007, 0.4297588, 0.499146, 0.5457723, 
    0.8744599, 1.634933, 5.208012, 10.96983, 7.812253, 4.479939, 3.738578, 
    4.423577, 5.955397,
  11.91618, 11.08157, 10.90409, 8.359364, 4.26669, 3.288913, 4.567597, 
    4.311891, 4.551157, 3.242229, 2.26896, 1.77285, 1.289031, 1.111883, 
    0.8554312, 0.835398, 0.8056557, 1.009362, 1.123106, 1.343839, 1.663274, 
    2.218811, 3.594744, 4.60871, 1.997598, 2.588714, 3.608673, 6.268638, 
    11.68186,
  6.696975, 5.189197, 4.619781, 8.883954, 6.542037, 5.546227, 6.188489, 
    7.474323, 8.293995, 5.538041, 3.820868, 2.779479, 2.428518, 2.873258, 
    3.032251, 2.725155, 2.083644, 1.920317, 1.753466, 2.248694, 3.000601, 
    4.324953, 2.296054, 2.063001, 1.819004, 2.111558, 3.07814, 4.458473, 
    4.944296,
  5.358634, 5.347701, 5.305471, 6.366942, 7.340802, 7.732112, 11.46079, 
    10.44122, 17.60733, 20.83975, 14.09571, 9.962207, 7.77075, 6.780212, 
    6.208395, 5.216723, 3.875997, 2.934543, 2.694544, 3.265342, 5.172385, 
    5.618476, 5.299451, 4.321221, 2.957787, 3.199229, 3.73034, 3.706909, 
    6.180785,
  5.977592, 6.529166, 7.669988, 8.624274, 13.1497, 10.50512, 14.89364, 
    17.08409, 16.16846, 15.07292, 13.21002, 11.05927, 9.933534, 8.327136, 
    7.149693, 6.037865, 5.178108, 4.234618, 3.543078, 3.705114, 6.276491, 
    8.814159, 7.654101, 7.760366, 6.892274, 5.991087, 4.953948, 4.370724, 
    4.510204,
  5.260959, 7.427051, 7.386576, 8.153484, 9.563104, 9.321963, 9.002777, 
    9.655906, 11.1051, 12.11073, 11.95998, 11.08745, 9.34289, 7.841994, 
    7.075999, 6.225314, 5.239411, 4.424889, 4.189902, 5.069248, 6.452775, 
    8.182209, 8.110361, 8.917301, 8.770969, 6.299463, 5.716386, 4.77071, 
    4.49317,
  4.963151, 5.966902, 6.847655, 7.327396, 7.982314, 8.619234, 8.673343, 
    9.164788, 9.300966, 8.799747, 9.670236, 9.497055, 8.223426, 7.028707, 
    6.246568, 5.603807, 5.139411, 4.718205, 4.724623, 5.574917, 6.167809, 
    5.982191, 6.160029, 7.368781, 7.42207, 6.438667, 5.500326, 4.997224, 
    4.681905,
  5.019511, 5.589746, 5.907118, 6.650708, 6.568672, 6.754752, 6.86503, 
    6.843895, 6.741898, 6.799544, 7.372096, 7.187245, 6.522538, 5.971663, 
    5.494614, 4.936649, 5.052636, 4.745072, 4.381207, 4.308669, 4.47867, 
    4.831729, 5.300239, 5.658435, 5.749367, 4.985647, 4.673476, 4.787138, 
    4.65831,
  4.712903, 4.713703, 4.84224, 4.936086, 5.158194, 5.357385, 5.350399, 
    5.49746, 5.617131, 5.609337, 5.543673, 5.558936, 5.431035, 5.130193, 
    4.841757, 4.519231, 4.374754, 4.259281, 4.238707, 4.308121, 4.326588, 
    4.38295, 4.424768, 4.709711, 4.965761, 4.550707, 4.468385, 4.820172, 
    4.807682,
  0.422201, 0.422201, 0.422201, 0.422201, 0.422201, 0.422201, 0.422201, 
    0.4153799, 0.4153799, 0.4153799, 0.4153799, 0.4153799, 0.4153799, 
    0.4153799, 0.4358175, 0.4358175, 0.4358175, 0.4358175, 0.4358175, 
    0.4358175, 0.4358175, 0.4382435, 0.4382435, 0.4382435, 0.4382435, 
    0.4382435, 0.4382435, 0.4382435, 0.422201,
  0.5396417, 0.5166984, 0.4949176, 0.4686637, 0.4620216, 0.436177, 0.4141854, 
    0.4143952, 0.4288028, 0.438999, 0.4503074, 0.4695933, 0.4582317, 
    0.3256658, 0.3280679, 0.3425202, 0.3575713, 0.4037128, 0.4552437, 
    0.4800135, 0.5037284, 0.5050967, 0.5166811, 0.4717281, 0.4709797, 
    0.4466813, 0.4195999, 0.4698704, 0.5417879,
  0.6222394, 0.6070442, 0.5586631, 0.5746126, 0.6913928, 0.6330594, 0.460942, 
    0.5423606, 0.4973672, 0.4659756, 0.5140303, 0.6260799, 0.6314629, 
    0.7043722, 0.7917068, 0.882282, 0.8722698, 0.7820233, 0.6306342, 
    0.5426329, 0.5138301, 0.5122885, 0.4903864, 0.6113013, 0.6978735, 
    0.7030692, 0.7513611, 0.7346159, 0.6696401,
  1.130131, 1.011918, 0.9639743, 0.9903185, 1.039952, 0.9726974, 0.7932405, 
    0.6809173, 0.5660404, 0.4879263, 0.483977, 0.7299343, 1.272265, 1.356744, 
    1.464241, 1.526034, 1.428223, 1.319208, 1.117286, 0.9428564, 0.7236208, 
    0.6350176, 0.6031497, 0.5982482, 1.045716, 1.288032, 1.491464, 1.333966, 
    1.227677,
  1.559357, 1.431251, 1.307014, 1.445425, 1.483069, 1.368485, 1.29047, 
    1.139005, 0.9623064, 0.8423779, 0.8264484, 1.143004, 1.885986, 2.275335, 
    2.246109, 2.002321, 1.693538, 1.616535, 1.456264, 1.218399, 1.062611, 
    0.9515331, 0.8196194, 0.954924, 1.583543, 2.078137, 1.988721, 1.917584, 
    1.724325,
  1.716971, 1.524672, 1.847669, 2.976717, 2.831978, 2.220216, 1.841259, 
    1.618934, 1.493076, 1.422031, 1.800308, 2.425164, 3.321371, 3.245917, 
    2.854721, 2.30045, 1.998562, 1.837837, 1.591597, 1.332078, 1.171094, 
    0.9591963, 0.9158268, 1.007814, 4.330112, 3.409727, 2.379594, 1.968235, 
    1.815021,
  2.182167, 2.694879, 6.33064, 6.052653, 3.38738, 2.716713, 2.33483, 2.26916, 
    2.211156, 2.569715, 5.404548, 5.854051, 5.26606, 3.41179, 2.691488, 
    2.534992, 2.220807, 1.761607, 1.3453, 1.116685, 0.8492827, 0.7525206, 
    0.703116, 1.080327, 8.272486, 5.434963, 3.42513, 2.562685, 2.259004,
  2.876342, 7.289421, 8.684439, 5.558702, 4.034698, 2.512774, 2.362023, 
    2.09862, 2.316746, 3.314503, 7.107865, 5.307982, 3.516088, 2.502909, 
    1.962608, 1.673885, 1.341314, 0.9925347, 0.7497688, 0.5596669, 0.4983103, 
    0.5858061, 0.9877203, 4.28679, 10.80539, 8.232718, 3.805631, 2.809447, 
    2.703176,
  5.028776, 11.51879, 10.79039, 5.407426, 2.335625, 1.786319, 1.586511, 
    1.602277, 2.141746, 2.74149, 2.864215, 3.109175, 2.210244, 1.173597, 
    0.6151419, 0.4492225, 0.4992974, 0.497488, 0.3958354, 0.3989694, 
    0.7326111, 1.699651, 5.731009, 12.87393, 11.26628, 8.448075, 2.408434, 
    2.322911, 3.19188,
  11.1414, 19.53128, 18.96892, 4.643572, 2.115223, 1.779477, 1.968068, 
    2.334266, 4.621789, 7.230543, 3.073791, 2.138183, 1.091242, 0.453858, 
    0.3477579, 0.3729907, 0.3944002, 0.4490445, 0.5413742, 0.6766378, 
    1.132279, 2.23228, 7.906651, 13.03254, 9.266685, 4.141261, 3.593157, 
    4.763458, 6.607039,
  12.49452, 12.38421, 12.86446, 11.16024, 5.190011, 3.543722, 4.99495, 
    4.998531, 4.719877, 3.273442, 2.22882, 1.766113, 1.245325, 1.064204, 
    0.8156128, 0.8097067, 0.8327226, 1.054056, 1.163124, 1.455718, 1.772574, 
    2.461455, 3.975625, 4.61583, 2.035338, 2.731457, 3.940603, 7.011693, 
    12.13184,
  10.46556, 7.626664, 6.212755, 11.49518, 8.697038, 6.756638, 6.60305, 
    8.630671, 8.916993, 6.130147, 3.801515, 2.622576, 2.401021, 2.85433, 
    3.034057, 2.678625, 2.017499, 1.803689, 1.898768, 2.459776, 3.436586, 
    5.103041, 2.337862, 2.067127, 1.81559, 2.251461, 3.649036, 6.085769, 
    8.469297,
  6.313296, 6.520682, 5.980338, 8.213882, 8.878246, 9.480556, 13.79578, 
    11.64729, 19.20183, 22.13269, 14.37177, 10.14791, 8.006044, 6.995897, 
    6.13848, 5.220359, 3.79, 2.870825, 2.685888, 3.379495, 5.904315, 
    6.469068, 5.769128, 4.48436, 2.985853, 3.164558, 3.68042, 3.977916, 
    7.584461,
  6.352198, 7.071095, 8.173812, 9.105913, 14.92999, 11.3853, 16.00791, 
    18.22509, 17.44188, 15.34707, 13.41362, 11.17571, 9.873379, 8.278228, 
    7.07072, 5.925046, 5.071661, 4.06995, 3.445087, 3.809483, 7.466981, 
    10.12538, 8.505663, 8.310048, 7.222537, 6.054366, 4.998078, 4.421699, 
    4.60625,
  5.373535, 7.74966, 7.602589, 8.496441, 9.939557, 9.8794, 9.503038, 
    9.911647, 11.7106, 12.89409, 12.41043, 11.7267, 9.680846, 7.962805, 
    7.110279, 6.201485, 5.166747, 4.40027, 4.054518, 5.166869, 7.172553, 
    9.022318, 8.882177, 9.770814, 9.539816, 6.571889, 5.821634, 4.788642, 
    4.513183,
  5.146191, 6.177919, 7.200531, 7.661706, 8.291861, 8.94287, 9.038209, 
    9.685389, 9.920354, 9.243078, 10.15154, 9.988005, 8.458743, 7.245403, 
    6.367535, 5.64791, 5.200042, 4.79294, 4.868264, 6.175256, 6.878348, 
    6.660987, 6.650882, 7.886792, 7.911841, 6.780308, 5.61394, 5.061311, 
    4.785237,
  5.251488, 5.811729, 6.157922, 7.00059, 6.957948, 7.130335, 7.37722, 
    7.204622, 7.132786, 7.140299, 7.638323, 7.47152, 6.652973, 6.118165, 
    5.662624, 5.040814, 5.216999, 4.936801, 4.570227, 4.508616, 4.839351, 
    5.198215, 5.646109, 5.986827, 6.057902, 5.206463, 4.919448, 4.91229, 
    4.755561,
  4.946179, 4.901503, 4.979996, 5.014976, 5.276876, 5.495563, 5.472912, 
    5.673965, 5.802153, 5.791982, 5.728997, 5.665944, 5.574175, 5.216418, 
    4.916191, 4.622755, 4.513306, 4.442266, 4.424323, 4.42187, 4.514665, 
    4.584603, 4.740288, 5.070077, 5.33653, 4.866573, 4.745408, 5.10942, 
    5.061909,
  0.4085007, 0.4085007, 0.4085007, 0.4085007, 0.4085007, 0.4085007, 
    0.4085007, 0.4025953, 0.4025953, 0.4025953, 0.4025953, 0.4025953, 
    0.4025953, 0.4025953, 0.4207416, 0.4207416, 0.4207416, 0.4207416, 
    0.4207416, 0.4207416, 0.4207416, 0.4239167, 0.4239167, 0.4239167, 
    0.4239167, 0.4239167, 0.4239167, 0.4239167, 0.4085007,
  0.5178865, 0.4952067, 0.4719208, 0.4446789, 0.4443918, 0.4201009, 
    0.4022813, 0.4040679, 0.4176518, 0.4251699, 0.4261926, 0.4263141, 
    0.4013544, 0.2826695, 0.282661, 0.2943943, 0.3100562, 0.3609417, 
    0.4146357, 0.4438801, 0.4717794, 0.4800691, 0.4905145, 0.4601744, 
    0.4591856, 0.4231157, 0.3996142, 0.449747, 0.5103241,
  0.5854673, 0.5377709, 0.4905567, 0.5133541, 0.6502429, 0.5868708, 
    0.3974669, 0.493475, 0.4486746, 0.4224141, 0.4582591, 0.5758483, 
    0.5702977, 0.6279431, 0.7041332, 0.7857108, 0.7816647, 0.6950992, 
    0.575071, 0.4918195, 0.459661, 0.4629921, 0.4482715, 0.5834113, 
    0.6748348, 0.6899661, 0.7376934, 0.7148767, 0.6349729,
  1.083838, 0.9729016, 0.9103451, 0.9496826, 0.9935474, 0.900965, 0.7267334, 
    0.6250674, 0.5125477, 0.4445347, 0.4389457, 0.6601321, 1.236635, 
    1.269136, 1.344147, 1.396411, 1.293928, 1.161872, 1.007508, 0.8323194, 
    0.6491666, 0.55835, 0.5568988, 0.563101, 1.037375, 1.330773, 1.530387, 
    1.357285, 1.214047,
  1.576121, 1.392368, 1.261735, 1.410142, 1.427376, 1.302441, 1.209655, 
    1.036952, 0.8574746, 0.7685022, 0.7593694, 1.106879, 1.866243, 2.232638, 
    2.175567, 1.873151, 1.5529, 1.490427, 1.329314, 1.11077, 0.9768289, 
    0.8642536, 0.7521284, 0.9200097, 1.746734, 2.248215, 2.022495, 1.952384, 
    1.713147,
  1.657063, 1.448026, 1.811552, 3.117473, 2.76112, 2.060162, 1.701016, 
    1.465502, 1.339107, 1.324163, 1.889058, 2.568473, 3.746917, 3.403244, 
    2.740799, 2.175376, 1.879223, 1.676296, 1.462974, 1.242674, 1.09901, 
    0.8789531, 0.8662632, 1.03009, 5.313493, 3.680618, 2.393399, 1.953385, 
    1.772343,
  1.926104, 2.629132, 7.341014, 6.85968, 3.411253, 2.59425, 2.152327, 
    2.04335, 2.013447, 2.639838, 6.525577, 7.383804, 6.4665, 3.861833, 
    2.678456, 2.344095, 2.035825, 1.669234, 1.289236, 1.081687, 0.825924, 
    0.7455428, 0.6732551, 1.241314, 10.19787, 5.841956, 3.424361, 2.358335, 
    2.010806,
  2.878006, 9.135267, 9.757432, 6.303328, 4.096229, 2.312392, 2.162508, 
    1.993305, 2.371456, 3.965542, 9.229852, 6.604053, 3.650014, 2.407322, 
    1.846342, 1.634052, 1.229051, 0.9321774, 0.7030004, 0.5624092, 0.4920509, 
    0.6053295, 0.9704955, 4.582595, 12.6065, 8.841123, 3.695661, 2.554951, 
    2.440643,
  5.733972, 13.10889, 12.176, 5.866297, 2.388083, 1.670569, 1.481503, 
    1.52733, 2.122234, 2.960692, 3.004035, 3.189665, 2.269888, 1.134982, 
    0.5537133, 0.4119806, 0.4647304, 0.452564, 0.3802148, 0.478104, 1.008141, 
    2.287427, 7.51822, 14.44441, 12.56179, 9.416573, 2.261592, 2.188044, 
    3.165449,
  12.65036, 21.40991, 22.48511, 5.441207, 2.427013, 1.752241, 1.900383, 
    2.398619, 4.727294, 7.255778, 3.14032, 2.234562, 1.145368, 0.4439801, 
    0.3301685, 0.360096, 0.3938824, 0.4727516, 0.6248598, 0.9041242, 1.535, 
    3.351877, 11.16195, 15.11526, 10.15949, 3.764845, 3.616124, 5.214777, 
    7.62129,
  15.15291, 16.00085, 16.38928, 15.46259, 6.511304, 4.1182, 5.800113, 
    5.58042, 5.002998, 3.363351, 2.215693, 1.769192, 1.202015, 0.9974856, 
    0.7847748, 0.762325, 0.8557, 1.061285, 1.19223, 1.572682, 2.004011, 
    2.826579, 4.517325, 4.815728, 2.168135, 2.948451, 4.634333, 8.276731, 
    14.20634,
  14.25737, 11.35691, 8.501834, 13.83794, 11.20703, 7.988535, 7.342865, 
    10.15465, 10.05503, 7.117935, 4.1278, 2.5325, 2.429636, 2.889133, 
    2.999347, 2.616574, 1.915408, 1.814106, 2.079954, 2.6517, 4.011153, 
    6.254336, 2.478878, 2.175897, 1.882515, 2.688405, 4.585261, 7.942596, 
    12.41204,
  7.662095, 7.996233, 6.903494, 10.51807, 11.21674, 11.96964, 16.63029, 
    13.08563, 21.13773, 23.45951, 14.48596, 10.0716, 7.972322, 6.992015, 
    5.996451, 5.178723, 3.752561, 2.81302, 2.662016, 3.436779, 6.8268, 
    7.733213, 6.365531, 4.711733, 3.094453, 3.255763, 3.641943, 4.174583, 
    9.161661,
  7.010302, 7.826947, 8.959682, 9.962252, 16.90058, 12.79811, 17.37388, 
    19.80398, 19.14335, 15.86227, 13.94258, 11.60736, 9.845632, 8.231084, 
    6.920034, 5.786883, 4.924114, 3.909558, 3.376107, 3.959286, 8.882689, 
    11.80634, 9.611359, 9.078629, 7.806161, 6.265675, 5.089943, 4.564965, 
    4.847975,
  5.567079, 8.204716, 8.131557, 9.03103, 10.75931, 10.78774, 10.4134, 
    10.30567, 12.58707, 14.1032, 13.14912, 12.41857, 10.1495, 8.187666, 
    7.235732, 6.223372, 5.176535, 4.385185, 3.998873, 5.37366, 8.276681, 
    10.13764, 9.843697, 10.80315, 10.45115, 6.964316, 6.003477, 4.853985, 
    4.587971,
  5.375735, 6.489884, 7.773575, 8.263179, 8.815295, 9.485557, 9.601275, 
    10.48691, 10.72726, 9.909494, 10.94053, 10.5005, 8.721387, 7.495829, 
    6.518252, 5.676002, 5.380864, 4.942713, 5.127532, 7.064194, 7.703445, 
    7.515315, 7.32713, 8.550297, 8.406244, 7.177379, 5.729695, 5.178922, 
    4.924329,
  5.470695, 5.963122, 6.550839, 7.409849, 7.420152, 7.523644, 7.894755, 
    7.647454, 7.649834, 7.440273, 8.014024, 7.773956, 6.864933, 6.283387, 
    5.950289, 5.257502, 5.436222, 5.252913, 4.911655, 4.842297, 5.341891, 
    5.633408, 5.993402, 6.338379, 6.448245, 5.439291, 5.156918, 5.054216, 
    4.902549,
  5.167388, 5.119462, 5.193062, 5.189609, 5.440862, 5.632386, 5.66115, 
    5.867475, 5.976771, 5.961003, 5.983583, 5.830003, 5.697035, 5.30933, 
    5.002367, 4.696952, 4.657707, 4.628367, 4.594543, 4.508456, 4.665158, 
    4.742321, 5.042722, 5.442081, 5.724158, 5.223844, 5.041474, 5.37058, 
    5.292368,
  0.386014, 0.386014, 0.386014, 0.386014, 0.386014, 0.386014, 0.386014, 
    0.3830342, 0.3830342, 0.3830342, 0.3830342, 0.3830342, 0.3830342, 
    0.3830342, 0.401552, 0.401552, 0.401552, 0.401552, 0.401552, 0.401552, 
    0.401552, 0.4015134, 0.4015134, 0.4015134, 0.4015134, 0.4015134, 
    0.4015134, 0.4015134, 0.386014,
  0.4916043, 0.4708295, 0.4404637, 0.4188446, 0.4189212, 0.4014156, 
    0.3882928, 0.385456, 0.394096, 0.4036878, 0.3969638, 0.3766678, 
    0.3543891, 0.2487591, 0.2429411, 0.2497381, 0.2683475, 0.3212067, 
    0.3748664, 0.4123826, 0.4410431, 0.4556623, 0.465684, 0.446905, 0.447824, 
    0.4045849, 0.3831765, 0.430271, 0.4787789,
  0.5506598, 0.4650751, 0.4263449, 0.4480257, 0.6040003, 0.5420875, 
    0.3424127, 0.4464269, 0.4058186, 0.383694, 0.4154946, 0.522185, 
    0.5194613, 0.5613132, 0.6358685, 0.7113853, 0.7009028, 0.6234919, 
    0.5258039, 0.4482213, 0.4086617, 0.4157642, 0.4246732, 0.5667987, 
    0.6751621, 0.6926973, 0.7204195, 0.700236, 0.6044539,
  1.0401, 0.9266856, 0.8618289, 0.8930199, 0.9443891, 0.8243532, 0.6656476, 
    0.5720145, 0.4603932, 0.4075617, 0.3995584, 0.6034288, 1.205645, 
    1.185781, 1.240844, 1.272915, 1.169276, 1.036667, 0.9048151, 0.7394927, 
    0.5798562, 0.4950227, 0.5126013, 0.5349408, 1.048149, 1.39505, 1.604709, 
    1.391193, 1.197364,
  1.58677, 1.338758, 1.220271, 1.394009, 1.380713, 1.249544, 1.14586, 
    0.9314539, 0.7584853, 0.6948277, 0.702108, 1.0895, 1.85334, 2.222469, 
    2.129946, 1.759653, 1.450547, 1.358988, 1.214831, 0.9984766, 0.8813043, 
    0.7779297, 0.6845802, 0.9004177, 2.049775, 2.479788, 2.102053, 2.013136, 
    1.722473,
  1.599625, 1.422771, 1.836078, 3.297168, 2.62628, 1.874534, 1.559741, 
    1.333121, 1.185052, 1.243197, 1.965535, 2.724534, 4.284273, 3.633725, 
    2.68896, 2.087752, 1.773894, 1.526362, 1.310964, 1.158372, 1.024011, 
    0.8189529, 0.8265727, 1.094708, 6.38239, 3.998225, 2.381033, 2.013583, 
    1.739837,
  1.739973, 2.696682, 8.746685, 7.644805, 3.460996, 2.50772, 2.02963, 
    1.868342, 1.786925, 2.834172, 7.987703, 9.102013, 7.969521, 4.397571, 
    2.657378, 2.142466, 1.851154, 1.570716, 1.211855, 1.025812, 0.7894882, 
    0.7196169, 0.6533027, 1.578876, 12.20948, 6.348591, 3.473634, 2.178874, 
    1.743895,
  2.980038, 10.87679, 11.66725, 7.024571, 4.284504, 2.162306, 1.996759, 
    1.916327, 2.54829, 4.906534, 12.01634, 8.102642, 4.083969, 2.457218, 
    1.752808, 1.592566, 1.166787, 0.8954374, 0.6665742, 0.5554736, 0.5003049, 
    0.6160262, 0.948887, 4.66363, 14.82086, 9.707255, 3.585842, 2.349146, 
    2.305006,
  6.733028, 14.74518, 14.36307, 6.537492, 2.523408, 1.591638, 1.397973, 
    1.522694, 2.160167, 3.224741, 3.254379, 3.357115, 2.321369, 1.074453, 
    0.500952, 0.3871958, 0.4393167, 0.4317013, 0.3889903, 0.6110874, 
    1.266945, 2.962965, 9.105339, 15.86286, 13.93409, 11.10744, 2.230859, 
    2.164061, 3.481225,
  14.54674, 23.83436, 26.07857, 6.834761, 3.028037, 1.778256, 1.902703, 
    2.545148, 4.930189, 7.315205, 3.229786, 2.301886, 1.17961, 0.4375384, 
    0.3186407, 0.3506802, 0.4116109, 0.5273649, 0.7420083, 1.153094, 
    2.168866, 4.865694, 13.93444, 16.90498, 11.40959, 3.603854, 3.910183, 
    5.90994, 9.385674,
  19.74921, 20.07997, 20.72582, 20.33154, 7.824087, 4.993701, 6.964091, 
    6.053187, 5.433716, 3.510124, 2.246131, 1.7733, 1.201076, 0.917092, 
    0.7474464, 0.7117423, 0.8411539, 1.043512, 1.2539, 1.729297, 2.342953, 
    3.219156, 5.036291, 5.366856, 2.373295, 3.266048, 5.608731, 10.4106, 
    18.85046,
  16.59542, 15.55372, 10.99593, 15.50974, 14.98792, 8.99147, 8.596321, 
    11.78421, 11.55481, 8.550052, 4.665978, 2.625885, 2.52107, 2.973607, 
    2.984877, 2.49862, 1.923262, 1.859848, 2.143517, 2.785295, 4.610756, 
    7.740342, 2.717589, 2.41936, 2.129325, 3.1786, 5.369482, 9.206231, 
    15.08452,
  9.542372, 9.675598, 8.009172, 12.86524, 13.9561, 14.75342, 19.86579, 
    14.65578, 23.55725, 24.70598, 14.49007, 9.912906, 7.805354, 6.850552, 
    5.882484, 5.069831, 3.69663, 2.769198, 2.630056, 3.479846, 7.970852, 
    9.41915, 7.18258, 4.97342, 3.278705, 3.379791, 3.614964, 4.38204, 10.69407,
  8.040668, 8.760389, 10.20903, 11.20384, 19.06792, 14.58714, 19.11154, 
    22.00142, 21.43536, 16.872, 14.99541, 12.38645, 10.07528, 8.182185, 
    6.768749, 5.659452, 4.721403, 3.73766, 3.289271, 4.227012, 10.36442, 
    13.95394, 11.00732, 10.17562, 8.721286, 6.629236, 5.184361, 4.775175, 
    5.222241,
  5.865205, 8.762828, 9.065492, 9.997684, 12.06332, 12.18645, 11.61605, 
    10.92828, 13.83514, 15.70537, 14.41628, 13.2212, 10.87754, 8.635732, 
    7.420787, 6.235508, 5.192486, 4.43733, 4.029924, 5.70355, 9.892266, 
    11.46633, 10.9859, 12.2056, 11.51183, 7.571972, 6.318246, 5.048354, 
    4.656279,
  5.755693, 6.953564, 8.629956, 9.159878, 9.840661, 10.36504, 10.55446, 
    11.66584, 11.94622, 11.0542, 12.00478, 11.15517, 9.158191, 7.754143, 
    6.730337, 5.797534, 5.623931, 5.274483, 5.555952, 8.129274, 8.686009, 
    8.405701, 8.056548, 9.3703, 9.112658, 7.580389, 5.911492, 5.360667, 
    5.182347,
  5.731811, 6.241568, 7.084182, 7.998657, 7.856518, 7.986168, 8.471828, 
    8.273198, 8.407713, 7.902462, 8.460793, 8.171296, 7.195158, 6.530008, 
    6.246881, 5.610616, 5.687343, 5.675488, 5.372723, 5.349068, 5.918868, 
    6.126933, 6.393237, 6.733722, 6.944304, 5.710747, 5.372824, 5.249614, 
    5.107621,
  5.375138, 5.293825, 5.525606, 5.542349, 5.837532, 5.95204, 6.001205, 
    6.140661, 6.226977, 6.132669, 6.207244, 6.026155, 5.838483, 5.485769, 
    5.226771, 4.855654, 4.791479, 4.834975, 4.790953, 4.570291, 4.737272, 
    4.871879, 5.321206, 5.790784, 6.097824, 5.591469, 5.380283, 5.630061, 
    5.516533,
  0.3577868, 0.3577868, 0.3577868, 0.3577868, 0.3577868, 0.3577868, 
    0.3577868, 0.3595785, 0.3595785, 0.3595785, 0.3595785, 0.3595785, 
    0.3595785, 0.3595785, 0.3793937, 0.3793937, 0.3793937, 0.3793937, 
    0.3793937, 0.3793937, 0.3793937, 0.3737674, 0.3737674, 0.3737674, 
    0.3737674, 0.3737674, 0.3737674, 0.3737674, 0.3577868,
  0.4621152, 0.4425593, 0.4075545, 0.3912147, 0.3872158, 0.3793467, 
    0.3720371, 0.3638122, 0.3684734, 0.3792154, 0.3628754, 0.335804, 
    0.3172847, 0.2213806, 0.2095009, 0.2143663, 0.2336375, 0.2835575, 
    0.3374804, 0.3821969, 0.4108911, 0.4321919, 0.4440573, 0.422275, 
    0.431178, 0.3883352, 0.3682009, 0.4121437, 0.4477853,
  0.5135285, 0.3972056, 0.3747752, 0.3900538, 0.5547303, 0.49357, 0.2972864, 
    0.4042055, 0.3711668, 0.3483461, 0.3824038, 0.4761887, 0.470999, 
    0.4975251, 0.5922672, 0.6547085, 0.6307587, 0.568052, 0.4775018, 
    0.4065716, 0.3595491, 0.3737726, 0.3958505, 0.5659656, 0.6899595, 
    0.7117273, 0.7289334, 0.6891961, 0.5826855,
  0.9984945, 0.8755718, 0.8113584, 0.8257257, 0.8878483, 0.7511522, 
    0.6100084, 0.5161628, 0.4106474, 0.374864, 0.3643626, 0.5546753, 
    1.162654, 1.109022, 1.159776, 1.169568, 1.064526, 0.9307426, 0.817423, 
    0.6601735, 0.511801, 0.4357206, 0.4719939, 0.5207644, 1.086937, 1.500477, 
    1.70061, 1.438472, 1.178898,
  1.58914, 1.296246, 1.185556, 1.390983, 1.343958, 1.212417, 1.078007, 
    0.8302355, 0.6660163, 0.6153575, 0.6601291, 1.073194, 1.85231, 2.207075, 
    2.100458, 1.678368, 1.361323, 1.249611, 1.119394, 0.8945985, 0.7884684, 
    0.6994275, 0.6147751, 0.9136242, 2.529721, 2.715071, 2.280047, 2.095911, 
    1.769615,
  1.568499, 1.403091, 1.908261, 3.506229, 2.486282, 1.708029, 1.419128, 
    1.215822, 1.052658, 1.132549, 2.065155, 2.912438, 4.946997, 3.926001, 
    2.717625, 2.024386, 1.661132, 1.397155, 1.165009, 1.062635, 0.9336925, 
    0.7628322, 0.7771778, 1.208556, 7.50268, 4.270973, 2.411995, 2.095499, 
    1.742175,
  1.575328, 2.686958, 10.60588, 8.156214, 3.435246, 2.412279, 1.879996, 
    1.720024, 1.564537, 3.223666, 9.681874, 10.94058, 9.681306, 4.890268, 
    2.6472, 1.977858, 1.662989, 1.44125, 1.095193, 0.9674371, 0.7468223, 
    0.6696823, 0.6242568, 2.13555, 14.33309, 7.013193, 3.465991, 1.998886, 
    1.513772,
  2.85318, 12.12838, 14.00944, 7.628555, 4.56813, 2.075727, 1.852334, 
    1.967404, 2.834832, 6.380524, 15.1788, 10.1697, 4.68844, 2.478406, 
    1.664788, 1.499651, 1.161308, 0.8462805, 0.6420256, 0.5531222, 0.5270361, 
    0.6242578, 0.8183963, 4.601675, 17.41826, 10.92691, 3.56691, 2.087685, 
    2.183079,
  7.331345, 16.15655, 16.86195, 7.418595, 2.571653, 1.577271, 1.36382, 
    1.641644, 2.296813, 3.582144, 3.729985, 3.664105, 2.38983, 0.9983396, 
    0.4597539, 0.3811181, 0.4331723, 0.394558, 0.4548983, 0.7638806, 
    1.585839, 3.776247, 9.869789, 17.57279, 15.70627, 12.77052, 2.314155, 
    2.184293, 3.86025,
  16.7887, 26.40076, 29.34356, 8.499919, 3.533456, 1.907966, 2.0033, 
    2.587203, 5.36577, 7.668701, 3.383436, 2.327813, 1.188104, 0.4341869, 
    0.3098183, 0.3449872, 0.4297146, 0.6021509, 0.9058422, 1.453673, 
    2.937604, 6.726599, 15.96726, 18.55647, 13.36374, 3.901952, 4.433115, 
    7.036042, 11.8323,
  24.69301, 24.64498, 24.75267, 24.70407, 9.22546, 5.976706, 8.412181, 
    6.618783, 5.961825, 3.838469, 2.386973, 1.806071, 1.229897, 0.8456407, 
    0.6788554, 0.6664755, 0.8009912, 1.039566, 1.343314, 1.91869, 2.725571, 
    3.657526, 5.477835, 6.37036, 2.653505, 3.791264, 6.629488, 13.59436, 
    23.81636,
  18.15504, 18.7805, 13.46883, 16.774, 19.20833, 10.2148, 10.62656, 13.55903, 
    13.52152, 10.12945, 5.413561, 2.943255, 2.724312, 3.137978, 3.014012, 
    2.401267, 1.965469, 1.840395, 2.167859, 2.835049, 5.279309, 9.468008, 
    3.013271, 2.777852, 2.436518, 3.551137, 5.764651, 9.838005, 17.15692,
  12.00575, 11.56741, 9.49785, 15.33572, 16.98326, 17.48139, 23.19144, 
    16.4981, 26.239, 25.78434, 14.35931, 9.720002, 7.689239, 6.634391, 
    5.802736, 4.901485, 3.643173, 2.706789, 2.606884, 3.594208, 9.187654, 
    11.56088, 8.302844, 5.372352, 3.637206, 3.506068, 3.550413, 4.588746, 
    12.12108,
  9.374531, 9.758392, 11.95661, 12.82915, 21.33667, 16.79852, 21.13767, 
    24.19665, 24.09283, 18.44169, 16.64661, 13.64163, 10.6202, 8.204003, 
    6.733275, 5.539207, 4.557349, 3.569892, 3.205585, 4.678806, 11.83634, 
    16.3805, 12.75873, 11.64714, 9.917389, 7.102674, 5.402394, 5.016577, 
    5.823049,
  6.342595, 9.452209, 10.32368, 11.4183, 13.95693, 14.21024, 13.19123, 
    11.84682, 15.407, 17.69206, 16.36497, 14.30107, 11.86751, 9.402524, 
    7.64706, 6.284827, 5.234653, 4.575281, 4.09865, 6.171132, 12.0544, 
    13.3494, 12.42595, 14.01606, 13.05674, 8.434604, 6.793062, 5.356889, 
    4.834651,
  6.266198, 7.717208, 9.824766, 10.38107, 11.15088, 11.58399, 11.92878, 
    13.25989, 13.58702, 12.44086, 13.46331, 12.05295, 9.778989, 8.173794, 
    7.115692, 6.065775, 5.990602, 5.78584, 6.185392, 9.540585, 10.17593, 
    9.49236, 8.874978, 10.42885, 9.971107, 8.037108, 6.164961, 5.622756, 
    5.567425,
  6.069885, 6.651186, 7.683175, 8.703354, 8.527191, 8.618951, 9.166674, 
    9.092841, 9.475831, 8.66279, 9.074577, 8.794359, 7.718733, 6.944767, 
    6.625087, 6.032003, 6.029583, 6.24219, 5.948531, 6.175092, 6.584741, 
    6.693428, 6.886294, 7.16985, 7.415013, 5.998874, 5.562516, 5.447266, 
    5.376709,
  5.526995, 5.435729, 5.816034, 5.988952, 6.333632, 6.514092, 6.50246, 
    6.612515, 6.679512, 6.543686, 6.523313, 6.367948, 6.106547, 5.838532, 
    5.575667, 5.091429, 5.047163, 5.10196, 5.056419, 4.744507, 4.853909, 
    5.096746, 5.622617, 6.132305, 6.44678, 5.953058, 5.723473, 5.84987, 
    5.72502,
  0.3326207, 0.3326207, 0.3326207, 0.3326207, 0.3326207, 0.3326207, 
    0.3326207, 0.3342404, 0.3342404, 0.3342404, 0.3342404, 0.3342404, 
    0.3342404, 0.3342404, 0.3538899, 0.3538899, 0.3538899, 0.3538899, 
    0.3538899, 0.3538899, 0.3538899, 0.3456289, 0.3456289, 0.3456289, 
    0.3456289, 0.3456289, 0.3456289, 0.3456289, 0.3326207,
  0.432183, 0.4118441, 0.3793661, 0.3662605, 0.3563295, 0.3532245, 0.3518472, 
    0.3419802, 0.3443062, 0.3509765, 0.3294756, 0.3014341, 0.2867844, 
    0.2002295, 0.1849979, 0.1902862, 0.2076301, 0.2517448, 0.3019792, 
    0.3521689, 0.3820268, 0.4119865, 0.424049, 0.3922689, 0.405971, 
    0.3694567, 0.3518106, 0.3943675, 0.417764,
  0.4682986, 0.3393969, 0.3316727, 0.3416774, 0.5036536, 0.4425448, 
    0.2588435, 0.3665715, 0.3435279, 0.3211982, 0.3551404, 0.4396911, 
    0.4261993, 0.4399126, 0.5589776, 0.6094783, 0.5642729, 0.5173516, 
    0.4329465, 0.374484, 0.3231242, 0.3481743, 0.3784904, 0.5824266, 
    0.7120097, 0.7288107, 0.745435, 0.683933, 0.5642129,
  0.9631189, 0.8206059, 0.7629514, 0.757503, 0.8204271, 0.6816905, 0.554069, 
    0.4630088, 0.3649595, 0.3406985, 0.3344384, 0.5251477, 1.104862, 
    1.040543, 1.082356, 1.07601, 0.9694422, 0.8415248, 0.737057, 0.5862724, 
    0.4562699, 0.3906625, 0.4279428, 0.5257705, 1.168334, 1.666375, 1.807984, 
    1.482689, 1.178445,
  1.57598, 1.25908, 1.169961, 1.402462, 1.297657, 1.173851, 1.011669, 
    0.7531738, 0.5904865, 0.5407007, 0.6195559, 1.061969, 1.863931, 2.184549, 
    2.104008, 1.628421, 1.298345, 1.149686, 1.021699, 0.7939112, 0.6970042, 
    0.6171115, 0.5512077, 0.9810577, 3.155931, 2.997403, 2.558931, 2.192266, 
    1.813643,
  1.550659, 1.383609, 2.000563, 3.663587, 2.344079, 1.577258, 1.293459, 
    1.115098, 0.9570969, 1.019388, 2.158909, 3.09289, 5.680274, 4.146613, 
    2.801975, 1.974612, 1.538662, 1.257467, 1.030509, 0.9595098, 0.841924, 
    0.7040387, 0.7187905, 1.399749, 8.572908, 4.474637, 2.506349, 2.126166, 
    1.769662,
  1.436017, 2.60629, 12.77791, 8.366887, 3.411251, 2.241537, 1.694247, 
    1.566914, 1.375473, 3.745356, 11.50945, 13.03197, 11.70771, 5.254215, 
    2.660142, 1.780192, 1.480093, 1.284204, 0.9855334, 0.8887178, 0.6936936, 
    0.6364708, 0.6026437, 2.696293, 16.45351, 7.777997, 3.392865, 1.792721, 
    1.321216,
  2.583278, 13.33637, 17.0301, 8.193953, 4.818723, 1.936141, 1.739769, 
    2.031457, 3.192549, 8.555649, 19.37386, 13.31595, 5.225355, 2.540392, 
    1.576877, 1.348109, 1.124004, 0.7897964, 0.5728529, 0.5304452, 0.5456712, 
    0.5948945, 0.7331609, 4.517885, 20.79429, 12.59955, 3.492125, 1.783479, 
    2.04045,
  7.067732, 17.59692, 19.36902, 8.768515, 2.556671, 1.507043, 1.355292, 
    1.861194, 2.667509, 4.295358, 4.655681, 4.106831, 2.467562, 0.9279485, 
    0.4384148, 0.3526246, 0.4355804, 0.3983923, 0.5717857, 0.9461907, 
    1.954609, 4.325752, 9.557686, 19.79542, 17.86095, 14.2259, 2.356148, 
    2.218385, 3.964425,
  18.63166, 29.23258, 32.61956, 10.46144, 3.788923, 2.126274, 2.174945, 
    2.569672, 6.154706, 8.481604, 3.536264, 2.346076, 1.185528, 0.4290014, 
    0.3084539, 0.3603823, 0.4729608, 0.6926748, 1.079644, 1.884566, 3.923146, 
    8.301534, 17.06477, 20.64576, 15.92218, 4.683109, 5.116963, 8.323365, 
    13.92214,
  29.48943, 28.70185, 28.62796, 28.12488, 10.80742, 6.861437, 10.11266, 
    7.2941, 6.690565, 4.341392, 2.673907, 1.88516, 1.241314, 0.8066381, 
    0.6238084, 0.6439293, 0.786463, 1.076429, 1.462234, 2.154159, 3.133757, 
    4.310938, 5.994026, 7.975487, 2.980314, 4.192974, 7.499698, 17.27044, 
    28.54628,
  19.90008, 21.33663, 15.83748, 18.13738, 22.51963, 11.71377, 13.73624, 
    15.64869, 16.08646, 11.70947, 6.187667, 3.349791, 3.087202, 3.403272, 
    3.144082, 2.367933, 1.981249, 1.822758, 2.120688, 2.877769, 5.861704, 
    11.32762, 3.473439, 3.360561, 2.623927, 3.722178, 6.011337, 10.16253, 
    18.9528,
  14.9304, 13.73322, 11.36128, 18.08123, 20.00519, 20.32267, 26.3177, 
    18.49464, 28.87523, 26.68645, 14.08636, 9.727609, 7.678439, 6.442278, 
    5.692255, 4.718297, 3.558086, 2.673314, 2.647877, 3.805799, 10.57777, 
    14.09147, 9.575438, 5.978464, 4.090816, 3.679265, 3.54278, 4.822485, 
    13.53388,
  11.02217, 10.98313, 14.15526, 14.91146, 23.97664, 19.62215, 23.4639, 
    26.75547, 27.02871, 20.68734, 18.97766, 15.41738, 11.58395, 8.402224, 
    6.774495, 5.429474, 4.500171, 3.478561, 3.177764, 5.534088, 13.43634, 
    19.1659, 15.10409, 13.70077, 11.41332, 7.659076, 5.730975, 5.382191, 
    6.5722,
  7.052025, 10.4278, 12.02876, 13.49007, 16.35554, 17.17268, 15.5322, 
    13.06652, 17.38842, 20.08398, 19.34436, 15.97333, 13.10491, 10.32931, 
    7.940414, 6.424524, 5.329937, 4.795416, 4.312059, 6.918139, 14.8136, 
    15.72757, 14.31437, 16.19739, 14.81749, 9.452079, 7.396464, 5.744777, 
    5.171534,
  6.974178, 8.7914, 11.43868, 11.9663, 12.84739, 13.35057, 13.76736, 
    15.43374, 15.69164, 14.06473, 15.24736, 13.32362, 10.49825, 8.72414, 
    7.732598, 6.505746, 6.415236, 6.535479, 7.082987, 11.45292, 12.1308, 
    10.89771, 9.875382, 11.77002, 10.98646, 8.535945, 6.475324, 5.897233, 
    5.974955,
  6.560389, 7.317565, 8.479062, 9.520387, 9.481074, 9.53187, 9.973522, 
    10.26442, 10.76093, 9.824098, 9.973387, 9.668852, 8.474718, 7.51317, 
    7.076726, 6.577693, 6.62678, 6.999592, 6.792582, 7.174347, 7.450513, 
    7.331534, 7.478308, 7.631031, 7.794359, 6.263442, 5.721426, 5.633676, 
    5.679035,
  5.672016, 5.689579, 6.106973, 6.543521, 6.944693, 7.279668, 7.246957, 
    7.329135, 7.336554, 7.203969, 7.02449, 6.843297, 6.597921, 6.309377, 
    6.024082, 5.516025, 5.442975, 5.475163, 5.404041, 5.066904, 5.123554, 
    5.456636, 5.920841, 6.47606, 6.756511, 6.289413, 6.038975, 6.06457, 
    5.885837,
  0.3141891, 0.3141891, 0.3141891, 0.3141891, 0.3141891, 0.3141891, 
    0.3141891, 0.3133451, 0.3133451, 0.3133451, 0.3133451, 0.3133451, 
    0.3133451, 0.3133451, 0.3310637, 0.3310637, 0.3310637, 0.3310637, 
    0.3310637, 0.3310637, 0.3310637, 0.3248012, 0.3248012, 0.3248012, 
    0.3248012, 0.3248012, 0.3248012, 0.3248012, 0.3141891,
  0.4043238, 0.3821345, 0.3562676, 0.3480269, 0.3264943, 0.3261846, 
    0.3297152, 0.3214499, 0.3206889, 0.3209597, 0.2981658, 0.2722267, 
    0.2599746, 0.1856776, 0.1688999, 0.1746962, 0.1879235, 0.227186, 
    0.2703045, 0.3227807, 0.3575906, 0.3926541, 0.4062383, 0.356951, 
    0.3832273, 0.3527659, 0.333094, 0.3752245, 0.3955382,
  0.4124414, 0.2919462, 0.2903674, 0.3006163, 0.4508547, 0.3917387, 
    0.2271082, 0.3323115, 0.3207025, 0.3002974, 0.332868, 0.4087169, 
    0.3845711, 0.3857533, 0.5148599, 0.5561337, 0.5128297, 0.4705262, 
    0.3961415, 0.348511, 0.2956603, 0.3318829, 0.3668692, 0.6051595, 
    0.7183058, 0.7497523, 0.7523414, 0.6739088, 0.5415813,
  0.9259799, 0.7642347, 0.7103467, 0.6964974, 0.7544551, 0.6149823, 
    0.4990429, 0.417933, 0.3273261, 0.3134174, 0.3100398, 0.4895061, 
    1.052216, 0.9935879, 1.022023, 1.020013, 0.8999429, 0.7647614, 0.6642144, 
    0.5264824, 0.4096563, 0.3511035, 0.3905554, 0.5337487, 1.279386, 
    1.808987, 1.895239, 1.508447, 1.193873,
  1.540464, 1.225595, 1.160095, 1.389137, 1.244034, 1.139116, 0.9473259, 
    0.6820261, 0.529213, 0.4760045, 0.5818937, 1.030873, 1.876259, 2.168595, 
    2.107407, 1.606039, 1.230268, 1.080678, 0.9230027, 0.71333, 0.6075619, 
    0.5352368, 0.4925869, 1.153492, 3.947908, 3.36704, 2.847662, 2.272657, 
    1.843152,
  1.553338, 1.378231, 2.078479, 3.606371, 2.142649, 1.442056, 1.182558, 
    1.017918, 0.8766025, 0.9120506, 2.260875, 3.257392, 6.407698, 4.231384, 
    3.005481, 1.961103, 1.412143, 1.121171, 0.9018645, 0.8641638, 0.767226, 
    0.6489313, 0.6794383, 1.76678, 9.634652, 4.634138, 2.642349, 2.141187, 
    1.790335,
  1.344231, 2.646756, 15.15038, 8.147523, 3.308192, 2.01959, 1.489762, 
    1.39431, 1.222132, 4.343234, 13.60446, 14.83629, 13.61248, 5.354979, 
    2.61159, 1.62033, 1.301033, 1.10575, 0.8614949, 0.7724336, 0.6316273, 
    0.5964534, 0.5684513, 3.25112, 18.41408, 8.509464, 3.207131, 1.600623, 
    1.219337,
  2.472952, 14.89827, 20.72622, 8.688679, 4.840539, 1.742574, 1.60459, 
    2.053518, 3.685723, 11.00723, 23.7486, 17.17923, 5.668155, 2.557147, 
    1.49079, 1.198635, 1.050246, 0.7044977, 0.5246773, 0.4948629, 0.5576551, 
    0.5360993, 0.6968706, 4.613519, 24.34445, 14.60716, 3.13864, 1.492566, 
    1.823762,
  6.42875, 18.76912, 22.24078, 10.48147, 2.39456, 1.399178, 1.385494, 
    2.103833, 3.259803, 5.508416, 6.151264, 4.498104, 2.55251, 0.8679014, 
    0.4250869, 0.3454378, 0.4258737, 0.4351785, 0.6903651, 1.15543, 2.22402, 
    4.374835, 8.189422, 22.51671, 20.96322, 15.77774, 2.394017, 2.242861, 
    3.732141,
  19.80203, 32.26421, 35.91308, 13.2245, 3.709595, 2.341053, 2.332423, 
    2.671166, 7.345254, 9.90032, 3.678992, 2.427442, 1.180614, 0.424693, 
    0.3184368, 0.4016238, 0.551599, 0.825692, 1.31696, 2.487421, 4.900678, 
    9.350656, 17.4181, 23.21645, 18.49309, 5.835291, 5.826652, 9.36684, 
    15.27281,
  34.17523, 32.04915, 31.36699, 30.49985, 12.34155, 7.528187, 12.03026, 
    8.075918, 7.864016, 4.988306, 3.119113, 2.049792, 1.275753, 0.8274334, 
    0.5993829, 0.6558725, 0.81436, 1.148577, 1.608962, 2.399221, 3.649952, 
    5.213066, 6.597746, 9.905416, 3.187158, 4.337492, 8.597584, 20.32112, 
    33.73159,
  22.25683, 23.7877, 18.15446, 19.69978, 25.06741, 13.22767, 16.9684, 
    17.75799, 19.09029, 13.18487, 6.859272, 3.850619, 3.666955, 3.71783, 
    3.311999, 2.365121, 1.995238, 1.849338, 2.108473, 2.89715, 6.261796, 
    13.26826, 4.178957, 4.195512, 2.711157, 3.80386, 6.089437, 10.40413, 
    20.57803,
  18.14904, 16.09904, 13.69685, 21.28767, 22.73487, 23.15167, 29.13702, 
    20.77517, 31.49061, 27.86576, 14.10108, 10.06324, 7.809581, 6.326763, 
    5.589664, 4.558803, 3.413965, 2.669034, 2.741291, 4.165518, 12.15309, 
    16.76005, 10.97557, 7.020956, 4.589012, 3.858871, 3.5625, 5.014575, 
    14.95627,
  12.99197, 12.38115, 16.58363, 17.3449, 27.05569, 22.42281, 25.8613, 
    29.58266, 30.24482, 23.71635, 22.00528, 17.76134, 12.67977, 8.747373, 
    6.935437, 5.388694, 4.516201, 3.470422, 3.21847, 6.937133, 15.1522, 
    22.3233, 18.14536, 16.62381, 13.20255, 8.258942, 6.136657, 5.766225, 
    7.451026,
  8.039016, 11.79911, 14.15095, 16.05512, 19.01669, 20.37052, 18.368, 
    14.73614, 19.84023, 23.01449, 23.02519, 18.3945, 14.71878, 11.3931, 
    8.349963, 6.671067, 5.521569, 5.042399, 4.561929, 7.927204, 17.93193, 
    18.86878, 16.84904, 19.19691, 16.86593, 10.66466, 8.092819, 6.240869, 
    5.695092,
  7.831084, 10.19897, 13.30391, 14.01179, 14.95597, 15.57871, 16.18685, 
    18.04422, 18.06336, 16.12319, 17.15767, 14.72208, 11.43336, 9.476033, 
    8.608068, 7.172544, 7.103455, 7.425115, 8.068835, 13.81286, 14.66338, 
    12.70794, 11.25565, 13.06559, 12.17747, 8.999932, 6.901917, 6.273988, 
    6.411841,
  7.062912, 8.021914, 9.257833, 10.44017, 10.66504, 10.75985, 10.99366, 
    11.70968, 12.20951, 11.1093, 11.01311, 10.77439, 9.296811, 8.152157, 
    7.710881, 7.194204, 7.504001, 8.031941, 7.927028, 8.283611, 8.385488, 
    7.986227, 8.021174, 8.114985, 8.137836, 6.50913, 5.891754, 5.767591, 
    5.938109,
  5.884809, 6.058145, 6.462124, 7.154435, 7.620001, 8.074273, 8.092852, 
    8.173054, 8.165791, 7.986963, 7.648643, 7.490717, 7.288277, 6.906931, 
    6.627526, 6.142787, 5.953024, 5.988512, 5.883817, 5.507158, 5.50049, 
    5.958723, 6.328794, 6.808258, 7.037171, 6.618635, 6.323128, 6.342176, 
    6.106665,
  0.2990493, 0.2990493, 0.2990493, 0.2990493, 0.2990493, 0.2990493, 
    0.2990493, 0.2971749, 0.2971749, 0.2971749, 0.2971749, 0.2971749, 
    0.2971749, 0.2971749, 0.3113742, 0.3113742, 0.3113742, 0.3113742, 
    0.3113742, 0.3113742, 0.3113742, 0.3110233, 0.3110233, 0.3110233, 
    0.3110233, 0.3110233, 0.3110233, 0.3110233, 0.2990493,
  0.3825701, 0.354023, 0.3352614, 0.3331631, 0.2984086, 0.3010359, 0.3068528, 
    0.3011803, 0.2970305, 0.2920082, 0.2721946, 0.2493206, 0.2386916, 
    0.1771485, 0.1581355, 0.1644888, 0.1755156, 0.2064283, 0.2438451, 
    0.2958391, 0.3390072, 0.3767769, 0.387423, 0.3255202, 0.3619894, 
    0.3408173, 0.3108852, 0.3554581, 0.3819218,
  0.3656503, 0.2536117, 0.2557227, 0.2652448, 0.4013685, 0.3440868, 
    0.2017763, 0.3014389, 0.3017407, 0.2846109, 0.3149809, 0.3786195, 
    0.3465651, 0.3295949, 0.4647798, 0.5031633, 0.4628187, 0.4226803, 
    0.3678931, 0.3270571, 0.2765586, 0.316481, 0.3692326, 0.6206207, 
    0.7214739, 0.7702122, 0.7577399, 0.658246, 0.5255492,
  0.8944967, 0.7218501, 0.6522789, 0.6382866, 0.6866418, 0.5548621, 
    0.4517966, 0.3773546, 0.2969324, 0.2899988, 0.2904931, 0.4544898, 
    1.003552, 0.9588338, 0.9651436, 0.9833712, 0.8666608, 0.7069955, 
    0.6064271, 0.4758947, 0.372784, 0.3186247, 0.3617896, 0.5508676, 
    1.420447, 1.967524, 1.936546, 1.479757, 1.171214,
  1.480507, 1.174986, 1.130041, 1.352988, 1.194709, 1.089111, 0.8923802, 
    0.6119223, 0.4797904, 0.4308539, 0.5571089, 0.9915191, 1.908921, 
    2.175294, 2.133072, 1.622441, 1.179293, 1.018267, 0.8316183, 0.649109, 
    0.5407079, 0.4719338, 0.4482258, 1.466945, 4.850534, 3.784184, 3.081509, 
    2.343787, 1.849848,
  1.51111, 1.349176, 2.233587, 3.453643, 1.898038, 1.299959, 1.083916, 
    0.9082735, 0.7968531, 0.8510156, 2.304929, 3.356328, 7.124082, 4.307992, 
    3.413406, 1.985355, 1.302096, 1.005901, 0.7948411, 0.7663751, 0.7008489, 
    0.5943245, 0.6476589, 2.430688, 10.95503, 4.834943, 2.654318, 2.16365, 
    1.762995,
  1.294172, 2.981643, 18.0116, 7.587829, 3.081714, 1.772978, 1.288943, 
    1.20842, 1.067614, 5.245986, 15.76, 17.21394, 15.44567, 5.348175, 
    2.471733, 1.466038, 1.153015, 0.9584416, 0.7498757, 0.661429, 0.5687481, 
    0.5442173, 0.5374265, 3.968967, 20.47781, 9.159015, 2.947823, 1.470154, 
    1.184374,
  2.4868, 16.84328, 24.78878, 9.220135, 4.682009, 1.524686, 1.452211, 
    2.068917, 4.219191, 12.91142, 28.26579, 21.03305, 6.11842, 2.530603, 
    1.435164, 1.092863, 0.897174, 0.6350996, 0.4925435, 0.4511582, 0.5136086, 
    0.5288684, 0.6719244, 5.072219, 27.5482, 17.37659, 2.673561, 1.249219, 
    1.589492,
  5.877928, 20.11379, 25.43835, 12.19078, 2.20068, 1.317856, 1.41796, 
    2.332356, 4.029373, 6.822755, 7.938746, 4.883009, 2.696108, 0.842081, 
    0.4173524, 0.347813, 0.4149177, 0.4819202, 0.7860335, 1.346086, 2.398318, 
    4.00296, 6.777039, 25.50431, 24.47729, 17.80489, 2.267529, 2.11595, 
    3.32241,
  20.18858, 35.46019, 38.98978, 16.27707, 3.335058, 2.435157, 2.518137, 
    2.859231, 8.685114, 11.87876, 3.834611, 2.571417, 1.159223, 0.4155422, 
    0.3319809, 0.4448908, 0.6337553, 1.011396, 1.689632, 3.184367, 5.614921, 
    9.736381, 17.23756, 26.00025, 20.76244, 6.894566, 6.342106, 10.03281, 
    16.1947,
  38.34431, 35.43719, 32.77482, 32.07778, 13.61116, 8.1235, 13.77217, 
    8.897931, 9.358263, 5.648719, 3.572789, 2.290384, 1.412016, 0.8989564, 
    0.6275512, 0.6829064, 0.8721015, 1.254521, 1.755287, 2.660373, 4.236442, 
    6.235478, 7.174972, 11.77142, 3.293612, 4.539906, 9.220257, 21.96533, 
    38.68513,
  25.85565, 26.33642, 20.3201, 21.49055, 27.23074, 14.78788, 20.57626, 
    19.89351, 22.69788, 14.48823, 7.511169, 4.325292, 4.145705, 3.915152, 
    3.315957, 2.263101, 2.018477, 1.985073, 2.135602, 2.911337, 6.565655, 
    15.19202, 5.055014, 5.187411, 2.750202, 3.848535, 6.134109, 10.57619, 
    22.75213,
  21.31797, 19.00454, 16.63799, 24.68817, 25.21179, 26.22834, 31.88884, 
    23.21807, 33.95829, 30.33351, 14.813, 10.67719, 8.020176, 6.312846, 
    5.502434, 4.418649, 3.258846, 2.666816, 2.859369, 4.872088, 14.22378, 
    19.76894, 12.77841, 8.388692, 5.157394, 4.094907, 3.767609, 5.258105, 
    16.37041,
  15.19054, 14.14921, 19.39559, 20.20809, 30.31492, 25.39545, 28.61729, 
    32.79892, 33.92443, 27.59783, 25.68748, 20.61987, 13.84915, 9.22766, 
    7.118275, 5.405971, 4.559148, 3.492479, 3.333118, 8.986459, 17.26908, 
    26.0599, 22.08733, 20.31694, 15.00151, 8.974498, 6.510892, 6.211424, 
    8.70154,
  9.295711, 13.70506, 17.09926, 19.42832, 22.16, 23.53147, 21.6366, 16.82883, 
    23.04443, 26.64367, 27.35459, 21.61029, 16.5913, 12.43911, 8.88055, 
    7.118305, 5.803191, 5.397613, 4.942393, 9.23107, 21.69902, 22.88197, 
    20.2511, 22.83668, 19.47694, 12.03713, 8.683719, 6.622472, 6.365243,
  8.804612, 12.11683, 15.40809, 16.45987, 17.86456, 18.32682, 18.8956, 
    21.07412, 21.24582, 19.29679, 19.7531, 16.28632, 12.72463, 10.38854, 
    9.686273, 7.939917, 8.116419, 8.548525, 9.418964, 16.70202, 17.38174, 
    14.77178, 13.09761, 14.57527, 13.55283, 9.438924, 7.307325, 6.694681, 
    6.87514,
  7.429345, 8.7639, 10.16886, 11.48064, 12.09122, 12.17643, 12.46988, 
    13.6844, 13.98518, 12.54449, 12.33364, 12.33532, 10.30803, 8.994902, 
    8.535055, 8.00637, 8.650227, 9.418283, 9.344234, 9.758239, 9.409531, 
    8.81354, 8.668581, 8.644058, 8.561033, 6.72879, 6.065496, 5.854684, 
    6.161591,
  6.183407, 6.478043, 6.970573, 7.820632, 8.337979, 9.002526, 9.072468, 
    9.234627, 9.204309, 8.992249, 8.585729, 8.423381, 8.119756, 7.674732, 
    7.297405, 6.784788, 6.538764, 6.646362, 6.46863, 6.063922, 5.922051, 
    6.478015, 6.696134, 7.155434, 7.289748, 6.914669, 6.583482, 6.66081, 
    6.437249,
  0.2843398, 0.2843398, 0.2843398, 0.2843398, 0.2843398, 0.2843398, 
    0.2843398, 0.2861641, 0.2861641, 0.2861641, 0.2861641, 0.2861641, 
    0.2861641, 0.2861641, 0.2963867, 0.2963867, 0.2963867, 0.2963867, 
    0.2963867, 0.2963867, 0.2963867, 0.2989272, 0.2989272, 0.2989272, 
    0.2989272, 0.2989272, 0.2989272, 0.2989272, 0.2843398,
  0.363676, 0.3297343, 0.3174675, 0.3180227, 0.2747826, 0.2795744, 0.2857454, 
    0.282168, 0.2751657, 0.2673869, 0.250599, 0.2319114, 0.2220674, 
    0.1729754, 0.150125, 0.1549878, 0.1657069, 0.1881282, 0.2237448, 
    0.2747176, 0.3256456, 0.3639873, 0.3676159, 0.2843213, 0.3311221, 
    0.3258395, 0.2880622, 0.3364189, 0.369875,
  0.3231106, 0.223414, 0.2259121, 0.2358201, 0.3568701, 0.3010482, 0.182407, 
    0.2751589, 0.2845421, 0.2672542, 0.2990027, 0.3472113, 0.3141037, 
    0.2817432, 0.4109708, 0.4568604, 0.4189886, 0.3787999, 0.3389116, 
    0.3064405, 0.2593336, 0.2989667, 0.3850076, 0.6173314, 0.7033888, 
    0.7932942, 0.7546177, 0.6525851, 0.511556,
  0.8810792, 0.6862349, 0.6027118, 0.5868939, 0.6213807, 0.5073436, 
    0.4116665, 0.3420145, 0.2762339, 0.2674545, 0.271995, 0.4248824, 
    0.930819, 0.9294913, 0.9155474, 0.9400565, 0.8431318, 0.6600235, 
    0.5496988, 0.4270049, 0.3412397, 0.2905822, 0.3431478, 0.5617098, 
    1.634403, 2.189899, 1.955251, 1.443191, 1.152344,
  1.435008, 1.14886, 1.095082, 1.309136, 1.142863, 1.027092, 0.8198633, 
    0.5446299, 0.4358392, 0.3960707, 0.5203366, 0.9409563, 1.971276, 
    2.165886, 2.166947, 1.639305, 1.144685, 0.9653095, 0.7499828, 0.5927477, 
    0.4866289, 0.4270401, 0.4131572, 2.028345, 5.772911, 4.237988, 3.281641, 
    2.412915, 1.837259,
  1.44781, 1.324143, 2.411414, 3.23353, 1.665792, 1.150545, 0.9718634, 
    0.7955191, 0.7043514, 0.7896169, 2.312003, 3.469235, 7.881898, 4.392642, 
    4.07748, 2.05588, 1.220377, 0.9267258, 0.7308241, 0.6777779, 0.6444502, 
    0.5655961, 0.6464247, 3.42067, 12.53866, 5.009211, 2.639461, 2.176543, 
    1.695823,
  1.202739, 3.540309, 21.34131, 6.880089, 2.725516, 1.526064, 1.078001, 
    1.007111, 0.9842018, 6.457189, 18.12206, 20.20575, 17.38207, 5.233265, 
    2.290729, 1.363015, 1.037037, 0.860933, 0.657104, 0.5811583, 0.5095204, 
    0.4845533, 0.5251701, 5.133357, 22.83886, 9.606769, 2.613795, 1.319734, 
    1.122656,
  2.591202, 18.76666, 28.70206, 9.421081, 4.276315, 1.341519, 1.277386, 
    2.035877, 4.769808, 14.90575, 31.42006, 24.24593, 6.505034, 2.418469, 
    1.36144, 1.019494, 0.7674428, 0.585878, 0.4864149, 0.4210232, 0.4251962, 
    0.5055617, 0.6181068, 5.748434, 30.85908, 20.16369, 2.182087, 1.021083, 
    1.414371,
  5.43414, 21.30937, 28.86953, 13.26074, 2.021635, 1.298753, 1.436488, 
    2.503186, 4.634144, 7.936133, 9.461168, 5.255292, 2.834494, 0.8355262, 
    0.4189768, 0.3556581, 0.4160037, 0.5152364, 0.7899187, 1.324921, 
    2.381479, 3.139225, 5.401128, 29.10067, 28.23389, 20.04543, 2.084253, 
    1.887534, 2.93714,
  19.7466, 38.59562, 41.76822, 18.29058, 3.441077, 2.623247, 2.739788, 
    3.10834, 10.06112, 14.28786, 4.001438, 2.794432, 1.105728, 0.3996986, 
    0.3450851, 0.4771375, 0.6961549, 1.128594, 1.941727, 3.473515, 5.815841, 
    9.295584, 16.34498, 28.88361, 22.61824, 7.710786, 6.66355, 10.22763, 
    16.49062,
  41.14019, 38.75451, 33.78275, 33.04678, 14.79872, 8.890121, 15.05417, 
    9.37681, 11.07918, 6.095754, 3.921096, 2.489775, 1.577601, 1.016013, 
    0.6900475, 0.7263814, 0.9431343, 1.356071, 1.886482, 2.899346, 4.815918, 
    7.38012, 7.670706, 13.33527, 3.258578, 4.932137, 9.537843, 22.14848, 
    41.65372,
  30.60749, 29.62272, 22.85616, 23.34759, 29.32575, 16.9523, 24.22923, 
    22.22051, 26.73858, 15.77911, 7.975129, 4.64444, 4.257494, 3.884085, 
    3.139216, 2.188138, 2.085069, 2.23592, 2.344307, 3.032485, 6.953249, 
    17.08756, 6.190028, 5.809456, 2.814665, 3.782611, 6.126548, 11.04051, 
    26.45618,
  24.59972, 22.28807, 19.81108, 28.23923, 27.48706, 29.62587, 34.68635, 
    25.60027, 36.4097, 35.07773, 16.42525, 11.51982, 8.197167, 6.314696, 
    5.373242, 4.313176, 3.162079, 2.669553, 3.129423, 5.931499, 16.62624, 
    22.85231, 15.65795, 10.24256, 5.868859, 4.462021, 3.975688, 5.585057, 
    17.88615,
  17.51308, 16.4567, 22.89686, 23.26633, 33.65165, 29.26093, 31.56299, 
    36.1461, 37.9573, 32.20425, 30.20445, 23.42745, 15.04822, 9.687998, 
    7.394521, 5.431438, 4.618068, 3.590087, 3.468758, 11.20776, 19.68907, 
    30.40818, 27.36696, 25.2114, 16.69245, 9.723692, 6.92428, 6.583556, 
    10.41422,
  11.01931, 16.31708, 20.69535, 23.55502, 25.72029, 26.90325, 25.54778, 
    19.31544, 26.67495, 31.19834, 32.47297, 25.73658, 18.81787, 13.27951, 
    9.309443, 7.692425, 6.234173, 5.770047, 5.42693, 11.08304, 25.80123, 
    28.42566, 25.23914, 27.03861, 22.34942, 13.56424, 9.231513, 7.01663, 
    7.305234,
  9.921772, 14.30255, 17.9693, 19.79033, 21.60994, 22.31794, 22.66637, 
    24.74709, 25.57405, 23.78682, 23.86769, 18.32681, 14.31401, 11.83686, 
    10.96151, 8.971134, 9.482587, 9.84549, 11.19822, 20.01926, 20.64291, 
    17.63213, 15.15003, 16.54568, 15.02429, 9.788063, 7.67285, 7.16388, 
    7.424049,
  7.750371, 9.564883, 11.38895, 13.00028, 13.82789, 13.93916, 14.25915, 
    16.20633, 16.22078, 14.32853, 14.24714, 14.36405, 11.51004, 10.18824, 
    9.679282, 9.113441, 10.1294, 11.06029, 11.13201, 11.65605, 10.44695, 
    9.878273, 9.736784, 9.231435, 9.080626, 6.960367, 6.236952, 5.867185, 
    6.402864,
  6.495965, 6.939672, 7.43204, 8.441461, 9.136636, 10.00921, 10.29299, 
    10.53886, 10.58307, 10.34356, 10.00446, 9.729712, 9.170202, 8.61409, 
    7.980806, 7.445165, 7.255861, 7.30532, 7.07376, 6.70609, 6.380611, 6.91, 
    7.086012, 7.458575, 7.447979, 7.133189, 6.817133, 6.934138, 6.756274,
  0.2687275, 0.2687275, 0.2687275, 0.2687275, 0.2687275, 0.2687275, 
    0.2687275, 0.2754089, 0.2754089, 0.2754089, 0.2754089, 0.2754089, 
    0.2754089, 0.2754089, 0.2845536, 0.2845536, 0.2845536, 0.2845536, 
    0.2845536, 0.2845536, 0.2845536, 0.2856445, 0.2856445, 0.2856445, 
    0.2856445, 0.2856445, 0.2856445, 0.2856445, 0.2687275,
  0.3479453, 0.3093624, 0.3011045, 0.3039462, 0.2562994, 0.260901, 0.2660033, 
    0.2631235, 0.2554973, 0.247283, 0.2337672, 0.2182372, 0.2094817, 
    0.172107, 0.1450515, 0.146036, 0.1566134, 0.1737535, 0.2090131, 
    0.2582762, 0.3147454, 0.3525748, 0.3452002, 0.2345979, 0.2912801, 
    0.3082741, 0.2669687, 0.3204782, 0.3602282,
  0.2876714, 0.1987722, 0.1997417, 0.213966, 0.3175634, 0.2621026, 0.1690124, 
    0.254731, 0.2663315, 0.2494681, 0.2824357, 0.3157665, 0.2853966, 
    0.2457648, 0.3619657, 0.4213515, 0.3828472, 0.3384673, 0.310992, 
    0.2836064, 0.2451782, 0.2814873, 0.4039566, 0.5980667, 0.678642, 
    0.8174949, 0.7536567, 0.6534032, 0.4857502,
  0.8518418, 0.6573772, 0.5563975, 0.5345141, 0.5624182, 0.4619969, 
    0.3766563, 0.3130571, 0.2586974, 0.2485677, 0.2536921, 0.394994, 
    0.8488244, 0.9032817, 0.864994, 0.9001041, 0.797565, 0.622815, 0.4940907, 
    0.3847333, 0.3129373, 0.2698056, 0.3433288, 0.588424, 1.94591, 2.389619, 
    1.97019, 1.40958, 1.137544,
  1.41487, 1.111054, 1.042458, 1.235359, 1.074929, 0.9701834, 0.7423533, 
    0.4976695, 0.3969902, 0.3672568, 0.4816322, 0.8898536, 2.010664, 
    2.118959, 2.246004, 1.63872, 1.112546, 0.9080339, 0.6957475, 0.5385507, 
    0.4480202, 0.3959748, 0.3872613, 2.935012, 6.643823, 4.762277, 3.428838, 
    2.46757, 1.81263,
  1.368598, 1.291002, 2.617868, 3.00006, 1.481193, 1.013299, 0.8552387, 
    0.696519, 0.627158, 0.7411468, 2.304153, 3.67549, 8.626563, 4.407376, 
    4.958845, 2.118927, 1.169379, 0.8690842, 0.6931748, 0.6150893, 0.5766585, 
    0.5554669, 0.6872588, 4.827305, 14.3672, 5.049482, 2.709871, 2.161219, 
    1.618916,
  1.14134, 4.276403, 24.87384, 6.085731, 2.308145, 1.289638, 0.8898614, 
    0.8088861, 0.9626297, 7.657077, 20.73699, 22.99523, 19.25747, 4.903491, 
    2.144292, 1.311522, 0.9673856, 0.7960009, 0.588094, 0.5243694, 0.4601173, 
    0.4457464, 0.5288464, 7.136859, 25.67422, 9.840184, 2.307389, 1.198478, 
    1.059357,
  2.763466, 20.71124, 31.90475, 9.382594, 3.767755, 1.184198, 1.141957, 
    1.918334, 5.105091, 16.61927, 33.75927, 26.75241, 6.504213, 2.25736, 
    1.30432, 0.9047952, 0.6497427, 0.5315772, 0.4551353, 0.3839243, 
    0.3791175, 0.452397, 0.6531561, 6.297855, 34.46746, 23.15367, 1.801219, 
    0.901469, 1.301822,
  5.08613, 22.15813, 31.98842, 14.02282, 1.888524, 1.279181, 1.443254, 
    2.667555, 5.044423, 8.731775, 10.65352, 5.512383, 2.962222, 0.8357103, 
    0.425798, 0.3653543, 0.4240624, 0.5442702, 0.7663411, 1.077448, 1.767047, 
    2.143524, 4.096879, 32.76171, 31.332, 22.2331, 1.895152, 1.582999, 
    2.568171,
  18.85352, 42.05167, 44.61063, 19.52223, 3.590635, 2.956293, 3.080556, 
    3.382021, 11.49322, 16.82398, 4.149704, 3.080608, 1.035713, 0.3843222, 
    0.3560222, 0.5000356, 0.7402034, 1.183954, 1.976215, 3.270911, 5.434183, 
    8.514749, 14.82246, 31.81113, 24.25986, 8.336017, 6.82572, 10.03132, 
    15.58742,
  42.8835, 41.56568, 35.46364, 33.64735, 16.2248, 9.788512, 15.84804, 
    9.964705, 13.12737, 6.440232, 4.257641, 2.615225, 1.683738, 1.090493, 
    0.7481893, 0.7951223, 1.024348, 1.462103, 2.001922, 3.111388, 5.353076, 
    8.58357, 8.04726, 14.45034, 3.177261, 4.999735, 9.318697, 21.4506, 
    43.45099,
  35.79327, 34.01204, 26.76542, 25.03722, 31.60429, 19.83449, 27.96959, 
    25.12712, 31.26694, 17.58761, 8.288644, 4.748306, 4.148841, 3.646394, 
    2.944316, 2.178144, 2.177906, 2.393817, 2.880906, 3.585065, 7.828329, 
    18.84622, 7.556993, 6.21163, 2.802126, 3.69354, 6.130964, 12.77506, 
    32.37706,
  27.82725, 25.90248, 23.10047, 31.52121, 29.72894, 33.4449, 37.96108, 
    28.02401, 38.75617, 40.70332, 19.37613, 12.47692, 8.39743, 6.314065, 
    5.327087, 4.279474, 3.181785, 2.749575, 3.506315, 7.387977, 19.4064, 
    26.16796, 19.78828, 11.87619, 6.541607, 4.843598, 4.150869, 6.020236, 
    19.83472,
  19.8543, 19.30888, 26.70615, 26.29173, 37.39678, 33.48264, 34.8728, 
    39.81469, 42.56393, 37.27365, 35.31606, 25.94982, 16.16221, 10.19027, 
    7.672401, 5.579011, 4.701001, 3.716818, 3.613341, 13.66917, 22.57807, 
    35.79047, 33.85115, 31.02125, 18.41674, 10.53032, 7.313816, 6.854661, 
    12.48337,
  13.19627, 19.74742, 25.06448, 28.11891, 30.03303, 30.76165, 30.41832, 
    22.1956, 30.56443, 36.66918, 39.07541, 30.97594, 21.61699, 14.10165, 
    9.729695, 8.217316, 6.994309, 6.318615, 6.273479, 13.68885, 30.31472, 
    35.18689, 31.76508, 32.22545, 25.92709, 15.27916, 9.765356, 7.399515, 
    8.722329,
  11.1712, 16.42697, 21.30842, 24.27605, 26.49331, 27.28054, 27.57357, 
    29.90257, 30.86144, 29.28509, 29.30891, 21.10403, 16.10117, 13.83587, 
    12.71436, 10.11371, 11.12614, 11.52436, 13.74578, 23.95716, 24.89047, 
    21.24921, 17.38337, 19.06363, 16.78047, 10.02734, 8.03503, 7.503171, 
    7.91543,
  7.92724, 10.16975, 12.71049, 14.96153, 15.91736, 16.34086, 16.85816, 
    19.44331, 18.74605, 16.40553, 16.69157, 16.77881, 13.12526, 11.92872, 
    11.39362, 10.5151, 11.83173, 12.92796, 12.8889, 13.53045, 11.53859, 
    11.37149, 11.05609, 9.873787, 9.582034, 7.188984, 6.379082, 5.81023, 
    6.609983,
  6.757342, 7.319344, 7.888938, 9.068604, 9.929606, 11.12249, 11.61886, 
    12.13894, 12.28209, 12.12003, 11.74951, 11.10231, 10.34798, 9.594935, 
    8.822229, 8.216036, 8.009921, 8.037846, 7.802186, 7.519916, 6.983832, 
    7.416598, 7.456749, 7.654363, 7.477963, 7.249768, 7.014091, 7.067791, 
    6.953017,
  0.2555091, 0.2555091, 0.2555091, 0.2555091, 0.2555091, 0.2555091, 
    0.2555091, 0.2621664, 0.2621664, 0.2621664, 0.2621664, 0.2621664, 
    0.2621664, 0.2621664, 0.2736266, 0.2736266, 0.2736266, 0.2736266, 
    0.2736266, 0.2736266, 0.2736266, 0.2721828, 0.2721828, 0.2721828, 
    0.2721828, 0.2721828, 0.2721828, 0.2721828, 0.2555091,
  0.3332098, 0.2909473, 0.2868015, 0.2899759, 0.242202, 0.2451533, 0.2476065, 
    0.2450356, 0.2387917, 0.2315809, 0.2214003, 0.2065923, 0.1998931, 
    0.1727896, 0.1421203, 0.1379069, 0.1469377, 0.1616628, 0.1982282, 
    0.247664, 0.3061936, 0.3413741, 0.3213387, 0.1977027, 0.2429286, 
    0.2828912, 0.2497413, 0.3084668, 0.3507191,
  0.2576542, 0.181776, 0.1825655, 0.1987673, 0.2848707, 0.2299245, 0.1609614, 
    0.2379207, 0.2461116, 0.2312427, 0.2630936, 0.2878277, 0.2604485, 
    0.2207106, 0.3190266, 0.3822934, 0.3448559, 0.3067397, 0.2849994, 
    0.2648847, 0.2318019, 0.2638715, 0.4139797, 0.5823188, 0.6549275, 
    0.828566, 0.7621222, 0.650187, 0.4527743,
  0.8156695, 0.6349842, 0.5153666, 0.5024285, 0.5167669, 0.4248594, 
    0.3490572, 0.2887028, 0.2408271, 0.2318384, 0.2404332, 0.3691703, 
    0.7769674, 0.857356, 0.8275741, 0.8620675, 0.7453287, 0.5821254, 
    0.4468713, 0.3530559, 0.2845674, 0.257127, 0.3582637, 0.6499015, 2.29835, 
    2.574073, 1.963594, 1.368544, 1.10879,
  1.404398, 1.064858, 0.9951029, 1.162354, 1.003628, 0.9076484, 0.6719416, 
    0.4613456, 0.3722944, 0.3446777, 0.4512075, 0.8160525, 1.986641, 
    2.101165, 2.29795, 1.63362, 1.091587, 0.8684328, 0.6604029, 0.5031974, 
    0.4180173, 0.3733076, 0.369869, 4.324761, 7.556637, 5.274325, 3.554323, 
    2.508214, 1.804048,
  1.284918, 1.259773, 2.747526, 2.705317, 1.299292, 0.8931254, 0.7313226, 
    0.6054085, 0.5639638, 0.7047538, 2.295476, 3.961341, 9.230262, 4.383079, 
    5.97435, 2.14451, 1.12982, 0.8284443, 0.6617109, 0.5678599, 0.5241535, 
    0.5513767, 0.7640932, 6.65885, 16.4084, 5.061016, 2.712382, 2.101345, 
    1.546027,
  1.120664, 4.947349, 28.06816, 5.312283, 1.928401, 1.075724, 0.7712404, 
    0.6568611, 0.9510142, 8.833773, 22.70903, 25.08, 20.84095, 4.531604, 
    2.08259, 1.27746, 0.9325497, 0.7420626, 0.5502962, 0.4899655, 0.4275382, 
    0.429282, 0.5628517, 9.971706, 29.42046, 9.765859, 2.056707, 1.138204, 
    1.048471,
  2.839825, 22.73735, 34.39952, 9.261024, 3.228284, 1.057912, 1.011396, 
    1.773245, 5.19054, 17.65404, 35.22852, 28.53794, 6.073923, 2.155481, 
    1.268661, 0.8333306, 0.6263855, 0.5079481, 0.4434846, 0.3733123, 
    0.3692653, 0.428715, 0.7571179, 6.599907, 38.2128, 26.24142, 1.5514, 
    0.8345939, 1.179774,
  4.693958, 22.59717, 34.62894, 14.70605, 1.804388, 1.268997, 1.454784, 
    2.801694, 5.360919, 9.436922, 11.81265, 5.715101, 3.103755, 0.8296898, 
    0.4390494, 0.37666, 0.4371001, 0.5631105, 0.736655, 0.8890523, 1.129057, 
    1.413913, 3.122509, 37.32267, 34.32925, 24.34112, 1.762505, 1.415433, 
    2.40286,
  17.66986, 44.41589, 46.67401, 20.44996, 3.733689, 3.32953, 3.571985, 
    3.651301, 12.89833, 19.4743, 4.351407, 3.349386, 0.9634926, 0.3717136, 
    0.3639968, 0.513459, 0.7671538, 1.217767, 1.956089, 3.029936, 4.542068, 
    7.461402, 13.1628, 34.41151, 25.78381, 8.746934, 7.027672, 9.77346, 
    14.27948,
  44.15864, 43.47303, 38.96325, 34.12915, 17.52991, 10.6336, 16.32077, 
    10.7563, 15.68706, 6.783856, 4.613023, 2.736865, 1.779392, 1.156224, 
    0.7920964, 0.8604506, 1.104472, 1.562549, 2.109267, 3.311422, 5.832511, 
    9.748972, 8.323095, 15.44559, 3.126047, 4.869083, 9.279019, 20.76792, 
    44.51447,
  39.85163, 39.31818, 31.81919, 26.35634, 35.13963, 22.62103, 31.20715, 
    30.25289, 35.20369, 20.39842, 8.510159, 4.901515, 4.134681, 3.607025, 
    2.917708, 2.241441, 2.324135, 2.53838, 3.497522, 5.094298, 9.506528, 
    20.45775, 8.91952, 6.353048, 2.867544, 3.663118, 6.295133, 14.47286, 
    38.13097,
  31.21271, 29.53498, 25.85627, 34.36658, 32.18757, 37.61874, 41.4231, 
    30.49337, 41.14282, 46.79691, 21.27167, 13.23505, 8.5252, 6.386826, 
    5.370107, 4.301341, 3.214222, 2.827227, 3.934952, 9.304761, 22.42983, 
    29.45852, 24.78481, 12.51775, 6.92691, 5.101887, 4.30833, 6.48616, 
    22.23276,
  22.17645, 22.25251, 30.37139, 29.39584, 41.46554, 38.82522, 38.28992, 
    43.98185, 47.57669, 42.65413, 40.60368, 27.87266, 17.00153, 10.51686, 
    7.775785, 5.804147, 4.73781, 3.819511, 3.811823, 16.31043, 25.8193, 
    41.46323, 40.8582, 36.87252, 20.20727, 11.15561, 7.560823, 7.063392, 
    14.67454,
  15.7006, 23.50718, 30.43958, 33.16998, 35.04547, 35.38855, 35.9565, 
    25.29665, 34.79008, 43.14539, 46.32125, 37.35803, 24.13138, 14.7063, 
    10.30468, 8.59783, 7.472197, 6.839998, 7.15629, 16.67833, 35.2842, 
    42.51002, 38.44846, 37.79896, 30.15084, 16.88906, 10.18314, 7.670363, 
    10.22917,
  12.29358, 18.68296, 25.16866, 29.76369, 32.3349, 33.09345, 33.37443, 
    36.43488, 36.73749, 35.81429, 34.80353, 24.66342, 18.34753, 16.2834, 
    14.98426, 11.46917, 13.01492, 13.44494, 16.82639, 28.34237, 30.60524, 
    25.61109, 20.40005, 22.07027, 18.80411, 10.14397, 8.336499, 7.785648, 
    8.454614,
  7.912992, 10.75924, 13.88052, 17.07657, 18.5695, 19.36699, 20.22735, 
    23.71262, 21.79493, 18.90563, 19.65562, 19.70669, 15.26488, 14.45134, 
    13.59613, 12.03508, 13.75038, 14.99531, 14.93289, 15.72297, 12.85895, 
    13.00091, 12.36562, 10.69145, 9.984112, 7.342838, 6.48902, 5.732481, 
    6.720255,
  6.983796, 7.697377, 8.421252, 9.728044, 10.79689, 12.3454, 12.97057, 
    13.75862, 14.04776, 13.99587, 13.59803, 12.61022, 11.75851, 10.86075, 
    9.85208, 9.145173, 8.940885, 8.933352, 8.717065, 8.389482, 7.712662, 
    7.921227, 7.761354, 7.750506, 7.424536, 7.257544, 7.128934, 7.017962, 
    7.112415,
  0.2406541, 0.2406541, 0.2406541, 0.2406541, 0.2406541, 0.2406541, 
    0.2406541, 0.2487088, 0.2487088, 0.2487088, 0.2487088, 0.2487088, 
    0.2487088, 0.2487088, 0.2609453, 0.2609453, 0.2609453, 0.2609453, 
    0.2609453, 0.2609453, 0.2609453, 0.2547974, 0.2547974, 0.2547974, 
    0.2547974, 0.2547974, 0.2547974, 0.2547974, 0.2406541,
  0.3152442, 0.2749273, 0.2749184, 0.2784969, 0.2313534, 0.2316616, 
    0.2312679, 0.2287757, 0.2240928, 0.2179321, 0.2104342, 0.1976401, 
    0.1931963, 0.1739921, 0.1404116, 0.1316987, 0.1385211, 0.1528425, 
    0.1903075, 0.2398342, 0.2953101, 0.3302951, 0.2949161, 0.1841697, 
    0.2137241, 0.2527169, 0.2372937, 0.2989912, 0.3361188,
  0.2336108, 0.1721284, 0.1724055, 0.1889929, 0.2590373, 0.2056679, 
    0.1574798, 0.2242652, 0.2259023, 0.2147702, 0.2445718, 0.2624925, 
    0.2397024, 0.2021618, 0.2832258, 0.3437741, 0.3127106, 0.2747032, 
    0.2634161, 0.2448565, 0.2190577, 0.2498578, 0.4223393, 0.5651522, 
    0.633326, 0.8417046, 0.7659869, 0.6444019, 0.4131697,
  0.7879763, 0.6110783, 0.4820262, 0.4808373, 0.4833869, 0.3959151, 
    0.3269384, 0.2699987, 0.2233608, 0.2167949, 0.224575, 0.3418054, 
    0.7019718, 0.8073213, 0.7943768, 0.8180402, 0.6891295, 0.5452574, 
    0.4084206, 0.3255129, 0.2705944, 0.2480586, 0.3650125, 0.7318103, 
    2.647163, 2.723922, 1.958084, 1.300871, 1.068461,
  1.37141, 1.031995, 0.955687, 1.092464, 0.9441747, 0.8474289, 0.6114483, 
    0.4362102, 0.3571222, 0.3312094, 0.4252899, 0.7492974, 1.953853, 
    2.063613, 2.373294, 1.635647, 1.080691, 0.8367375, 0.6245356, 0.4742435, 
    0.3958354, 0.3548836, 0.3571841, 6.184701, 8.602274, 5.691222, 3.655237, 
    2.499898, 1.793686,
  1.201945, 1.182971, 2.803708, 2.429783, 1.140102, 0.7982652, 0.6533562, 
    0.5513501, 0.5261596, 0.6780486, 2.199124, 4.202044, 9.726505, 4.279876, 
    7.156804, 2.13512, 1.094127, 0.8013155, 0.6367949, 0.5391038, 0.4947426, 
    0.556627, 0.8278857, 9.080991, 18.44654, 5.065032, 2.679878, 2.021101, 
    1.498616,
  1.110152, 5.353672, 30.8152, 4.667676, 1.645221, 0.9660497, 0.7038665, 
    0.5836928, 0.9269657, 9.772548, 24.45147, 26.73391, 22.25801, 4.098508, 
    2.018789, 1.255542, 0.9186657, 0.7171113, 0.5401067, 0.4703636, 
    0.4174033, 0.4313459, 0.5764383, 13.44651, 33.6523, 9.458438, 1.920344, 
    1.09203, 1.026906,
  2.792313, 25.27164, 36.52031, 9.22397, 2.780669, 0.9686337, 0.9494882, 
    1.684564, 5.114912, 18.51036, 36.50622, 29.8712, 5.539056, 2.066261, 
    1.27592, 0.8079693, 0.6194535, 0.512156, 0.439864, 0.3694658, 0.3654271, 
    0.4147994, 0.851321, 6.780877, 42.38766, 29.27513, 1.401328, 0.7897366, 
    1.110419,
  4.611792, 22.85933, 36.4763, 15.45014, 1.743538, 1.260311, 1.466661, 
    2.913417, 5.682425, 9.993044, 12.4885, 5.999394, 3.279755, 0.8220256, 
    0.4451985, 0.3868598, 0.449222, 0.567246, 0.6996185, 0.7774609, 
    0.7980633, 0.9319016, 2.585043, 41.02449, 36.45627, 26.02828, 1.660148, 
    1.314506, 2.335785,
  15.77576, 45.09292, 47.16542, 21.64048, 3.876715, 3.655979, 4.036498, 
    3.970913, 14.08969, 21.58933, 4.640563, 3.678928, 0.9313592, 0.3642681, 
    0.3683051, 0.5201839, 0.7829519, 1.232319, 1.913215, 2.855775, 3.927823, 
    5.840368, 11.61758, 36.26664, 26.99056, 9.025648, 7.177109, 9.440448, 
    12.49503,
  45.26125, 45.11354, 41.78677, 34.5613, 18.68433, 11.56771, 16.92014, 
    11.36145, 18.29474, 7.122463, 5.018014, 2.887063, 1.895087, 1.239213, 
    0.845256, 0.9125754, 1.177417, 1.6478, 2.200679, 3.490748, 6.242664, 
    10.94479, 8.527595, 16.37865, 3.082811, 4.865874, 8.96294, 20.40565, 
    45.46419,
  42.70404, 43.93698, 37.39948, 27.21728, 38.21938, 23.49604, 33.61959, 
    35.30167, 38.64563, 23.58579, 8.772184, 5.058591, 4.205277, 3.663695, 
    2.969243, 2.334264, 2.495073, 2.674211, 4.010714, 6.829283, 11.3508, 
    22.06664, 9.749897, 6.446459, 2.945104, 3.67765, 6.364323, 15.04451, 
    41.94544,
  34.88103, 32.95064, 28.22223, 36.7893, 34.81575, 41.79934, 44.97136, 
    32.92364, 43.72127, 52.90019, 22.1633, 13.51058, 8.703155, 6.480554, 
    5.393868, 4.320969, 3.274886, 2.942801, 4.367424, 11.46318, 25.78026, 
    32.62109, 29.08237, 12.77303, 7.120324, 5.242965, 4.456874, 6.729471, 
    24.90104,
  24.59532, 24.38208, 33.71397, 32.5671, 45.76873, 45.54496, 41.67558, 
    49.34583, 53.09797, 48.07786, 45.12975, 29.06492, 17.35346, 10.62291, 
    7.815907, 5.938464, 4.724005, 3.975065, 3.970688, 19.39363, 29.29253, 
    46.86195, 47.76657, 42.14864, 21.18077, 11.60911, 7.776028, 7.168334, 
    16.73268,
  18.95437, 28.15601, 36.16409, 39.33776, 41.75703, 41.98747, 42.97971, 
    28.84192, 39.48494, 50.03738, 54.22924, 44.66062, 25.634, 15.04091, 
    10.58761, 8.802453, 7.864009, 7.230102, 7.927874, 20.02436, 40.25793, 
    50.48598, 45.44022, 43.59793, 34.37114, 17.82649, 10.40957, 7.856347, 
    11.66665,
  13.23457, 21.23746, 29.33388, 35.95981, 38.66679, 39.22611, 40.11907, 
    44.13675, 43.65362, 43.04144, 41.18779, 29.03333, 20.92114, 19.13235, 
    17.67627, 12.87235, 15.48308, 15.58062, 20.66952, 33.06432, 36.75272, 
    31.33673, 24.26183, 25.64058, 20.93239, 10.17377, 8.535556, 7.951367, 
    8.939139,
  7.81625, 11.18758, 14.98651, 18.97418, 21.27134, 22.48368, 23.93791, 
    28.81874, 25.68627, 21.68051, 23.33186, 23.13567, 17.94429, 17.78999, 
    16.40158, 13.904, 16.0628, 17.18924, 17.23397, 18.50687, 14.79468, 
    14.90706, 13.67148, 11.58791, 10.34012, 7.396251, 6.541937, 5.649925, 
    6.693912,
  7.137356, 8.037487, 8.989552, 10.42834, 11.80638, 13.66231, 14.51941, 
    15.63913, 15.95418, 15.86079, 15.31169, 14.17818, 13.19746, 12.16042, 
    10.9276, 10.13345, 9.9278, 9.958167, 9.800444, 9.338352, 8.421479, 
    8.365955, 7.961207, 7.771192, 7.340245, 7.209704, 7.152281, 6.877131, 
    7.204244,
  0.2266015, 0.2266015, 0.2266015, 0.2266015, 0.2266015, 0.2266015, 
    0.2266015, 0.2338538, 0.2338538, 0.2338538, 0.2338538, 0.2338538, 
    0.2338538, 0.2338538, 0.2457233, 0.2457233, 0.2457233, 0.2457233, 
    0.2457233, 0.2457233, 0.2457233, 0.2350092, 0.2350092, 0.2350092, 
    0.2350092, 0.2350092, 0.2350092, 0.2350092, 0.2266015,
  0.2942939, 0.2590224, 0.2593313, 0.2647382, 0.2221366, 0.2207597, 
    0.2182656, 0.2149413, 0.2105658, 0.2053609, 0.2008042, 0.1917366, 
    0.1882525, 0.1753933, 0.1396763, 0.1290338, 0.1316793, 0.1467994, 
    0.1839653, 0.2303774, 0.2839442, 0.3197635, 0.2692691, 0.1828515, 
    0.199644, 0.2277151, 0.2287359, 0.2892972, 0.314227,
  0.2166543, 0.1673619, 0.1669387, 0.1843538, 0.2388967, 0.1885775, 
    0.1573867, 0.2133105, 0.2074421, 0.2013936, 0.2285277, 0.2385962, 
    0.2226438, 0.1893539, 0.2551593, 0.3120398, 0.2884859, 0.2522981, 
    0.2453857, 0.227032, 0.2101335, 0.241933, 0.4298913, 0.544476, 0.6122949, 
    0.8255862, 0.7644207, 0.6310945, 0.3648591,
  0.7565339, 0.587281, 0.4550153, 0.4635709, 0.4558422, 0.3831306, 0.3139653, 
    0.2561671, 0.2105167, 0.2058155, 0.212854, 0.3169695, 0.6368816, 
    0.7476831, 0.7517293, 0.7819054, 0.6597085, 0.5093775, 0.3827181, 
    0.3095843, 0.2615388, 0.2429174, 0.3708766, 0.8409622, 2.980339, 
    2.781775, 1.95478, 1.230006, 1.005873,
  1.323371, 1.009927, 0.9219798, 1.040261, 0.8937065, 0.7878225, 0.5660625, 
    0.4216118, 0.3496276, 0.3236803, 0.4057295, 0.6958906, 1.934378, 
    2.021839, 2.459384, 1.64939, 1.071645, 0.8104174, 0.5989395, 0.4545611, 
    0.3829457, 0.3443579, 0.3571723, 8.384976, 9.695794, 6.004473, 3.608607, 
    2.459139, 1.776353,
  1.154799, 1.129216, 2.799378, 2.194623, 1.034491, 0.736441, 0.6143628, 
    0.5256384, 0.5033202, 0.6667122, 2.082507, 4.326686, 10.03811, 4.142851, 
    8.480131, 2.118382, 1.067472, 0.7890128, 0.6191257, 0.5195956, 0.4815067, 
    0.5561917, 0.8861129, 11.82994, 20.36097, 4.999855, 2.626222, 1.953635, 
    1.463578,
  1.085427, 5.493469, 32.94056, 4.221551, 1.4794, 0.8912227, 0.6697752, 
    0.5526655, 0.907894, 10.31259, 26.10748, 28.42219, 23.76384, 3.813558, 
    1.968834, 1.241055, 0.906076, 0.707232, 0.5356287, 0.4638508, 0.4143825, 
    0.4278885, 0.5701579, 17.4282, 37.46937, 9.073395, 1.81756, 1.069671, 
    1.014627,
  2.663268, 28.24445, 38.52528, 9.229617, 2.517752, 0.9298616, 0.921799, 
    1.628027, 5.013583, 19.44479, 37.94589, 31.14793, 5.276794, 2.046558, 
    1.295115, 0.8037074, 0.6212416, 0.5153877, 0.4361453, 0.3668096, 
    0.3592893, 0.4104355, 0.923547, 7.407237, 45.70504, 31.79953, 1.320019, 
    0.7662137, 1.089209,
  4.759985, 23.06463, 37.90148, 16.63243, 1.722279, 1.259841, 1.468505, 
    2.969314, 5.893988, 10.33739, 12.73953, 6.30401, 3.513716, 0.8222026, 
    0.4540763, 0.3941346, 0.455264, 0.5628431, 0.6599459, 0.689079, 
    0.6636467, 0.7306214, 2.22665, 42.47094, 37.35363, 27.44389, 1.618387, 
    1.247338, 2.282561,
  14.65849, 44.64545, 46.54307, 23.03556, 3.978271, 3.822756, 4.295541, 
    4.190718, 14.59461, 22.61761, 4.876502, 3.803984, 0.9282818, 0.3623472, 
    0.3691901, 0.52198, 0.785924, 1.228039, 1.855285, 2.707646, 3.531593, 
    4.510461, 9.677018, 37.08067, 27.96339, 9.007564, 7.254722, 9.141612, 
    11.47964,
  46.06445, 46.5294, 43.74965, 35.16559, 19.67435, 11.72973, 17.65917, 
    11.57395, 20.35664, 7.471319, 5.389327, 3.012612, 1.967965, 1.302659, 
    0.8833761, 0.9529556, 1.222996, 1.712849, 2.266773, 3.625734, 6.573338, 
    11.95208, 8.88249, 17.28155, 3.029157, 4.769705, 8.651968, 20.57189, 
    46.15695,
  44.9274, 47.03259, 41.89862, 27.95202, 40.17459, 22.96036, 35.52294, 
    37.82108, 41.72372, 25.74968, 8.954253, 5.174289, 4.241837, 3.70428, 
    3.014185, 2.40635, 2.587631, 2.75642, 4.189323, 7.985758, 12.68044, 
    23.58759, 10.13976, 6.755657, 2.951254, 3.612915, 6.206734, 14.8348, 
    44.47807,
  38.71736, 35.64634, 30.22731, 38.90229, 37.32778, 45.53873, 48.54768, 
    35.42207, 46.43203, 58.16311, 22.60768, 13.66908, 8.801521, 6.562729, 
    5.430595, 4.344669, 3.333298, 2.996655, 4.656348, 13.56293, 29.03911, 
    35.53107, 32.22464, 12.76546, 7.203958, 5.29784, 4.51502, 6.658809, 
    27.45471,
  26.86596, 25.59284, 36.70307, 35.83273, 50.50413, 53.08842, 44.90922, 
    55.43269, 58.79503, 53.03225, 49.00933, 29.83819, 17.43068, 10.6451, 
    7.841006, 5.98493, 4.722697, 4.075233, 4.079265, 22.80876, 32.93505, 
    51.59288, 53.50788, 45.35264, 21.57551, 11.74029, 7.865088, 7.237274, 
    18.63917,
  22.34307, 33.77787, 42.73988, 47.02584, 50.0713, 51.00076, 50.06722, 
    32.47762, 44.42091, 57.25926, 63.43726, 52.58194, 26.29333, 15.2568, 
    10.78118, 8.895558, 8.050209, 7.554502, 8.525399, 24.01155, 45.89151, 
    57.61418, 52.54882, 49.67369, 38.74896, 18.36773, 10.43626, 7.907604, 
    12.56011,
  13.91591, 24.11717, 33.95396, 42.79527, 45.26741, 45.61855, 47.63085, 
    53.3106, 51.10802, 51.43363, 49.34699, 34.17583, 23.76194, 22.6583, 
    19.52681, 14.16817, 18.56748, 17.98029, 25.04168, 37.83854, 44.07181, 
    37.34154, 27.64768, 29.48845, 22.30828, 10.19172, 8.641829, 8.013843, 
    9.289974,
  7.777571, 11.48786, 16.02697, 20.8125, 23.75225, 25.65305, 28.32633, 
    34.95976, 29.98731, 24.84573, 27.81907, 26.93987, 21.39478, 21.44866, 
    19.64598, 15.59365, 18.01782, 19.70613, 20.02184, 21.76837, 17.1351, 
    17.13493, 15.1611, 12.66395, 10.62456, 7.377668, 6.53191, 5.553197, 
    6.62282,
  7.262084, 8.368874, 9.655175, 11.16686, 12.84065, 15.057, 16.33612, 
    17.54413, 17.9068, 17.65327, 17.10889, 15.95687, 14.78685, 13.52915, 
    12.23675, 11.12766, 10.83533, 10.92738, 10.82649, 10.25439, 9.174309, 
    8.708855, 8.001207, 7.743292, 7.22006, 7.121406, 7.103294, 6.671535, 
    7.051307,
  0.2121684, 0.2121684, 0.2121684, 0.2121684, 0.2121684, 0.2121684, 
    0.2121684, 0.2211976, 0.2211976, 0.2211976, 0.2211976, 0.2211976, 
    0.2211976, 0.2211976, 0.2298353, 0.2298353, 0.2298353, 0.2298353, 
    0.2298353, 0.2298353, 0.2298353, 0.2156998, 0.2156998, 0.2156998, 
    0.2156998, 0.2156998, 0.2156998, 0.2156998, 0.2121684,
  0.275326, 0.2455239, 0.2430588, 0.2483182, 0.2143765, 0.2111904, 0.2082938, 
    0.2040882, 0.1993012, 0.1945066, 0.1905111, 0.1840114, 0.1844856, 
    0.1766085, 0.1396889, 0.1281355, 0.1268771, 0.1430555, 0.1789336, 
    0.2214995, 0.2725159, 0.3061523, 0.2501554, 0.182193, 0.1881934, 
    0.2101838, 0.2228265, 0.2791847, 0.2921259,
  0.2043765, 0.1664654, 0.1651296, 0.1829219, 0.2231341, 0.1770311, 
    0.1591114, 0.2038256, 0.191384, 0.191544, 0.214398, 0.2177341, 0.2113422, 
    0.1826495, 0.2348853, 0.284482, 0.2659336, 0.2335105, 0.2292778, 
    0.2132672, 0.20491, 0.2358717, 0.428776, 0.516064, 0.5949415, 0.7860578, 
    0.7418979, 0.601243, 0.3249059,
  0.7222602, 0.5609685, 0.4359986, 0.4554656, 0.4379613, 0.3786412, 
    0.3069429, 0.2494773, 0.1996553, 0.1973155, 0.2073658, 0.293654, 
    0.5829603, 0.7020718, 0.729664, 0.7487649, 0.62971, 0.4831213, 0.3650751, 
    0.3003282, 0.255899, 0.240589, 0.3741917, 0.9305108, 3.23508, 2.822839, 
    1.947993, 1.182039, 0.9325101,
  1.293008, 0.9929271, 0.9026502, 1.007656, 0.8627341, 0.7455295, 0.5448422, 
    0.4163254, 0.3464801, 0.3191228, 0.3950456, 0.6550367, 1.911555, 
    2.021106, 2.595744, 1.642089, 1.065524, 0.7947049, 0.5846204, 0.444443, 
    0.375902, 0.3401252, 0.3641621, 10.7682, 10.69139, 6.228361, 3.528667, 
    2.363497, 1.723215,
  1.135818, 1.107546, 2.787409, 2.026124, 0.9811168, 0.7085916, 0.5917847, 
    0.5111827, 0.4914318, 0.6669035, 1.976481, 4.438077, 10.1752, 4.056872, 
    9.844956, 2.08917, 1.053183, 0.7808672, 0.6110412, 0.5109298, 0.4746803, 
    0.5607571, 0.9228639, 14.86992, 22.39325, 4.91537, 2.59214, 1.911237, 
    1.437259,
  1.070807, 5.474974, 35.34364, 4.013284, 1.403315, 0.8422814, 0.6547639, 
    0.5416721, 0.9008455, 10.58767, 28.07999, 30.55401, 25.77362, 3.687989, 
    1.954634, 1.232214, 0.8996706, 0.7029512, 0.5330108, 0.4609279, 
    0.4139309, 0.4275807, 0.5677394, 21.2404, 40.91842, 8.825224, 1.761693, 
    1.05734, 1.010485,
  2.613705, 31.94802, 40.90599, 9.243153, 2.422944, 0.9148062, 0.9141067, 
    1.583997, 4.924589, 20.37357, 39.87851, 32.65453, 5.17833, 2.054279, 
    1.305645, 0.8045096, 0.6225275, 0.5169068, 0.4354219, 0.3676674, 
    0.3583539, 0.4087081, 0.9392521, 8.131169, 48.40033, 34.12795, 1.294314, 
    0.758707, 1.08413,
  4.800344, 23.97169, 39.23547, 18.3575, 1.726291, 1.259019, 1.460229, 
    2.996279, 5.941132, 10.48227, 12.87367, 6.460266, 3.80707, 0.8238528, 
    0.4565932, 0.395889, 0.4574282, 0.5626879, 0.6513517, 0.6740649, 
    0.6364015, 0.7056729, 2.19715, 43.175, 38.01282, 29.24312, 1.633437, 
    1.227601, 2.270739,
  14.48907, 43.6334, 45.76482, 24.55988, 4.022579, 3.862811, 4.368524, 
    4.238746, 15.00961, 23.19883, 4.975522, 3.847567, 0.9322844, 0.3614912, 
    0.3679597, 0.5217429, 0.7877872, 1.215981, 1.809066, 2.574406, 3.273599, 
    3.88101, 8.349621, 37.75962, 29.33364, 9.044528, 7.279744, 8.886703, 
    10.98727,
  47.09783, 48.12553, 45.55158, 36.34564, 20.69247, 11.76855, 18.40115, 
    11.55697, 21.37372, 7.603295, 5.643266, 3.074064, 1.981736, 1.331475, 
    0.9032318, 0.9724611, 1.240787, 1.741416, 2.31111, 3.668315, 6.647932, 
    12.40697, 9.598971, 18.39653, 3.003652, 4.743378, 8.537838, 20.64628, 
    47.13638,
  47.00815, 49.87823, 45.29858, 28.81287, 42.18431, 22.04566, 37.85503, 
    37.8883, 44.85072, 27.14042, 9.051709, 5.238094, 4.25355, 3.718469, 
    3.033005, 2.428618, 2.615391, 2.780641, 4.247148, 8.407842, 13.59703, 
    24.99298, 10.23584, 7.087601, 2.953665, 3.566, 6.108559, 14.36561, 
    46.56471,
  42.14116, 38.12627, 32.08921, 41.25736, 39.87299, 49.26427, 52.32122, 
    38.32299, 49.47882, 63.20845, 22.902, 13.74733, 8.838875, 6.607987, 
    5.445612, 4.352273, 3.36282, 3.0191, 4.734205, 15.19507, 32.3665, 
    38.37357, 34.93692, 12.74416, 7.231593, 5.326924, 4.528205, 6.514729, 
    30.18548,
  29.19647, 26.50309, 39.35647, 39.3191, 56.63214, 59.81326, 48.22999, 
    62.22655, 64.51469, 57.66348, 52.62439, 30.4178, 17.40402, 10.61633, 
    7.829302, 5.986796, 4.720626, 4.098568, 4.227117, 26.6615, 36.97337, 
    56.36802, 58.25502, 47.25101, 21.70003, 11.78336, 7.894668, 7.280598, 
    20.66666,
  25.84244, 39.41565, 49.61137, 55.87584, 59.7959, 60.95244, 57.35936, 
    36.45903, 49.9564, 64.44161, 72.68729, 61.02437, 26.63696, 15.32889, 
    10.8635, 8.902562, 8.101133, 7.84994, 8.920084, 28.45563, 51.72504, 
    64.48637, 59.12078, 56.09322, 42.76602, 18.6003, 10.38626, 7.887611, 
    13.11056,
  14.50769, 27.16378, 38.75932, 50.12393, 52.30812, 52.81951, 55.98282, 
    62.78484, 59.70288, 60.95259, 58.5201, 40.27714, 27.40008, 26.95479, 
    20.61497, 15.4989, 22.22117, 20.6624, 30.34105, 43.05768, 52.35533, 
    43.25941, 30.9087, 33.44934, 22.92673, 10.21195, 8.682396, 8.042104, 
    9.55768,
  7.702012, 11.71786, 17.30605, 22.15807, 25.73183, 28.88001, 33.28051, 
    42.17609, 34.06222, 28.41252, 32.75702, 31.43505, 25.92082, 26.48115, 
    23.46069, 17.42136, 20.04946, 22.51772, 22.95665, 25.30235, 19.46322, 
    19.6003, 16.83591, 14.05661, 10.79448, 7.306567, 6.491508, 5.458089, 
    6.500249,
  7.260473, 8.600894, 10.08791, 11.91739, 13.85673, 16.14276, 17.88238, 
    19.36809, 19.83593, 19.2913, 18.78264, 17.58838, 16.22276, 14.65668, 
    13.28467, 11.99564, 11.48015, 11.77722, 11.73307, 11.03591, 9.989864, 
    8.930477, 7.889748, 7.627321, 7.110322, 7.035539, 7.017481, 6.505445, 
    6.775091,
  0.195764, 0.195764, 0.195764, 0.195764, 0.195764, 0.195764, 0.195764, 
    0.2043555, 0.2043555, 0.2043555, 0.2043555, 0.2043555, 0.2043555, 
    0.2043555, 0.2107716, 0.2107716, 0.2107716, 0.2107716, 0.2107716, 
    0.2107716, 0.2107716, 0.1983764, 0.1983764, 0.1983764, 0.1983764, 
    0.1983764, 0.1983764, 0.1983764, 0.195764,
  0.2611513, 0.2370166, 0.2305889, 0.2299524, 0.2080239, 0.203764, 0.200634, 
    0.1962758, 0.1897181, 0.1860653, 0.181326, 0.1775193, 0.1818507, 0.1774, 
    0.1400097, 0.1276894, 0.124663, 0.1407733, 0.1761979, 0.2122974, 
    0.2616779, 0.289562, 0.23667, 0.1809869, 0.1759436, 0.1979714, 0.2198165, 
    0.2721188, 0.2767511,
  0.1962656, 0.1674542, 0.1654752, 0.182507, 0.2101007, 0.1694916, 0.161252, 
    0.1930094, 0.1790545, 0.1838403, 0.1996603, 0.2052872, 0.2031964, 
    0.1799374, 0.2210182, 0.2626783, 0.2496312, 0.2203103, 0.2195387, 
    0.2019244, 0.2016264, 0.2301341, 0.4212892, 0.4883763, 0.581776, 
    0.7453459, 0.7093021, 0.5542116, 0.2926745,
  0.6942412, 0.5417504, 0.4258201, 0.4500644, 0.4301654, 0.3748413, 
    0.3028273, 0.2464243, 0.1938362, 0.1903535, 0.2041537, 0.278611, 
    0.5429095, 0.6741519, 0.7152815, 0.7279339, 0.5998979, 0.4665461, 
    0.3532391, 0.2952192, 0.2531216, 0.2392961, 0.3764728, 0.9808582, 
    3.414662, 2.856965, 1.940078, 1.151042, 0.897864,
  1.280673, 0.9846819, 0.8882395, 0.9810452, 0.8514594, 0.7137513, 0.5329982, 
    0.4147837, 0.3449349, 0.3146295, 0.3911304, 0.6340643, 1.88626, 2.023787, 
    2.753528, 1.636008, 1.057727, 0.7838089, 0.5772471, 0.4393377, 0.3717802, 
    0.3378355, 0.3674813, 13.45672, 11.3589, 6.388869, 3.483057, 2.303645, 
    1.694863,
  1.129584, 1.098608, 2.770511, 1.946599, 0.9603832, 0.6975251, 0.5831634, 
    0.5041894, 0.4859666, 0.6667458, 1.896353, 4.558115, 10.21559, 4.004609, 
    11.32012, 2.0721, 1.045369, 0.7764171, 0.607924, 0.5075554, 0.4717408, 
    0.5646879, 0.9163234, 18.11405, 24.60431, 4.857249, 2.571036, 1.886602, 
    1.423395,
  1.068525, 5.49917, 38.28203, 3.927137, 1.364771, 0.8119534, 0.6490895, 
    0.5370944, 0.899968, 10.78746, 30.78601, 33.15181, 28.39949, 3.630659, 
    1.947277, 1.229216, 0.8967509, 0.7010406, 0.5318517, 0.4602844, 
    0.4136883, 0.4278758, 0.5684248, 24.03648, 44.56504, 8.710939, 1.730878, 
    1.05333, 1.008035,
  2.599302, 36.02434, 43.97667, 9.233204, 2.406974, 0.9098226, 0.9123706, 
    1.577813, 4.910471, 20.80041, 42.47845, 34.80716, 5.134535, 2.056073, 
    1.309512, 0.8046656, 0.6224453, 0.5173114, 0.4354357, 0.3678566, 
    0.357946, 0.4085094, 0.9459483, 8.502193, 50.87075, 36.78303, 1.285071, 
    0.7561007, 1.083562,
  4.804586, 25.07329, 41.01508, 20.67373, 1.72755, 1.260449, 1.458021, 
    3.001771, 5.94753, 10.50856, 12.94488, 6.506135, 4.090027, 0.8236834, 
    0.457845, 0.3961606, 0.4577336, 0.5625899, 0.6496847, 0.6694801, 
    0.6289841, 0.6994231, 2.195022, 43.35966, 38.92494, 31.6103, 1.653672, 
    1.225557, 2.26811,
  14.46666, 43.19961, 45.12115, 25.90226, 4.029648, 3.870651, 4.388427, 
    4.250419, 15.48625, 23.96176, 4.998051, 3.855317, 0.9334015, 0.3615482, 
    0.3679188, 0.5218325, 0.7878162, 1.214887, 1.795351, 2.534538, 3.156162, 
    3.652349, 8.07533, 38.40601, 31.1296, 9.055709, 7.271106, 8.822683, 
    10.90136,
  48.77173, 50.12035, 47.66673, 38.16347, 21.89359, 11.79002, 19.09182, 
    11.55525, 21.75874, 7.634747, 5.770342, 3.083613, 1.987126, 1.337466, 
    0.9081188, 0.9751826, 1.244417, 1.745775, 2.318366, 3.673357, 6.657397, 
    12.50163, 10.70638, 19.63947, 3.002066, 4.738377, 8.522297, 20.68167, 
    48.60423,
  49.46647, 53.20917, 48.39312, 29.69054, 44.93978, 21.4803, 40.59826, 
    37.64338, 48.5958, 27.81733, 9.093001, 5.256363, 4.254266, 3.721743, 
    3.039614, 2.435754, 2.622834, 2.790165, 4.273513, 8.486026, 13.90797, 
    26.3844, 10.26145, 7.313838, 2.956017, 3.557861, 6.091661, 14.22158, 
    49.30745,
  45.82119, 40.78819, 34.13701, 44.19228, 42.65784, 53.23024, 56.75504, 
    41.65401, 52.96112, 68.04729, 23.07446, 13.76461, 8.852608, 6.621539, 
    5.45148, 4.358914, 3.370574, 3.026951, 4.744162, 15.93316, 35.86044, 
    41.48547, 37.86736, 12.74802, 7.240216, 5.337346, 4.530416, 6.464262, 
    33.23998,
  31.78845, 27.31449, 41.85855, 42.88332, 62.93739, 66.3722, 51.76861, 
    70.0228, 70.20433, 62.2962, 56.33536, 30.81623, 17.35469, 10.57629, 
    7.8074, 5.977814, 4.712821, 4.10868, 4.314877, 30.73436, 41.578, 
    61.15531, 62.79827, 48.73385, 21.73528, 11.76964, 7.89087, 7.281248, 
    22.99314,
  29.03808, 45.26522, 55.76379, 64.66347, 70.88466, 71.45867, 64.23087, 
    40.70045, 56.08872, 71.55356, 80.89432, 69.88081, 26.76277, 15.37046, 
    10.83151, 8.860952, 8.113016, 7.942384, 9.207063, 33.48481, 57.92752, 
    70.48018, 64.86586, 62.97461, 46.17809, 18.64217, 10.34604, 7.872706, 
    13.5359,
  14.98536, 30.65819, 43.17519, 57.48373, 60.8425, 61.24574, 66.14278, 
    73.45976, 70.06905, 72.34147, 68.19557, 46.63331, 32.46106, 32.28476, 
    21.24172, 16.41578, 26.731, 23.65375, 36.41852, 49.1644, 60.35355, 
    49.53646, 33.58229, 37.67405, 23.20782, 10.269, 8.688784, 8.038992, 
    9.733064,
  7.679257, 11.845, 18.96325, 22.90652, 27.45417, 31.86518, 38.72274, 
    49.17467, 38.17368, 32.87269, 38.02326, 37.43887, 31.82724, 32.90553, 
    27.9642, 19.52426, 22.34661, 25.93785, 26.00523, 29.06587, 22.41787, 
    22.32015, 18.92415, 15.72639, 10.95178, 7.211775, 6.433012, 5.403213, 
    6.429934,
  7.239048, 8.617623, 10.41571, 12.48708, 14.59139, 16.79046, 19.17505, 
    20.89267, 20.83559, 20.28587, 19.79056, 18.78233, 17.54317, 15.72068, 
    14.19119, 12.80561, 12.07206, 12.29873, 12.13819, 11.40176, 10.47393, 
    8.910903, 7.816611, 7.5334, 7.063246, 6.957053, 6.924455, 6.410952, 
    6.557846,
  0.1867052, 0.1867052, 0.1867052, 0.1867052, 0.1867052, 0.1867052, 
    0.1867052, 0.1893054, 0.1893054, 0.1893054, 0.1893054, 0.1893054, 
    0.1893054, 0.1893054, 0.1935619, 0.1935619, 0.1935619, 0.1935619, 
    0.1935619, 0.1935619, 0.1935619, 0.1879463, 0.1879463, 0.1879463, 
    0.1879463, 0.1879463, 0.1879463, 0.1879463, 0.1867052,
  0.2500449, 0.2307612, 0.2198764, 0.2145719, 0.2027036, 0.1980734, 
    0.1953363, 0.1909217, 0.1845458, 0.1812636, 0.1758073, 0.1728161, 
    0.1782444, 0.1775847, 0.1413715, 0.1275861, 0.1241487, 0.139655, 
    0.1770186, 0.2051513, 0.2516343, 0.2719839, 0.2285404, 0.1797423, 
    0.1697517, 0.1914527, 0.2186254, 0.2677292, 0.2657917,
  0.1910064, 0.1693244, 0.1663672, 0.1825181, 0.1992918, 0.1647302, 
    0.1630526, 0.1824051, 0.1724635, 0.1774581, 0.187796, 0.1953025, 
    0.1973228, 0.1787373, 0.2111252, 0.2490548, 0.2387944, 0.2119059, 
    0.2133378, 0.1965547, 0.1984813, 0.2263266, 0.4165221, 0.4668813, 
    0.5731247, 0.7160949, 0.6723729, 0.5237899, 0.2711837,
  0.6797754, 0.5321198, 0.420503, 0.445086, 0.4248545, 0.3721754, 0.2999102, 
    0.2449481, 0.1916342, 0.1860887, 0.201698, 0.267336, 0.5213138, 
    0.6519991, 0.7077314, 0.7128854, 0.5848143, 0.454929, 0.3480155, 
    0.2926254, 0.2516883, 0.2386, 0.3774142, 1.013312, 3.498182, 2.887146, 
    1.922171, 1.129272, 0.8791083,
  1.272847, 0.9806931, 0.8777222, 0.9592381, 0.8377293, 0.689424, 0.5260914, 
    0.4140604, 0.3442505, 0.3121245, 0.3899424, 0.6262205, 1.860621, 
    2.015262, 2.850809, 1.630151, 1.053925, 0.7787705, 0.5742834, 0.4373533, 
    0.370098, 0.3369881, 0.3688741, 16.68666, 11.67084, 6.442644, 3.452917, 
    2.275736, 1.679859,
  1.127208, 1.094425, 2.755901, 1.91774, 0.9519091, 0.6933822, 0.5801195, 
    0.5012026, 0.4836093, 0.665244, 1.859211, 4.671752, 10.23715, 3.970969, 
    13.13378, 2.062603, 1.041849, 0.7741466, 0.6062357, 0.5059522, 0.4704908, 
    0.5662143, 0.8976187, 21.94486, 26.91518, 4.821564, 2.559227, 1.876912, 
    1.417125,
  1.067589, 5.548201, 42.88445, 3.888777, 1.345818, 0.79978, 0.6471738, 
    0.5352955, 0.8991517, 10.92076, 34.63051, 37.00253, 32.10093, 3.606786, 
    1.943526, 1.228183, 0.8954831, 0.7001292, 0.5314704, 0.4601965, 
    0.4134983, 0.4282122, 0.5688039, 26.26876, 49.25433, 8.670573, 1.718588, 
    1.051597, 1.007031,
  2.591822, 40.89777, 48.36079, 9.189458, 2.415803, 0.9089587, 0.9118194, 
    1.575513, 4.908525, 20.90507, 47.09244, 38.45109, 5.124647, 2.056438, 
    1.310562, 0.8050019, 0.6223341, 0.517481, 0.4355338, 0.3679273, 
    0.3578693, 0.4083922, 0.9472308, 8.497594, 54.72517, 40.45848, 1.282061, 
    0.7556199, 1.083106,
  4.804395, 26.7767, 44.53823, 23.79728, 1.727944, 1.260697, 1.457722, 
    3.003271, 5.94907, 10.51983, 12.98494, 6.521163, 4.397038, 0.8231829, 
    0.4581558, 0.3962502, 0.4578476, 0.5625429, 0.6491777, 0.6681923, 
    0.6265399, 0.6974167, 2.191362, 45.00033, 40.89997, 35.57382, 1.660215, 
    1.2248, 2.267285,
  14.45673, 44.24976, 46.18502, 27.58977, 4.03104, 3.873757, 4.39433, 
    4.254692, 17.08376, 25.77821, 5.005329, 3.857808, 0.9340573, 0.3616026, 
    0.3679526, 0.5218638, 0.7878243, 1.21447, 1.791432, 2.520246, 3.119374, 
    3.584282, 7.995908, 39.95953, 34.43647, 9.059086, 7.269742, 8.809716, 
    10.87865,
  52.43768, 53.2168, 51.06952, 41.68251, 23.36385, 11.7964, 19.98894, 
    11.55801, 21.9743, 7.642304, 5.836987, 3.086072, 1.988994, 1.338942, 
    0.9092814, 0.9759701, 1.245442, 1.747068, 2.320508, 3.675125, 6.660601, 
    12.527, 12.27075, 21.74222, 3.00158, 4.736437, 8.518579, 20.68565, 
    51.96306,
  53.81883, 58.21296, 53.02913, 30.5582, 49.42389, 21.30037, 44.8419, 
    37.65874, 53.32299, 28.09521, 9.103786, 5.262394, 4.254794, 3.722752, 
    3.041495, 2.43796, 2.625238, 2.792964, 4.282369, 8.508824, 13.98468, 
    28.17405, 10.27203, 7.480675, 2.956948, 3.556372, 6.091595, 14.24818, 
    53.75571,
  50.69237, 44.61756, 37.14478, 48.87573, 46.3351, 58.356, 63.29585, 
    45.86584, 57.17307, 74.20384, 23.18259, 13.77229, 8.855392, 6.626689, 
    5.451811, 4.362412, 3.37323, 3.028405, 4.750277, 16.6368, 40.36232, 
    45.50519, 41.74606, 12.7541, 7.24524, 5.341165, 4.53177, 6.43579, 37.07895,
  34.88197, 28.26084, 44.58963, 46.69896, 72.27171, 73.06049, 56.39895, 
    79.22845, 76.69729, 67.29247, 60.62931, 31.05644, 17.29705, 10.54953, 
    7.7858, 5.964715, 4.703483, 4.114715, 4.31671, 35.70296, 47.63676, 
    66.91745, 67.77468, 49.97493, 21.73852, 11.76299, 7.88819, 7.27971, 
    25.65241,
  32.40907, 51.08319, 62.56683, 73.06059, 83.87714, 84.3652, 71.30239, 
    45.99367, 63.7015, 78.53375, 88.29085, 78.28038, 26.76658, 15.29309, 
    10.75474, 8.820501, 8.127961, 7.922163, 9.384232, 39.9307, 64.50861, 
    76.01182, 70.57733, 69.84995, 48.89018, 18.58285, 10.32343, 7.864083, 
    13.84569,
  15.29571, 34.98876, 47.27845, 64.11396, 69.39729, 70.14425, 77.21525, 
    83.97734, 82.61196, 85.52794, 78.13716, 53.90767, 39.49162, 38.00174, 
    21.6481, 17.1606, 32.17857, 27.1318, 43.65988, 56.17321, 67.52496, 
    56.37355, 34.68335, 42.81758, 23.36034, 10.33718, 8.690552, 8.039106, 
    9.8059,
  7.649647, 11.89977, 21.20312, 23.37815, 29.10966, 34.80414, 44.53082, 
    55.59069, 42.90729, 38.83072, 43.66844, 45.16835, 38.75761, 40.49028, 
    32.74329, 21.75126, 25.237, 29.3591, 29.30426, 32.95084, 26.17994, 
    25.44525, 21.14864, 17.65637, 11.15607, 7.130839, 6.361743, 5.371073, 
    6.392998,
  7.130416, 8.546899, 10.28519, 12.40856, 14.51229, 16.68701, 19.51777, 
    21.54721, 21.18429, 20.58559, 20.33407, 19.77964, 18.62097, 16.81156, 
    14.97784, 13.37198, 12.51611, 12.49946, 12.17888, 11.5442, 10.5963, 
    8.776625, 7.695233, 7.47488, 7.032848, 6.912582, 6.841928, 6.369389, 
    6.406349,
  0.1845552, 0.1845552, 0.1845552, 0.1845552, 0.1845552, 0.1845552, 
    0.1845552, 0.1828895, 0.1828895, 0.1828895, 0.1828895, 0.1828895, 
    0.1828895, 0.1828895, 0.1845149, 0.1845149, 0.1845149, 0.1845149, 
    0.1845149, 0.1845149, 0.1845149, 0.1837774, 0.1837774, 0.1837774, 
    0.1837774, 0.1837774, 0.1837774, 0.1837774, 0.1845552,
  0.2397681, 0.2250075, 0.2104963, 0.2013103, 0.199289, 0.1946204, 0.1921776, 
    0.188555, 0.1817753, 0.1777173, 0.1730631, 0.1695651, 0.1745418, 
    0.1775456, 0.1432465, 0.1269255, 0.1234704, 0.1396185, 0.1805927, 
    0.2025109, 0.2455323, 0.2576008, 0.2244135, 0.1780916, 0.1656251, 
    0.1887873, 0.2183464, 0.2646837, 0.2560225,
  0.1881869, 0.1710618, 0.166899, 0.1829061, 0.1904972, 0.1623828, 0.1644562, 
    0.1775724, 0.1695806, 0.1740866, 0.1827623, 0.1874391, 0.1946867, 
    0.1780111, 0.2045175, 0.2418015, 0.2331291, 0.2070241, 0.2096896, 
    0.194564, 0.1956645, 0.2243773, 0.411575, 0.4555787, 0.568494, 0.6965212, 
    0.6502396, 0.5099524, 0.2605556,
  0.6726427, 0.5277817, 0.4176444, 0.4433385, 0.4215862, 0.3705168, 
    0.2979971, 0.2440869, 0.1906692, 0.1841103, 0.2000821, 0.2608142, 
    0.50725, 0.6383215, 0.7035049, 0.7026245, 0.5755251, 0.4485439, 
    0.3457421, 0.2914527, 0.2510441, 0.2382343, 0.3778683, 1.029963, 
    3.523914, 2.891545, 1.902837, 1.118525, 0.8693191,
  1.268146, 0.9783456, 0.870056, 0.9435769, 0.8208601, 0.6758505, 0.5219946, 
    0.4135914, 0.3438983, 0.3110952, 0.3889126, 0.6230808, 1.840206, 
    2.006521, 2.882354, 1.627042, 1.051872, 0.7763708, 0.5731888, 0.4365072, 
    0.3693286, 0.3364354, 0.3695155, 20.87469, 11.71763, 6.446299, 3.427727, 
    2.262058, 1.670725,
  1.125914, 1.092101, 2.743991, 1.905465, 0.9474032, 0.6915993, 0.5784665, 
    0.4999328, 0.482563, 0.662756, 1.844346, 4.74862, 10.25518, 3.95339, 
    15.57555, 2.05722, 1.040247, 0.7729503, 0.605381, 0.5049847, 0.4701181, 
    0.5669353, 0.8949122, 26.93799, 29.13792, 4.801504, 2.552644, 1.871998, 
    1.414665,
  1.067205, 5.604344, 50.72953, 3.869162, 1.337974, 0.795091, 0.6464919, 
    0.5344356, 0.8985594, 11.00226, 40.33926, 42.91748, 37.50831, 3.596719, 
    1.942062, 1.227666, 0.894893, 0.6997467, 0.5312957, 0.46014, 0.4134173, 
    0.4282407, 0.5689083, 28.45717, 55.56522, 8.65313, 1.714538, 1.050685, 
    1.006636,
  2.589266, 46.81869, 54.93798, 9.165668, 2.422075, 0.9086167, 0.9115017, 
    1.574368, 4.906776, 20.91386, 54.88425, 44.60778, 5.123438, 2.056486, 
    1.310873, 0.8051016, 0.6222708, 0.5175461, 0.4355734, 0.3679446, 
    0.3578337, 0.4083354, 0.9473932, 8.463987, 61.63586, 46.47627, 1.280939, 
    0.7554066, 1.082741,
  4.804418, 29.44862, 52.03605, 27.99464, 1.728094, 1.260764, 1.457595, 
    3.003698, 5.949598, 10.52548, 13.00278, 6.527547, 4.76335, 0.8229759, 
    0.4582883, 0.3962836, 0.457893, 0.5625123, 0.6489339, 0.6675755, 
    0.625425, 0.6965777, 2.189941, 50.77832, 46.87601, 42.71595, 1.661739, 
    1.224478, 2.266927,
  14.45173, 49.76954, 52.36669, 29.94906, 4.031525, 3.875176, 4.396851, 
    4.256516, 21.6397, 31.08896, 5.008983, 3.858869, 0.9342227, 0.361617, 
    0.3679736, 0.5218629, 0.7878124, 1.214288, 1.790111, 2.515454, 3.10917, 
    3.564449, 7.965623, 45.49673, 40.60741, 9.058471, 7.26975, 8.805715, 
    10.87099,
  59.97418, 58.8932, 56.61495, 48.24759, 25.68839, 11.79975, 21.25548, 
    11.55948, 22.07857, 7.645186, 5.866838, 3.087037, 1.989859, 1.339618, 
    0.9098313, 0.9762926, 1.245848, 1.747602, 2.321338, 3.675802, 6.661912, 
    12.53778, 14.63148, 25.43095, 3.001256, 4.735564, 8.517083, 20.68551, 
    59.40228,
  61.89168, 65.51559, 60.15525, 31.14913, 57.1203, 21.25211, 50.97587, 
    37.72766, 60.70229, 28.22816, 9.107894, 5.264795, 4.254961, 3.723117, 
    3.042229, 2.438946, 2.626245, 2.793805, 4.285938, 8.518045, 14.0044, 
    30.9957, 10.27744, 7.600688, 2.957366, 3.555892, 6.091552, 14.26972, 
    61.7774,
  58.35569, 51.02323, 42.43321, 56.23833, 52.10713, 65.57144, 73.51981, 
    51.47336, 62.66194, 82.35292, 23.23916, 13.77341, 8.856837, 6.628286, 
    5.450861, 4.363534, 3.374472, 3.028928, 4.752496, 17.06978, 47.20175, 
    51.56445, 47.93272, 12.75747, 7.247174, 5.342814, 4.53264, 6.424783, 
    42.8965,
  38.77036, 29.25283, 47.64825, 51.62401, 87.15549, 81.49844, 63.41759, 
    89.89162, 85.12155, 73.87016, 66.35784, 31.20949, 17.24053, 10.53871, 
    7.775557, 5.952922, 4.696519, 4.116264, 4.318249, 42.985, 55.98639, 
    74.23471, 74.06078, 51.01447, 21.73991, 11.76076, 7.885429, 7.279345, 
    28.55933,
  35.09585, 57.54869, 70.64131, 82.79121, 97.78465, 99.76031, 79.85188, 
    53.40354, 73.67348, 86.71268, 96.64599, 86.36521, 26.69184, 15.18844, 
    10.72396, 8.797892, 8.133154, 7.919512, 9.442423, 48.73418, 72.20205, 
    82.18509, 77.18464, 76.94688, 51.20487, 18.52412, 10.3116, 7.861915, 
    14.02471,
  15.41194, 40.99143, 50.71993, 69.65706, 76.83022, 78.812, 86.83138, 
    93.13291, 95.55847, 98.1207, 87.90301, 63.05593, 48.77492, 43.6333, 
    21.92811, 17.53808, 39.16222, 31.2341, 51.61818, 64.39787, 73.9232, 
    63.71401, 35.01596, 49.03832, 23.4367, 10.392, 8.690084, 8.03912, 9.826776,
  7.628272, 11.90363, 23.85019, 23.72729, 30.14043, 37.53691, 50.08922, 
    61.08013, 48.64536, 46.11203, 48.81365, 53.78066, 47.98763, 47.92721, 
    37.18465, 23.6, 28.54797, 32.19622, 32.22576, 36.06083, 31.13611, 
    28.62473, 22.86014, 20.49327, 11.27639, 7.060326, 6.289242, 5.338724, 
    6.382876,
  7.089921, 8.489287, 10.05322, 12.2933, 14.3477, 16.41586, 19.30546, 
    21.47076, 21.09914, 20.49807, 20.52957, 20.2022, 19.36539, 17.70084, 
    15.70968, 13.8146, 12.83927, 12.65027, 12.1785, 11.48137, 10.54172, 
    8.615923, 7.568262, 7.415557, 7.01511, 6.875118, 6.778393, 6.323478, 
    6.347658,
  0.1836565, 0.1836565, 0.1836565, 0.1836565, 0.1836565, 0.1836565, 
    0.1836565, 0.1807598, 0.1807598, 0.1807598, 0.1807598, 0.1807598, 
    0.1807598, 0.1807598, 0.1807906, 0.1807906, 0.1807906, 0.1807906, 
    0.1807906, 0.1807906, 0.1807906, 0.1815091, 0.1815091, 0.1815091, 
    0.1815091, 0.1815091, 0.1815091, 0.1815091, 0.1836565,
  0.2343223, 0.2209795, 0.2043144, 0.1929999, 0.196169, 0.1922857, 0.1902238, 
    0.1871262, 0.1794737, 0.1754618, 0.1716341, 0.168156, 0.1719578, 
    0.1771545, 0.1443741, 0.1261234, 0.1229006, 0.1411362, 0.1843873, 
    0.2022168, 0.2420906, 0.2492415, 0.2225556, 0.1764602, 0.162214, 
    0.1870906, 0.2181509, 0.2639144, 0.2490561,
  0.187228, 0.1723244, 0.1671597, 0.183319, 0.1845763, 0.161212, 0.1654558, 
    0.1764194, 0.1688847, 0.1726112, 0.1811739, 0.1847244, 0.193287, 
    0.1778324, 0.200062, 0.2383002, 0.2304534, 0.2043, 0.2079306, 0.1936612, 
    0.1943502, 0.2235549, 0.4095752, 0.4505627, 0.5675382, 0.6857195, 
    0.6385227, 0.5033849, 0.2565751,
  0.6692104, 0.5255449, 0.4162678, 0.4427462, 0.4198182, 0.3694432, 
    0.2970594, 0.2435003, 0.1901297, 0.183154, 0.1991171, 0.2583236, 
    0.496224, 0.6298807, 0.7018982, 0.695527, 0.5687647, 0.4444426, 
    0.3446104, 0.2908211, 0.2506852, 0.2380324, 0.3780979, 1.039287, 
    3.533101, 2.884131, 1.890347, 1.113117, 0.8638209,
  1.265332, 0.9765645, 0.8644835, 0.9311904, 0.8076512, 0.667938, 0.5196292, 
    0.4131946, 0.3436314, 0.3104378, 0.3878539, 0.6208835, 1.825306, 
    1.999833, 2.889953, 1.625039, 1.050875, 0.7753155, 0.5727338, 0.4360855, 
    0.368906, 0.3360259, 0.3699007, 26.46751, 11.67662, 6.427775, 3.409189, 
    2.25289, 1.665016,
  1.125143, 1.090926, 2.735896, 1.899451, 0.9444568, 0.6904944, 0.577505, 
    0.4992432, 0.4820609, 0.6605859, 1.838848, 4.785595, 10.25125, 3.942703, 
    19.70147, 2.054244, 1.039447, 0.772244, 0.6049566, 0.5044069, 0.4700631, 
    0.5672522, 0.8942916, 35.10328, 30.76228, 4.789558, 2.549204, 1.869313, 
    1.413412,
  1.066987, 5.616731, 65.2174, 3.859627, 1.33377, 0.7929817, 0.646174, 
    0.5340014, 0.8981586, 11.03702, 49.63142, 53.18906, 47.08826, 3.591935, 
    1.941287, 1.227369, 0.8945679, 0.6995367, 0.5312002, 0.4600841, 
    0.4133792, 0.4282277, 0.5689552, 30.72219, 64.7382, 8.63851, 1.7128, 
    1.050262, 1.006442,
  2.587937, 55.26173, 66.61246, 9.156287, 2.427219, 0.9084311, 0.9113001, 
    1.573689, 4.90568, 20.91534, 69.32765, 55.59047, 5.123151, 2.056499, 
    1.310961, 0.805125, 0.6222373, 0.5175669, 0.4355883, 0.3679458, 
    0.3578088, 0.4082975, 0.9474543, 8.447308, 75.0431, 57.63905, 1.280465, 
    0.7552859, 1.082506,
  4.804389, 35.53048, 68.88678, 34.17503, 1.728119, 1.260759, 1.457487, 
    3.003799, 5.949768, 10.52855, 13.01329, 6.531019, 5.159082, 0.8229438, 
    0.4583569, 0.396302, 0.4579116, 0.5624893, 0.6487924, 0.6672221, 
    0.6248209, 0.6961494, 2.189254, 67.65474, 62.13598, 56.54036, 1.662983, 
    1.224285, 2.266722,
  14.44894, 68.66165, 71.60869, 33.77109, 4.031725, 3.87579, 4.397975, 
    4.25724, 36.1696, 46.90523, 5.011384, 3.85936, 0.9342781, 0.3616183, 
    0.3679781, 0.521856, 0.7877957, 1.214173, 1.789536, 2.513306, 3.10559, 
    3.557343, 7.952315, 61.11032, 54.76284, 9.056561, 7.269518, 8.803885, 
    10.86757,
  75.88767, 72.41269, 67.49055, 62.37434, 29.94206, 11.80157, 23.35758, 
    11.56019, 22.14093, 7.646518, 5.886144, 3.087468, 1.990319, 1.339994, 
    0.9100928, 0.976455, 1.246033, 1.747849, 2.321726, 3.676073, 6.662572, 
    12.54361, 19.68689, 30.72467, 3.001044, 4.735106, 8.516404, 20.68588, 
    77.35792,
  78.41781, 78.34711, 74.31876, 31.43154, 72.3616, 21.23942, 60.89283, 
    37.78557, 74.44736, 28.2912, 9.109962, 5.266012, 4.255089, 3.723299, 
    3.042576, 2.439414, 2.626636, 2.794168, 4.287537, 8.522753, 14.01115, 
    36.19541, 10.28058, 7.673872, 2.957584, 3.555638, 6.091353, 14.27055, 
    79.01308,
  73.45344, 63.06799, 52.82583, 69.74151, 63.70716, 78.69741, 89.39156, 
    60.41645, 71.33209, 95.98394, 23.26324, 13.77409, 8.857118, 6.628799, 
    5.450278, 4.363347, 3.375047, 3.02917, 4.753617, 17.2068, 59.40361, 
    61.07218, 59.12729, 12.75884, 7.247752, 5.343589, 4.533027, 6.421901, 
    53.74182,
  44.01929, 30.27309, 51.28828, 60.28422, 117.4128, 94.04648, 77.82687, 
    104.5106, 99.07629, 84.50882, 75.98818, 31.28512, 17.21382, 10.53013, 
    7.771493, 5.945718, 4.692236, 4.11666, 4.318878, 55.29141, 69.23284, 
    84.80025, 83.27959, 51.86977, 21.73946, 11.75972, 7.88328, 7.278702, 
    31.52883,
  37.11136, 65.40439, 80.59516, 94.685, 113.1168, 117.2172, 91.47063, 
    69.19384, 87.52202, 98.12813, 108.4864, 96.41669, 26.63271, 15.13416, 
    10.71245, 8.787526, 8.136562, 7.920138, 9.458996, 61.05651, 83.08198, 
    90.49181, 86.02306, 85.06693, 53.52443, 18.4789, 10.30646, 7.859756, 
    14.09122,
  15.4431, 48.98676, 54.23183, 75.017, 83.01718, 87.06475, 95.00419, 
    100.8271, 106.7053, 108.4566, 98.32821, 74.93463, 59.67374, 48.74986, 
    22.0565, 17.64916, 46.65129, 36.67875, 59.98475, 73.91439, 80.26309, 
    71.776, 35.03218, 57.17186, 23.45749, 10.42999, 8.689426, 8.038771, 
    9.834986,
  7.625116, 11.87654, 26.48655, 23.92744, 30.4024, 39.14312, 53.89163, 
    66.36544, 54.58265, 51.35251, 52.30616, 59.72591, 54.59047, 52.34892, 
    40.18656, 24.31417, 31.86068, 34.1584, 33.9488, 38.11263, 36.68829, 
    31.12383, 24.02641, 25.56618, 11.26998, 7.006742, 6.220743, 5.321117, 
    6.377306,
  7.075942, 8.490022, 9.955416, 12.26578, 14.30707, 16.26779, 19.18691, 
    21.37566, 21.00982, 20.41423, 20.52216, 20.20891, 19.47036, 17.92389, 
    15.99089, 13.97516, 12.93176, 12.62361, 12.11427, 11.42475, 10.46203, 
    8.503734, 7.480387, 7.335333, 6.998674, 6.825962, 6.726771, 6.299751, 
    6.327248,
  0.1830172, 0.1830172, 0.1830172, 0.1830172, 0.1830172, 0.1830172, 
    0.1830172, 0.1800378, 0.1800378, 0.1800378, 0.1800378, 0.1800378, 
    0.1800378, 0.1800378, 0.1797999, 0.1797999, 0.1797999, 0.1797999, 
    0.1797999, 0.1797999, 0.1797999, 0.1809472, 0.1809472, 0.1809472, 
    0.1809472, 0.1809472, 0.1809472, 0.1809472, 0.1830172,
  0.2321628, 0.2189483, 0.2018014, 0.1904988, 0.1947195, 0.191612, 0.1895826, 
    0.1863981, 0.1786638, 0.1745263, 0.1710492, 0.1676851, 0.1707922, 
    0.1766776, 0.1446727, 0.1256107, 0.122343, 0.1417824, 0.1855617, 
    0.2022805, 0.2406474, 0.2465921, 0.2213084, 0.1755888, 0.1603592, 
    0.1860067, 0.2172446, 0.2634422, 0.2457712,
  0.1867602, 0.1726869, 0.1672785, 0.183544, 0.182448, 0.1605894, 0.1659336, 
    0.1760402, 0.168776, 0.172488, 0.1808398, 0.1840364, 0.1928882, 
    0.1775319, 0.196972, 0.2368892, 0.2292691, 0.2028779, 0.2072551, 
    0.1932683, 0.193972, 0.2231889, 0.4087738, 0.4489911, 0.5688769, 
    0.6792787, 0.6331583, 0.5003545, 0.2550911,
  0.6675171, 0.5245636, 0.4155932, 0.4423693, 0.4190683, 0.3689176, 
    0.2966548, 0.2432142, 0.1897729, 0.1827032, 0.1985791, 0.2572365, 
    0.4894466, 0.6252253, 0.7012065, 0.6900014, 0.564952, 0.4414373, 
    0.3438663, 0.2904543, 0.2504925, 0.2379246, 0.378119, 1.044761, 3.537332, 
    2.871844, 1.878893, 1.109964, 0.8610432,
  1.263211, 0.9750137, 0.8631408, 0.9233932, 0.8011606, 0.6642553, 0.5183473, 
    0.4129584, 0.343445, 0.3099774, 0.3865496, 0.6194767, 1.812166, 1.993407, 
    2.889472, 1.623603, 1.050326, 0.7747726, 0.572476, 0.4358628, 0.368777, 
    0.3357699, 0.3702446, 35.64325, 11.63918, 6.400451, 3.394313, 2.246086, 
    1.66126,
  1.124637, 1.090405, 2.72992, 1.896371, 0.9423411, 0.6897693, 0.5768511, 
    0.4988052, 0.481804, 0.659327, 1.836756, 4.79586, 10.23618, 3.935667, 
    26.66829, 2.052795, 1.038963, 0.77184, 0.6047231, 0.5040893, 0.470017, 
    0.5673311, 0.8940023, 49.52427, 31.49985, 4.781196, 2.54718, 1.86758, 
    1.412739,
  1.066847, 5.610649, 95.4231, 3.854683, 1.331165, 0.7920783, 0.6459973, 
    0.5337813, 0.8979549, 11.03432, 66.72967, 70.55579, 65.66341, 3.589753, 
    1.940846, 1.227177, 0.8943897, 0.699414, 0.5311333, 0.4600443, 0.4133559, 
    0.4282141, 0.5689664, 32.5528, 80.69199, 8.629315, 1.711867, 1.05005, 
    1.006337,
  2.587434, 67.78394, 90.20565, 9.151943, 2.42884, 0.9083194, 0.9111699, 
    1.573273, 4.904991, 20.91595, 96.18049, 77.11339, 5.123066, 2.056493, 
    1.310971, 0.8051205, 0.6222165, 0.5175743, 0.4355918, 0.3679433, 
    0.3577901, 0.4082721, 0.947472, 8.43866, 106.6334, 81.71753, 1.280231, 
    0.7552118, 1.082368,
  4.804335, 48.30406, 110.2506, 44.51353, 1.728109, 1.260731, 1.457399, 
    3.003777, 5.949725, 10.53098, 13.0199, 6.532798, 5.717745, 0.8229315, 
    0.4583899, 0.3963081, 0.4579161, 0.562469, 0.6487076, 0.6670259, 
    0.6245047, 0.6959379, 2.188928, 120.4041, 102.1439, 84.88774, 1.663718, 
    1.224161, 2.266579,
  14.44728, 123.6215, 126.3112, 39.79053, 4.031743, 3.876026, 4.398426, 
    4.257525, 76.76659, 89.82708, 5.013388, 3.859617, 0.9342878, 0.3616148, 
    0.3679737, 0.5218433, 0.7877705, 1.214084, 1.789225, 2.512375, 3.104146, 
    3.55487, 7.947061, 102.6705, 86.51524, 9.054829, 7.269166, 8.802851, 
    10.86563,
  113.2795, 98.66676, 85.21989, 93.10471, 36.3805, 11.80242, 27.82697, 
    11.56033, 22.18229, 7.647018, 5.900556, 3.087621, 1.990525, 1.340179, 
    0.9102095, 0.9765242, 1.246101, 1.747941, 2.321887, 3.676137, 6.662781, 
    12.54657, 32.90568, 38.4539, 3.000876, 4.734792, 8.515959, 20.6861, 
    118.0746,
  97.53346, 102.4282, 92.7276, 31.52845, 98.72373, 21.23565, 75.36081, 
    37.81243, 102.1569, 28.3223, 9.111006, 5.266669, 4.255156, 3.723375, 
    3.042743, 2.439646, 2.626757, 2.794273, 4.288209, 8.525073, 14.01415, 
    45.10903, 10.28232, 7.711299, 2.957678, 3.555452, 6.091117, 14.26911, 
    103.9206,
  101.2534, 83.46094, 71.27958, 88.89589, 87.33348, 101.676, 114.8962, 
    72.02972, 85.7618, 121.2348, 23.26675, 13.77406, 8.856251, 6.628633, 
    5.449748, 4.362847, 3.375314, 3.029182, 4.754155, 17.22709, 82.45274, 
    81.17115, 81.51618, 12.75913, 7.247625, 5.343802, 4.533104, 6.420838, 
    71.07201,
  51.91103, 30.85057, 56.52483, 78.98534, 158.5402, 114.5219, 100.4564, 
    129.3025, 122.0926, 102.8396, 93.43543, 31.30679, 17.1978, 10.52232, 
    7.768935, 5.941621, 4.689216, 4.116649, 4.319179, 76.63359, 91.09911, 
    104.2968, 100.7001, 52.88546, 21.73624, 11.75871, 7.882007, 7.277975, 
    34.97157,
  39.0601, 79.06976, 98.03624, 116.2615, 133.3574, 142.6494, 111.994, 
    95.76788, 107.5593, 120.7536, 130.1772, 113.3673, 26.6072, 15.11478, 
    10.70878, 8.783196, 8.137673, 7.919577, 9.46513, 81.66874, 102.8623, 
    105.6434, 102.1064, 98.4668, 56.60724, 18.44585, 10.30405, 7.857541, 
    14.11692,
  15.45422, 60.46137, 59.71362, 82.46527, 91.8737, 99.06068, 107.0777, 
    111.8517, 123.196, 123.2894, 112.8761, 90.47037, 72.81858, 56.09212, 
    22.07834, 17.66465, 57.48666, 41.069, 72.15166, 88.21484, 89.91603, 
    84.13793, 34.99161, 68.28332, 23.44573, 10.45828, 8.688264, 8.038462, 
    9.837646,
  7.620437, 11.85673, 28.40279, 23.97136, 30.45284, 39.53924, 56.07699, 
    72.81481, 59.78307, 54.14567, 54.07816, 62.64185, 57.79655, 53.77367, 
    41.71376, 24.38621, 34.30349, 35.54052, 34.45811, 39.24881, 44.72125, 
    32.03192, 24.59001, 33.40801, 11.24519, 6.97137, 6.191442, 5.318031, 
    6.370452,
  7.069119, 8.491707, 9.932939, 12.2496, 14.27919, 16.21104, 19.11423, 
    21.33723, 20.96618, 20.35874, 20.48543, 20.19796, 19.48082, 17.95564, 
    16.01758, 14.00328, 12.9283, 12.60122, 12.08921, 11.39805, 10.42944, 
    8.467238, 7.462381, 7.30438, 6.982195, 6.795946, 6.68722, 6.269146, 
    6.312067 ;

 time = 912.5 ;

 time_bnds =
  730, 1095 ;
}
