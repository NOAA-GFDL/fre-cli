netcdf atmos.1980-1981.alb_sfc.03 {
dimensions:
	time = UNLIMITED ; // (1 currently)
	lat = 18 ;
	lon = 29 ;
	bnds = 2 ;
variables:
	float alb_sfc(time, lat, lon) ;
		alb_sfc:long_name = "Surface Albedo for  Flux" ;
		alb_sfc:units = "percent" ;
		alb_sfc:_FillValue = 1.e+20f ;
		alb_sfc:missing_value = 1.e+20f ;
		alb_sfc:cell_measures = "area: area" ;
		alb_sfc:interp_method = "conserve_order1" ;
		alb_sfc:cell_methods = "time: mean within months time: mean over years" ;
		alb_sfc:time_avg_info = "average_T1,average_T2,average_DT" ;
	double average_DT(time) ;
		average_DT:long_name = "Length of average period" ;
		average_DT:units = "days" ;
	double average_T1(time) ;
		average_T1:long_name = "Start time for average period" ;
		average_T1:units = "days since 1979-01-01 00:00:00" ;
	double average_T2(time) ;
		average_T2:long_name = "End time for average period" ;
		average_T2:units = "days since 1979-01-01 00:00:00" ;
	double climatology_bounds(time, bnds) ;
	double lat(lat) ;
		lat:standard_name = "latitude" ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_N" ;
		lat:axis = "Y" ;
		lat:bounds = "lat_bnds" ;
	double lat_bnds(lat, bnds) ;
	double lon(lon) ;
		lon:standard_name = "longitude" ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_E" ;
		lon:axis = "X" ;
		lon:bounds = "lon_bnds" ;
	double lon_bnds(lon, bnds) ;
	double time(time) ;
		time:standard_name = "time" ;
		time:long_name = "time" ;
		time:climatology = "climatology_bounds" ;
		time:units = "days since 1979-01-01 00:00:00" ;
		time:calendar = "standard" ;
		time:axis = "T" ;

// global attributes:
		:CDI = "Climate Data Interface version 2.4.4 (https://mpimet.mpg.de/cdi)" ;
		:Conventions = "CF-1.6" ;
		:title = "c96L65_am5f9d8r0_amip" ;
		:associated_files = "area: 19800101.grid_spec.nc" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
		:code_release_version = "2024.05" ;
		:git_hash = "5d306c05d9fe755cab04eedc8fd3de0d3c8355a0" ;
		:creationtime = "Mon Aug 25 14:09:46 2025" ;
		:hostname = "pp050" ;
		:history = "Mon Aug 25 13:32:16 2025: ncks -d lat,,,10 -d lon,,,10 atmos.1980-1981.alb_sfc.03.nc reduced/atmos.1980-1981.alb_sfc.03.nc\n",
			"Mon Aug 25 14:40:04 2025: cdo -O -s -select,month=3 merged_output.nc monthly_nc_files/all_years.3.nc\n",
			"Mon Aug 25 14:40:01 2025: cdo -O -s -mergetime /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/shards/ts/regrid-xy/180_288.conserve_order2/atmos_month/P1M/P1Y/atmos_month.198001-198012.alb_sfc.nc /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/shards/ts/regrid-xy/180_288.conserve_order2/atmos_month/P1M/P1Y/atmos_month.198101-198112.alb_sfc.nc merged_output.nc\n",
			"Mon Aug 25 14:12:17 2025: cdo --history splitname 19800101.atmos_month.nc /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/cycle/19800101T0000Z/split/regrid-xy/180_288.conserve_order2/19800101.atmos_month.\n",
			"fregrid --debug --standard_dimension --input_mosaic C96_mosaic.nc --input_dir /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/cycle/19800101T0000Z/history/native --input_file 19800101.atmos_month --associated_file_dir /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/cycle/19800101T0000Z/history/native --interp_method conserve_order2 --remap_file fregrid_remap_file_288_by_180.nc --nlon 288 --nlat 180 --scalar_field (**please see the field list in this file**) --output_file 19800101.atmos_month.nc" ;
		:CDO = "Climate Data Operators version 2.4.4 (https://mpimet.mpg.de/cdo)" ;
		:comment = "FMS time averaging, version 3.0, precision=double" ;
		:NCO = "netCDF Operators version 5.2.4 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco, Citation = 10.1016/j.envsoft.2008.03.004)" ;
data:

 alb_sfc =
  47.43417, 47.43417, 47.43417, 47.43417, 47.43417, 47.43417, 47.43417, 
    47.59669, 47.59669, 47.59669, 47.59669, 47.59669, 47.59669, 47.59669, 
    47.61921, 47.61921, 47.61921, 47.61921, 47.61921, 47.61921, 47.61921, 
    47.46468, 47.46468, 47.46468, 47.46468, 47.46468, 47.46468, 47.46468, 
    47.43417,
  43.5118, 43.41313, 43.37036, 43.4233, 43.34738, 43.27142, 43.21986, 
    43.16364, 43.16291, 43.08019, 43.10503, 43.17345, 43.27472, 43.73903, 
    43.99079, 44.35541, 44.28147, 44.11162, 43.8757, 44.02043, 44.13496, 
    43.95731, 43.94007, 44.31731, 44.26321, 43.96834, 44.14059, 43.97385, 
    43.53454,
  26.7236, 16.41761, 7.966278, 35.78895, 41.79649, 41.75282, 43.79784, 
    41.65121, 41.46552, 41.64182, 41.6374, 41.627, 41.87435, 10.6217, 
    4.606793, 4.578598, 4.524013, 4.308167, 4.425159, 5.285616, 8.286122, 
    11.52913, 33.27543, 39.1891, 43.22599, 22.12953, 4.541925, 4.264524, 
    14.46985,
  4.410142, 4.518198, 4.669731, 4.199453, 4.158391, 4.037917, 3.989242, 
    3.818337, 3.904713, 4.22206, 4.473274, 4.074083, 3.690371, 3.926199, 
    4.158232, 4.037803, 3.922801, 3.802495, 3.853079, 4.105456, 4.215384, 
    4.275981, 4.060549, 4.061829, 3.773694, 3.679171, 3.764771, 3.856111, 
    4.230276,
  3.639926, 3.829758, 3.834495, 3.892229, 3.764282, 3.857962, 3.818746, 
    3.830472, 3.901062, 3.877645, 3.794396, 3.887465, 3.775724, 3.71369, 
    3.934788, 3.721147, 3.769408, 3.764766, 3.870242, 3.926732, 3.939211, 
    4.013168, 3.882056, 7.232795, 4.353914, 3.982586, 3.670774, 3.511096, 
    3.600022,
  3.641325, 3.7892, 3.976749, 3.814518, 3.792114, 3.882679, 3.715187, 
    3.557861, 3.673491, 3.769892, 3.782632, 3.852752, 3.977583, 3.584382, 
    8.780268, 3.861363, 3.809021, 3.78386, 3.718145, 3.767006, 3.676623, 
    3.580771, 3.905207, 8.803297, 4.328143, 3.777349, 3.70266, 3.604915, 
    3.652615,
  3.74546, 3.983719, 11.5186, 3.707229, 3.711147, 3.527759, 3.522706, 
    3.630677, 3.642393, 3.822381, 9.471046, 14.07704, 9.842587, 3.749553, 
    3.701789, 3.781526, 3.580466, 3.497125, 3.467586, 3.74583, 3.706888, 
    3.886431, 3.735367, 4.319248, 8.952963, 3.731999, 3.575386, 3.728696, 
    3.899436,
  3.50742, 9.670603, 11.71459, 3.609141, 3.36628, 3.433098, 3.624848, 
    3.502537, 3.482238, 3.632973, 12.03836, 11.295, 3.631648, 3.437924, 
    3.306992, 3.447149, 3.424329, 3.450294, 3.522445, 3.708003, 3.617065, 
    3.817372, 3.467546, 3.322013, 8.883327, 8.742012, 3.49592, 3.572309, 
    3.86863,
  3.321374, 6.202157, 8.453776, 8.980318, 3.309302, 3.440564, 3.390748, 
    3.255559, 3.234333, 3.279746, 4.651907, 3.258299, 4.239234, 3.25945, 
    3.327178, 3.426277, 3.244133, 3.416974, 3.374014, 3.537418, 3.556986, 
    3.694318, 3.44858, 8.366242, 8.293596, 8.593252, 3.467623, 3.540089, 
    3.613626,
  3.036963, 8.607241, 8.298052, 9.843227, 3.318223, 3.289852, 3.23226, 
    3.240616, 8.473204, 8.144125, 3.288433, 3.230237, 3.280407, 3.248574, 
    3.241026, 3.32691, 3.378343, 3.641906, 3.528069, 3.57112, 3.4649, 
    3.46364, 3.23815, 8.437507, 8.380023, 3.148606, 3.217084, 3.254031, 
    3.045958,
  9.98345, 10.37729, 10.50356, 9.571718, 14.96064, 3.358743, 5.22686, 
    3.389226, 3.681864, 3.390008, 4.284321, 3.42228, 3.335911, 3.433167, 
    3.410778, 3.364733, 3.463377, 3.435695, 3.362568, 3.423584, 3.275271, 
    3.405106, 8.768454, 7.381003, 3.384129, 3.268433, 3.178878, 3.176008, 
    8.986258,
  17.55748, 20.01732, 22.10609, 3.499441, 22.11784, 3.705402, 10.63408, 
    3.748679, 9.675865, 3.28196, 3.534585, 3.588541, 3.653285, 3.752709, 
    3.74703, 3.717777, 3.606305, 3.748666, 3.402335, 3.480055, 3.695015, 
    6.224007, 3.706169, 4.433354, 3.690275, 3.629511, 3.392702, 3.345877, 
    22.87215,
  22.73115, 18.50284, 19.72854, 18.40043, 12.29249, 13.97918, 12.22011, 
    25.39712, 9.471245, 10.2568, 3.425316, 3.529753, 3.550213, 3.490078, 
    3.517384, 3.513832, 3.588286, 3.55178, 3.560022, 3.891266, 12.58634, 
    11.28694, 9.027315, 3.553791, 3.525265, 3.598995, 3.457394, 3.584906, 
    11.05108,
  6.862658, 4.24641, 6.099311, 21.99548, 1.907975, 13.77354, 27.28526, 
    14.25956, 12.25579, 9.852301, 9.669758, 3.805349, 3.762033, 3.801228, 
    3.806376, 3.713762, 3.686108, 3.516, 3.564968, 11.78414, 21.65573, 
    15.0246, 15.5598, 4.605766, 3.59783, 3.544308, 3.631895, 3.681892, 
    5.572101,
  5.710312, 14.32593, 15.17859, 14.85682, 20.07127, 32.8579, 11.70861, 
    34.25611, 14.14958, 7.993164, 7.885602, 23.5869, 18.52461, 3.999243, 
    4.003437, 4.027384, 3.780671, 3.724721, 3.877232, 26.05449, 15.99785, 
    28.24509, 27.0799, 31.89691, 18.29533, 3.741544, 3.660026, 3.855, 3.832637,
  4.235409, 20.35779, 19.5347, 27.41287, 27.35172, 26.15433, 27.5785, 
    28.89903, 24.97812, 25.73755, 23.16117, 37.04792, 38.28573, 34.68979, 
    4.64973, 40.23306, 32.64667, 15.88013, 35.85291, 25.77517, 27.16916, 
    37.32644, 45.4029, 38.35985, 3.857375, 12.98213, 4.63226, 4.31885, 
    4.353382,
  4.95221, 4.941158, 25.73737, 4.007228, 29.15009, 42.70691, 37.38919, 
    37.44806, 37.39031, 37.21919, 26.11864, 22.41674, 37.10708, 43.86335, 
    43.59488, 44.62059, 39.81145, 39.8255, 43.22331, 43.07043, 36.97938, 
    41.05639, 38.20845, 37.84148, 44.72926, 37.89758, 37.7412, 41.86723, 
    4.748385,
  40.04799, 41.25996, 39.19645, 41.5205, 40.40662, 40.06661, 41.54838, 
    41.28444, 41.52411, 41.66435, 41.79435, 41.83583, 41.79807, 41.85226, 
    41.77138, 41.59155, 41.57026, 41.60006, 41.64032, 41.6435, 41.67337, 
    39.35219, 36.38178, 37.18844, 35.34088, 35.16234, 35.18691, 35.81013, 
    41.71321 ;

 average_DT = 730 ;

 average_T1 = 75.5 ;

 average_T2 = 805.5 ;

 climatology_bounds =
  75.5, 805.5 ;

 lat = -89.5, -79.5, -69.5, -59.5, -49.5, -39.5, -29.5, -19.5, -9.5, 0.5, 
    10.5, 20.5, 30.5, 40.5, 50.5, 60.5, 70.5, 80.5 ;

 lat_bnds =
  -90, -89,
  -80, -79,
  -70, -69,
  -60, -59,
  -50, -49,
  -40, -39,
  -30, -29,
  -20, -19,
  -10, -9,
  0, 1,
  10, 11,
  20, 21,
  30, 31,
  40, 41,
  50, 51,
  60, 61,
  70, 71,
  80, 81 ;

 lon = 0.625, 13.125, 25.625, 38.125, 50.625, 63.125, 75.625, 88.125, 
    100.625, 113.125, 125.625, 138.125, 150.625, 163.125, 175.625, 188.125, 
    200.625, 213.125, 225.625, 238.125, 250.625, 263.125, 275.625, 288.125, 
    300.625, 313.125, 325.625, 338.125, 350.625 ;

 lon_bnds =
  0, 1.25,
  12.5, 13.75,
  25, 26.25,
  37.5, 38.75,
  50, 51.25,
  62.5, 63.75,
  75, 76.25,
  87.5, 88.75,
  100, 101.25,
  112.5, 113.75,
  125, 126.25,
  137.5, 138.75,
  150, 151.25,
  162.5, 163.75,
  175, 176.25,
  187.5, 188.75,
  200, 201.25,
  212.5, 213.75,
  225, 226.25,
  237.5, 238.75,
  250, 251.25,
  262.5, 263.75,
  275, 276.25,
  287.5, 288.75,
  300, 301.25,
  312.5, 313.75,
  325, 326.25,
  337.5, 338.75,
  350, 351.25 ;

 time = 0 ;
}
