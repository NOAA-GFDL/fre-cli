netcdf atmos.1980-1981.alb_sfc.06 {
dimensions:
	time = UNLIMITED ; // (1 currently)
	lat = 18 ;
	lon = 29 ;
	bnds = 2 ;
variables:
	float alb_sfc(time, lat, lon) ;
		alb_sfc:long_name = "Surface Albedo for  Flux" ;
		alb_sfc:units = "percent" ;
		alb_sfc:_FillValue = 1.e+20f ;
		alb_sfc:missing_value = 1.e+20f ;
		alb_sfc:cell_measures = "area: area" ;
		alb_sfc:interp_method = "conserve_order1" ;
		alb_sfc:cell_methods = "time: mean within months time: mean over years" ;
		alb_sfc:time_avg_info = "average_T1,average_T2,average_DT" ;
	double average_DT(time) ;
		average_DT:long_name = "Length of average period" ;
		average_DT:units = "days" ;
	double average_T1(time) ;
		average_T1:long_name = "Start time for average period" ;
		average_T1:units = "days since 1979-01-01 00:00:00" ;
	double average_T2(time) ;
		average_T2:long_name = "End time for average period" ;
		average_T2:units = "days since 1979-01-01 00:00:00" ;
	double climatology_bounds(time, bnds) ;
	double lat(lat) ;
		lat:standard_name = "latitude" ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_N" ;
		lat:axis = "Y" ;
		lat:bounds = "lat_bnds" ;
	double lat_bnds(lat, bnds) ;
	double lon(lon) ;
		lon:standard_name = "longitude" ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_E" ;
		lon:axis = "X" ;
		lon:bounds = "lon_bnds" ;
	double lon_bnds(lon, bnds) ;
	double time(time) ;
		time:standard_name = "time" ;
		time:long_name = "time" ;
		time:climatology = "climatology_bounds" ;
		time:units = "days since 1979-01-01 00:00:00" ;
		time:calendar = "standard" ;
		time:axis = "T" ;

// global attributes:
		:CDI = "Climate Data Interface version 2.4.4 (https://mpimet.mpg.de/cdi)" ;
		:Conventions = "CF-1.6" ;
		:title = "c96L65_am5f9d8r0_amip" ;
		:associated_files = "area: 19800101.grid_spec.nc" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
		:code_release_version = "2024.05" ;
		:git_hash = "5d306c05d9fe755cab04eedc8fd3de0d3c8355a0" ;
		:creationtime = "Mon Aug 25 14:09:46 2025" ;
		:hostname = "pp050" ;
		:history = "Mon Aug 25 13:32:19 2025: ncks -d lat,,,10 -d lon,,,10 atmos.1980-1981.alb_sfc.06.nc reduced/atmos.1980-1981.alb_sfc.06.nc\n",
			"Mon Aug 25 14:40:06 2025: cdo -O -s -select,month=6 merged_output.nc monthly_nc_files/all_years.6.nc\n",
			"Mon Aug 25 14:40:01 2025: cdo -O -s -mergetime /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/shards/ts/regrid-xy/180_288.conserve_order2/atmos_month/P1M/P1Y/atmos_month.198001-198012.alb_sfc.nc /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/shards/ts/regrid-xy/180_288.conserve_order2/atmos_month/P1M/P1Y/atmos_month.198101-198112.alb_sfc.nc merged_output.nc\n",
			"Mon Aug 25 14:12:17 2025: cdo --history splitname 19800101.atmos_month.nc /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/cycle/19800101T0000Z/split/regrid-xy/180_288.conserve_order2/19800101.atmos_month.\n",
			"fregrid --debug --standard_dimension --input_mosaic C96_mosaic.nc --input_dir /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/cycle/19800101T0000Z/history/native --input_file 19800101.atmos_month --associated_file_dir /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/cycle/19800101T0000Z/history/native --interp_method conserve_order2 --remap_file fregrid_remap_file_288_by_180.nc --nlon 288 --nlat 180 --scalar_field (**please see the field list in this file**) --output_file 19800101.atmos_month.nc" ;
		:CDO = "Climate Data Operators version 2.4.4 (https://mpimet.mpg.de/cdo)" ;
		:comment = "FMS time averaging, version 3.0, precision=double" ;
		:NCO = "netCDF Operators version 5.2.4 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco, Citation = 10.1016/j.envsoft.2008.03.004)" ;
data:

 alb_sfc =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  6.10913, 2.472299, 2.821715, 2.640081, 2.49383, 2.439744, 2.064852, 
    2.271052, 2.550112, 2.157125, 2.364811, 2.38126, 2.13951, 2.103727, 
    2.316686, 2.330638, 2.17626, 2.630388, 2.752551, 2.662262, 2.696767, 
    2.792917, 2.893465, 2.750311, 2.416049, 12.22941, 15.65005, 10.34081, 
    13.9831,
  3.227399, 3.566913, 3.501629, 3.672955, 3.543805, 3.578784, 3.365438, 
    3.531744, 3.62255, 3.486609, 3.486244, 3.616765, 3.598236, 3.408287, 
    3.211436, 3.196608, 3.135719, 3.021747, 3.144073, 3.177851, 3.407255, 
    3.508275, 3.624202, 7.784444, 4.128461, 3.603603, 2.985872, 3.295046, 
    3.35557,
  3.882885, 3.998829, 3.78594, 3.958253, 3.573961, 3.819581, 4.017222, 
    3.588875, 3.628383, 4.052907, 3.963184, 3.756925, 4.385285, 4.080914, 
    10.40794, 4.140424, 3.815361, 3.643842, 3.755473, 3.643792, 3.513572, 
    3.693882, 3.850002, 9.394314, 4.243852, 3.859491, 3.620617, 3.699072, 
    3.843531,
  3.936741, 4.360675, 11.45523, 4.24957, 3.956027, 3.867745, 4.202823, 
    3.977661, 4.262262, 4.388114, 8.481571, 12.33008, 9.58466, 4.193267, 
    3.96261, 3.976026, 3.932655, 3.925729, 3.634832, 3.57807, 3.766159, 
    4.081422, 3.855513, 4.145562, 8.333965, 3.768728, 4.045858, 4.185052, 
    4.097891,
  3.549889, 9.438309, 9.558647, 3.902886, 4.081747, 4.242013, 3.880852, 
    3.978007, 3.843688, 4.178564, 11.46663, 11.92268, 3.910018, 3.888362, 
    3.767899, 3.632597, 3.831578, 3.711967, 3.842808, 3.871082, 4.120521, 
    3.745393, 3.686062, 3.9026, 8.390615, 8.940468, 3.915594, 3.801316, 
    3.691058,
  3.491963, 6.487567, 9.229486, 9.060808, 3.634311, 3.630728, 3.595816, 
    3.578713, 3.30456, 3.750729, 4.638881, 3.677724, 4.266951, 3.472409, 
    3.426909, 3.490531, 3.751797, 3.710634, 4.114725, 3.879488, 3.933003, 
    3.565532, 3.334886, 8.584091, 8.868982, 9.069365, 3.779548, 4.025764, 
    3.455439,
  3.217942, 8.751482, 8.470738, 10.12177, 3.573646, 3.424278, 3.224331, 
    3.285343, 8.661646, 8.59764, 3.472167, 3.371392, 3.352608, 3.486397, 
    3.448731, 3.553501, 3.595276, 3.751022, 3.68049, 3.796342, 3.646607, 
    3.633111, 3.294773, 8.281111, 8.507886, 3.549616, 3.552839, 3.471088, 
    3.308708,
  9.806553, 10.2914, 10.54464, 10.00444, 15.20477, 3.351101, 5.060882, 
    3.055056, 3.557211, 3.206537, 4.279098, 3.329697, 3.252438, 3.378843, 
    3.510272, 3.442339, 3.289331, 3.675989, 3.370578, 3.524721, 3.499994, 
    3.34456, 8.99514, 7.75107, 3.391173, 3.243975, 3.40188, 3.11311, 8.907709,
  19.44018, 21.78009, 23.58921, 3.558252, 24.28801, 3.184416, 11.16966, 
    3.207238, 9.231133, 3.395174, 3.477529, 3.468552, 3.864067, 3.771709, 
    3.686505, 3.949712, 3.816407, 3.873244, 3.670712, 3.745437, 3.720231, 
    6.931602, 3.477043, 4.056266, 3.800932, 3.669249, 3.650343, 3.469378, 
    24.63101,
  25.87786, 21.85138, 22.7486, 20.91747, 13.92895, 15.91502, 13.16095, 
    10.83539, 8.459892, 11.03952, 3.625111, 3.643754, 3.634988, 3.747644, 
    3.687321, 3.762459, 4.016238, 3.95763, 3.847518, 3.838506, 11.63663, 
    12.42416, 9.90737, 3.742181, 3.645398, 4.102548, 3.92161, 3.961878, 
    11.98179,
  8.264321, 4.211575, 6.782467, 11.05632, 2.353259, 16.72853, 9.819856, 
    17.30908, 14.99815, 11.67514, 8.188787, 3.989883, 3.779939, 3.841346, 
    3.915041, 3.75757, 3.873854, 3.862718, 3.849194, 13.64296, 12.80821, 
    14.70553, 14.10074, 4.936634, 3.882792, 4.015848, 4.066926, 3.992003, 
    5.436654,
  6.884028, 14.11233, 15.28396, 16.58824, 15.39645, 13.47851, 9.54277, 
    12.88732, 8.883905, 8.166033, 7.933316, 7.611247, 4.264384, 4.285189, 
    4.124409, 4.230452, 4.181227, 4.26473, 4.434647, 10.29861, 11.61545, 
    11.33044, 8.018856, 7.64455, 6.040251, 4.502963, 4.432994, 4.406594, 
    4.685765,
  5.425042, 9.156954, 10.88309, 8.931665, 9.364049, 9.234555, 9.374854, 
    9.407482, 9.809399, 9.519079, 9.161164, 17.04486, 25.16867, 8.731203, 
    5.489271, 5.986596, 12.17577, 17.24231, 14.02074, 9.358944, 8.427878, 
    21.62209, 45.21049, 23.24934, 5.620914, 10.04432, 5.119761, 5.17194, 
    5.255353,
  6.312997, 7.03748, 12.17826, 7.056308, 10.77177, 59.7938, 43.33971, 
    44.12855, 35.48384, 34.78027, 17.22225, 15.04599, 31.56168, 58.9479, 
    58.23514, 57.21755, 35.97139, 34.61705, 52.02171, 36.98507, 32.3983, 
    49.13464, 36.09002, 53.41291, 37.01002, 68.90591, 74.33415, 39.78078, 
    6.757262,
  60.45778, 58.45857, 57.89606, 60.52255, 48.92993, 59.73045, 60.41017, 
    59.18221, 60.1264, 60.40049, 60.53784, 60.60666, 60.55488, 60.59946, 
    60.51875, 60.42652, 60.39294, 60.5252, 60.69265, 60.43377, 60.52378, 
    56.54607, 58.05941, 64.68721, 66.17075, 69.03517, 69.42293, 64.27591, 
    60.87678 ;

 average_DT = 730 ;

 average_T1 = 167 ;

 average_T2 = 897 ;

 climatology_bounds =
  167, 897 ;

 lat = -89.5, -79.5, -69.5, -59.5, -49.5, -39.5, -29.5, -19.5, -9.5, 0.5, 
    10.5, 20.5, 30.5, 40.5, 50.5, 60.5, 70.5, 80.5 ;

 lat_bnds =
  -90, -89,
  -80, -79,
  -70, -69,
  -60, -59,
  -50, -49,
  -40, -39,
  -30, -29,
  -20, -19,
  -10, -9,
  0, 1,
  10, 11,
  20, 21,
  30, 31,
  40, 41,
  50, 51,
  60, 61,
  70, 71,
  80, 81 ;

 lon = 0.625, 13.125, 25.625, 38.125, 50.625, 63.125, 75.625, 88.125, 
    100.625, 113.125, 125.625, 138.125, 150.625, 163.125, 175.625, 188.125, 
    200.625, 213.125, 225.625, 238.125, 250.625, 263.125, 275.625, 288.125, 
    300.625, 313.125, 325.625, 338.125, 350.625 ;

 lon_bnds =
  0, 1.25,
  12.5, 13.75,
  25, 26.25,
  37.5, 38.75,
  50, 51.25,
  62.5, 63.75,
  75, 76.25,
  87.5, 88.75,
  100, 101.25,
  112.5, 113.75,
  125, 126.25,
  137.5, 138.75,
  150, 151.25,
  162.5, 163.75,
  175, 176.25,
  187.5, 188.75,
  200, 201.25,
  212.5, 213.75,
  225, 226.25,
  237.5, 238.75,
  250, 251.25,
  262.5, 263.75,
  275, 276.25,
  287.5, 288.75,
  300, 301.25,
  312.5, 313.75,
  325, 326.25,
  337.5, 338.75,
  350, 351.25 ;

 time = 0 ;
}
